VERSION 5.7 ;
NOWIREEXTENSIONATPIN ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
MACRO tdc_inline_3
  CLASS BLOCK ;
  FOREIGN tdc_inline_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 460.000 BY 408.000 ;
  PIN bus_in[0]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 2.850 404.000 3.130 408.000 ;
    END
  END bus_in[0]
  PIN bus_in[10]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 121.990 404.000 122.270 408.000 ;
    END
  END bus_in[10]
  PIN bus_in[11]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 133.950 404.000 134.230 408.000 ;
    END
  END bus_in[11]
  PIN bus_in[12]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 145.910 404.000 146.190 408.000 ;
    END
  END bus_in[12]
  PIN bus_in[13]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 157.870 404.000 158.150 408.000 ;
    END
  END bus_in[13]
  PIN bus_in[14]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 169.830 404.000 170.110 408.000 ;
    END
  END bus_in[14]
  PIN bus_in[15]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 181.790 404.000 182.070 408.000 ;
    END
  END bus_in[15]
  PIN bus_in[16]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 193.750 404.000 194.030 408.000 ;
    END
  END bus_in[16]
  PIN bus_in[17]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 205.710 404.000 205.990 408.000 ;
    END
  END bus_in[17]
  PIN bus_in[18]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 217.670 404.000 217.950 408.000 ;
    END
  END bus_in[18]
  PIN bus_in[19]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 229.630 404.000 229.910 408.000 ;
    END
  END bus_in[19]
  PIN bus_in[1]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 14.350 404.000 14.630 408.000 ;
    END
  END bus_in[1]
  PIN bus_in[20]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 241.590 404.000 241.870 408.000 ;
    END
  END bus_in[20]
  PIN bus_in[21]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 253.550 404.000 253.830 408.000 ;
    END
  END bus_in[21]
  PIN bus_in[22]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 265.510 404.000 265.790 408.000 ;
    END
  END bus_in[22]
  PIN bus_in[23]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 277.470 404.000 277.750 408.000 ;
    END
  END bus_in[23]
  PIN bus_in[24]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 289.430 404.000 289.710 408.000 ;
    END
  END bus_in[24]
  PIN bus_in[25]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 301.390 404.000 301.670 408.000 ;
    END
  END bus_in[25]
  PIN bus_in[26]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 313.350 404.000 313.630 408.000 ;
    END
  END bus_in[26]
  PIN bus_in[27]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 325.310 404.000 325.590 408.000 ;
    END
  END bus_in[27]
  PIN bus_in[28]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 337.270 404.000 337.550 408.000 ;
    END
  END bus_in[28]
  PIN bus_in[29]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 349.230 404.000 349.510 408.000 ;
    END
  END bus_in[29]
  PIN bus_in[2]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 26.310 404.000 26.590 408.000 ;
    END
  END bus_in[2]
  PIN bus_in[30]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 361.190 404.000 361.470 408.000 ;
    END
  END bus_in[30]
  PIN bus_in[31]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 373.150 404.000 373.430 408.000 ;
    END
  END bus_in[31]
  PIN bus_in[32]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 385.110 404.000 385.390 408.000 ;
    END
  END bus_in[32]
  PIN bus_in[33]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 397.070 404.000 397.350 408.000 ;
    END
  END bus_in[33]
  PIN bus_in[34]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 409.030 404.000 409.310 408.000 ;
    END
  END bus_in[34]
  PIN bus_in[35]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 420.990 404.000 421.270 408.000 ;
    END
  END bus_in[35]
  PIN bus_in[36]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 426.970 404.000 427.250 408.000 ;
    END
  END bus_in[36]
  PIN bus_in[37]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 432.950 404.000 433.230 408.000 ;
    END
  END bus_in[37]
  PIN bus_in[38]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 438.930 404.000 439.210 408.000 ;
    END
  END bus_in[38]
  PIN bus_in[39]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 444.910 404.000 445.190 408.000 ;
    END
  END bus_in[39]
  PIN bus_in[3]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 38.270 404.000 38.550 408.000 ;
    END
  END bus_in[3]
  PIN bus_in[40]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 450.890 404.000 451.170 408.000 ;
    END
  END bus_in[40]
  PIN bus_in[41]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 456.870 404.000 457.150 408.000 ;
    END
  END bus_in[41]
  PIN bus_in[4]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 50.230 404.000 50.510 408.000 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 62.190 404.000 62.470 408.000 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 74.150 404.000 74.430 408.000 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 86.110 404.000 86.390 408.000 ;
    END
  END bus_in[7]
  PIN bus_in[8]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 98.070 404.000 98.350 408.000 ;
    END
  END bus_in[8]
  PIN bus_in[9]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 110.030 404.000 110.310 408.000 ;
    END
  END bus_in[9]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 8.370 404.000 8.650 408.000 ;
    END
  END bus_out[0]
  PIN bus_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 127.970 404.000 128.250 408.000 ;
    END
  END bus_out[10]
  PIN bus_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 139.930 404.000 140.210 408.000 ;
    END
  END bus_out[11]
  PIN bus_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 151.890 404.000 152.170 408.000 ;
    END
  END bus_out[12]
  PIN bus_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 163.850 404.000 164.130 408.000 ;
    END
  END bus_out[13]
  PIN bus_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 175.810 404.000 176.090 408.000 ;
    END
  END bus_out[14]
  PIN bus_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 187.770 404.000 188.050 408.000 ;
    END
  END bus_out[15]
  PIN bus_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 199.730 404.000 200.010 408.000 ;
    END
  END bus_out[16]
  PIN bus_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 211.690 404.000 211.970 408.000 ;
    END
  END bus_out[17]
  PIN bus_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 223.650 404.000 223.930 408.000 ;
    END
  END bus_out[18]
  PIN bus_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 235.610 404.000 235.890 408.000 ;
    END
  END bus_out[19]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 20.330 404.000 20.610 408.000 ;
    END
  END bus_out[1]
  PIN bus_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 247.570 404.000 247.850 408.000 ;
    END
  END bus_out[20]
  PIN bus_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 259.530 404.000 259.810 408.000 ;
    END
  END bus_out[21]
  PIN bus_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 271.490 404.000 271.770 408.000 ;
    END
  END bus_out[22]
  PIN bus_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 283.450 404.000 283.730 408.000 ;
    END
  END bus_out[23]
  PIN bus_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 295.410 404.000 295.690 408.000 ;
    END
  END bus_out[24]
  PIN bus_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 307.370 404.000 307.650 408.000 ;
    END
  END bus_out[25]
  PIN bus_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 319.330 404.000 319.610 408.000 ;
    END
  END bus_out[26]
  PIN bus_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 331.290 404.000 331.570 408.000 ;
    END
  END bus_out[27]
  PIN bus_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 343.250 404.000 343.530 408.000 ;
    END
  END bus_out[28]
  PIN bus_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 355.210 404.000 355.490 408.000 ;
    END
  END bus_out[29]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 32.290 404.000 32.570 408.000 ;
    END
  END bus_out[2]
  PIN bus_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 367.170 404.000 367.450 408.000 ;
    END
  END bus_out[30]
  PIN bus_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 379.130 404.000 379.410 408.000 ;
    END
  END bus_out[31]
  PIN bus_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 391.090 404.000 391.370 408.000 ;
    END
  END bus_out[32]
  PIN bus_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 403.050 404.000 403.330 408.000 ;
    END
  END bus_out[33]
  PIN bus_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 415.010 404.000 415.290 408.000 ;
    END
  END bus_out[34]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 44.250 404.000 44.530 408.000 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 56.210 404.000 56.490 408.000 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 68.170 404.000 68.450 408.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 80.130 404.000 80.410 408.000 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 92.090 404.000 92.370 408.000 ;
    END
  END bus_out[7]
  PIN bus_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 104.050 404.000 104.330 408.000 ;
    END
  END bus_out[8]
  PIN bus_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 116.010 404.000 116.290 408.000 ;
    END
  END bus_out[9]
  PIN clk_i
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 102.040 460.000 102.640 ;
    END
  END clk_i
  PIN inp_i
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 0.000 204.040 4.000 204.640 ;
    END
  END inp_i
  PIN rst_n_i
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 306.040 460.000 306.640 ;
    END
  END rst_n_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT 
      LAYER met4 ;
      RECT 174.64 10.64 176.24 397.36 ;
      RECT 328.24 10.64 329.84 397.36 ;
      RECT 21.040 10.640 22.640 397.360 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT 
      LAYER met4 ;
      RECT 251.44 10.64 253.04 397.36 ;
      RECT 405.04 10.64 406.64 397.36 ;
      RECT 97.840 10.640 99.440 397.360 ;
    END
  END VGND
  OBS 
    LAYER li1 ;
    RECT 5.520 10.795 454.480 397.205 ;
    LAYER met1 ;
    RECT 5.520 10.640 457.170 397.360 ;
    LAYER met2 ;
    RECT 3.410 403.720 8.090 404.000 ;
    RECT 8.930 403.720 14.070 404.000 ;
    RECT 14.910 403.720 20.050 404.000 ;
    RECT 20.890 403.720 26.030 404.000 ;
    RECT 26.870 403.720 32.010 404.000 ;
    RECT 32.850 403.720 37.990 404.000 ;
    RECT 38.830 403.720 43.970 404.000 ;
    RECT 44.810 403.720 49.950 404.000 ;
    RECT 50.790 403.720 55.930 404.000 ;
    RECT 56.770 403.720 61.910 404.000 ;
    RECT 62.750 403.720 67.890 404.000 ;
    RECT 68.730 403.720 73.870 404.000 ;
    RECT 74.710 403.720 79.850 404.000 ;
    RECT 80.690 403.720 85.830 404.000 ;
    RECT 86.670 403.720 91.810 404.000 ;
    RECT 92.650 403.720 97.790 404.000 ;
    RECT 98.630 403.720 103.770 404.000 ;
    RECT 104.610 403.720 109.750 404.000 ;
    RECT 110.590 403.720 115.730 404.000 ;
    RECT 116.570 403.720 121.710 404.000 ;
    RECT 122.550 403.720 127.690 404.000 ;
    RECT 128.530 403.720 133.670 404.000 ;
    RECT 134.510 403.720 139.650 404.000 ;
    RECT 140.490 403.720 145.630 404.000 ;
    RECT 146.470 403.720 151.610 404.000 ;
    RECT 152.450 403.720 157.590 404.000 ;
    RECT 158.430 403.720 163.570 404.000 ;
    RECT 164.410 403.720 169.550 404.000 ;
    RECT 170.390 403.720 175.530 404.000 ;
    RECT 176.370 403.720 181.510 404.000 ;
    RECT 182.350 403.720 187.490 404.000 ;
    RECT 188.330 403.720 193.470 404.000 ;
    RECT 194.310 403.720 199.450 404.000 ;
    RECT 200.290 403.720 205.430 404.000 ;
    RECT 206.270 403.720 211.410 404.000 ;
    RECT 212.250 403.720 217.390 404.000 ;
    RECT 218.230 403.720 223.370 404.000 ;
    RECT 224.210 403.720 229.350 404.000 ;
    RECT 230.190 403.720 235.330 404.000 ;
    RECT 236.170 403.720 241.310 404.000 ;
    RECT 242.150 403.720 247.290 404.000 ;
    RECT 248.130 403.720 253.270 404.000 ;
    RECT 254.110 403.720 259.250 404.000 ;
    RECT 260.090 403.720 265.230 404.000 ;
    RECT 266.070 403.720 271.210 404.000 ;
    RECT 272.050 403.720 277.190 404.000 ;
    RECT 278.030 403.720 283.170 404.000 ;
    RECT 284.010 403.720 289.150 404.000 ;
    RECT 289.990 403.720 295.130 404.000 ;
    RECT 295.970 403.720 301.110 404.000 ;
    RECT 301.950 403.720 307.090 404.000 ;
    RECT 307.930 403.720 313.070 404.000 ;
    RECT 313.910 403.720 319.050 404.000 ;
    RECT 319.890 403.720 325.030 404.000 ;
    RECT 325.870 403.720 331.010 404.000 ;
    RECT 331.850 403.720 336.990 404.000 ;
    RECT 337.830 403.720 342.970 404.000 ;
    RECT 343.810 403.720 348.950 404.000 ;
    RECT 349.790 403.720 354.930 404.000 ;
    RECT 355.770 403.720 360.910 404.000 ;
    RECT 361.750 403.720 366.890 404.000 ;
    RECT 367.730 403.720 372.870 404.000 ;
    RECT 373.710 403.720 378.850 404.000 ;
    RECT 379.690 403.720 384.830 404.000 ;
    RECT 385.670 403.720 390.810 404.000 ;
    RECT 391.650 403.720 396.790 404.000 ;
    RECT 397.630 403.720 402.770 404.000 ;
    RECT 403.610 403.720 408.750 404.000 ;
    RECT 409.590 403.720 414.730 404.000 ;
    RECT 415.570 403.720 420.710 404.000 ;
    RECT 421.550 403.720 426.690 404.000 ;
    RECT 427.530 403.720 432.670 404.000 ;
    RECT 433.510 403.720 438.650 404.000 ;
    RECT 439.490 403.720 444.630 404.000 ;
    RECT 445.470 403.720 450.610 404.000 ;
    RECT 451.450 403.720 456.590 404.000 ;
    RECT 2.850 10.640 457.140 403.720 ;
    LAYER met3 ;
    RECT 2.825 307.040 456.000 397.285 ;
    RECT 2.825 305.640 455.600 307.040 ;
    RECT 2.825 205.040 456.000 305.640 ;
    RECT 4.400 203.640 456.000 205.040 ;
    RECT 2.825 103.040 456.000 203.640 ;
    RECT 2.825 101.640 455.600 103.040 ;
    RECT 2.825 10.715 456.000 101.640 ;
    LAYER met4 ;
    RECT 174.640 10.640 406.640 397.360 ;
  END
END tdc_inline_3
END LIBRARY
