VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2902.210 2846.040 2902.530 2846.100 ;
        RECT 2866.000 2845.900 2902.530 2846.040 ;
        RECT 2902.210 2845.840 2902.530 2845.900 ;
      LAYER via ;
        RECT 2902.240 2845.840 2902.500 2846.100 ;
      LAYER met2 ;
        RECT 2902.230 2962.235 2902.510 2962.605 ;
        RECT 2902.300 2846.130 2902.440 2962.235 ;
        RECT 2902.240 2845.810 2902.500 2846.130 ;
      LAYER via2 ;
        RECT 2902.230 2962.280 2902.510 2962.560 ;
      LAYER met3 ;
        RECT 2902.205 2962.570 2902.535 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2902.205 2962.270 2924.800 2962.570 ;
        RECT 2902.205 2962.255 2902.535 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2901.750 2514.880 2902.070 2514.940 ;
        RECT 2866.000 2514.740 2902.070 2514.880 ;
        RECT 2901.750 2514.680 2902.070 2514.740 ;
      LAYER via ;
        RECT 2901.780 2514.680 2902.040 2514.940 ;
      LAYER met2 ;
        RECT 2901.770 3196.835 2902.050 3197.205 ;
        RECT 2901.840 2514.970 2901.980 3196.835 ;
        RECT 2901.780 2514.650 2902.040 2514.970 ;
      LAYER via2 ;
        RECT 2901.770 3196.880 2902.050 3197.160 ;
      LAYER met3 ;
        RECT 2901.745 3197.170 2902.075 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.745 3196.870 2924.800 3197.170 ;
        RECT 2901.745 3196.855 2902.075 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2901.290 417.420 2901.610 417.480 ;
        RECT 2866.000 417.280 2901.610 417.420 ;
        RECT 2901.290 417.220 2901.610 417.280 ;
      LAYER via ;
        RECT 2901.320 417.220 2901.580 417.480 ;
      LAYER met2 ;
        RECT 2901.310 3431.435 2901.590 3431.805 ;
        RECT 2901.380 417.510 2901.520 3431.435 ;
        RECT 2901.320 417.190 2901.580 417.510 ;
      LAYER via2 ;
        RECT 2901.310 3431.480 2901.590 3431.760 ;
      LAYER met3 ;
        RECT 2901.285 3431.770 2901.615 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2901.285 3431.470 2924.800 3431.770 ;
        RECT 2901.285 3431.455 2901.615 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.845 2717.520 3517.600 ;
        RECT 2717.310 3501.475 2717.590 3501.845 ;
      LAYER via2 ;
        RECT 2717.310 3501.520 2717.590 3501.800 ;
      LAYER met3 ;
        RECT 1584.510 3501.810 1584.890 3501.820 ;
        RECT 2717.285 3501.810 2717.615 3501.825 ;
        RECT 1584.510 3501.510 2717.615 3501.810 ;
        RECT 1584.510 3501.500 1584.890 3501.510 ;
        RECT 2717.285 3501.495 2717.615 3501.510 ;
      LAYER via3 ;
        RECT 1584.540 3501.500 1584.860 3501.820 ;
      LAYER met4 ;
        RECT 1584.535 3501.495 1584.865 3501.825 ;
        RECT 1584.550 3466.000 1584.850 3501.495 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3502.525 2392.760 3517.600 ;
        RECT 2392.550 3502.155 2392.830 3502.525 ;
      LAYER via2 ;
        RECT 2392.550 3502.200 2392.830 3502.480 ;
      LAYER met3 ;
        RECT 1586.350 3502.490 1586.730 3502.500 ;
        RECT 2392.525 3502.490 2392.855 3502.505 ;
        RECT 1586.350 3502.190 2392.855 3502.490 ;
        RECT 1586.350 3502.180 1586.730 3502.190 ;
        RECT 2392.525 3502.175 2392.855 3502.190 ;
      LAYER via3 ;
        RECT 1586.380 3502.180 1586.700 3502.500 ;
      LAYER met4 ;
        RECT 1586.375 3502.175 1586.705 3502.505 ;
        RECT 1586.390 3466.000 1586.690 3502.175 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1569.590 3502.240 1569.910 3502.300 ;
        RECT 2068.230 3502.240 2068.550 3502.300 ;
        RECT 1569.590 3502.100 2068.550 3502.240 ;
        RECT 1569.590 3502.040 1569.910 3502.100 ;
        RECT 2068.230 3502.040 2068.550 3502.100 ;
      LAYER via ;
        RECT 1569.620 3502.040 1569.880 3502.300 ;
        RECT 2068.260 3502.040 2068.520 3502.300 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3502.330 2068.460 3517.600 ;
        RECT 1569.620 3502.010 1569.880 3502.330 ;
        RECT 2068.260 3502.010 2068.520 3502.330 ;
        RECT 1569.680 3466.000 1569.820 3502.010 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3503.205 1744.160 3517.600 ;
        RECT 1743.950 3502.835 1744.230 3503.205 ;
      LAYER via2 ;
        RECT 1743.950 3502.880 1744.230 3503.160 ;
      LAYER met3 ;
        RECT 1585.430 3503.170 1585.810 3503.180 ;
        RECT 1743.925 3503.170 1744.255 3503.185 ;
        RECT 1585.430 3502.870 1744.255 3503.170 ;
        RECT 1585.430 3502.860 1585.810 3502.870 ;
        RECT 1743.925 3502.855 1744.255 3502.870 ;
      LAYER via3 ;
        RECT 1585.460 3502.860 1585.780 3503.180 ;
      LAYER met4 ;
        RECT 1585.455 3502.855 1585.785 3503.185 ;
        RECT 1585.470 3466.000 1585.770 3502.855 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1416.410 3491.360 1416.730 3491.420 ;
        RECT 1419.630 3491.360 1419.950 3491.420 ;
        RECT 1416.410 3491.220 1419.950 3491.360 ;
        RECT 1416.410 3491.160 1416.730 3491.220 ;
        RECT 1419.630 3491.160 1419.950 3491.220 ;
        RECT 1415.490 3470.620 1415.810 3470.680 ;
        RECT 1416.410 3470.620 1416.730 3470.680 ;
        RECT 1415.490 3470.480 1416.730 3470.620 ;
        RECT 1415.490 3470.420 1415.810 3470.480 ;
        RECT 1416.410 3470.420 1416.730 3470.480 ;
      LAYER via ;
        RECT 1416.440 3491.160 1416.700 3491.420 ;
        RECT 1419.660 3491.160 1419.920 3491.420 ;
        RECT 1415.520 3470.420 1415.780 3470.680 ;
        RECT 1416.440 3470.420 1416.700 3470.680 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3517.370 1419.400 3517.600 ;
        RECT 1419.260 3517.230 1419.860 3517.370 ;
        RECT 1419.720 3491.450 1419.860 3517.230 ;
        RECT 1416.440 3491.130 1416.700 3491.450 ;
        RECT 1419.660 3491.130 1419.920 3491.450 ;
        RECT 1416.500 3470.710 1416.640 3491.130 ;
        RECT 1415.520 3470.390 1415.780 3470.710 ;
        RECT 1416.440 3470.390 1416.700 3470.710 ;
        RECT 1415.580 3466.000 1415.720 3470.390 ;
    END
  END io_out[19]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3502.240 1095.190 3502.300 ;
        RECT 1412.270 3502.240 1412.590 3502.300 ;
        RECT 1094.870 3502.100 1412.590 3502.240 ;
        RECT 1094.870 3502.040 1095.190 3502.100 ;
        RECT 1412.270 3502.040 1412.590 3502.100 ;
      LAYER via ;
        RECT 1094.900 3502.040 1095.160 3502.300 ;
        RECT 1412.300 3502.040 1412.560 3502.300 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3502.330 1095.100 3517.600 ;
        RECT 1094.900 3502.010 1095.160 3502.330 ;
        RECT 1412.300 3502.010 1412.560 3502.330 ;
        RECT 1412.360 3466.000 1412.500 3502.010 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 693.290 3502.580 693.610 3502.640 ;
        RECT 770.570 3502.580 770.890 3502.640 ;
        RECT 693.290 3502.440 770.890 3502.580 ;
        RECT 693.290 3502.380 693.610 3502.440 ;
        RECT 770.570 3502.380 770.890 3502.440 ;
      LAYER via ;
        RECT 693.320 3502.380 693.580 3502.640 ;
        RECT 770.600 3502.380 770.860 3502.640 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3502.670 770.800 3517.600 ;
        RECT 693.320 3502.350 693.580 3502.670 ;
        RECT 770.600 3502.350 770.860 3502.670 ;
        RECT 693.380 3466.000 693.520 3502.350 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3502.240 446.130 3502.300 ;
        RECT 693.750 3502.240 694.070 3502.300 ;
        RECT 445.810 3502.100 694.070 3502.240 ;
        RECT 445.810 3502.040 446.130 3502.100 ;
        RECT 693.750 3502.040 694.070 3502.100 ;
      LAYER via ;
        RECT 445.840 3502.040 446.100 3502.300 ;
        RECT 693.780 3502.040 694.040 3502.300 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3502.330 446.040 3517.600 ;
        RECT 445.840 3502.010 446.100 3502.330 ;
        RECT 693.780 3502.010 694.040 3502.330 ;
        RECT 693.840 3466.000 693.980 3502.010 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1411.350 3501.560 1411.670 3501.620 ;
        RECT 121.510 3501.420 1411.670 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1411.350 3501.360 1411.670 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1411.380 3501.360 1411.640 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1411.380 3501.330 1411.640 3501.650 ;
        RECT 1411.440 3466.000 1411.580 3501.330 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 17.090 3339.580 54.000 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 3050.040 16.950 3050.100 ;
        RECT 16.630 3049.900 54.000 3050.040 ;
        RECT 16.630 3049.840 16.950 3049.900 ;
      LAYER via ;
        RECT 16.660 3049.840 16.920 3050.100 ;
      LAYER met2 ;
        RECT 16.650 3051.995 16.930 3052.365 ;
        RECT 16.720 3050.130 16.860 3051.995 ;
        RECT 16.660 3049.810 16.920 3050.130 ;
      LAYER via2 ;
        RECT 16.650 3052.040 16.930 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 16.625 3052.330 16.955 3052.345 ;
        RECT -4.800 3052.030 16.955 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 16.625 3052.015 16.955 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 15.710 2760.220 54.000 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
    END
  END io_out[26]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 137.940 17.410 138.000 ;
        RECT 17.090 137.800 54.000 137.940 ;
        RECT 17.090 137.740 17.410 137.800 ;
      LAYER via ;
        RECT 17.120 137.740 17.380 138.000 ;
      LAYER met2 ;
        RECT 17.110 2189.755 17.390 2190.125 ;
        RECT 17.180 138.030 17.320 2189.755 ;
        RECT 17.120 137.710 17.380 138.030 ;
      LAYER via2 ;
        RECT 17.110 2189.800 17.390 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 17.085 2190.090 17.415 2190.105 ;
        RECT -4.800 2189.790 17.415 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 17.085 2189.775 17.415 2189.790 ;
    END
  END io_out[28]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2118.440 17.870 2118.500 ;
        RECT 17.550 2118.300 54.000 2118.440 ;
        RECT 17.550 2118.240 17.870 2118.300 ;
      LAYER via ;
        RECT 17.580 2118.240 17.840 2118.500 ;
      LAYER met2 ;
        RECT 17.570 2118.355 17.850 2118.725 ;
        RECT 17.580 2118.210 17.840 2118.355 ;
      LAYER via2 ;
        RECT 17.570 2118.400 17.850 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 17.545 2118.690 17.875 2118.705 ;
        RECT -4.800 2118.390 17.875 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 17.545 2118.375 17.875 2118.390 ;
    END
  END io_oeb[28]
  PIN analog_io[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2477.480 17.870 2477.540 ;
        RECT 17.550 2477.340 54.000 2477.480 ;
        RECT 17.550 2477.280 17.870 2477.340 ;
      LAYER via ;
        RECT 17.580 2477.280 17.840 2477.540 ;
      LAYER met2 ;
        RECT 17.570 2477.395 17.850 2477.765 ;
        RECT 17.580 2477.250 17.840 2477.395 ;
      LAYER via2 ;
        RECT 17.570 2477.440 17.850 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.545 2477.730 17.875 2477.745 ;
        RECT -4.800 2477.430 17.875 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.545 2477.415 17.875 2477.430 ;
    END
  END io_out[27]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2901.750 1518.000 2902.070 1518.060 ;
        RECT 2866.000 1517.860 2902.070 1518.000 ;
        RECT 2901.750 1517.800 2902.070 1517.860 ;
      LAYER via ;
        RECT 2901.780 1517.800 2902.040 1518.060 ;
      LAYER met2 ;
        RECT 2904.530 2727.635 2904.810 2728.005 ;
        RECT 2904.600 2493.405 2904.740 2727.635 ;
        RECT 2904.530 2493.035 2904.810 2493.405 ;
        RECT 2904.600 2258.805 2904.740 2493.035 ;
        RECT 2904.530 2258.435 2904.810 2258.805 ;
        RECT 2904.600 2024.205 2904.740 2258.435 ;
        RECT 2904.530 2023.835 2904.810 2024.205 ;
        RECT 2904.600 1789.605 2904.740 2023.835 ;
        RECT 2904.530 1789.235 2904.810 1789.605 ;
        RECT 2904.600 1554.325 2904.740 1789.235 ;
        RECT 2901.770 1553.955 2902.050 1554.325 ;
        RECT 2904.530 1553.955 2904.810 1554.325 ;
        RECT 2901.840 1518.090 2901.980 1553.955 ;
        RECT 2901.780 1517.770 2902.040 1518.090 ;
        RECT 2901.840 1319.725 2901.980 1517.770 ;
        RECT 2901.770 1319.355 2902.050 1319.725 ;
        RECT 2904.530 1319.355 2904.810 1319.725 ;
        RECT 2904.600 1085.125 2904.740 1319.355 ;
        RECT 2904.530 1084.755 2904.810 1085.125 ;
        RECT 2904.600 850.525 2904.740 1084.755 ;
        RECT 2904.530 850.155 2904.810 850.525 ;
        RECT 2904.600 615.925 2904.740 850.155 ;
        RECT 2904.530 615.555 2904.810 615.925 ;
        RECT 2904.600 381.325 2904.740 615.555 ;
        RECT 2904.530 380.955 2904.810 381.325 ;
        RECT 2904.600 146.725 2904.740 380.955 ;
        RECT 2904.530 146.355 2904.810 146.725 ;
      LAYER via2 ;
        RECT 2904.530 2727.680 2904.810 2727.960 ;
        RECT 2904.530 2493.080 2904.810 2493.360 ;
        RECT 2904.530 2258.480 2904.810 2258.760 ;
        RECT 2904.530 2023.880 2904.810 2024.160 ;
        RECT 2904.530 1789.280 2904.810 1789.560 ;
        RECT 2901.770 1554.000 2902.050 1554.280 ;
        RECT 2904.530 1554.000 2904.810 1554.280 ;
        RECT 2901.770 1319.400 2902.050 1319.680 ;
        RECT 2904.530 1319.400 2904.810 1319.680 ;
        RECT 2904.530 1084.800 2904.810 1085.080 ;
        RECT 2904.530 850.200 2904.810 850.480 ;
        RECT 2904.530 615.600 2904.810 615.880 ;
        RECT 2904.530 381.000 2904.810 381.280 ;
        RECT 2904.530 146.400 2904.810 146.680 ;
      LAYER met3 ;
        RECT 2904.505 2727.970 2904.835 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2904.505 2727.670 2924.800 2727.970 ;
        RECT 2904.505 2727.655 2904.835 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2904.505 2493.370 2904.835 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2904.505 2493.070 2924.800 2493.370 ;
        RECT 2904.505 2493.055 2904.835 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2904.505 2258.770 2904.835 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2904.505 2258.470 2924.800 2258.770 ;
        RECT 2904.505 2258.455 2904.835 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2904.505 2024.170 2904.835 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2904.505 2023.870 2924.800 2024.170 ;
        RECT 2904.505 2023.855 2904.835 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2904.505 1789.570 2904.835 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2904.505 1789.270 2924.800 1789.570 ;
        RECT 2904.505 1789.255 2904.835 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2901.745 1554.290 2902.075 1554.305 ;
        RECT 2904.505 1554.290 2904.835 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2901.745 1553.990 2924.800 1554.290 ;
        RECT 2901.745 1553.975 2902.075 1553.990 ;
        RECT 2904.505 1553.975 2904.835 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 2901.745 1319.690 2902.075 1319.705 ;
        RECT 2904.505 1319.690 2904.835 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2901.745 1319.390 2924.800 1319.690 ;
        RECT 2901.745 1319.375 2902.075 1319.390 ;
        RECT 2904.505 1319.375 2904.835 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 2904.505 1085.090 2904.835 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2904.505 1084.790 2924.800 1085.090 ;
        RECT 2904.505 1084.775 2904.835 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 2904.505 850.490 2904.835 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2904.505 850.190 2924.800 850.490 ;
        RECT 2904.505 850.175 2904.835 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 2904.505 615.890 2904.835 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2904.505 615.590 2924.800 615.890 ;
        RECT 2904.505 615.575 2904.835 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 2904.505 381.290 2904.835 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2904.505 380.990 2924.800 381.290 ;
        RECT 2904.505 380.975 2904.835 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2904.505 146.690 2904.835 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2904.505 146.390 2924.800 146.690 ;
        RECT 2904.505 146.375 2904.835 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 1583.620 14.190 1583.680 ;
        RECT 17.550 1583.620 17.870 1583.680 ;
        RECT 13.870 1583.480 54.000 1583.620 ;
        RECT 13.870 1583.420 14.190 1583.480 ;
        RECT 17.550 1583.420 17.870 1583.480 ;
      LAYER via ;
        RECT 13.900 1583.420 14.160 1583.680 ;
        RECT 17.580 1583.420 17.840 1583.680 ;
      LAYER met2 ;
        RECT 13.890 1902.795 14.170 1903.165 ;
        RECT 13.960 1831.085 14.100 1902.795 ;
        RECT 13.890 1830.715 14.170 1831.085 ;
        RECT 13.960 1615.525 14.100 1830.715 ;
        RECT 13.890 1615.155 14.170 1615.525 ;
        RECT 13.960 1583.710 14.100 1615.155 ;
        RECT 13.900 1583.390 14.160 1583.710 ;
        RECT 17.580 1583.390 17.840 1583.710 ;
        RECT 17.640 1545.485 17.780 1583.390 ;
        RECT 13.890 1545.115 14.170 1545.485 ;
        RECT 17.570 1545.115 17.850 1545.485 ;
        RECT 13.960 1544.125 14.100 1545.115 ;
        RECT 13.890 1543.755 14.170 1544.125 ;
        RECT 13.960 1400.645 14.100 1543.755 ;
        RECT 13.890 1400.275 14.170 1400.645 ;
        RECT 13.960 1328.565 14.100 1400.275 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
        RECT 13.960 1185.085 14.100 1328.195 ;
        RECT 13.890 1184.715 14.170 1185.085 ;
        RECT 13.960 1113.005 14.100 1184.715 ;
        RECT 13.890 1112.635 14.170 1113.005 ;
        RECT 13.960 969.525 14.100 1112.635 ;
        RECT 13.890 969.155 14.170 969.525 ;
        RECT 13.960 897.445 14.100 969.155 ;
        RECT 13.890 897.075 14.170 897.445 ;
        RECT 13.960 753.965 14.100 897.075 ;
        RECT 13.890 753.595 14.170 753.965 ;
        RECT 13.960 681.885 14.100 753.595 ;
        RECT 13.890 681.515 14.170 681.885 ;
        RECT 13.960 538.405 14.100 681.515 ;
        RECT 13.890 538.035 14.170 538.405 ;
        RECT 13.960 466.325 14.100 538.035 ;
        RECT 13.890 465.955 14.170 466.325 ;
        RECT 13.960 322.845 14.100 465.955 ;
        RECT 13.890 322.475 14.170 322.845 ;
        RECT 13.960 250.765 14.100 322.475 ;
        RECT 13.890 250.395 14.170 250.765 ;
        RECT 13.960 107.285 14.100 250.395 ;
        RECT 13.890 106.915 14.170 107.285 ;
        RECT 13.960 35.885 14.100 106.915 ;
        RECT 13.890 35.515 14.170 35.885 ;
      LAYER via2 ;
        RECT 13.890 1902.840 14.170 1903.120 ;
        RECT 13.890 1830.760 14.170 1831.040 ;
        RECT 13.890 1615.200 14.170 1615.480 ;
        RECT 13.890 1545.160 14.170 1545.440 ;
        RECT 17.570 1545.160 17.850 1545.440 ;
        RECT 13.890 1543.800 14.170 1544.080 ;
        RECT 13.890 1400.320 14.170 1400.600 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
        RECT 13.890 1184.760 14.170 1185.040 ;
        RECT 13.890 1112.680 14.170 1112.960 ;
        RECT 13.890 969.200 14.170 969.480 ;
        RECT 13.890 897.120 14.170 897.400 ;
        RECT 13.890 753.640 14.170 753.920 ;
        RECT 13.890 681.560 14.170 681.840 ;
        RECT 13.890 538.080 14.170 538.360 ;
        RECT 13.890 466.000 14.170 466.280 ;
        RECT 13.890 322.520 14.170 322.800 ;
        RECT 13.890 250.440 14.170 250.720 ;
        RECT 13.890 106.960 14.170 107.240 ;
        RECT 13.890 35.560 14.170 35.840 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 13.865 1903.130 14.195 1903.145 ;
        RECT -4.800 1902.830 14.195 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 13.865 1902.815 14.195 1902.830 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 13.865 1831.050 14.195 1831.065 ;
        RECT -4.800 1830.750 14.195 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 13.865 1830.735 14.195 1830.750 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 13.865 1615.490 14.195 1615.505 ;
        RECT -4.800 1615.190 14.195 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 13.865 1615.175 14.195 1615.190 ;
        RECT 13.865 1545.450 14.195 1545.465 ;
        RECT 17.545 1545.450 17.875 1545.465 ;
        RECT 13.865 1545.150 17.875 1545.450 ;
        RECT 13.865 1545.135 14.195 1545.150 ;
        RECT 17.545 1545.135 17.875 1545.150 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 13.865 1544.090 14.195 1544.105 ;
        RECT -4.800 1543.790 14.195 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 13.865 1543.775 14.195 1543.790 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 13.865 1400.610 14.195 1400.625 ;
        RECT -4.800 1400.310 14.195 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 13.865 1400.295 14.195 1400.310 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.800 1328.230 14.195 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 13.865 1185.050 14.195 1185.065 ;
        RECT -4.800 1184.750 14.195 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 13.865 1184.735 14.195 1184.750 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 13.865 1112.970 14.195 1112.985 ;
        RECT -4.800 1112.670 14.195 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 13.865 1112.655 14.195 1112.670 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 13.865 969.490 14.195 969.505 ;
        RECT -4.800 969.190 14.195 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 13.865 969.175 14.195 969.190 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 13.865 753.930 14.195 753.945 ;
        RECT -4.800 753.630 14.195 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 13.865 753.615 14.195 753.630 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 13.865 681.850 14.195 681.865 ;
        RECT -4.800 681.550 14.195 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 13.865 681.535 14.195 681.550 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 13.865 538.370 14.195 538.385 ;
        RECT -4.800 538.070 14.195 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 13.865 538.055 14.195 538.070 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 13.865 466.290 14.195 466.305 ;
        RECT -4.800 465.990 14.195 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 13.865 465.975 14.195 465.990 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 13.865 322.810 14.195 322.825 ;
        RECT -4.800 322.510 14.195 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 13.865 322.495 14.195 322.510 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 13.865 250.730 14.195 250.745 ;
        RECT -4.800 250.430 14.195 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 13.865 250.415 14.195 250.430 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 13.865 107.250 14.195 107.265 ;
        RECT -4.800 106.950 14.195 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 13.865 106.935 14.195 106.950 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 13.865 35.850 14.195 35.865 ;
        RECT -4.800 35.550 14.195 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 13.865 35.535 14.195 35.550 ;
    END
  END io_oeb[29]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2881.050 2898.400 2881.370 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2881.050 2898.260 2901.150 2898.400 ;
        RECT 2881.050 2898.200 2881.370 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2881.050 314.060 2881.370 314.120 ;
        RECT 2866.000 313.920 2881.370 314.060 ;
        RECT 2881.050 313.860 2881.370 313.920 ;
      LAYER via ;
        RECT 2881.080 2898.200 2881.340 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2881.080 313.860 2881.340 314.120 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2881.080 2898.170 2881.340 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2881.140 314.150 2881.280 2898.170 ;
        RECT 2881.080 313.830 2881.340 314.150 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 1411.810 3501.900 1412.130 3501.960 ;
        RECT 202.470 3501.760 1412.130 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 1411.810 3501.700 1412.130 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 1411.840 3501.700 1412.100 3501.960 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 1411.840 3501.670 1412.100 3501.990 ;
        RECT 1411.900 3466.000 1412.040 3501.670 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 17.550 3408.600 54.000 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2425.460 17.410 2425.520 ;
        RECT 17.090 2425.320 54.000 2425.460 ;
        RECT 17.090 2425.260 17.410 2425.320 ;
      LAYER via ;
        RECT 17.120 2425.260 17.380 2425.520 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 2425.550 17.320 3124.075 ;
        RECT 17.120 2425.230 17.380 2425.550 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2836.180 17.870 2836.240 ;
        RECT 45.610 2836.180 45.930 2836.240 ;
        RECT 17.550 2836.040 45.930 2836.180 ;
        RECT 17.550 2835.980 17.870 2836.040 ;
        RECT 45.610 2835.980 45.930 2836.040 ;
        RECT 45.610 2221.800 45.930 2221.860 ;
        RECT 45.610 2221.660 54.000 2221.800 ;
        RECT 45.610 2221.600 45.930 2221.660 ;
      LAYER via ;
        RECT 17.580 2835.980 17.840 2836.240 ;
        RECT 45.640 2835.980 45.900 2836.240 ;
        RECT 45.640 2221.600 45.900 2221.860 ;
      LAYER met2 ;
        RECT 17.570 2836.435 17.850 2836.805 ;
        RECT 17.640 2836.270 17.780 2836.435 ;
        RECT 17.580 2835.950 17.840 2836.270 ;
        RECT 45.640 2835.950 45.900 2836.270 ;
        RECT 45.700 2221.890 45.840 2835.950 ;
        RECT 45.640 2221.570 45.900 2221.890 ;
      LAYER via2 ;
        RECT 17.570 2836.480 17.850 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.545 2836.770 17.875 2836.785 ;
        RECT -4.800 2836.470 17.875 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.545 2836.455 17.875 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.330 2546.500 14.650 2546.560 ;
        RECT 14.330 2546.360 54.000 2546.500 ;
        RECT 14.330 2546.300 14.650 2546.360 ;
      LAYER via ;
        RECT 14.360 2546.300 14.620 2546.560 ;
      LAYER met2 ;
        RECT 14.350 2549.475 14.630 2549.845 ;
        RECT 14.420 2546.590 14.560 2549.475 ;
        RECT 14.360 2546.270 14.620 2546.590 ;
      LAYER via2 ;
        RECT 14.350 2549.520 14.630 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 14.325 2549.810 14.655 2549.825 ;
        RECT -4.800 2549.510 14.655 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 14.325 2549.495 14.655 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2256.480 17.410 2256.540 ;
        RECT 17.090 2256.340 54.000 2256.480 ;
        RECT 17.090 2256.280 17.410 2256.340 ;
      LAYER via ;
        RECT 17.120 2256.280 17.380 2256.540 ;
      LAYER met2 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
        RECT 17.180 2256.570 17.320 2261.835 ;
        RECT 17.120 2256.250 17.380 2256.570 ;
      LAYER via2 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 1974.875 24.290 1975.245 ;
        RECT 24.080 868.885 24.220 1974.875 ;
        RECT 24.010 868.515 24.290 868.885 ;
      LAYER via2 ;
        RECT 24.010 1974.920 24.290 1975.200 ;
        RECT 24.010 868.560 24.290 868.840 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 23.985 1975.210 24.315 1975.225 ;
        RECT -4.800 1974.910 24.315 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 23.985 1974.895 24.315 1974.910 ;
        RECT 23.985 868.850 24.315 868.865 ;
        RECT 23.985 868.550 46.610 868.850 ;
        RECT 23.985 868.535 24.315 868.550 ;
        RECT 46.310 867.980 46.610 868.550 ;
        RECT 46.000 867.380 50.000 867.980 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1683.920 16.030 1683.980 ;
        RECT 30.890 1683.920 31.210 1683.980 ;
        RECT 15.710 1683.780 31.210 1683.920 ;
        RECT 15.710 1683.720 16.030 1683.780 ;
        RECT 30.890 1683.720 31.210 1683.780 ;
      LAYER via ;
        RECT 15.740 1683.720 16.000 1683.980 ;
        RECT 30.920 1683.720 31.180 1683.980 ;
      LAYER met2 ;
        RECT 15.730 1687.235 16.010 1687.605 ;
        RECT 15.800 1684.010 15.940 1687.235 ;
        RECT 15.740 1683.690 16.000 1684.010 ;
        RECT 30.920 1683.690 31.180 1684.010 ;
        RECT 30.980 327.605 31.120 1683.690 ;
        RECT 30.910 327.235 31.190 327.605 ;
      LAYER via2 ;
        RECT 15.730 1687.280 16.010 1687.560 ;
        RECT 30.910 327.280 31.190 327.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 15.705 1687.570 16.035 1687.585 ;
        RECT -4.800 1687.270 16.035 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 15.705 1687.255 16.035 1687.270 ;
        RECT 30.885 327.570 31.215 327.585 ;
        RECT 46.000 327.570 50.000 327.840 ;
        RECT 30.885 327.270 50.000 327.570 ;
        RECT 30.885 327.255 31.215 327.270 ;
        RECT 46.000 327.240 50.000 327.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 1121.220 18.330 1121.280 ;
        RECT 18.010 1121.080 54.000 1121.220 ;
        RECT 18.010 1121.020 18.330 1121.080 ;
      LAYER via ;
        RECT 18.040 1121.020 18.300 1121.280 ;
      LAYER met2 ;
        RECT 18.030 1471.675 18.310 1472.045 ;
        RECT 18.100 1121.310 18.240 1471.675 ;
        RECT 18.040 1120.990 18.300 1121.310 ;
      LAYER via2 ;
        RECT 18.030 1471.720 18.310 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 18.005 1472.010 18.335 1472.025 ;
        RECT -4.800 1471.710 18.335 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 18.005 1471.695 18.335 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 1118.160 17.870 1118.220 ;
        RECT 17.550 1118.020 54.000 1118.160 ;
        RECT 17.550 1117.960 17.870 1118.020 ;
      LAYER via ;
        RECT 17.580 1117.960 17.840 1118.220 ;
      LAYER met2 ;
        RECT 17.580 1117.930 17.840 1118.250 ;
        RECT 17.640 179.365 17.780 1117.930 ;
        RECT 17.570 178.995 17.850 179.365 ;
      LAYER via2 ;
        RECT 17.570 179.040 17.850 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.545 179.330 17.875 179.345 ;
        RECT -4.800 179.030 17.875 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.545 179.015 17.875 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2866.000 206.820 2901.150 206.960 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2887.950 2548.200 2888.270 2548.260 ;
        RECT 2898.070 2548.200 2898.390 2548.260 ;
        RECT 2887.950 2548.060 2898.390 2548.200 ;
        RECT 2887.950 2548.000 2888.270 2548.060 ;
        RECT 2898.070 2548.000 2898.390 2548.060 ;
        RECT 2887.950 1635.300 2888.270 1635.360 ;
        RECT 2866.000 1635.160 2888.270 1635.300 ;
        RECT 2887.950 1635.100 2888.270 1635.160 ;
      LAYER via ;
        RECT 2887.980 2548.000 2888.240 2548.260 ;
        RECT 2898.100 2548.000 2898.360 2548.260 ;
        RECT 2887.980 1635.100 2888.240 1635.360 ;
      LAYER met2 ;
        RECT 2898.090 2551.515 2898.370 2551.885 ;
        RECT 2898.160 2548.290 2898.300 2551.515 ;
        RECT 2887.980 2547.970 2888.240 2548.290 ;
        RECT 2898.100 2547.970 2898.360 2548.290 ;
        RECT 2888.040 1635.390 2888.180 2547.970 ;
        RECT 2887.980 1635.070 2888.240 1635.390 ;
      LAYER via2 ;
        RECT 2898.090 2551.560 2898.370 2551.840 ;
      LAYER met3 ;
        RECT 2898.065 2551.850 2898.395 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2898.065 2551.550 2924.800 2551.850 ;
        RECT 2898.065 2551.535 2898.395 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2866.000 2780.960 2901.150 2781.100 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2894.390 469.100 2894.710 469.160 ;
        RECT 2866.000 468.960 2894.710 469.100 ;
        RECT 2894.390 468.900 2894.710 468.960 ;
      LAYER via ;
        RECT 2894.420 468.900 2894.680 469.160 ;
      LAYER met2 ;
        RECT 2894.410 3020.715 2894.690 3021.085 ;
        RECT 2894.480 469.190 2894.620 3020.715 ;
        RECT 2894.420 468.870 2894.680 469.190 ;
      LAYER via2 ;
        RECT 2894.410 3020.760 2894.690 3021.040 ;
      LAYER met3 ;
        RECT 2894.385 3021.050 2894.715 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2894.385 3020.750 2924.800 3021.050 ;
        RECT 2894.385 3020.735 2894.715 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2887.490 3250.300 2887.810 3250.360 ;
        RECT 2898.070 3250.300 2898.390 3250.360 ;
        RECT 2887.490 3250.160 2898.390 3250.300 ;
        RECT 2887.490 3250.100 2887.810 3250.160 ;
        RECT 2898.070 3250.100 2898.390 3250.160 ;
        RECT 2887.490 468.760 2887.810 468.820 ;
        RECT 2866.000 468.620 2887.810 468.760 ;
        RECT 2887.490 468.560 2887.810 468.620 ;
      LAYER via ;
        RECT 2887.520 3250.100 2887.780 3250.360 ;
        RECT 2898.100 3250.100 2898.360 3250.360 ;
        RECT 2887.520 468.560 2887.780 468.820 ;
      LAYER met2 ;
        RECT 2898.090 3255.315 2898.370 3255.685 ;
        RECT 2898.160 3250.390 2898.300 3255.315 ;
        RECT 2887.520 3250.070 2887.780 3250.390 ;
        RECT 2898.100 3250.070 2898.360 3250.390 ;
        RECT 2887.580 468.850 2887.720 3250.070 ;
        RECT 2887.520 468.530 2887.780 468.850 ;
      LAYER via2 ;
        RECT 2898.090 3255.360 2898.370 3255.640 ;
      LAYER met3 ;
        RECT 2898.065 3255.650 2898.395 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2898.065 3255.350 2924.800 3255.650 ;
        RECT 2898.065 3255.335 2898.395 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2880.590 3484.900 2880.910 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2880.590 3484.760 2901.150 3484.900 ;
        RECT 2880.590 3484.700 2880.910 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 2880.590 475.900 2880.910 475.960 ;
        RECT 2866.000 475.760 2880.910 475.900 ;
        RECT 2880.590 475.700 2880.910 475.760 ;
      LAYER via ;
        RECT 2880.620 3484.700 2880.880 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 2880.620 475.700 2880.880 475.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2880.620 3484.670 2880.880 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2880.680 475.990 2880.820 3484.670 ;
        RECT 2880.620 475.670 2880.880 475.990 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1576.490 3501.560 1576.810 3501.620 ;
        RECT 2635.870 3501.560 2636.190 3501.620 ;
        RECT 1576.490 3501.420 2636.190 3501.560 ;
        RECT 1576.490 3501.360 1576.810 3501.420 ;
        RECT 2635.870 3501.360 2636.190 3501.420 ;
      LAYER via ;
        RECT 1576.520 3501.360 1576.780 3501.620 ;
        RECT 2635.900 3501.360 2636.160 3501.620 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.650 2636.100 3517.600 ;
        RECT 1576.520 3501.330 1576.780 3501.650 ;
        RECT 2635.900 3501.330 2636.160 3501.650 ;
        RECT 1576.580 3466.000 1576.720 3501.330 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1562.690 3501.900 1563.010 3501.960 ;
        RECT 2311.570 3501.900 2311.890 3501.960 ;
        RECT 1562.690 3501.760 2311.890 3501.900 ;
        RECT 1562.690 3501.700 1563.010 3501.760 ;
        RECT 2311.570 3501.700 2311.890 3501.760 ;
      LAYER via ;
        RECT 1562.720 3501.700 1562.980 3501.960 ;
        RECT 2311.600 3501.700 2311.860 3501.960 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.990 2311.800 3517.600 ;
        RECT 1562.720 3501.670 1562.980 3501.990 ;
        RECT 2311.600 3501.670 2311.860 3501.990 ;
        RECT 1562.780 3466.000 1562.920 3501.670 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1507.490 3502.580 1507.810 3502.640 ;
        RECT 1987.270 3502.580 1987.590 3502.640 ;
        RECT 1507.490 3502.440 1987.590 3502.580 ;
        RECT 1507.490 3502.380 1507.810 3502.440 ;
        RECT 1987.270 3502.380 1987.590 3502.440 ;
      LAYER via ;
        RECT 1507.520 3502.380 1507.780 3502.640 ;
        RECT 1987.300 3502.380 1987.560 3502.640 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3502.670 1987.500 3517.600 ;
        RECT 1507.520 3502.350 1507.780 3502.670 ;
        RECT 1987.300 3502.350 1987.560 3502.670 ;
        RECT 1507.580 3466.000 1507.720 3502.350 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1528.190 3502.920 1528.510 3502.980 ;
        RECT 1662.510 3502.920 1662.830 3502.980 ;
        RECT 1528.190 3502.780 1662.830 3502.920 ;
        RECT 1528.190 3502.720 1528.510 3502.780 ;
        RECT 1662.510 3502.720 1662.830 3502.780 ;
      LAYER via ;
        RECT 1528.220 3502.720 1528.480 3502.980 ;
        RECT 1662.540 3502.720 1662.800 3502.980 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.010 1662.740 3517.600 ;
        RECT 1528.220 3502.690 1528.480 3503.010 ;
        RECT 1662.540 3502.690 1662.800 3503.010 ;
        RECT 1528.280 3466.000 1528.420 3502.690 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3502.580 1338.530 3502.640 ;
        RECT 1410.890 3502.580 1411.210 3502.640 ;
        RECT 1338.210 3502.440 1411.210 3502.580 ;
        RECT 1338.210 3502.380 1338.530 3502.440 ;
        RECT 1410.890 3502.380 1411.210 3502.440 ;
      LAYER via ;
        RECT 1338.240 3502.380 1338.500 3502.640 ;
        RECT 1410.920 3502.380 1411.180 3502.640 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3502.670 1338.440 3517.600 ;
        RECT 1338.240 3502.350 1338.500 3502.670 ;
        RECT 1410.920 3502.350 1411.180 3502.670 ;
        RECT 1410.980 3466.000 1411.120 3502.350 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2866.000 441.420 2901.150 441.560 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3502.580 1014.230 3502.640 ;
        RECT 1253.110 3502.580 1253.430 3502.640 ;
        RECT 1013.910 3502.440 1253.430 3502.580 ;
        RECT 1013.910 3502.380 1014.230 3502.440 ;
        RECT 1253.110 3502.380 1253.430 3502.440 ;
        RECT 1253.110 3493.400 1253.430 3493.460 ;
        RECT 1262.770 3493.400 1263.090 3493.460 ;
        RECT 1253.110 3493.260 1263.090 3493.400 ;
        RECT 1253.110 3493.200 1253.430 3493.260 ;
        RECT 1262.770 3493.200 1263.090 3493.260 ;
        RECT 1262.770 3484.560 1263.090 3484.620 ;
        RECT 1300.030 3484.560 1300.350 3484.620 ;
        RECT 1262.770 3484.420 1300.350 3484.560 ;
        RECT 1262.770 3484.360 1263.090 3484.420 ;
        RECT 1300.030 3484.360 1300.350 3484.420 ;
        RECT 1300.030 3474.020 1300.350 3474.080 ;
        RECT 1334.990 3474.020 1335.310 3474.080 ;
        RECT 1300.030 3473.880 1335.310 3474.020 ;
        RECT 1300.030 3473.820 1300.350 3473.880 ;
        RECT 1334.990 3473.820 1335.310 3473.880 ;
      LAYER via ;
        RECT 1013.940 3502.380 1014.200 3502.640 ;
        RECT 1253.140 3502.380 1253.400 3502.640 ;
        RECT 1253.140 3493.200 1253.400 3493.460 ;
        RECT 1262.800 3493.200 1263.060 3493.460 ;
        RECT 1262.800 3484.360 1263.060 3484.620 ;
        RECT 1300.060 3484.360 1300.320 3484.620 ;
        RECT 1300.060 3473.820 1300.320 3474.080 ;
        RECT 1335.020 3473.820 1335.280 3474.080 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3502.670 1014.140 3517.600 ;
        RECT 1013.940 3502.350 1014.200 3502.670 ;
        RECT 1253.140 3502.350 1253.400 3502.670 ;
        RECT 1253.200 3493.490 1253.340 3502.350 ;
        RECT 1253.140 3493.170 1253.400 3493.490 ;
        RECT 1262.800 3493.170 1263.060 3493.490 ;
        RECT 1262.860 3484.650 1263.000 3493.170 ;
        RECT 1262.800 3484.330 1263.060 3484.650 ;
        RECT 1300.060 3484.330 1300.320 3484.650 ;
        RECT 1300.120 3474.110 1300.260 3484.330 ;
        RECT 1300.060 3473.790 1300.320 3474.110 ;
        RECT 1335.020 3473.790 1335.280 3474.110 ;
        RECT 1335.080 3466.000 1335.220 3473.790 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 683.170 3487.960 683.490 3488.020 ;
        RECT 689.150 3487.960 689.470 3488.020 ;
        RECT 683.170 3487.820 689.470 3487.960 ;
        RECT 683.170 3487.760 683.490 3487.820 ;
        RECT 689.150 3487.760 689.470 3487.820 ;
      LAYER via ;
        RECT 683.200 3487.760 683.460 3488.020 ;
        RECT 689.180 3487.760 689.440 3488.020 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3488.050 689.380 3517.600 ;
        RECT 683.200 3487.730 683.460 3488.050 ;
        RECT 689.180 3487.730 689.440 3488.050 ;
        RECT 683.260 3466.000 683.400 3487.730 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 258.590 3502.240 258.910 3502.300 ;
        RECT 364.850 3502.240 365.170 3502.300 ;
        RECT 258.590 3502.100 365.170 3502.240 ;
        RECT 258.590 3502.040 258.910 3502.100 ;
        RECT 364.850 3502.040 365.170 3502.100 ;
      LAYER via ;
        RECT 258.620 3502.040 258.880 3502.300 ;
        RECT 364.880 3502.040 365.140 3502.300 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 258.620 3502.010 258.880 3502.330 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 258.680 3466.000 258.820 3502.010 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.560 40.870 3501.620 ;
        RECT 44.690 3501.560 45.010 3501.620 ;
        RECT 40.550 3501.420 45.010 3501.560 ;
        RECT 40.550 3501.360 40.870 3501.420 ;
        RECT 44.690 3501.360 45.010 3501.420 ;
        RECT 44.690 627.880 45.010 627.940 ;
        RECT 44.690 627.740 54.000 627.880 ;
        RECT 44.690 627.680 45.010 627.740 ;
      LAYER via ;
        RECT 40.580 3501.360 40.840 3501.620 ;
        RECT 44.720 3501.360 44.980 3501.620 ;
        RECT 44.720 627.680 44.980 627.940 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.650 40.780 3517.600 ;
        RECT 40.580 3501.330 40.840 3501.650 ;
        RECT 44.720 3501.330 44.980 3501.650 ;
        RECT 44.780 627.970 44.920 3501.330 ;
        RECT 44.720 627.650 44.980 627.970 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 51.590 3263.900 51.910 3263.960 ;
        RECT 15.250 3263.760 51.910 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 51.590 3263.700 51.910 3263.760 ;
        RECT 51.590 634.680 51.910 634.740 ;
        RECT 51.590 634.540 54.000 634.680 ;
        RECT 51.590 634.480 51.910 634.540 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 51.620 3263.700 51.880 3263.960 ;
        RECT 51.620 634.480 51.880 634.740 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 51.620 3263.670 51.880 3263.990 ;
        RECT 51.680 634.770 51.820 3263.670 ;
        RECT 51.620 634.450 51.880 634.770 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2974.220 17.870 2974.280 ;
        RECT 45.150 2974.220 45.470 2974.280 ;
        RECT 17.550 2974.080 45.470 2974.220 ;
        RECT 17.550 2974.020 17.870 2974.080 ;
        RECT 45.150 2974.020 45.470 2974.080 ;
        RECT 45.150 641.480 45.470 641.540 ;
        RECT 45.150 641.340 54.000 641.480 ;
        RECT 45.150 641.280 45.470 641.340 ;
      LAYER via ;
        RECT 17.580 2974.020 17.840 2974.280 ;
        RECT 45.180 2974.020 45.440 2974.280 ;
        RECT 45.180 641.280 45.440 641.540 ;
      LAYER met2 ;
        RECT 17.570 2979.915 17.850 2980.285 ;
        RECT 17.640 2974.310 17.780 2979.915 ;
        RECT 17.580 2973.990 17.840 2974.310 ;
        RECT 45.180 2973.990 45.440 2974.310 ;
        RECT 45.240 641.570 45.380 2973.990 ;
        RECT 45.180 641.250 45.440 641.570 ;
      LAYER via2 ;
        RECT 17.570 2979.960 17.850 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 17.545 2980.250 17.875 2980.265 ;
        RECT -4.800 2979.950 17.875 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 17.545 2979.935 17.875 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2691.340 17.870 2691.400 ;
        RECT 52.050 2691.340 52.370 2691.400 ;
        RECT 17.550 2691.200 52.370 2691.340 ;
        RECT 17.550 2691.140 17.870 2691.200 ;
        RECT 52.050 2691.140 52.370 2691.200 ;
        RECT 52.140 646.440 54.000 646.580 ;
        RECT 52.140 646.300 52.280 646.440 ;
        RECT 52.050 646.040 52.370 646.300 ;
      LAYER via ;
        RECT 17.580 2691.140 17.840 2691.400 ;
        RECT 52.080 2691.140 52.340 2691.400 ;
        RECT 52.080 646.040 52.340 646.300 ;
      LAYER met2 ;
        RECT 17.570 2692.955 17.850 2693.325 ;
        RECT 17.640 2691.430 17.780 2692.955 ;
        RECT 17.580 2691.110 17.840 2691.430 ;
        RECT 52.080 2691.110 52.340 2691.430 ;
        RECT 52.140 646.330 52.280 2691.110 ;
        RECT 52.080 646.010 52.340 646.330 ;
      LAYER via2 ;
        RECT 17.570 2693.000 17.850 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.545 2693.290 17.875 2693.305 ;
        RECT -4.800 2692.990 17.875 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.545 2692.975 17.875 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2401.320 16.030 2401.380 ;
        RECT 15.710 2401.180 54.000 2401.320 ;
        RECT 15.710 2401.120 16.030 2401.180 ;
      LAYER via ;
        RECT 15.740 2401.120 16.000 2401.380 ;
      LAYER met2 ;
        RECT 15.730 2405.315 16.010 2405.685 ;
        RECT 15.800 2401.410 15.940 2405.315 ;
        RECT 15.740 2401.090 16.000 2401.410 ;
      LAYER via2 ;
        RECT 15.730 2405.360 16.010 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.705 2405.650 16.035 2405.665 ;
        RECT -4.800 2405.350 16.035 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.705 2405.335 16.035 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2866.000 676.020 2901.150 676.160 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.910 910.760 2900.230 910.820 ;
        RECT 2866.000 910.620 2900.230 910.760 ;
        RECT 2899.910 910.560 2900.230 910.620 ;
      LAYER via ;
        RECT 2899.940 910.560 2900.200 910.820 ;
      LAYER met2 ;
        RECT 2899.940 910.530 2900.200 910.850 ;
        RECT 2900.000 909.685 2900.140 910.530 ;
        RECT 2899.930 909.315 2900.210 909.685 ;
      LAYER via2 ;
        RECT 2899.930 909.360 2900.210 909.640 ;
      LAYER met3 ;
        RECT 2899.905 909.650 2900.235 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2899.905 909.350 2924.800 909.650 ;
        RECT 2899.905 909.335 2900.235 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2899.910 1145.360 2900.230 1145.420 ;
        RECT 2866.000 1145.220 2900.230 1145.360 ;
        RECT 2899.910 1145.160 2900.230 1145.220 ;
      LAYER via ;
        RECT 2899.940 1145.160 2900.200 1145.420 ;
      LAYER met2 ;
        RECT 2899.940 1145.130 2900.200 1145.450 ;
        RECT 2900.000 1144.285 2900.140 1145.130 ;
        RECT 2899.930 1143.915 2900.210 1144.285 ;
      LAYER via2 ;
        RECT 2899.930 1143.960 2900.210 1144.240 ;
      LAYER met3 ;
        RECT 2899.905 1144.250 2900.235 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2899.905 1143.950 2924.800 1144.250 ;
        RECT 2899.905 1143.935 2900.235 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 2866.000 1379.820 2901.150 1379.960 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 1608.100 2901.150 1608.160 ;
        RECT 2866.000 1607.960 2901.150 1608.100 ;
        RECT 2900.830 1607.900 2901.150 1607.960 ;
      LAYER via ;
        RECT 2900.860 1607.900 2901.120 1608.160 ;
      LAYER met2 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
        RECT 2900.920 1608.190 2901.060 1613.115 ;
        RECT 2900.860 1607.870 2901.120 1608.190 ;
      LAYER via2 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
      LAYER met3 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 1842.700 2901.150 1842.760 ;
        RECT 2866.000 1842.560 2901.150 1842.700 ;
        RECT 2900.830 1842.500 2901.150 1842.560 ;
      LAYER via ;
        RECT 2900.860 1842.500 2901.120 1842.760 ;
      LAYER met2 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
        RECT 2900.920 1842.790 2901.060 1847.715 ;
        RECT 2900.860 1842.470 2901.120 1842.790 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 2866.000 2077.160 2901.150 2077.300 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
      LAYER via ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2866.000 2311.760 2901.150 2311.900 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
      LAYER via ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 633.105 2.805 633.275 48.195 ;
      LAYER mcon ;
        RECT 633.105 48.025 633.275 48.195 ;
      LAYER met1 ;
        RECT 633.045 48.180 633.335 48.225 ;
        RECT 634.410 48.180 634.730 48.240 ;
        RECT 633.045 48.040 634.730 48.180 ;
        RECT 633.045 47.995 633.335 48.040 ;
        RECT 634.410 47.980 634.730 48.040 ;
        RECT 633.030 2.960 633.350 3.020 ;
        RECT 632.835 2.820 633.350 2.960 ;
        RECT 633.030 2.760 633.350 2.820 ;
      LAYER via ;
        RECT 634.440 47.980 634.700 48.240 ;
        RECT 633.060 2.760 633.320 3.020 ;
      LAYER met2 ;
        RECT 634.500 48.270 634.640 54.000 ;
        RECT 634.440 47.950 634.700 48.270 ;
        RECT 633.060 2.730 633.320 3.050 ;
        RECT 633.120 2.400 633.260 2.730 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2417.370 46.480 2417.690 46.540 ;
        RECT 2645.990 46.480 2646.310 46.540 ;
        RECT 2417.370 46.340 2646.310 46.480 ;
        RECT 2417.370 46.280 2417.690 46.340 ;
        RECT 2645.990 46.280 2646.310 46.340 ;
      LAYER via ;
        RECT 2417.400 46.280 2417.660 46.540 ;
        RECT 2646.020 46.280 2646.280 46.540 ;
      LAYER met2 ;
        RECT 2646.080 46.570 2646.220 54.000 ;
        RECT 2417.400 46.250 2417.660 46.570 ;
        RECT 2646.020 46.250 2646.280 46.570 ;
        RECT 2417.460 2.400 2417.600 46.250 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2434.850 51.920 2435.170 51.980 ;
        RECT 2651.510 51.920 2651.830 51.980 ;
        RECT 2434.850 51.780 2651.830 51.920 ;
        RECT 2434.850 51.720 2435.170 51.780 ;
        RECT 2651.510 51.720 2651.830 51.780 ;
      LAYER via ;
        RECT 2434.880 51.720 2435.140 51.980 ;
        RECT 2651.540 51.720 2651.800 51.980 ;
      LAYER met2 ;
        RECT 2651.600 52.010 2651.740 54.000 ;
        RECT 2434.880 51.690 2435.140 52.010 ;
        RECT 2651.540 51.690 2651.800 52.010 ;
        RECT 2434.940 2.400 2435.080 51.690 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2452.790 16.900 2453.110 16.960 ;
        RECT 2456.010 16.900 2456.330 16.960 ;
        RECT 2452.790 16.760 2456.330 16.900 ;
        RECT 2452.790 16.700 2453.110 16.760 ;
        RECT 2456.010 16.700 2456.330 16.760 ;
      LAYER via ;
        RECT 2452.820 16.700 2453.080 16.960 ;
        RECT 2456.040 16.700 2456.300 16.960 ;
      LAYER met2 ;
        RECT 2456.100 16.990 2456.240 54.000 ;
        RECT 2452.820 16.670 2453.080 16.990 ;
        RECT 2456.040 16.670 2456.300 16.990 ;
        RECT 2452.880 2.400 2453.020 16.670 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2471.190 47.160 2471.510 47.220 ;
        RECT 2661.630 47.160 2661.950 47.220 ;
        RECT 2471.190 47.020 2661.950 47.160 ;
        RECT 2471.190 46.960 2471.510 47.020 ;
        RECT 2661.630 46.960 2661.950 47.020 ;
      LAYER via ;
        RECT 2471.220 46.960 2471.480 47.220 ;
        RECT 2661.660 46.960 2661.920 47.220 ;
      LAYER met2 ;
        RECT 2661.720 47.250 2661.860 54.000 ;
        RECT 2471.220 46.930 2471.480 47.250 ;
        RECT 2661.660 46.930 2661.920 47.250 ;
        RECT 2471.280 3.130 2471.420 46.930 ;
        RECT 2470.820 2.990 2471.420 3.130 ;
        RECT 2470.820 2.400 2470.960 2.990 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2490.510 52.260 2490.830 52.320 ;
        RECT 2668.990 52.260 2669.310 52.320 ;
        RECT 2490.510 52.120 2669.310 52.260 ;
        RECT 2490.510 52.060 2490.830 52.120 ;
        RECT 2668.990 52.060 2669.310 52.120 ;
      LAYER via ;
        RECT 2490.540 52.060 2490.800 52.320 ;
        RECT 2669.020 52.060 2669.280 52.320 ;
      LAYER met2 ;
        RECT 2669.080 52.350 2669.220 54.000 ;
        RECT 2490.540 52.030 2490.800 52.350 ;
        RECT 2669.020 52.030 2669.280 52.350 ;
        RECT 2490.600 3.130 2490.740 52.030 ;
        RECT 2488.760 2.990 2490.740 3.130 ;
        RECT 2488.760 2.400 2488.900 2.990 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2506.150 17.580 2506.470 17.640 ;
        RECT 2511.210 17.580 2511.530 17.640 ;
        RECT 2506.150 17.440 2511.530 17.580 ;
        RECT 2506.150 17.380 2506.470 17.440 ;
        RECT 2511.210 17.380 2511.530 17.440 ;
      LAYER via ;
        RECT 2506.180 17.380 2506.440 17.640 ;
        RECT 2511.240 17.380 2511.500 17.640 ;
      LAYER met2 ;
        RECT 2511.300 17.670 2511.440 54.000 ;
        RECT 2506.180 17.350 2506.440 17.670 ;
        RECT 2511.240 17.350 2511.500 17.670 ;
        RECT 2506.240 2.400 2506.380 17.350 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2524.090 32.200 2524.410 32.260 ;
        RECT 2677.730 32.200 2678.050 32.260 ;
        RECT 2524.090 32.060 2678.050 32.200 ;
        RECT 2524.090 32.000 2524.410 32.060 ;
        RECT 2677.730 32.000 2678.050 32.060 ;
      LAYER via ;
        RECT 2524.120 32.000 2524.380 32.260 ;
        RECT 2677.760 32.000 2678.020 32.260 ;
      LAYER met2 ;
        RECT 2677.820 32.290 2677.960 54.000 ;
        RECT 2524.120 31.970 2524.380 32.290 ;
        RECT 2677.760 31.970 2678.020 32.290 ;
        RECT 2524.180 2.400 2524.320 31.970 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2542.030 21.660 2542.350 21.720 ;
        RECT 2685.090 21.660 2685.410 21.720 ;
        RECT 2542.030 21.520 2685.410 21.660 ;
        RECT 2542.030 21.460 2542.350 21.520 ;
        RECT 2685.090 21.460 2685.410 21.520 ;
      LAYER via ;
        RECT 2542.060 21.460 2542.320 21.720 ;
        RECT 2685.120 21.460 2685.380 21.720 ;
      LAYER met2 ;
        RECT 2685.180 21.750 2685.320 54.000 ;
        RECT 2542.060 21.430 2542.320 21.750 ;
        RECT 2685.120 21.430 2685.380 21.750 ;
        RECT 2542.120 2.400 2542.260 21.430 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2559.970 37.980 2560.290 38.040 ;
        RECT 2691.990 37.980 2692.310 38.040 ;
        RECT 2559.970 37.840 2692.310 37.980 ;
        RECT 2559.970 37.780 2560.290 37.840 ;
        RECT 2691.990 37.780 2692.310 37.840 ;
      LAYER via ;
        RECT 2560.000 37.780 2560.260 38.040 ;
        RECT 2692.020 37.780 2692.280 38.040 ;
      LAYER met2 ;
        RECT 2692.080 38.070 2692.220 54.000 ;
        RECT 2560.000 37.750 2560.260 38.070 ;
        RECT 2692.020 37.750 2692.280 38.070 ;
        RECT 2560.060 2.400 2560.200 37.750 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2577.910 20.640 2578.230 20.700 ;
        RECT 2580.210 20.640 2580.530 20.700 ;
        RECT 2577.910 20.500 2580.530 20.640 ;
        RECT 2577.910 20.440 2578.230 20.500 ;
        RECT 2580.210 20.440 2580.530 20.500 ;
      LAYER via ;
        RECT 2577.940 20.440 2578.200 20.700 ;
        RECT 2580.240 20.440 2580.500 20.700 ;
      LAYER met2 ;
        RECT 2580.300 20.730 2580.440 54.000 ;
        RECT 2577.940 20.410 2578.200 20.730 ;
        RECT 2580.240 20.410 2580.500 20.730 ;
        RECT 2578.000 2.400 2578.140 20.410 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 911.405 17.425 912.035 17.595 ;
      LAYER mcon ;
        RECT 911.865 17.425 912.035 17.595 ;
      LAYER met1 ;
        RECT 811.510 17.580 811.830 17.640 ;
        RECT 911.345 17.580 911.635 17.625 ;
        RECT 811.510 17.440 911.635 17.580 ;
        RECT 811.510 17.380 811.830 17.440 ;
        RECT 911.345 17.395 911.635 17.440 ;
        RECT 911.805 17.580 912.095 17.625 ;
        RECT 1196.990 17.580 1197.310 17.640 ;
        RECT 911.805 17.440 1197.310 17.580 ;
        RECT 911.805 17.395 912.095 17.440 ;
        RECT 1196.990 17.380 1197.310 17.440 ;
      LAYER via ;
        RECT 811.540 17.380 811.800 17.640 ;
        RECT 1197.020 17.380 1197.280 17.640 ;
      LAYER met2 ;
        RECT 1197.080 17.670 1197.220 54.000 ;
        RECT 811.540 17.350 811.800 17.670 ;
        RECT 1197.020 17.350 1197.280 17.670 ;
        RECT 811.600 2.400 811.740 17.350 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2697.970 34.580 2698.290 34.640 ;
        RECT 2702.570 34.580 2702.890 34.640 ;
        RECT 2697.970 34.440 2702.890 34.580 ;
        RECT 2697.970 34.380 2698.290 34.440 ;
        RECT 2702.570 34.380 2702.890 34.440 ;
        RECT 2595.390 30.840 2595.710 30.900 ;
        RECT 2697.970 30.840 2698.290 30.900 ;
        RECT 2595.390 30.700 2698.290 30.840 ;
        RECT 2595.390 30.640 2595.710 30.700 ;
        RECT 2697.970 30.640 2698.290 30.700 ;
      LAYER via ;
        RECT 2698.000 34.380 2698.260 34.640 ;
        RECT 2702.600 34.380 2702.860 34.640 ;
        RECT 2595.420 30.640 2595.680 30.900 ;
        RECT 2698.000 30.640 2698.260 30.900 ;
      LAYER met2 ;
        RECT 2702.660 34.670 2702.800 54.000 ;
        RECT 2698.000 34.350 2698.260 34.670 ;
        RECT 2702.600 34.350 2702.860 34.670 ;
        RECT 2698.060 30.930 2698.200 34.350 ;
        RECT 2595.420 30.610 2595.680 30.930 ;
        RECT 2698.000 30.610 2698.260 30.930 ;
        RECT 2595.480 2.400 2595.620 30.610 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2632.740 17.440 2643.000 17.580 ;
        RECT 2613.330 17.240 2613.650 17.300 ;
        RECT 2632.740 17.240 2632.880 17.440 ;
        RECT 2613.330 17.100 2632.880 17.240 ;
        RECT 2613.330 17.040 2613.650 17.100 ;
        RECT 2642.860 16.560 2643.000 17.440 ;
        RECT 2673.590 16.560 2673.910 16.620 ;
        RECT 2642.860 16.420 2673.910 16.560 ;
        RECT 2673.590 16.360 2673.910 16.420 ;
      LAYER via ;
        RECT 2613.360 17.040 2613.620 17.300 ;
        RECT 2673.620 16.360 2673.880 16.620 ;
      LAYER met2 ;
        RECT 2613.360 17.010 2613.620 17.330 ;
        RECT 2613.420 2.400 2613.560 17.010 ;
        RECT 2673.680 16.650 2673.820 54.000 ;
        RECT 2673.620 16.330 2673.880 16.650 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2666.230 44.780 2666.550 44.840 ;
        RECT 2714.990 44.780 2715.310 44.840 ;
        RECT 2666.230 44.640 2715.310 44.780 ;
        RECT 2666.230 44.580 2666.550 44.640 ;
        RECT 2714.990 44.580 2715.310 44.640 ;
        RECT 2631.270 17.920 2631.590 17.980 ;
        RECT 2666.230 17.920 2666.550 17.980 ;
        RECT 2631.270 17.780 2666.550 17.920 ;
        RECT 2631.270 17.720 2631.590 17.780 ;
        RECT 2666.230 17.720 2666.550 17.780 ;
      LAYER via ;
        RECT 2666.260 44.580 2666.520 44.840 ;
        RECT 2715.020 44.580 2715.280 44.840 ;
        RECT 2631.300 17.720 2631.560 17.980 ;
        RECT 2666.260 17.720 2666.520 17.980 ;
      LAYER met2 ;
        RECT 2715.080 44.870 2715.220 54.000 ;
        RECT 2666.260 44.550 2666.520 44.870 ;
        RECT 2715.020 44.550 2715.280 44.870 ;
        RECT 2666.320 18.010 2666.460 44.550 ;
        RECT 2631.300 17.690 2631.560 18.010 ;
        RECT 2666.260 17.690 2666.520 18.010 ;
        RECT 2631.360 2.400 2631.500 17.690 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2719.590 17.580 2719.910 17.640 ;
        RECT 2693.000 17.440 2719.910 17.580 ;
        RECT 2693.000 17.240 2693.140 17.440 ;
        RECT 2719.590 17.380 2719.910 17.440 ;
        RECT 2649.300 17.100 2693.140 17.240 ;
        RECT 2649.300 16.960 2649.440 17.100 ;
        RECT 2649.210 16.700 2649.530 16.960 ;
      LAYER via ;
        RECT 2719.620 17.380 2719.880 17.640 ;
        RECT 2649.240 16.700 2649.500 16.960 ;
      LAYER met2 ;
        RECT 2719.680 17.670 2719.820 54.000 ;
        RECT 2719.620 17.350 2719.880 17.670 ;
        RECT 2649.240 16.670 2649.500 16.990 ;
        RECT 2649.300 2.400 2649.440 16.670 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2667.150 17.580 2667.470 17.640 ;
        RECT 2669.910 17.580 2670.230 17.640 ;
        RECT 2667.150 17.440 2670.230 17.580 ;
        RECT 2667.150 17.380 2667.470 17.440 ;
        RECT 2669.910 17.380 2670.230 17.440 ;
      LAYER via ;
        RECT 2667.180 17.380 2667.440 17.640 ;
        RECT 2669.940 17.380 2670.200 17.640 ;
      LAYER met2 ;
        RECT 2670.000 17.670 2670.140 54.000 ;
        RECT 2667.180 17.350 2667.440 17.670 ;
        RECT 2669.940 17.350 2670.200 17.670 ;
        RECT 2667.240 2.400 2667.380 17.350 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2684.630 17.920 2684.950 17.980 ;
        RECT 2721.890 17.920 2722.210 17.980 ;
        RECT 2684.630 17.780 2722.210 17.920 ;
        RECT 2684.630 17.720 2684.950 17.780 ;
        RECT 2721.890 17.720 2722.210 17.780 ;
      LAYER via ;
        RECT 2684.660 17.720 2684.920 17.980 ;
        RECT 2721.920 17.720 2722.180 17.980 ;
      LAYER met2 ;
        RECT 2721.980 18.010 2722.120 54.000 ;
        RECT 2684.660 17.690 2684.920 18.010 ;
        RECT 2721.920 17.690 2722.180 18.010 ;
        RECT 2684.720 2.400 2684.860 17.690 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2702.570 14.520 2702.890 14.580 ;
        RECT 2736.610 14.520 2736.930 14.580 ;
        RECT 2702.570 14.380 2736.930 14.520 ;
        RECT 2702.570 14.320 2702.890 14.380 ;
        RECT 2736.610 14.320 2736.930 14.380 ;
      LAYER via ;
        RECT 2702.600 14.320 2702.860 14.580 ;
        RECT 2736.640 14.320 2736.900 14.580 ;
      LAYER met2 ;
        RECT 2736.700 14.610 2736.840 54.000 ;
        RECT 2702.600 14.290 2702.860 14.610 ;
        RECT 2736.640 14.290 2736.900 14.610 ;
        RECT 2702.660 2.400 2702.800 14.290 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2720.510 18.600 2720.830 18.660 ;
        RECT 2725.110 18.600 2725.430 18.660 ;
        RECT 2720.510 18.460 2725.430 18.600 ;
        RECT 2720.510 18.400 2720.830 18.460 ;
        RECT 2725.110 18.400 2725.430 18.460 ;
      LAYER via ;
        RECT 2720.540 18.400 2720.800 18.660 ;
        RECT 2725.140 18.400 2725.400 18.660 ;
      LAYER met2 ;
        RECT 2725.200 18.690 2725.340 54.000 ;
        RECT 2720.540 18.370 2720.800 18.690 ;
        RECT 2725.140 18.370 2725.400 18.690 ;
        RECT 2720.600 2.400 2720.740 18.370 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2739.000 16.050 2739.140 54.000 ;
        RECT 2738.540 15.910 2739.140 16.050 ;
        RECT 2738.540 2.400 2738.680 15.910 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2754.090 14.180 2754.410 14.240 ;
        RECT 2754.090 14.040 2756.160 14.180 ;
        RECT 2754.090 13.980 2754.410 14.040 ;
        RECT 2756.020 13.900 2756.160 14.040 ;
        RECT 2755.930 13.640 2756.250 13.900 ;
      LAYER via ;
        RECT 2754.120 13.980 2754.380 14.240 ;
        RECT 2755.960 13.640 2756.220 13.900 ;
      LAYER met2 ;
        RECT 2754.180 14.270 2754.320 54.000 ;
        RECT 2754.120 13.950 2754.380 14.270 ;
        RECT 2755.960 13.610 2756.220 13.930 ;
        RECT 2756.020 2.400 2756.160 13.610 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 840.105 4.845 840.275 19.635 ;
      LAYER mcon ;
        RECT 840.105 19.465 840.275 19.635 ;
      LAYER met1 ;
        RECT 840.045 19.620 840.335 19.665 ;
        RECT 1162.490 19.620 1162.810 19.680 ;
        RECT 840.045 19.480 1162.810 19.620 ;
        RECT 840.045 19.435 840.335 19.480 ;
        RECT 1162.490 19.420 1162.810 19.480 ;
        RECT 829.450 5.000 829.770 5.060 ;
        RECT 840.045 5.000 840.335 5.045 ;
        RECT 829.450 4.860 840.335 5.000 ;
        RECT 829.450 4.800 829.770 4.860 ;
        RECT 840.045 4.815 840.335 4.860 ;
      LAYER via ;
        RECT 1162.520 19.420 1162.780 19.680 ;
        RECT 829.480 4.800 829.740 5.060 ;
      LAYER met2 ;
        RECT 1162.580 19.710 1162.720 54.000 ;
        RECT 1162.520 19.390 1162.780 19.710 ;
        RECT 829.480 4.770 829.740 5.090 ;
        RECT 829.540 2.400 829.680 4.770 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2773.870 2.960 2774.190 3.020 ;
        RECT 2774.790 2.960 2775.110 3.020 ;
        RECT 2773.870 2.820 2775.110 2.960 ;
        RECT 2773.870 2.760 2774.190 2.820 ;
        RECT 2774.790 2.760 2775.110 2.820 ;
      LAYER via ;
        RECT 2773.900 2.760 2774.160 3.020 ;
        RECT 2774.820 2.760 2775.080 3.020 ;
      LAYER met2 ;
        RECT 2774.880 3.050 2775.020 54.000 ;
        RECT 2773.900 2.730 2774.160 3.050 ;
        RECT 2774.820 2.730 2775.080 3.050 ;
        RECT 2773.960 2.400 2774.100 2.730 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2777.550 19.960 2777.870 20.020 ;
        RECT 2791.810 19.960 2792.130 20.020 ;
        RECT 2777.550 19.820 2792.130 19.960 ;
        RECT 2777.550 19.760 2777.870 19.820 ;
        RECT 2791.810 19.760 2792.130 19.820 ;
      LAYER via ;
        RECT 2777.580 19.760 2777.840 20.020 ;
        RECT 2791.840 19.760 2792.100 20.020 ;
      LAYER met2 ;
        RECT 2777.640 20.050 2777.780 54.000 ;
        RECT 2777.580 19.730 2777.840 20.050 ;
        RECT 2791.840 19.730 2792.100 20.050 ;
        RECT 2791.900 2.400 2792.040 19.730 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2783.530 17.920 2783.850 17.980 ;
        RECT 2809.750 17.920 2810.070 17.980 ;
        RECT 2783.530 17.780 2810.070 17.920 ;
        RECT 2783.530 17.720 2783.850 17.780 ;
        RECT 2809.750 17.720 2810.070 17.780 ;
      LAYER via ;
        RECT 2783.560 17.720 2783.820 17.980 ;
        RECT 2809.780 17.720 2810.040 17.980 ;
      LAYER met2 ;
        RECT 2783.620 18.010 2783.760 54.000 ;
        RECT 2783.560 17.690 2783.820 18.010 ;
        RECT 2809.780 17.690 2810.040 18.010 ;
        RECT 2809.840 2.400 2809.980 17.690 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2779.850 15.540 2780.170 15.600 ;
        RECT 2827.690 15.540 2828.010 15.600 ;
        RECT 2779.850 15.400 2828.010 15.540 ;
        RECT 2779.850 15.340 2780.170 15.400 ;
        RECT 2827.690 15.340 2828.010 15.400 ;
      LAYER via ;
        RECT 2779.880 15.340 2780.140 15.600 ;
        RECT 2827.720 15.340 2827.980 15.600 ;
      LAYER met2 ;
        RECT 2779.940 15.630 2780.080 54.000 ;
        RECT 2779.880 15.310 2780.140 15.630 ;
        RECT 2827.720 15.310 2827.980 15.630 ;
        RECT 2827.780 2.400 2827.920 15.310 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2787.210 16.560 2787.530 16.620 ;
        RECT 2845.170 16.560 2845.490 16.620 ;
        RECT 2787.210 16.420 2845.490 16.560 ;
        RECT 2787.210 16.360 2787.530 16.420 ;
        RECT 2845.170 16.360 2845.490 16.420 ;
      LAYER via ;
        RECT 2787.240 16.360 2787.500 16.620 ;
        RECT 2845.200 16.360 2845.460 16.620 ;
      LAYER met2 ;
        RECT 2787.300 16.650 2787.440 54.000 ;
        RECT 2787.240 16.330 2787.500 16.650 ;
        RECT 2845.200 16.330 2845.460 16.650 ;
        RECT 2845.260 2.400 2845.400 16.330 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2793.190 20.640 2793.510 20.700 ;
        RECT 2863.110 20.640 2863.430 20.700 ;
        RECT 2793.190 20.500 2863.430 20.640 ;
        RECT 2793.190 20.440 2793.510 20.500 ;
        RECT 2863.110 20.440 2863.430 20.500 ;
      LAYER via ;
        RECT 2793.220 20.440 2793.480 20.700 ;
        RECT 2863.140 20.440 2863.400 20.700 ;
      LAYER met2 ;
        RECT 2793.280 20.730 2793.420 54.000 ;
        RECT 2793.220 20.410 2793.480 20.730 ;
        RECT 2863.140 20.410 2863.400 20.730 ;
        RECT 2863.200 2.400 2863.340 20.410 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2800.550 19.620 2800.870 19.680 ;
        RECT 2881.050 19.620 2881.370 19.680 ;
        RECT 2800.550 19.480 2881.370 19.620 ;
        RECT 2800.550 19.420 2800.870 19.480 ;
        RECT 2881.050 19.420 2881.370 19.480 ;
      LAYER via ;
        RECT 2800.580 19.420 2800.840 19.680 ;
        RECT 2881.080 19.420 2881.340 19.680 ;
      LAYER met2 ;
        RECT 2800.640 19.710 2800.780 54.000 ;
        RECT 2800.580 19.390 2800.840 19.710 ;
        RECT 2881.080 19.390 2881.340 19.710 ;
        RECT 2881.140 2.400 2881.280 19.390 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2898.990 17.240 2899.310 17.300 ;
        RECT 2822.720 17.100 2899.310 17.240 ;
        RECT 2800.090 16.900 2800.410 16.960 ;
        RECT 2822.720 16.900 2822.860 17.100 ;
        RECT 2898.990 17.040 2899.310 17.100 ;
        RECT 2800.090 16.760 2822.860 16.900 ;
        RECT 2800.090 16.700 2800.410 16.760 ;
      LAYER via ;
        RECT 2800.120 16.700 2800.380 16.960 ;
        RECT 2899.020 17.040 2899.280 17.300 ;
      LAYER met2 ;
        RECT 2800.180 16.990 2800.320 54.000 ;
        RECT 2899.020 17.010 2899.280 17.330 ;
        RECT 2800.120 16.670 2800.380 16.990 ;
        RECT 2899.080 2.400 2899.220 17.010 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 911.405 18.105 912.955 18.275 ;
      LAYER mcon ;
        RECT 912.785 18.105 912.955 18.275 ;
      LAYER met1 ;
        RECT 846.930 18.260 847.250 18.320 ;
        RECT 911.345 18.260 911.635 18.305 ;
        RECT 846.930 18.120 911.635 18.260 ;
        RECT 846.930 18.060 847.250 18.120 ;
        RECT 911.345 18.075 911.635 18.120 ;
        RECT 912.725 18.260 913.015 18.305 ;
        RECT 1217.690 18.260 1218.010 18.320 ;
        RECT 912.725 18.120 1218.010 18.260 ;
        RECT 912.725 18.075 913.015 18.120 ;
        RECT 1217.690 18.060 1218.010 18.120 ;
      LAYER via ;
        RECT 846.960 18.060 847.220 18.320 ;
        RECT 1217.720 18.060 1217.980 18.320 ;
      LAYER met2 ;
        RECT 1217.780 18.350 1217.920 54.000 ;
        RECT 846.960 18.030 847.220 18.350 ;
        RECT 1217.720 18.030 1217.980 18.350 ;
        RECT 847.020 2.400 847.160 18.030 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 864.870 20.640 865.190 20.700 ;
        RECT 869.010 20.640 869.330 20.700 ;
        RECT 864.870 20.500 869.330 20.640 ;
        RECT 864.870 20.440 865.190 20.500 ;
        RECT 869.010 20.440 869.330 20.500 ;
      LAYER via ;
        RECT 864.900 20.440 865.160 20.700 ;
        RECT 869.040 20.440 869.300 20.700 ;
      LAYER met2 ;
        RECT 869.100 20.730 869.240 54.000 ;
        RECT 864.900 20.410 865.160 20.730 ;
        RECT 869.040 20.410 869.300 20.730 ;
        RECT 864.960 2.400 865.100 20.410 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.350 18.600 882.670 18.660 ;
        RECT 1252.190 18.600 1252.510 18.660 ;
        RECT 882.350 18.460 1252.510 18.600 ;
        RECT 882.350 18.400 882.670 18.460 ;
        RECT 1252.190 18.400 1252.510 18.460 ;
      LAYER via ;
        RECT 882.380 18.400 882.640 18.660 ;
        RECT 1252.220 18.400 1252.480 18.660 ;
      LAYER met2 ;
        RECT 1252.280 18.690 1252.420 54.000 ;
        RECT 882.380 18.370 882.640 18.690 ;
        RECT 1252.220 18.370 1252.480 18.690 ;
        RECT 882.440 9.250 882.580 18.370 ;
        RECT 882.440 9.110 883.040 9.250 ;
        RECT 882.900 2.400 883.040 9.110 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.750 17.920 901.070 17.980 ;
        RECT 910.870 17.920 911.190 17.980 ;
        RECT 900.750 17.780 911.190 17.920 ;
        RECT 900.750 17.720 901.070 17.780 ;
        RECT 910.870 17.720 911.190 17.780 ;
        RECT 913.170 17.920 913.490 17.980 ;
        RECT 1286.690 17.920 1287.010 17.980 ;
        RECT 913.170 17.780 1287.010 17.920 ;
        RECT 913.170 17.720 913.490 17.780 ;
        RECT 1286.690 17.720 1287.010 17.780 ;
      LAYER via ;
        RECT 900.780 17.720 901.040 17.980 ;
        RECT 910.900 17.720 911.160 17.980 ;
        RECT 913.200 17.720 913.460 17.980 ;
        RECT 1286.720 17.720 1286.980 17.980 ;
      LAYER met2 ;
        RECT 900.780 17.690 901.040 18.010 ;
        RECT 910.890 17.835 911.170 18.205 ;
        RECT 913.190 17.835 913.470 18.205 ;
        RECT 1286.780 18.010 1286.920 54.000 ;
        RECT 910.900 17.690 911.160 17.835 ;
        RECT 913.200 17.690 913.460 17.835 ;
        RECT 1286.720 17.690 1286.980 18.010 ;
        RECT 900.840 2.400 900.980 17.690 ;
        RECT 900.630 -4.800 901.190 2.400 ;
      LAYER via2 ;
        RECT 910.890 17.880 911.170 18.160 ;
        RECT 913.190 17.880 913.470 18.160 ;
      LAYER met3 ;
        RECT 910.865 18.170 911.195 18.185 ;
        RECT 913.165 18.170 913.495 18.185 ;
        RECT 910.865 17.870 913.495 18.170 ;
        RECT 910.865 17.855 911.195 17.870 ;
        RECT 913.165 17.855 913.495 17.870 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 924.285 48.365 924.455 54.000 ;
      LAYER met1 ;
        RECT 924.210 48.520 924.530 48.580 ;
        RECT 924.015 48.380 924.530 48.520 ;
        RECT 924.210 48.320 924.530 48.380 ;
        RECT 918.690 12.480 919.010 12.540 ;
        RECT 924.210 12.480 924.530 12.540 ;
        RECT 918.690 12.340 924.530 12.480 ;
        RECT 918.690 12.280 919.010 12.340 ;
        RECT 924.210 12.280 924.530 12.340 ;
      LAYER via ;
        RECT 924.240 48.320 924.500 48.580 ;
        RECT 918.720 12.280 918.980 12.540 ;
        RECT 924.240 12.280 924.500 12.540 ;
      LAYER met2 ;
        RECT 924.240 48.290 924.500 48.610 ;
        RECT 924.300 12.570 924.440 48.290 ;
        RECT 918.720 12.250 918.980 12.570 ;
        RECT 924.240 12.250 924.500 12.570 ;
        RECT 918.780 2.400 918.920 12.250 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 936.170 18.940 936.490 19.000 ;
        RECT 1307.390 18.940 1307.710 19.000 ;
        RECT 936.170 18.800 1307.710 18.940 ;
        RECT 936.170 18.740 936.490 18.800 ;
        RECT 1307.390 18.740 1307.710 18.800 ;
      LAYER via ;
        RECT 936.200 18.740 936.460 19.000 ;
        RECT 1307.420 18.740 1307.680 19.000 ;
      LAYER met2 ;
        RECT 1307.480 19.030 1307.620 54.000 ;
        RECT 936.200 18.710 936.460 19.030 ;
        RECT 1307.420 18.710 1307.680 19.030 ;
        RECT 936.260 2.400 936.400 18.710 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 954.110 16.900 954.430 16.960 ;
        RECT 958.710 16.900 959.030 16.960 ;
        RECT 954.110 16.760 959.030 16.900 ;
        RECT 954.110 16.700 954.430 16.760 ;
        RECT 958.710 16.700 959.030 16.760 ;
      LAYER via ;
        RECT 954.140 16.700 954.400 16.960 ;
        RECT 958.740 16.700 959.000 16.960 ;
      LAYER met2 ;
        RECT 958.800 16.990 958.940 54.000 ;
        RECT 954.140 16.670 954.400 16.990 ;
        RECT 958.740 16.670 959.000 16.990 ;
        RECT 954.200 2.400 954.340 16.670 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 976.725 16.745 976.895 19.295 ;
      LAYER mcon ;
        RECT 976.725 19.125 976.895 19.295 ;
      LAYER met1 ;
        RECT 976.665 19.280 976.955 19.325 ;
        RECT 1341.890 19.280 1342.210 19.340 ;
        RECT 976.665 19.140 1342.210 19.280 ;
        RECT 976.665 19.095 976.955 19.140 ;
        RECT 1341.890 19.080 1342.210 19.140 ;
        RECT 972.050 16.900 972.370 16.960 ;
        RECT 976.665 16.900 976.955 16.945 ;
        RECT 972.050 16.760 976.955 16.900 ;
        RECT 972.050 16.700 972.370 16.760 ;
        RECT 976.665 16.715 976.955 16.760 ;
      LAYER via ;
        RECT 1341.920 19.080 1342.180 19.340 ;
        RECT 972.080 16.700 972.340 16.960 ;
      LAYER met2 ;
        RECT 1341.980 19.370 1342.120 54.000 ;
        RECT 1341.920 19.050 1342.180 19.370 ;
        RECT 972.080 16.670 972.340 16.990 ;
        RECT 972.140 2.400 972.280 16.670 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 19.280 651.290 19.340 ;
        RECT 655.110 19.280 655.430 19.340 ;
        RECT 650.970 19.140 655.430 19.280 ;
        RECT 650.970 19.080 651.290 19.140 ;
        RECT 655.110 19.080 655.430 19.140 ;
      LAYER via ;
        RECT 651.000 19.080 651.260 19.340 ;
        RECT 655.140 19.080 655.400 19.340 ;
      LAYER met2 ;
        RECT 655.200 19.370 655.340 54.000 ;
        RECT 651.000 19.050 651.260 19.370 ;
        RECT 655.140 19.050 655.400 19.370 ;
        RECT 651.060 2.400 651.200 19.050 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 989.990 24.040 990.310 24.100 ;
        RECT 2184.150 24.040 2184.470 24.100 ;
        RECT 989.990 23.900 2184.470 24.040 ;
        RECT 989.990 23.840 990.310 23.900 ;
        RECT 2184.150 23.840 2184.470 23.900 ;
      LAYER via ;
        RECT 990.020 23.840 990.280 24.100 ;
        RECT 2184.180 23.840 2184.440 24.100 ;
      LAYER met2 ;
        RECT 2184.240 24.130 2184.380 54.000 ;
        RECT 990.020 23.810 990.280 24.130 ;
        RECT 2184.180 23.810 2184.440 24.130 ;
        RECT 990.080 2.400 990.220 23.810 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2187.460 24.325 2187.600 54.000 ;
        RECT 1007.490 23.955 1007.770 24.325 ;
        RECT 2187.390 23.955 2187.670 24.325 ;
        RECT 1007.560 2.400 1007.700 23.955 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER via2 ;
        RECT 1007.490 24.000 1007.770 24.280 ;
        RECT 2187.390 24.000 2187.670 24.280 ;
      LAYER met3 ;
        RECT 1007.465 24.290 1007.795 24.305 ;
        RECT 2187.365 24.290 2187.695 24.305 ;
        RECT 1007.465 23.990 2187.695 24.290 ;
        RECT 1007.465 23.975 1007.795 23.990 ;
        RECT 2187.365 23.975 2187.695 23.990 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2194.360 25.005 2194.500 54.000 ;
        RECT 1025.430 24.635 1025.710 25.005 ;
        RECT 2194.290 24.635 2194.570 25.005 ;
        RECT 1025.500 2.400 1025.640 24.635 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
      LAYER via2 ;
        RECT 1025.430 24.680 1025.710 24.960 ;
        RECT 2194.290 24.680 2194.570 24.960 ;
      LAYER met3 ;
        RECT 1025.405 24.970 1025.735 24.985 ;
        RECT 2194.265 24.970 2194.595 24.985 ;
        RECT 1025.405 24.670 2194.595 24.970 ;
        RECT 1025.405 24.655 1025.735 24.670 ;
        RECT 2194.265 24.655 2194.595 24.670 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.350 24.380 1043.670 24.440 ;
        RECT 2202.090 24.380 2202.410 24.440 ;
        RECT 1043.350 24.240 2202.410 24.380 ;
        RECT 1043.350 24.180 1043.670 24.240 ;
        RECT 2202.090 24.180 2202.410 24.240 ;
      LAYER via ;
        RECT 1043.380 24.180 1043.640 24.440 ;
        RECT 2202.120 24.180 2202.380 24.440 ;
      LAYER met2 ;
        RECT 2202.180 24.470 2202.320 54.000 ;
        RECT 1043.380 24.150 1043.640 24.470 ;
        RECT 2202.120 24.150 2202.380 24.470 ;
        RECT 1043.440 2.400 1043.580 24.150 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2209.080 25.685 2209.220 54.000 ;
        RECT 1061.310 25.315 1061.590 25.685 ;
        RECT 2209.010 25.315 2209.290 25.685 ;
        RECT 1061.380 2.400 1061.520 25.315 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
      LAYER via2 ;
        RECT 1061.310 25.360 1061.590 25.640 ;
        RECT 2209.010 25.360 2209.290 25.640 ;
      LAYER met3 ;
        RECT 1061.285 25.650 1061.615 25.665 ;
        RECT 2208.985 25.650 2209.315 25.665 ;
        RECT 1061.285 25.350 2209.315 25.650 ;
        RECT 1061.285 25.335 1061.615 25.350 ;
        RECT 2208.985 25.335 2209.315 25.350 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.230 25.060 1079.550 25.120 ;
        RECT 2208.530 25.060 2208.850 25.120 ;
        RECT 1079.230 24.920 2208.850 25.060 ;
        RECT 1079.230 24.860 1079.550 24.920 ;
        RECT 2208.530 24.860 2208.850 24.920 ;
      LAYER via ;
        RECT 1079.260 24.860 1079.520 25.120 ;
        RECT 2208.560 24.860 2208.820 25.120 ;
      LAYER met2 ;
        RECT 2208.620 25.150 2208.760 54.000 ;
        RECT 1079.260 24.830 1079.520 25.150 ;
        RECT 2208.560 24.830 2208.820 25.150 ;
        RECT 1079.320 2.400 1079.460 24.830 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 25.400 1097.030 25.460 ;
        RECT 2215.890 25.400 2216.210 25.460 ;
        RECT 1096.710 25.260 2216.210 25.400 ;
        RECT 1096.710 25.200 1097.030 25.260 ;
        RECT 2215.890 25.200 2216.210 25.260 ;
      LAYER via ;
        RECT 1096.740 25.200 1097.000 25.460 ;
        RECT 2215.920 25.200 2216.180 25.460 ;
      LAYER met2 ;
        RECT 2215.980 25.490 2216.120 54.000 ;
        RECT 1096.740 25.170 1097.000 25.490 ;
        RECT 2215.920 25.170 2216.180 25.490 ;
        RECT 1096.800 2.400 1096.940 25.170 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.650 25.740 1114.970 25.800 ;
        RECT 2222.330 25.740 2222.650 25.800 ;
        RECT 1114.650 25.600 2222.650 25.740 ;
        RECT 1114.650 25.540 1114.970 25.600 ;
        RECT 2222.330 25.540 2222.650 25.600 ;
      LAYER via ;
        RECT 1114.680 25.540 1114.940 25.800 ;
        RECT 2222.360 25.540 2222.620 25.800 ;
      LAYER met2 ;
        RECT 2225.180 45.290 2225.320 54.000 ;
        RECT 2222.420 45.150 2225.320 45.290 ;
        RECT 2222.420 25.830 2222.560 45.150 ;
        RECT 1114.680 25.510 1114.940 25.830 ;
        RECT 2222.360 25.510 2222.620 25.830 ;
        RECT 1114.740 2.400 1114.880 25.510 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1132.590 26.080 1132.910 26.140 ;
        RECT 2229.230 26.080 2229.550 26.140 ;
        RECT 1132.590 25.940 2229.550 26.080 ;
        RECT 1132.590 25.880 1132.910 25.940 ;
        RECT 2229.230 25.880 2229.550 25.940 ;
      LAYER via ;
        RECT 1132.620 25.880 1132.880 26.140 ;
        RECT 2229.260 25.880 2229.520 26.140 ;
      LAYER met2 ;
        RECT 2229.320 26.170 2229.460 54.000 ;
        RECT 1132.620 25.850 1132.880 26.170 ;
        RECT 2229.260 25.850 2229.520 26.170 ;
        RECT 1132.680 2.400 1132.820 25.850 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1150.530 26.420 1150.850 26.480 ;
        RECT 2236.590 26.420 2236.910 26.480 ;
        RECT 1150.530 26.280 2236.910 26.420 ;
        RECT 1150.530 26.220 1150.850 26.280 ;
        RECT 2236.590 26.220 2236.910 26.280 ;
      LAYER via ;
        RECT 1150.560 26.220 1150.820 26.480 ;
        RECT 2236.620 26.220 2236.880 26.480 ;
      LAYER met2 ;
        RECT 2236.680 26.510 2236.820 54.000 ;
        RECT 1150.560 26.190 1150.820 26.510 ;
        RECT 2236.620 26.190 2236.880 26.510 ;
        RECT 1150.620 2.400 1150.760 26.190 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1640.045 10.285 1641.595 10.455 ;
        RECT 1736.645 10.285 1738.655 10.455 ;
      LAYER mcon ;
        RECT 1641.425 10.285 1641.595 10.455 ;
        RECT 1738.485 10.285 1738.655 10.455 ;
      LAYER met1 ;
        RECT 668.910 10.440 669.230 10.500 ;
        RECT 1639.985 10.440 1640.275 10.485 ;
        RECT 668.910 10.300 1640.275 10.440 ;
        RECT 668.910 10.240 669.230 10.300 ;
        RECT 1639.985 10.255 1640.275 10.300 ;
        RECT 1641.365 10.440 1641.655 10.485 ;
        RECT 1736.585 10.440 1736.875 10.485 ;
        RECT 1641.365 10.300 1736.875 10.440 ;
        RECT 1641.365 10.255 1641.655 10.300 ;
        RECT 1736.585 10.255 1736.875 10.300 ;
        RECT 1738.425 10.440 1738.715 10.485 ;
        RECT 1907.690 10.440 1908.010 10.500 ;
        RECT 1738.425 10.300 1908.010 10.440 ;
        RECT 1738.425 10.255 1738.715 10.300 ;
        RECT 1907.690 10.240 1908.010 10.300 ;
        RECT 1931.610 10.440 1931.930 10.500 ;
        RECT 2077.430 10.440 2077.750 10.500 ;
        RECT 1931.610 10.300 2077.750 10.440 ;
        RECT 1931.610 10.240 1931.930 10.300 ;
        RECT 2077.430 10.240 2077.750 10.300 ;
      LAYER via ;
        RECT 668.940 10.240 669.200 10.500 ;
        RECT 1907.720 10.240 1907.980 10.500 ;
        RECT 1931.640 10.240 1931.900 10.500 ;
        RECT 2077.460 10.240 2077.720 10.500 ;
      LAYER met2 ;
        RECT 668.940 10.210 669.200 10.530 ;
        RECT 1907.710 10.355 1907.990 10.725 ;
        RECT 1931.630 10.355 1931.910 10.725 ;
        RECT 2077.520 10.530 2077.660 54.000 ;
        RECT 1907.720 10.210 1907.980 10.355 ;
        RECT 1931.640 10.210 1931.900 10.355 ;
        RECT 2077.460 10.210 2077.720 10.530 ;
        RECT 669.000 2.400 669.140 10.210 ;
        RECT 668.790 -4.800 669.350 2.400 ;
      LAYER via2 ;
        RECT 1907.710 10.400 1907.990 10.680 ;
        RECT 1931.630 10.400 1931.910 10.680 ;
      LAYER met3 ;
        RECT 1907.685 10.690 1908.015 10.705 ;
        RECT 1931.605 10.690 1931.935 10.705 ;
        RECT 1907.685 10.390 1931.935 10.690 ;
        RECT 1907.685 10.375 1908.015 10.390 ;
        RECT 1931.605 10.375 1931.935 10.390 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.470 26.760 1168.790 26.820 ;
        RECT 2243.490 26.760 2243.810 26.820 ;
        RECT 1168.470 26.620 2243.810 26.760 ;
        RECT 1168.470 26.560 1168.790 26.620 ;
        RECT 2243.490 26.560 2243.810 26.620 ;
      LAYER via ;
        RECT 1168.500 26.560 1168.760 26.820 ;
        RECT 2243.520 26.560 2243.780 26.820 ;
      LAYER met2 ;
        RECT 2243.580 26.850 2243.720 54.000 ;
        RECT 1168.500 26.530 1168.760 26.850 ;
        RECT 2243.520 26.530 2243.780 26.850 ;
        RECT 1168.560 2.400 1168.700 26.530 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 27.100 1186.270 27.160 ;
        RECT 2247.630 27.100 2247.950 27.160 ;
        RECT 1185.950 26.960 2247.950 27.100 ;
        RECT 1185.950 26.900 1186.270 26.960 ;
        RECT 2247.630 26.900 2247.950 26.960 ;
      LAYER via ;
        RECT 1185.980 26.900 1186.240 27.160 ;
        RECT 2247.660 26.900 2247.920 27.160 ;
      LAYER met2 ;
        RECT 2247.720 27.190 2247.860 54.000 ;
        RECT 1185.980 26.870 1186.240 27.190 ;
        RECT 2247.660 26.870 2247.920 27.190 ;
        RECT 1186.040 2.400 1186.180 26.870 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 27.440 1204.210 27.500 ;
        RECT 2253.150 27.440 2253.470 27.500 ;
        RECT 1203.890 27.300 2253.470 27.440 ;
        RECT 1203.890 27.240 1204.210 27.300 ;
        RECT 2253.150 27.240 2253.470 27.300 ;
      LAYER via ;
        RECT 1203.920 27.240 1204.180 27.500 ;
        RECT 2253.180 27.240 2253.440 27.500 ;
      LAYER met2 ;
        RECT 2253.240 27.530 2253.380 54.000 ;
        RECT 1203.920 27.210 1204.180 27.530 ;
        RECT 2253.180 27.210 2253.440 27.530 ;
        RECT 1203.980 2.400 1204.120 27.210 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.830 23.700 1222.150 23.760 ;
        RECT 2259.130 23.700 2259.450 23.760 ;
        RECT 1221.830 23.560 2259.450 23.700 ;
        RECT 1221.830 23.500 1222.150 23.560 ;
        RECT 2259.130 23.500 2259.450 23.560 ;
      LAYER via ;
        RECT 1221.860 23.500 1222.120 23.760 ;
        RECT 2259.160 23.500 2259.420 23.760 ;
      LAYER met2 ;
        RECT 2259.220 23.790 2259.360 54.000 ;
        RECT 1221.860 23.470 1222.120 23.790 ;
        RECT 2259.160 23.470 2259.420 23.790 ;
        RECT 1221.920 2.400 1222.060 23.470 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1239.770 23.360 1240.090 23.420 ;
        RECT 2264.650 23.360 2264.970 23.420 ;
        RECT 1239.770 23.220 2264.970 23.360 ;
        RECT 1239.770 23.160 1240.090 23.220 ;
        RECT 2264.650 23.160 2264.970 23.220 ;
      LAYER via ;
        RECT 1239.800 23.160 1240.060 23.420 ;
        RECT 2264.680 23.160 2264.940 23.420 ;
      LAYER met2 ;
        RECT 2264.740 23.450 2264.880 54.000 ;
        RECT 1239.800 23.130 1240.060 23.450 ;
        RECT 2264.680 23.130 2264.940 23.450 ;
        RECT 1239.860 2.400 1240.000 23.130 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1257.250 23.020 1257.570 23.080 ;
        RECT 2270.630 23.020 2270.950 23.080 ;
        RECT 1257.250 22.880 2270.950 23.020 ;
        RECT 1257.250 22.820 1257.570 22.880 ;
        RECT 2270.630 22.820 2270.950 22.880 ;
      LAYER via ;
        RECT 1257.280 22.820 1257.540 23.080 ;
        RECT 2270.660 22.820 2270.920 23.080 ;
      LAYER met2 ;
        RECT 2270.720 23.110 2270.860 54.000 ;
        RECT 1257.280 22.790 1257.540 23.110 ;
        RECT 2270.660 22.790 2270.920 23.110 ;
        RECT 1257.340 2.400 1257.480 22.790 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1275.190 22.680 1275.510 22.740 ;
        RECT 2277.070 22.680 2277.390 22.740 ;
        RECT 1275.190 22.540 2277.390 22.680 ;
        RECT 1275.190 22.480 1275.510 22.540 ;
        RECT 2277.070 22.480 2277.390 22.540 ;
      LAYER via ;
        RECT 1275.220 22.480 1275.480 22.740 ;
        RECT 2277.100 22.480 2277.360 22.740 ;
      LAYER met2 ;
        RECT 2277.160 22.770 2277.300 54.000 ;
        RECT 1275.220 22.450 1275.480 22.770 ;
        RECT 2277.100 22.450 2277.360 22.770 ;
        RECT 1275.280 2.400 1275.420 22.450 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1293.130 17.580 1293.450 17.640 ;
        RECT 1296.810 17.580 1297.130 17.640 ;
        RECT 1293.130 17.440 1297.130 17.580 ;
        RECT 1293.130 17.380 1293.450 17.440 ;
        RECT 1296.810 17.380 1297.130 17.440 ;
      LAYER via ;
        RECT 1293.160 17.380 1293.420 17.640 ;
        RECT 1296.840 17.380 1297.100 17.640 ;
      LAYER met2 ;
        RECT 1296.900 17.670 1297.040 54.000 ;
        RECT 1293.160 17.350 1293.420 17.670 ;
        RECT 1296.840 17.350 1297.100 17.670 ;
        RECT 1293.220 2.400 1293.360 17.350 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.070 13.160 1311.390 13.220 ;
        RECT 2284.430 13.160 2284.750 13.220 ;
        RECT 1311.070 13.020 2284.750 13.160 ;
        RECT 1311.070 12.960 1311.390 13.020 ;
        RECT 2284.430 12.960 2284.750 13.020 ;
      LAYER via ;
        RECT 1311.100 12.960 1311.360 13.220 ;
        RECT 2284.460 12.960 2284.720 13.220 ;
      LAYER met2 ;
        RECT 2284.520 13.250 2284.660 54.000 ;
        RECT 1311.100 12.930 1311.360 13.250 ;
        RECT 2284.460 12.930 2284.720 13.250 ;
        RECT 1311.160 2.400 1311.300 12.930 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1329.010 17.440 1331.630 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
      LAYER via ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1331.340 17.380 1331.600 17.640 ;
      LAYER met2 ;
        RECT 1331.400 17.670 1331.540 54.000 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 714.065 18.105 714.235 19.295 ;
        RECT 738.445 19.125 738.615 20.655 ;
        RECT 814.345 19.125 814.515 19.975 ;
        RECT 834.585 19.125 835.215 19.295 ;
        RECT 919.225 18.785 919.395 24.735 ;
      LAYER mcon ;
        RECT 919.225 24.565 919.395 24.735 ;
        RECT 738.445 20.485 738.615 20.655 ;
        RECT 714.065 19.125 714.235 19.295 ;
        RECT 814.345 19.805 814.515 19.975 ;
        RECT 835.045 19.125 835.215 19.295 ;
      LAYER met1 ;
        RECT 919.165 24.720 919.455 24.765 ;
        RECT 2083.870 24.720 2084.190 24.780 ;
        RECT 919.165 24.580 2084.190 24.720 ;
        RECT 919.165 24.535 919.455 24.580 ;
        RECT 2083.870 24.520 2084.190 24.580 ;
        RECT 738.385 20.640 738.675 20.685 ;
        RECT 738.385 20.500 786.900 20.640 ;
        RECT 738.385 20.455 738.675 20.500 ;
        RECT 786.760 19.960 786.900 20.500 ;
        RECT 814.285 19.960 814.575 20.005 ;
        RECT 786.760 19.820 814.575 19.960 ;
        RECT 814.285 19.775 814.575 19.820 ;
        RECT 714.005 19.280 714.295 19.325 ;
        RECT 738.385 19.280 738.675 19.325 ;
        RECT 714.005 19.140 738.675 19.280 ;
        RECT 714.005 19.095 714.295 19.140 ;
        RECT 738.385 19.095 738.675 19.140 ;
        RECT 814.285 19.280 814.575 19.325 ;
        RECT 834.525 19.280 834.815 19.325 ;
        RECT 814.285 19.140 834.815 19.280 ;
        RECT 814.285 19.095 814.575 19.140 ;
        RECT 834.525 19.095 834.815 19.140 ;
        RECT 834.985 19.280 835.275 19.325 ;
        RECT 834.985 19.140 903.280 19.280 ;
        RECT 834.985 19.095 835.275 19.140 ;
        RECT 903.140 18.940 903.280 19.140 ;
        RECT 919.165 18.940 919.455 18.985 ;
        RECT 903.140 18.800 919.455 18.940 ;
        RECT 919.165 18.755 919.455 18.800 ;
        RECT 686.390 18.260 686.710 18.320 ;
        RECT 714.005 18.260 714.295 18.305 ;
        RECT 686.390 18.120 714.295 18.260 ;
        RECT 686.390 18.060 686.710 18.120 ;
        RECT 714.005 18.075 714.295 18.120 ;
      LAYER via ;
        RECT 2083.900 24.520 2084.160 24.780 ;
        RECT 686.420 18.060 686.680 18.320 ;
      LAYER met2 ;
        RECT 2087.180 43.930 2087.320 54.000 ;
        RECT 2083.960 43.790 2087.320 43.930 ;
        RECT 2083.960 24.810 2084.100 43.790 ;
        RECT 2083.900 24.490 2084.160 24.810 ;
        RECT 686.420 18.030 686.680 18.350 ;
        RECT 686.480 2.400 686.620 18.030 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.490 13.500 1346.810 13.560 ;
        RECT 2299.150 13.500 2299.470 13.560 ;
        RECT 1346.490 13.360 2299.470 13.500 ;
        RECT 1346.490 13.300 1346.810 13.360 ;
        RECT 2299.150 13.300 2299.470 13.360 ;
      LAYER via ;
        RECT 1346.520 13.300 1346.780 13.560 ;
        RECT 2299.180 13.300 2299.440 13.560 ;
      LAYER met2 ;
        RECT 2299.240 13.590 2299.380 54.000 ;
        RECT 1346.520 13.270 1346.780 13.590 ;
        RECT 2299.180 13.270 2299.440 13.590 ;
        RECT 1346.580 2.400 1346.720 13.270 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1365.900 17.410 1366.040 54.000 ;
        RECT 1364.520 17.270 1366.040 17.410 ;
        RECT 1364.520 2.400 1364.660 17.270 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1382.370 10.100 1382.690 10.160 ;
        RECT 2312.030 10.100 2312.350 10.160 ;
        RECT 1382.370 9.960 2312.350 10.100 ;
        RECT 1382.370 9.900 1382.690 9.960 ;
        RECT 2312.030 9.900 2312.350 9.960 ;
      LAYER via ;
        RECT 1382.400 9.900 1382.660 10.160 ;
        RECT 2312.060 9.900 2312.320 10.160 ;
      LAYER met2 ;
        RECT 2312.120 10.190 2312.260 54.000 ;
        RECT 1382.400 9.870 1382.660 10.190 ;
        RECT 2312.060 9.870 2312.320 10.190 ;
        RECT 1382.460 2.400 1382.600 9.870 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.400 2.400 1400.540 54.000 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2319.020 31.805 2319.160 54.000 ;
        RECT 1418.270 31.435 1418.550 31.805 ;
        RECT 2318.950 31.435 2319.230 31.805 ;
        RECT 1418.340 2.400 1418.480 31.435 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
      LAYER via2 ;
        RECT 1418.270 31.480 1418.550 31.760 ;
        RECT 2318.950 31.480 2319.230 31.760 ;
      LAYER met3 ;
        RECT 1418.245 31.770 1418.575 31.785 ;
        RECT 2318.925 31.770 2319.255 31.785 ;
        RECT 1418.245 31.470 2319.255 31.770 ;
        RECT 1418.245 31.455 1418.575 31.470 ;
        RECT 2318.925 31.455 2319.255 31.470 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1435.730 31.520 1436.050 31.580 ;
        RECT 2325.830 31.520 2326.150 31.580 ;
        RECT 1435.730 31.380 2326.150 31.520 ;
        RECT 1435.730 31.320 1436.050 31.380 ;
        RECT 2325.830 31.320 2326.150 31.380 ;
      LAYER via ;
        RECT 1435.760 31.320 1436.020 31.580 ;
        RECT 2325.860 31.320 2326.120 31.580 ;
      LAYER met2 ;
        RECT 2325.920 31.610 2326.060 54.000 ;
        RECT 1435.760 31.290 1436.020 31.610 ;
        RECT 2325.860 31.290 2326.120 31.610 ;
        RECT 1435.820 2.400 1435.960 31.290 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1453.670 31.860 1453.990 31.920 ;
        RECT 2332.730 31.860 2333.050 31.920 ;
        RECT 1453.670 31.720 2333.050 31.860 ;
        RECT 1453.670 31.660 1453.990 31.720 ;
        RECT 2332.730 31.660 2333.050 31.720 ;
      LAYER via ;
        RECT 1453.700 31.660 1453.960 31.920 ;
        RECT 2332.760 31.660 2333.020 31.920 ;
      LAYER met2 ;
        RECT 2332.820 31.950 2332.960 54.000 ;
        RECT 1453.700 31.630 1453.960 31.950 ;
        RECT 2332.760 31.630 2333.020 31.950 ;
        RECT 1453.760 2.400 1453.900 31.630 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.610 32.200 1471.930 32.260 ;
        RECT 2340.090 32.200 2340.410 32.260 ;
        RECT 1471.610 32.060 2340.410 32.200 ;
        RECT 1471.610 32.000 1471.930 32.060 ;
        RECT 2340.090 32.000 2340.410 32.060 ;
      LAYER via ;
        RECT 1471.640 32.000 1471.900 32.260 ;
        RECT 2340.120 32.000 2340.380 32.260 ;
      LAYER met2 ;
        RECT 2340.180 32.290 2340.320 54.000 ;
        RECT 1471.640 31.970 1471.900 32.290 ;
        RECT 2340.120 31.970 2340.380 32.290 ;
        RECT 1471.700 2.400 1471.840 31.970 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1489.550 32.540 1489.870 32.600 ;
        RECT 2346.530 32.540 2346.850 32.600 ;
        RECT 1489.550 32.400 2346.850 32.540 ;
        RECT 1489.550 32.340 1489.870 32.400 ;
        RECT 2346.530 32.340 2346.850 32.400 ;
      LAYER via ;
        RECT 1489.580 32.340 1489.840 32.600 ;
        RECT 2346.560 32.340 2346.820 32.600 ;
      LAYER met2 ;
        RECT 2346.620 32.630 2346.760 54.000 ;
        RECT 1489.580 32.310 1489.840 32.630 ;
        RECT 2346.560 32.310 2346.820 32.630 ;
        RECT 1489.640 2.400 1489.780 32.310 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1507.030 32.880 1507.350 32.940 ;
        RECT 2346.990 32.880 2347.310 32.940 ;
        RECT 1507.030 32.740 2347.310 32.880 ;
        RECT 1507.030 32.680 1507.350 32.740 ;
        RECT 2346.990 32.680 2347.310 32.740 ;
      LAYER via ;
        RECT 1507.060 32.680 1507.320 32.940 ;
        RECT 2347.020 32.680 2347.280 32.940 ;
      LAYER met2 ;
        RECT 2347.080 32.970 2347.220 54.000 ;
        RECT 1507.060 32.650 1507.320 32.970 ;
        RECT 2347.020 32.650 2347.280 32.970 ;
        RECT 1507.120 2.400 1507.260 32.650 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2092.700 31.125 2092.840 54.000 ;
        RECT 704.810 30.755 705.090 31.125 ;
        RECT 2092.630 30.755 2092.910 31.125 ;
        RECT 704.880 14.010 705.020 30.755 ;
        RECT 704.420 13.870 705.020 14.010 ;
        RECT 704.420 2.400 704.560 13.870 ;
        RECT 704.210 -4.800 704.770 2.400 ;
      LAYER via2 ;
        RECT 704.810 30.800 705.090 31.080 ;
        RECT 2092.630 30.800 2092.910 31.080 ;
      LAYER met3 ;
        RECT 704.785 31.090 705.115 31.105 ;
        RECT 2092.605 31.090 2092.935 31.105 ;
        RECT 704.785 30.790 2092.935 31.090 ;
        RECT 704.785 30.775 705.115 30.790 ;
        RECT 2092.605 30.775 2092.935 30.790 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.970 33.220 1525.290 33.280 ;
        RECT 2353.430 33.220 2353.750 33.280 ;
        RECT 1524.970 33.080 2353.750 33.220 ;
        RECT 1524.970 33.020 1525.290 33.080 ;
        RECT 2353.430 33.020 2353.750 33.080 ;
      LAYER via ;
        RECT 1525.000 33.020 1525.260 33.280 ;
        RECT 2353.460 33.020 2353.720 33.280 ;
      LAYER met2 ;
        RECT 2353.520 33.310 2353.660 54.000 ;
        RECT 1525.000 32.990 1525.260 33.310 ;
        RECT 2353.460 32.990 2353.720 33.310 ;
        RECT 1525.060 2.400 1525.200 32.990 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1542.910 33.560 1543.230 33.620 ;
        RECT 2360.790 33.560 2361.110 33.620 ;
        RECT 1542.910 33.420 2361.110 33.560 ;
        RECT 1542.910 33.360 1543.230 33.420 ;
        RECT 2360.790 33.360 2361.110 33.420 ;
      LAYER via ;
        RECT 1542.940 33.360 1543.200 33.620 ;
        RECT 2360.820 33.360 2361.080 33.620 ;
      LAYER met2 ;
        RECT 2360.880 33.650 2361.020 54.000 ;
        RECT 1542.940 33.330 1543.200 33.650 ;
        RECT 2360.820 33.330 2361.080 33.650 ;
        RECT 1543.000 2.400 1543.140 33.330 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1560.850 33.900 1561.170 33.960 ;
        RECT 2367.230 33.900 2367.550 33.960 ;
        RECT 1560.850 33.760 2367.550 33.900 ;
        RECT 1560.850 33.700 1561.170 33.760 ;
        RECT 2367.230 33.700 2367.550 33.760 ;
      LAYER via ;
        RECT 1560.880 33.700 1561.140 33.960 ;
        RECT 2367.260 33.700 2367.520 33.960 ;
      LAYER met2 ;
        RECT 2367.320 33.990 2367.460 54.000 ;
        RECT 1560.880 33.670 1561.140 33.990 ;
        RECT 2367.260 33.670 2367.520 33.990 ;
        RECT 1560.940 2.400 1561.080 33.670 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1578.790 34.240 1579.110 34.300 ;
        RECT 2374.590 34.240 2374.910 34.300 ;
        RECT 1578.790 34.100 2374.910 34.240 ;
        RECT 1578.790 34.040 1579.110 34.100 ;
        RECT 2374.590 34.040 2374.910 34.100 ;
      LAYER via ;
        RECT 1578.820 34.040 1579.080 34.300 ;
        RECT 2374.620 34.040 2374.880 34.300 ;
      LAYER met2 ;
        RECT 2374.680 34.330 2374.820 54.000 ;
        RECT 1578.820 34.010 1579.080 34.330 ;
        RECT 2374.620 34.010 2374.880 34.330 ;
        RECT 1578.880 2.400 1579.020 34.010 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1596.270 30.500 1596.590 30.560 ;
        RECT 2381.030 30.500 2381.350 30.560 ;
        RECT 1596.270 30.360 2381.350 30.500 ;
        RECT 1596.270 30.300 1596.590 30.360 ;
        RECT 2381.030 30.300 2381.350 30.360 ;
      LAYER via ;
        RECT 1596.300 30.300 1596.560 30.560 ;
        RECT 2381.060 30.300 2381.320 30.560 ;
      LAYER met2 ;
        RECT 2381.120 30.590 2381.260 54.000 ;
        RECT 1596.300 30.270 1596.560 30.590 ;
        RECT 2381.060 30.270 2381.320 30.590 ;
        RECT 1596.360 2.400 1596.500 30.270 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 30.160 1614.530 30.220 ;
        RECT 2381.490 30.160 2381.810 30.220 ;
        RECT 1614.210 30.020 2381.810 30.160 ;
        RECT 1614.210 29.960 1614.530 30.020 ;
        RECT 2381.490 29.960 2381.810 30.020 ;
      LAYER via ;
        RECT 1614.240 29.960 1614.500 30.220 ;
        RECT 2381.520 29.960 2381.780 30.220 ;
      LAYER met2 ;
        RECT 2386.180 47.330 2386.320 54.000 ;
        RECT 2381.580 47.190 2386.320 47.330 ;
        RECT 2381.580 30.250 2381.720 47.190 ;
        RECT 1614.240 29.930 1614.500 30.250 ;
        RECT 2381.520 29.930 2381.780 30.250 ;
        RECT 1614.300 2.400 1614.440 29.930 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1632.150 29.820 1632.470 29.880 ;
        RECT 2387.470 29.820 2387.790 29.880 ;
        RECT 1632.150 29.680 2387.790 29.820 ;
        RECT 1632.150 29.620 1632.470 29.680 ;
        RECT 2387.470 29.620 2387.790 29.680 ;
      LAYER via ;
        RECT 1632.180 29.620 1632.440 29.880 ;
        RECT 2387.500 29.620 2387.760 29.880 ;
      LAYER met2 ;
        RECT 2391.700 53.450 2391.840 54.000 ;
        RECT 2387.560 53.310 2391.840 53.450 ;
        RECT 2387.560 29.910 2387.700 53.310 ;
        RECT 1632.180 29.590 1632.440 29.910 ;
        RECT 2387.500 29.590 2387.760 29.910 ;
        RECT 1632.240 2.400 1632.380 29.590 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1650.090 29.480 1650.410 29.540 ;
        RECT 2395.290 29.480 2395.610 29.540 ;
        RECT 1650.090 29.340 2395.610 29.480 ;
        RECT 1650.090 29.280 1650.410 29.340 ;
        RECT 2395.290 29.280 2395.610 29.340 ;
      LAYER via ;
        RECT 1650.120 29.280 1650.380 29.540 ;
        RECT 2395.320 29.280 2395.580 29.540 ;
      LAYER met2 ;
        RECT 2395.380 29.570 2395.520 54.000 ;
        RECT 1650.120 29.250 1650.380 29.570 ;
        RECT 2395.320 29.250 2395.580 29.570 ;
        RECT 1650.180 2.400 1650.320 29.250 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.030 29.140 1668.350 29.200 ;
        RECT 2401.730 29.140 2402.050 29.200 ;
        RECT 1668.030 29.000 2402.050 29.140 ;
        RECT 1668.030 28.940 1668.350 29.000 ;
        RECT 2401.730 28.940 2402.050 29.000 ;
      LAYER via ;
        RECT 1668.060 28.940 1668.320 29.200 ;
        RECT 2401.760 28.940 2402.020 29.200 ;
      LAYER met2 ;
        RECT 2401.820 29.230 2401.960 54.000 ;
        RECT 1668.060 28.910 1668.320 29.230 ;
        RECT 2401.760 28.910 2402.020 29.230 ;
        RECT 1668.120 2.400 1668.260 28.910 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.510 28.800 1685.830 28.860 ;
        RECT 2409.090 28.800 2409.410 28.860 ;
        RECT 1685.510 28.660 2409.410 28.800 ;
        RECT 1685.510 28.600 1685.830 28.660 ;
        RECT 2409.090 28.600 2409.410 28.660 ;
      LAYER via ;
        RECT 1685.540 28.600 1685.800 28.860 ;
        RECT 2409.120 28.600 2409.380 28.860 ;
      LAYER met2 ;
        RECT 2409.180 28.890 2409.320 54.000 ;
        RECT 1685.540 28.570 1685.800 28.890 ;
        RECT 2409.120 28.570 2409.380 28.890 ;
        RECT 1685.600 2.400 1685.740 28.570 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 722.270 30.840 722.590 30.900 ;
        RECT 2098.590 30.840 2098.910 30.900 ;
        RECT 722.270 30.700 2098.910 30.840 ;
        RECT 722.270 30.640 722.590 30.700 ;
        RECT 2098.590 30.640 2098.910 30.700 ;
      LAYER via ;
        RECT 722.300 30.640 722.560 30.900 ;
        RECT 2098.620 30.640 2098.880 30.900 ;
      LAYER met2 ;
        RECT 2098.680 30.930 2098.820 54.000 ;
        RECT 722.300 30.610 722.560 30.930 ;
        RECT 2098.620 30.610 2098.880 30.930 ;
        RECT 722.360 2.400 722.500 30.610 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.450 28.460 1703.770 28.520 ;
        RECT 2416.450 28.460 2416.770 28.520 ;
        RECT 1703.450 28.320 2416.770 28.460 ;
        RECT 1703.450 28.260 1703.770 28.320 ;
        RECT 2416.450 28.260 2416.770 28.320 ;
      LAYER via ;
        RECT 1703.480 28.260 1703.740 28.520 ;
        RECT 2416.480 28.260 2416.740 28.520 ;
      LAYER met2 ;
        RECT 2416.540 28.550 2416.680 54.000 ;
        RECT 1703.480 28.230 1703.740 28.550 ;
        RECT 2416.480 28.230 2416.740 28.550 ;
        RECT 1703.540 2.400 1703.680 28.230 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1721.390 28.120 1721.710 28.180 ;
        RECT 2415.530 28.120 2415.850 28.180 ;
        RECT 1721.390 27.980 2415.850 28.120 ;
        RECT 1721.390 27.920 1721.710 27.980 ;
        RECT 2415.530 27.920 2415.850 27.980 ;
      LAYER via ;
        RECT 1721.420 27.920 1721.680 28.180 ;
        RECT 2415.560 27.920 2415.820 28.180 ;
      LAYER met2 ;
        RECT 2415.620 28.210 2415.760 54.000 ;
        RECT 1721.420 27.890 1721.680 28.210 ;
        RECT 2415.560 27.890 2415.820 28.210 ;
        RECT 1721.480 2.400 1721.620 27.890 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.330 16.900 1739.650 16.960 ;
        RECT 1745.310 16.900 1745.630 16.960 ;
        RECT 1739.330 16.760 1745.630 16.900 ;
        RECT 1739.330 16.700 1739.650 16.760 ;
        RECT 1745.310 16.700 1745.630 16.760 ;
      LAYER via ;
        RECT 1739.360 16.700 1739.620 16.960 ;
        RECT 1745.340 16.700 1745.600 16.960 ;
      LAYER met2 ;
        RECT 1745.400 16.990 1745.540 54.000 ;
        RECT 1739.360 16.670 1739.620 16.990 ;
        RECT 1745.340 16.670 1745.600 16.990 ;
        RECT 1739.420 2.400 1739.560 16.670 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1756.810 16.900 1757.130 16.960 ;
        RECT 1759.110 16.900 1759.430 16.960 ;
        RECT 1756.810 16.760 1759.430 16.900 ;
        RECT 1756.810 16.700 1757.130 16.760 ;
        RECT 1759.110 16.700 1759.430 16.760 ;
      LAYER via ;
        RECT 1756.840 16.700 1757.100 16.960 ;
        RECT 1759.140 16.700 1759.400 16.960 ;
      LAYER met2 ;
        RECT 1759.200 16.990 1759.340 54.000 ;
        RECT 1756.840 16.670 1757.100 16.990 ;
        RECT 1759.140 16.670 1759.400 16.990 ;
        RECT 1756.900 2.400 1757.040 16.670 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1774.750 22.000 1775.070 22.060 ;
        RECT 2436.230 22.000 2436.550 22.060 ;
        RECT 1774.750 21.860 2436.550 22.000 ;
        RECT 1774.750 21.800 1775.070 21.860 ;
        RECT 2436.230 21.800 2436.550 21.860 ;
      LAYER via ;
        RECT 1774.780 21.800 1775.040 22.060 ;
        RECT 2436.260 21.800 2436.520 22.060 ;
      LAYER met2 ;
        RECT 2436.320 22.090 2436.460 54.000 ;
        RECT 1774.780 21.770 1775.040 22.090 ;
        RECT 2436.260 21.770 2436.520 22.090 ;
        RECT 1774.840 2.400 1774.980 21.770 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1793.700 17.410 1793.840 54.000 ;
        RECT 1792.780 17.270 1793.840 17.410 ;
        RECT 1792.780 2.400 1792.920 17.270 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1810.630 8.060 1810.950 8.120 ;
        RECT 2450.490 8.060 2450.810 8.120 ;
        RECT 1810.630 7.920 2450.810 8.060 ;
        RECT 1810.630 7.860 1810.950 7.920 ;
        RECT 2450.490 7.860 2450.810 7.920 ;
      LAYER via ;
        RECT 1810.660 7.860 1810.920 8.120 ;
        RECT 2450.520 7.860 2450.780 8.120 ;
      LAYER met2 ;
        RECT 2450.580 8.150 2450.720 54.000 ;
        RECT 1810.660 7.830 1810.920 8.150 ;
        RECT 2450.520 7.830 2450.780 8.150 ;
        RECT 1810.720 2.400 1810.860 7.830 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1828.570 40.700 1828.890 40.760 ;
        RECT 2454.630 40.700 2454.950 40.760 ;
        RECT 1828.570 40.560 2454.950 40.700 ;
        RECT 1828.570 40.500 1828.890 40.560 ;
        RECT 2454.630 40.500 2454.950 40.560 ;
      LAYER via ;
        RECT 1828.600 40.500 1828.860 40.760 ;
        RECT 2454.660 40.500 2454.920 40.760 ;
      LAYER met2 ;
        RECT 2454.720 40.790 2454.860 54.000 ;
        RECT 1828.600 40.470 1828.860 40.790 ;
        RECT 2454.660 40.470 2454.920 40.790 ;
        RECT 1828.660 2.400 1828.800 40.470 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1846.050 41.040 1846.370 41.100 ;
        RECT 2461.990 41.040 2462.310 41.100 ;
        RECT 1846.050 40.900 2462.310 41.040 ;
        RECT 1846.050 40.840 1846.370 40.900 ;
        RECT 2461.990 40.840 2462.310 40.900 ;
      LAYER via ;
        RECT 1846.080 40.840 1846.340 41.100 ;
        RECT 2462.020 40.840 2462.280 41.100 ;
      LAYER met2 ;
        RECT 2462.080 41.130 2462.220 54.000 ;
        RECT 1846.080 40.810 1846.340 41.130 ;
        RECT 2462.020 40.810 2462.280 41.130 ;
        RECT 1846.140 2.400 1846.280 40.810 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1863.990 41.380 1864.310 41.440 ;
        RECT 2467.510 41.380 2467.830 41.440 ;
        RECT 1863.990 41.240 2467.830 41.380 ;
        RECT 1863.990 41.180 1864.310 41.240 ;
        RECT 2467.510 41.180 2467.830 41.240 ;
      LAYER via ;
        RECT 1864.020 41.180 1864.280 41.440 ;
        RECT 2467.540 41.180 2467.800 41.440 ;
      LAYER met2 ;
        RECT 2467.600 41.470 2467.740 54.000 ;
        RECT 1864.020 41.150 1864.280 41.470 ;
        RECT 2467.540 41.150 2467.800 41.470 ;
        RECT 1864.080 2.400 1864.220 41.150 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2105.580 39.285 2105.720 54.000 ;
        RECT 740.230 38.915 740.510 39.285 ;
        RECT 2105.510 38.915 2105.790 39.285 ;
        RECT 740.300 2.400 740.440 38.915 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 740.230 38.960 740.510 39.240 ;
        RECT 2105.510 38.960 2105.790 39.240 ;
      LAYER met3 ;
        RECT 740.205 39.250 740.535 39.265 ;
        RECT 2105.485 39.250 2105.815 39.265 ;
        RECT 740.205 38.950 2105.815 39.250 ;
        RECT 740.205 38.935 740.535 38.950 ;
        RECT 2105.485 38.935 2105.815 38.950 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1881.930 37.640 1882.250 37.700 ;
        RECT 2473.490 37.640 2473.810 37.700 ;
        RECT 1881.930 37.500 2473.810 37.640 ;
        RECT 1881.930 37.440 1882.250 37.500 ;
        RECT 2473.490 37.440 2473.810 37.500 ;
      LAYER via ;
        RECT 1881.960 37.440 1882.220 37.700 ;
        RECT 2473.520 37.440 2473.780 37.700 ;
      LAYER met2 ;
        RECT 2473.580 37.730 2473.720 54.000 ;
        RECT 1881.960 37.410 1882.220 37.730 ;
        RECT 2473.520 37.410 2473.780 37.730 ;
        RECT 1882.020 2.400 1882.160 37.410 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1899.870 37.300 1900.190 37.360 ;
        RECT 2479.010 37.300 2479.330 37.360 ;
        RECT 1899.870 37.160 2479.330 37.300 ;
        RECT 1899.870 37.100 1900.190 37.160 ;
        RECT 2479.010 37.100 2479.330 37.160 ;
      LAYER via ;
        RECT 1899.900 37.100 1900.160 37.360 ;
        RECT 2479.040 37.100 2479.300 37.360 ;
      LAYER met2 ;
        RECT 2479.100 37.390 2479.240 54.000 ;
        RECT 1899.900 37.070 1900.160 37.390 ;
        RECT 2479.040 37.070 2479.300 37.390 ;
        RECT 1899.960 2.400 1900.100 37.070 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.350 36.960 1917.670 37.020 ;
        RECT 2484.990 36.960 2485.310 37.020 ;
        RECT 1917.350 36.820 2485.310 36.960 ;
        RECT 1917.350 36.760 1917.670 36.820 ;
        RECT 2484.990 36.760 2485.310 36.820 ;
      LAYER via ;
        RECT 1917.380 36.760 1917.640 37.020 ;
        RECT 2485.020 36.760 2485.280 37.020 ;
      LAYER met2 ;
        RECT 2485.080 37.050 2485.220 54.000 ;
        RECT 1917.380 36.730 1917.640 37.050 ;
        RECT 2485.020 36.730 2485.280 37.050 ;
        RECT 1917.440 17.410 1917.580 36.730 ;
        RECT 1917.440 17.270 1918.040 17.410 ;
        RECT 1917.900 2.400 1918.040 17.270 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1935.290 16.220 1935.610 16.280 ;
        RECT 1938.510 16.220 1938.830 16.280 ;
        RECT 1935.290 16.080 1938.830 16.220 ;
        RECT 1935.290 16.020 1935.610 16.080 ;
        RECT 1938.510 16.020 1938.830 16.080 ;
      LAYER via ;
        RECT 1935.320 16.020 1935.580 16.280 ;
        RECT 1938.540 16.020 1938.800 16.280 ;
      LAYER met2 ;
        RECT 1938.600 16.310 1938.740 54.000 ;
        RECT 1935.320 15.990 1935.580 16.310 ;
        RECT 1938.540 15.990 1938.800 16.310 ;
        RECT 1935.380 2.400 1935.520 15.990 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1953.230 36.620 1953.550 36.680 ;
        RECT 2496.490 36.620 2496.810 36.680 ;
        RECT 1953.230 36.480 2496.810 36.620 ;
        RECT 1953.230 36.420 1953.550 36.480 ;
        RECT 2496.490 36.420 2496.810 36.480 ;
      LAYER via ;
        RECT 1953.260 36.420 1953.520 36.680 ;
        RECT 2496.520 36.420 2496.780 36.680 ;
      LAYER met2 ;
        RECT 2496.580 36.710 2496.720 54.000 ;
        RECT 1953.260 36.390 1953.520 36.710 ;
        RECT 2496.520 36.390 2496.780 36.710 ;
        RECT 1953.320 2.400 1953.460 36.390 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1971.170 36.280 1971.490 36.340 ;
        RECT 2502.010 36.280 2502.330 36.340 ;
        RECT 1971.170 36.140 2502.330 36.280 ;
        RECT 1971.170 36.080 1971.490 36.140 ;
        RECT 2502.010 36.080 2502.330 36.140 ;
      LAYER via ;
        RECT 1971.200 36.080 1971.460 36.340 ;
        RECT 2502.040 36.080 2502.300 36.340 ;
      LAYER met2 ;
        RECT 2502.100 36.370 2502.240 54.000 ;
        RECT 1971.200 36.050 1971.460 36.370 ;
        RECT 2502.040 36.050 2502.300 36.370 ;
        RECT 1971.260 2.400 1971.400 36.050 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1989.110 35.940 1989.430 36.000 ;
        RECT 2507.990 35.940 2508.310 36.000 ;
        RECT 1989.110 35.800 2508.310 35.940 ;
        RECT 1989.110 35.740 1989.430 35.800 ;
        RECT 2507.990 35.740 2508.310 35.800 ;
      LAYER via ;
        RECT 1989.140 35.740 1989.400 36.000 ;
        RECT 2508.020 35.740 2508.280 36.000 ;
      LAYER met2 ;
        RECT 2508.080 36.030 2508.220 54.000 ;
        RECT 1989.140 35.710 1989.400 36.030 ;
        RECT 2508.020 35.710 2508.280 36.030 ;
        RECT 1989.200 2.400 1989.340 35.710 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2006.590 35.600 2006.910 35.660 ;
        RECT 2513.510 35.600 2513.830 35.660 ;
        RECT 2006.590 35.460 2513.830 35.600 ;
        RECT 2006.590 35.400 2006.910 35.460 ;
        RECT 2513.510 35.400 2513.830 35.460 ;
      LAYER via ;
        RECT 2006.620 35.400 2006.880 35.660 ;
        RECT 2513.540 35.400 2513.800 35.660 ;
      LAYER met2 ;
        RECT 2513.600 35.690 2513.740 54.000 ;
        RECT 2006.620 35.370 2006.880 35.690 ;
        RECT 2513.540 35.370 2513.800 35.690 ;
        RECT 2006.680 2.400 2006.820 35.370 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2024.530 35.260 2024.850 35.320 ;
        RECT 2519.490 35.260 2519.810 35.320 ;
        RECT 2024.530 35.120 2519.810 35.260 ;
        RECT 2024.530 35.060 2024.850 35.120 ;
        RECT 2519.490 35.060 2519.810 35.120 ;
      LAYER via ;
        RECT 2024.560 35.060 2024.820 35.320 ;
        RECT 2519.520 35.060 2519.780 35.320 ;
      LAYER met2 ;
        RECT 2519.580 35.350 2519.720 54.000 ;
        RECT 2024.560 35.030 2024.820 35.350 ;
        RECT 2519.520 35.030 2519.780 35.350 ;
        RECT 2024.620 2.400 2024.760 35.030 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.470 17.580 2042.790 17.640 ;
        RECT 2048.910 17.580 2049.230 17.640 ;
        RECT 2042.470 17.440 2049.230 17.580 ;
        RECT 2042.470 17.380 2042.790 17.440 ;
        RECT 2048.910 17.380 2049.230 17.440 ;
      LAYER via ;
        RECT 2042.500 17.380 2042.760 17.640 ;
        RECT 2048.940 17.380 2049.200 17.640 ;
      LAYER met2 ;
        RECT 2049.000 17.670 2049.140 54.000 ;
        RECT 2042.500 17.350 2042.760 17.670 ;
        RECT 2048.940 17.350 2049.200 17.670 ;
        RECT 2042.560 2.400 2042.700 17.350 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2111.100 39.965 2111.240 54.000 ;
        RECT 757.710 39.595 757.990 39.965 ;
        RECT 2111.030 39.595 2111.310 39.965 ;
        RECT 757.780 2.400 757.920 39.595 ;
        RECT 757.570 -4.800 758.130 2.400 ;
      LAYER via2 ;
        RECT 757.710 39.640 757.990 39.920 ;
        RECT 2111.030 39.640 2111.310 39.920 ;
      LAYER met3 ;
        RECT 757.685 39.930 758.015 39.945 ;
        RECT 2111.005 39.930 2111.335 39.945 ;
        RECT 757.685 39.630 2111.335 39.930 ;
        RECT 757.685 39.615 758.015 39.630 ;
        RECT 2111.005 39.615 2111.335 39.630 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2060.410 34.920 2060.730 34.980 ;
        RECT 2530.990 34.920 2531.310 34.980 ;
        RECT 2060.410 34.780 2531.310 34.920 ;
        RECT 2060.410 34.720 2060.730 34.780 ;
        RECT 2530.990 34.720 2531.310 34.780 ;
      LAYER via ;
        RECT 2060.440 34.720 2060.700 34.980 ;
        RECT 2531.020 34.720 2531.280 34.980 ;
      LAYER met2 ;
        RECT 2531.080 35.010 2531.220 54.000 ;
        RECT 2060.440 34.690 2060.700 35.010 ;
        RECT 2531.020 34.690 2531.280 35.010 ;
        RECT 2060.500 2.400 2060.640 34.690 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2078.350 17.580 2078.670 17.640 ;
        RECT 2083.410 17.580 2083.730 17.640 ;
        RECT 2078.350 17.440 2083.730 17.580 ;
        RECT 2078.350 17.380 2078.670 17.440 ;
        RECT 2083.410 17.380 2083.730 17.440 ;
      LAYER via ;
        RECT 2078.380 17.380 2078.640 17.640 ;
        RECT 2083.440 17.380 2083.700 17.640 ;
      LAYER met2 ;
        RECT 2083.500 17.670 2083.640 54.000 ;
        RECT 2078.380 17.350 2078.640 17.670 ;
        RECT 2083.440 17.350 2083.700 17.670 ;
        RECT 2078.440 2.400 2078.580 17.350 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2097.300 3.130 2097.440 54.000 ;
        RECT 2095.920 2.990 2097.440 3.130 ;
        RECT 2095.920 2.400 2096.060 2.990 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2113.770 17.580 2114.090 17.640 ;
        RECT 2117.910 17.580 2118.230 17.640 ;
        RECT 2113.770 17.440 2118.230 17.580 ;
        RECT 2113.770 17.380 2114.090 17.440 ;
        RECT 2117.910 17.380 2118.230 17.440 ;
      LAYER via ;
        RECT 2113.800 17.380 2114.060 17.640 ;
        RECT 2117.940 17.380 2118.200 17.640 ;
      LAYER met2 ;
        RECT 2118.000 17.670 2118.140 54.000 ;
        RECT 2113.800 17.350 2114.060 17.670 ;
        RECT 2117.940 17.350 2118.200 17.670 ;
        RECT 2113.860 2.400 2114.000 17.350 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 24.720 2132.030 24.780 ;
        RECT 2554.450 24.720 2554.770 24.780 ;
        RECT 2131.710 24.580 2554.770 24.720 ;
        RECT 2131.710 24.520 2132.030 24.580 ;
        RECT 2554.450 24.520 2554.770 24.580 ;
      LAYER via ;
        RECT 2131.740 24.520 2132.000 24.780 ;
        RECT 2554.480 24.520 2554.740 24.780 ;
      LAYER met2 ;
        RECT 2554.540 24.810 2554.680 54.000 ;
        RECT 2131.740 24.490 2132.000 24.810 ;
        RECT 2554.480 24.490 2554.740 24.810 ;
        RECT 2131.800 2.400 2131.940 24.490 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2149.650 21.320 2149.970 21.380 ;
        RECT 2553.530 21.320 2553.850 21.380 ;
        RECT 2149.650 21.180 2553.850 21.320 ;
        RECT 2149.650 21.120 2149.970 21.180 ;
        RECT 2553.530 21.120 2553.850 21.180 ;
      LAYER via ;
        RECT 2149.680 21.120 2149.940 21.380 ;
        RECT 2553.560 21.120 2553.820 21.380 ;
      LAYER met2 ;
        RECT 2553.620 21.410 2553.760 54.000 ;
        RECT 2149.680 21.090 2149.940 21.410 ;
        RECT 2553.560 21.090 2553.820 21.410 ;
        RECT 2149.740 2.400 2149.880 21.090 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2167.590 20.980 2167.910 21.040 ;
        RECT 2560.430 20.980 2560.750 21.040 ;
        RECT 2167.590 20.840 2560.750 20.980 ;
        RECT 2167.590 20.780 2167.910 20.840 ;
        RECT 2560.430 20.780 2560.750 20.840 ;
      LAYER via ;
        RECT 2167.620 20.780 2167.880 21.040 ;
        RECT 2560.460 20.780 2560.720 21.040 ;
      LAYER met2 ;
        RECT 2563.740 37.810 2563.880 54.000 ;
        RECT 2560.520 37.670 2563.880 37.810 ;
        RECT 2560.520 21.070 2560.660 37.670 ;
        RECT 2167.620 20.750 2167.880 21.070 ;
        RECT 2560.460 20.750 2560.720 21.070 ;
        RECT 2167.680 2.400 2167.820 20.750 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2185.070 24.040 2185.390 24.100 ;
        RECT 2567.790 24.040 2568.110 24.100 ;
        RECT 2185.070 23.900 2568.110 24.040 ;
        RECT 2185.070 23.840 2185.390 23.900 ;
        RECT 2567.790 23.840 2568.110 23.900 ;
      LAYER via ;
        RECT 2185.100 23.840 2185.360 24.100 ;
        RECT 2567.820 23.840 2568.080 24.100 ;
      LAYER met2 ;
        RECT 2567.880 24.130 2568.020 54.000 ;
        RECT 2185.100 23.810 2185.360 24.130 ;
        RECT 2567.820 23.810 2568.080 24.130 ;
        RECT 2185.160 2.400 2185.300 23.810 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2203.010 24.380 2203.330 24.440 ;
        RECT 2575.610 24.380 2575.930 24.440 ;
        RECT 2203.010 24.240 2575.930 24.380 ;
        RECT 2203.010 24.180 2203.330 24.240 ;
        RECT 2575.610 24.180 2575.930 24.240 ;
      LAYER via ;
        RECT 2203.040 24.180 2203.300 24.440 ;
        RECT 2575.640 24.180 2575.900 24.440 ;
      LAYER met2 ;
        RECT 2575.700 24.470 2575.840 54.000 ;
        RECT 2203.040 24.150 2203.300 24.470 ;
        RECT 2575.640 24.150 2575.900 24.470 ;
        RECT 2203.100 2.400 2203.240 24.150 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2220.950 25.060 2221.270 25.120 ;
        RECT 2581.590 25.060 2581.910 25.120 ;
        RECT 2220.950 24.920 2581.910 25.060 ;
        RECT 2220.950 24.860 2221.270 24.920 ;
        RECT 2581.590 24.860 2581.910 24.920 ;
      LAYER via ;
        RECT 2220.980 24.860 2221.240 25.120 ;
        RECT 2581.620 24.860 2581.880 25.120 ;
      LAYER met2 ;
        RECT 2581.680 25.150 2581.820 54.000 ;
        RECT 2220.980 24.830 2221.240 25.150 ;
        RECT 2581.620 24.830 2581.880 25.150 ;
        RECT 2221.040 2.400 2221.180 24.830 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2117.080 40.645 2117.220 54.000 ;
        RECT 775.650 40.275 775.930 40.645 ;
        RECT 2117.010 40.275 2117.290 40.645 ;
        RECT 775.720 2.400 775.860 40.275 ;
        RECT 775.510 -4.800 776.070 2.400 ;
      LAYER via2 ;
        RECT 775.650 40.320 775.930 40.600 ;
        RECT 2117.010 40.320 2117.290 40.600 ;
      LAYER met3 ;
        RECT 775.625 40.610 775.955 40.625 ;
        RECT 2116.985 40.610 2117.315 40.625 ;
        RECT 775.625 40.310 2117.315 40.610 ;
        RECT 775.625 40.295 775.955 40.310 ;
        RECT 2116.985 40.295 2117.315 40.310 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2239.350 25.400 2239.670 25.460 ;
        RECT 2588.490 25.400 2588.810 25.460 ;
        RECT 2239.350 25.260 2588.810 25.400 ;
        RECT 2239.350 25.200 2239.670 25.260 ;
        RECT 2588.490 25.200 2588.810 25.260 ;
      LAYER via ;
        RECT 2239.380 25.200 2239.640 25.460 ;
        RECT 2588.520 25.200 2588.780 25.460 ;
      LAYER met2 ;
        RECT 2588.580 25.490 2588.720 54.000 ;
        RECT 2239.380 25.170 2239.640 25.490 ;
        RECT 2588.520 25.170 2588.780 25.490 ;
        RECT 2239.440 12.820 2239.580 25.170 ;
        RECT 2238.980 12.680 2239.580 12.820 ;
        RECT 2238.980 2.400 2239.120 12.680 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2256.370 25.740 2256.690 25.800 ;
        RECT 2592.630 25.740 2592.950 25.800 ;
        RECT 2256.370 25.600 2592.950 25.740 ;
        RECT 2256.370 25.540 2256.690 25.600 ;
        RECT 2592.630 25.540 2592.950 25.600 ;
      LAYER via ;
        RECT 2256.400 25.540 2256.660 25.800 ;
        RECT 2592.660 25.540 2592.920 25.800 ;
      LAYER met2 ;
        RECT 2592.720 25.830 2592.860 54.000 ;
        RECT 2256.400 25.510 2256.660 25.830 ;
        RECT 2592.660 25.510 2592.920 25.830 ;
        RECT 2256.460 2.400 2256.600 25.510 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2274.310 26.080 2274.630 26.140 ;
        RECT 2598.150 26.080 2598.470 26.140 ;
        RECT 2274.310 25.940 2598.470 26.080 ;
        RECT 2274.310 25.880 2274.630 25.940 ;
        RECT 2598.150 25.880 2598.470 25.940 ;
      LAYER via ;
        RECT 2274.340 25.880 2274.600 26.140 ;
        RECT 2598.180 25.880 2598.440 26.140 ;
      LAYER met2 ;
        RECT 2598.240 26.170 2598.380 54.000 ;
        RECT 2274.340 25.850 2274.600 26.170 ;
        RECT 2598.180 25.850 2598.440 26.170 ;
        RECT 2274.400 2.400 2274.540 25.850 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2292.250 26.420 2292.570 26.480 ;
        RECT 2604.130 26.420 2604.450 26.480 ;
        RECT 2292.250 26.280 2604.450 26.420 ;
        RECT 2292.250 26.220 2292.570 26.280 ;
        RECT 2604.130 26.220 2604.450 26.280 ;
      LAYER via ;
        RECT 2292.280 26.220 2292.540 26.480 ;
        RECT 2604.160 26.220 2604.420 26.480 ;
      LAYER met2 ;
        RECT 2604.220 26.510 2604.360 54.000 ;
        RECT 2292.280 26.190 2292.540 26.510 ;
        RECT 2604.160 26.190 2604.420 26.510 ;
        RECT 2292.340 2.400 2292.480 26.190 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2310.190 26.760 2310.510 26.820 ;
        RECT 2609.650 26.760 2609.970 26.820 ;
        RECT 2310.190 26.620 2609.970 26.760 ;
        RECT 2310.190 26.560 2310.510 26.620 ;
        RECT 2609.650 26.560 2609.970 26.620 ;
      LAYER via ;
        RECT 2310.220 26.560 2310.480 26.820 ;
        RECT 2609.680 26.560 2609.940 26.820 ;
      LAYER met2 ;
        RECT 2609.740 26.850 2609.880 54.000 ;
        RECT 2310.220 26.530 2310.480 26.850 ;
        RECT 2609.680 26.530 2609.940 26.850 ;
        RECT 2310.280 2.400 2310.420 26.530 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2328.130 27.100 2328.450 27.160 ;
        RECT 2616.550 27.100 2616.870 27.160 ;
        RECT 2328.130 26.960 2616.870 27.100 ;
        RECT 2328.130 26.900 2328.450 26.960 ;
        RECT 2616.550 26.900 2616.870 26.960 ;
      LAYER via ;
        RECT 2328.160 26.900 2328.420 27.160 ;
        RECT 2616.580 26.900 2616.840 27.160 ;
      LAYER met2 ;
        RECT 2616.640 27.190 2616.780 54.000 ;
        RECT 2328.160 26.870 2328.420 27.190 ;
        RECT 2616.580 26.870 2616.840 27.190 ;
        RECT 2328.220 2.400 2328.360 26.870 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 27.440 2345.930 27.500 ;
        RECT 2622.530 27.440 2622.850 27.500 ;
        RECT 2345.610 27.300 2622.850 27.440 ;
        RECT 2345.610 27.240 2345.930 27.300 ;
        RECT 2622.530 27.240 2622.850 27.300 ;
      LAYER via ;
        RECT 2345.640 27.240 2345.900 27.500 ;
        RECT 2622.560 27.240 2622.820 27.500 ;
      LAYER met2 ;
        RECT 2622.620 27.530 2622.760 54.000 ;
        RECT 2345.640 27.210 2345.900 27.530 ;
        RECT 2622.560 27.210 2622.820 27.530 ;
        RECT 2345.700 2.400 2345.840 27.210 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2363.550 23.700 2363.870 23.760 ;
        RECT 2622.990 23.700 2623.310 23.760 ;
        RECT 2363.550 23.560 2623.310 23.700 ;
        RECT 2363.550 23.500 2363.870 23.560 ;
        RECT 2622.990 23.500 2623.310 23.560 ;
      LAYER via ;
        RECT 2363.580 23.500 2363.840 23.760 ;
        RECT 2623.020 23.500 2623.280 23.760 ;
      LAYER met2 ;
        RECT 2623.080 23.790 2623.220 54.000 ;
        RECT 2363.580 23.470 2363.840 23.790 ;
        RECT 2623.020 23.470 2623.280 23.790 ;
        RECT 2363.640 2.400 2363.780 23.470 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2381.490 23.360 2381.810 23.420 ;
        RECT 2629.890 23.360 2630.210 23.420 ;
        RECT 2381.490 23.220 2630.210 23.360 ;
        RECT 2381.490 23.160 2381.810 23.220 ;
        RECT 2629.890 23.160 2630.210 23.220 ;
      LAYER via ;
        RECT 2381.520 23.160 2381.780 23.420 ;
        RECT 2629.920 23.160 2630.180 23.420 ;
      LAYER met2 ;
        RECT 2629.980 23.450 2630.120 54.000 ;
        RECT 2381.520 23.130 2381.780 23.450 ;
        RECT 2629.920 23.130 2630.180 23.450 ;
        RECT 2381.580 2.400 2381.720 23.130 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2399.430 23.020 2399.750 23.080 ;
        RECT 2636.330 23.020 2636.650 23.080 ;
        RECT 2399.430 22.880 2636.650 23.020 ;
        RECT 2399.430 22.820 2399.750 22.880 ;
        RECT 2636.330 22.820 2636.650 22.880 ;
      LAYER via ;
        RECT 2399.460 22.820 2399.720 23.080 ;
        RECT 2636.360 22.820 2636.620 23.080 ;
      LAYER met2 ;
        RECT 2636.420 23.110 2636.560 54.000 ;
        RECT 2399.460 22.790 2399.720 23.110 ;
        RECT 2636.360 22.790 2636.620 23.110 ;
        RECT 2399.520 2.400 2399.660 22.790 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2122.600 41.325 2122.740 54.000 ;
        RECT 793.590 40.955 793.870 41.325 ;
        RECT 2122.530 40.955 2122.810 41.325 ;
        RECT 793.660 2.400 793.800 40.955 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 793.590 41.000 793.870 41.280 ;
        RECT 2122.530 41.000 2122.810 41.280 ;
      LAYER met3 ;
        RECT 793.565 41.290 793.895 41.305 ;
        RECT 2122.505 41.290 2122.835 41.305 ;
        RECT 793.565 40.990 2122.835 41.290 ;
        RECT 793.565 40.975 793.895 40.990 ;
        RECT 2122.505 40.975 2122.835 40.990 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2072.920 37.925 2073.060 54.000 ;
        RECT 639.030 37.555 639.310 37.925 ;
        RECT 2072.850 37.555 2073.130 37.925 ;
        RECT 639.100 2.400 639.240 37.555 ;
        RECT 638.890 -4.800 639.450 2.400 ;
      LAYER via2 ;
        RECT 639.030 37.600 639.310 37.880 ;
        RECT 2072.850 37.600 2073.130 37.880 ;
      LAYER met3 ;
        RECT 639.005 37.890 639.335 37.905 ;
        RECT 2072.825 37.890 2073.155 37.905 ;
        RECT 639.005 37.590 2073.155 37.890 ;
        RECT 639.005 37.575 639.335 37.590 ;
        RECT 2072.825 37.575 2073.155 37.590 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2422.890 22.680 2423.210 22.740 ;
        RECT 2643.690 22.680 2644.010 22.740 ;
        RECT 2422.890 22.540 2644.010 22.680 ;
        RECT 2422.890 22.480 2423.210 22.540 ;
        RECT 2643.690 22.480 2644.010 22.540 ;
      LAYER via ;
        RECT 2422.920 22.480 2423.180 22.740 ;
        RECT 2643.720 22.480 2643.980 22.740 ;
      LAYER met2 ;
        RECT 2643.780 22.770 2643.920 54.000 ;
        RECT 2422.920 22.450 2423.180 22.770 ;
        RECT 2643.720 22.450 2643.980 22.770 ;
        RECT 2422.980 2.400 2423.120 22.450 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2650.590 48.520 2650.910 48.580 ;
        RECT 2653.350 48.520 2653.670 48.580 ;
        RECT 2650.590 48.380 2653.670 48.520 ;
        RECT 2650.590 48.320 2650.910 48.380 ;
        RECT 2653.350 48.320 2653.670 48.380 ;
        RECT 2440.830 22.340 2441.150 22.400 ;
        RECT 2650.590 22.340 2650.910 22.400 ;
        RECT 2440.830 22.200 2650.910 22.340 ;
        RECT 2440.830 22.140 2441.150 22.200 ;
        RECT 2650.590 22.140 2650.910 22.200 ;
      LAYER via ;
        RECT 2650.620 48.320 2650.880 48.580 ;
        RECT 2653.380 48.320 2653.640 48.580 ;
        RECT 2440.860 22.140 2441.120 22.400 ;
        RECT 2650.620 22.140 2650.880 22.400 ;
      LAYER met2 ;
        RECT 2653.440 48.610 2653.580 54.000 ;
        RECT 2650.620 48.290 2650.880 48.610 ;
        RECT 2653.380 48.290 2653.640 48.610 ;
        RECT 2650.680 22.430 2650.820 48.290 ;
        RECT 2440.860 22.110 2441.120 22.430 ;
        RECT 2650.620 22.110 2650.880 22.430 ;
        RECT 2440.920 2.400 2441.060 22.110 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2458.770 22.000 2459.090 22.060 ;
        RECT 2657.490 22.000 2657.810 22.060 ;
        RECT 2458.770 21.860 2657.810 22.000 ;
        RECT 2458.770 21.800 2459.090 21.860 ;
        RECT 2657.490 21.800 2657.810 21.860 ;
      LAYER via ;
        RECT 2458.800 21.800 2459.060 22.060 ;
        RECT 2657.520 21.800 2657.780 22.060 ;
      LAYER met2 ;
        RECT 2657.580 22.090 2657.720 54.000 ;
        RECT 2458.800 21.770 2459.060 22.090 ;
        RECT 2657.520 21.770 2657.780 22.090 ;
        RECT 2458.860 2.400 2459.000 21.770 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2476.710 46.820 2477.030 46.880 ;
        RECT 2664.850 46.820 2665.170 46.880 ;
        RECT 2476.710 46.680 2665.170 46.820 ;
        RECT 2476.710 46.620 2477.030 46.680 ;
        RECT 2664.850 46.620 2665.170 46.680 ;
      LAYER via ;
        RECT 2476.740 46.620 2477.000 46.880 ;
        RECT 2664.880 46.620 2665.140 46.880 ;
      LAYER met2 ;
        RECT 2664.940 46.910 2665.080 54.000 ;
        RECT 2476.740 46.590 2477.000 46.910 ;
        RECT 2664.880 46.590 2665.140 46.910 ;
        RECT 2476.800 2.400 2476.940 46.590 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2497.410 52.600 2497.730 52.660 ;
        RECT 2670.830 52.600 2671.150 52.660 ;
        RECT 2497.410 52.460 2671.150 52.600 ;
        RECT 2497.410 52.400 2497.730 52.460 ;
        RECT 2670.830 52.400 2671.150 52.460 ;
        RECT 2494.650 16.900 2494.970 16.960 ;
        RECT 2497.410 16.900 2497.730 16.960 ;
        RECT 2494.650 16.760 2497.730 16.900 ;
        RECT 2494.650 16.700 2494.970 16.760 ;
        RECT 2497.410 16.700 2497.730 16.760 ;
      LAYER via ;
        RECT 2497.440 52.400 2497.700 52.660 ;
        RECT 2670.860 52.400 2671.120 52.660 ;
        RECT 2494.680 16.700 2494.940 16.960 ;
        RECT 2497.440 16.700 2497.700 16.960 ;
      LAYER met2 ;
        RECT 2670.920 52.690 2671.060 54.000 ;
        RECT 2497.440 52.370 2497.700 52.690 ;
        RECT 2670.860 52.370 2671.120 52.690 ;
        RECT 2497.500 16.990 2497.640 52.370 ;
        RECT 2494.680 16.670 2494.940 16.990 ;
        RECT 2497.440 16.670 2497.700 16.990 ;
        RECT 2494.740 2.400 2494.880 16.670 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2512.130 17.580 2512.450 17.640 ;
        RECT 2517.650 17.580 2517.970 17.640 ;
        RECT 2512.130 17.440 2517.970 17.580 ;
        RECT 2512.130 17.380 2512.450 17.440 ;
        RECT 2517.650 17.380 2517.970 17.440 ;
      LAYER via ;
        RECT 2512.160 17.380 2512.420 17.640 ;
        RECT 2517.680 17.380 2517.940 17.640 ;
      LAYER met2 ;
        RECT 2517.740 17.670 2517.880 54.000 ;
        RECT 2512.160 17.350 2512.420 17.670 ;
        RECT 2517.680 17.350 2517.940 17.670 ;
        RECT 2512.220 2.400 2512.360 17.350 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2530.070 32.540 2530.390 32.600 ;
        RECT 2678.190 32.540 2678.510 32.600 ;
        RECT 2530.070 32.400 2678.510 32.540 ;
        RECT 2530.070 32.340 2530.390 32.400 ;
        RECT 2678.190 32.340 2678.510 32.400 ;
      LAYER via ;
        RECT 2530.100 32.340 2530.360 32.600 ;
        RECT 2678.220 32.340 2678.480 32.600 ;
      LAYER met2 ;
        RECT 2678.280 32.630 2678.420 54.000 ;
        RECT 2530.100 32.310 2530.360 32.630 ;
        RECT 2678.220 32.310 2678.480 32.630 ;
        RECT 2530.160 2.400 2530.300 32.310 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2548.010 17.580 2548.330 17.640 ;
        RECT 2552.610 17.580 2552.930 17.640 ;
        RECT 2548.010 17.440 2552.930 17.580 ;
        RECT 2548.010 17.380 2548.330 17.440 ;
        RECT 2552.610 17.380 2552.930 17.440 ;
      LAYER via ;
        RECT 2548.040 17.380 2548.300 17.640 ;
        RECT 2552.640 17.380 2552.900 17.640 ;
      LAYER met2 ;
        RECT 2552.700 17.670 2552.840 54.000 ;
        RECT 2548.040 17.350 2548.300 17.670 ;
        RECT 2552.640 17.350 2552.900 17.670 ;
        RECT 2548.100 2.400 2548.240 17.350 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2565.950 38.320 2566.270 38.380 ;
        RECT 2693.830 38.320 2694.150 38.380 ;
        RECT 2565.950 38.180 2694.150 38.320 ;
        RECT 2565.950 38.120 2566.270 38.180 ;
        RECT 2693.830 38.120 2694.150 38.180 ;
      LAYER via ;
        RECT 2565.980 38.120 2566.240 38.380 ;
        RECT 2693.860 38.120 2694.120 38.380 ;
      LAYER met2 ;
        RECT 2693.920 38.410 2694.060 54.000 ;
        RECT 2565.980 38.090 2566.240 38.410 ;
        RECT 2693.860 38.090 2694.120 38.410 ;
        RECT 2566.040 2.400 2566.180 38.090 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2583.890 20.640 2584.210 20.700 ;
        RECT 2587.110 20.640 2587.430 20.700 ;
        RECT 2583.890 20.500 2587.430 20.640 ;
        RECT 2583.890 20.440 2584.210 20.500 ;
        RECT 2587.110 20.440 2587.430 20.500 ;
      LAYER via ;
        RECT 2583.920 20.440 2584.180 20.700 ;
        RECT 2587.140 20.440 2587.400 20.700 ;
      LAYER met2 ;
        RECT 2587.200 20.730 2587.340 54.000 ;
        RECT 2583.920 20.410 2584.180 20.730 ;
        RECT 2587.140 20.410 2587.400 20.730 ;
        RECT 2583.980 2.400 2584.120 20.410 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 37.980 817.810 38.040 ;
        RECT 2130.330 37.980 2130.650 38.040 ;
        RECT 817.490 37.840 2130.650 37.980 ;
        RECT 817.490 37.780 817.810 37.840 ;
        RECT 2130.330 37.780 2130.650 37.840 ;
      LAYER via ;
        RECT 817.520 37.780 817.780 38.040 ;
        RECT 2130.360 37.780 2130.620 38.040 ;
      LAYER met2 ;
        RECT 2130.420 38.070 2130.560 54.000 ;
        RECT 817.520 37.750 817.780 38.070 ;
        RECT 2130.360 37.750 2130.620 38.070 ;
        RECT 817.580 2.400 817.720 37.750 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2601.370 20.640 2601.690 20.700 ;
        RECT 2607.810 20.640 2608.130 20.700 ;
        RECT 2601.370 20.500 2608.130 20.640 ;
        RECT 2601.370 20.440 2601.690 20.500 ;
        RECT 2607.810 20.440 2608.130 20.500 ;
      LAYER via ;
        RECT 2601.400 20.440 2601.660 20.700 ;
        RECT 2607.840 20.440 2608.100 20.700 ;
      LAYER met2 ;
        RECT 2607.900 20.730 2608.040 54.000 ;
        RECT 2601.400 20.410 2601.660 20.730 ;
        RECT 2607.840 20.410 2608.100 20.730 ;
        RECT 2601.460 2.400 2601.600 20.410 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2619.310 20.640 2619.630 20.700 ;
        RECT 2621.610 20.640 2621.930 20.700 ;
        RECT 2619.310 20.500 2621.930 20.640 ;
        RECT 2619.310 20.440 2619.630 20.500 ;
        RECT 2621.610 20.440 2621.930 20.500 ;
      LAYER via ;
        RECT 2619.340 20.440 2619.600 20.700 ;
        RECT 2621.640 20.440 2621.900 20.700 ;
      LAYER met2 ;
        RECT 2621.700 20.730 2621.840 54.000 ;
        RECT 2619.340 20.410 2619.600 20.730 ;
        RECT 2621.640 20.410 2621.900 20.730 ;
        RECT 2619.400 2.400 2619.540 20.410 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2637.250 17.240 2637.570 17.300 ;
        RECT 2642.310 17.240 2642.630 17.300 ;
        RECT 2637.250 17.100 2642.630 17.240 ;
        RECT 2637.250 17.040 2637.570 17.100 ;
        RECT 2642.310 17.040 2642.630 17.100 ;
      LAYER via ;
        RECT 2637.280 17.040 2637.540 17.300 ;
        RECT 2642.340 17.040 2642.600 17.300 ;
      LAYER met2 ;
        RECT 2642.400 17.330 2642.540 54.000 ;
        RECT 2637.280 17.010 2637.540 17.330 ;
        RECT 2642.340 17.010 2642.600 17.330 ;
        RECT 2637.340 2.400 2637.480 17.010 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2656.200 17.410 2656.340 54.000 ;
        RECT 2655.280 17.270 2656.340 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2672.670 17.580 2672.990 17.640 ;
        RECT 2676.810 17.580 2677.130 17.640 ;
        RECT 2672.670 17.440 2677.130 17.580 ;
        RECT 2672.670 17.380 2672.990 17.440 ;
        RECT 2676.810 17.380 2677.130 17.440 ;
      LAYER via ;
        RECT 2672.700 17.380 2672.960 17.640 ;
        RECT 2676.840 17.380 2677.100 17.640 ;
      LAYER met2 ;
        RECT 2676.900 17.670 2677.040 54.000 ;
        RECT 2672.700 17.350 2672.960 17.670 ;
        RECT 2676.840 17.350 2677.100 17.670 ;
        RECT 2672.760 2.400 2672.900 17.350 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.700 2.400 2690.840 54.000 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2708.550 16.220 2708.870 16.280 ;
        RECT 2740.290 16.220 2740.610 16.280 ;
        RECT 2708.550 16.080 2740.610 16.220 ;
        RECT 2708.550 16.020 2708.870 16.080 ;
        RECT 2740.290 16.020 2740.610 16.080 ;
      LAYER via ;
        RECT 2708.580 16.020 2708.840 16.280 ;
        RECT 2740.320 16.020 2740.580 16.280 ;
      LAYER met2 ;
        RECT 2740.380 16.310 2740.520 54.000 ;
        RECT 2708.580 15.990 2708.840 16.310 ;
        RECT 2740.320 15.990 2740.580 16.310 ;
        RECT 2708.640 2.400 2708.780 15.990 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2726.490 19.280 2726.810 19.340 ;
        RECT 2731.550 19.280 2731.870 19.340 ;
        RECT 2726.490 19.140 2731.870 19.280 ;
        RECT 2726.490 19.080 2726.810 19.140 ;
        RECT 2731.550 19.080 2731.870 19.140 ;
      LAYER via ;
        RECT 2726.520 19.080 2726.780 19.340 ;
        RECT 2731.580 19.080 2731.840 19.340 ;
      LAYER met2 ;
        RECT 2731.640 19.370 2731.780 54.000 ;
        RECT 2726.520 19.050 2726.780 19.370 ;
        RECT 2731.580 19.050 2731.840 19.370 ;
        RECT 2726.580 2.400 2726.720 19.050 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2744.430 48.520 2744.750 48.580 ;
        RECT 2751.330 48.520 2751.650 48.580 ;
        RECT 2744.430 48.380 2751.650 48.520 ;
        RECT 2744.430 48.320 2744.750 48.380 ;
        RECT 2751.330 48.320 2751.650 48.380 ;
      LAYER via ;
        RECT 2744.460 48.320 2744.720 48.580 ;
        RECT 2751.360 48.320 2751.620 48.580 ;
      LAYER met2 ;
        RECT 2751.420 48.610 2751.560 54.000 ;
        RECT 2744.460 48.290 2744.720 48.610 ;
        RECT 2751.360 48.290 2751.620 48.610 ;
        RECT 2744.520 2.400 2744.660 48.290 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2759.610 20.640 2759.930 20.700 ;
        RECT 2761.910 20.640 2762.230 20.700 ;
        RECT 2759.610 20.500 2762.230 20.640 ;
        RECT 2759.610 20.440 2759.930 20.500 ;
        RECT 2761.910 20.440 2762.230 20.500 ;
      LAYER via ;
        RECT 2759.640 20.440 2759.900 20.700 ;
        RECT 2761.940 20.440 2762.200 20.700 ;
      LAYER met2 ;
        RECT 2759.700 20.730 2759.840 54.000 ;
        RECT 2759.640 20.410 2759.900 20.730 ;
        RECT 2761.940 20.410 2762.200 20.730 ;
        RECT 2762.000 2.400 2762.140 20.410 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 835.430 38.320 835.750 38.380 ;
        RECT 2135.850 38.320 2136.170 38.380 ;
        RECT 835.430 38.180 2136.170 38.320 ;
        RECT 835.430 38.120 835.750 38.180 ;
        RECT 2135.850 38.120 2136.170 38.180 ;
      LAYER via ;
        RECT 835.460 38.120 835.720 38.380 ;
        RECT 2135.880 38.120 2136.140 38.380 ;
      LAYER met2 ;
        RECT 2135.940 38.410 2136.080 54.000 ;
        RECT 835.460 38.090 835.720 38.410 ;
        RECT 2135.880 38.090 2136.140 38.410 ;
        RECT 835.520 2.400 835.660 38.090 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.480 14.690 2779.620 54.000 ;
        RECT 2779.480 14.550 2780.080 14.690 ;
        RECT 2779.940 2.400 2780.080 14.550 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2784.910 20.300 2785.230 20.360 ;
        RECT 2797.790 20.300 2798.110 20.360 ;
        RECT 2784.910 20.160 2798.110 20.300 ;
        RECT 2784.910 20.100 2785.230 20.160 ;
        RECT 2797.790 20.100 2798.110 20.160 ;
      LAYER via ;
        RECT 2784.940 20.100 2785.200 20.360 ;
        RECT 2797.820 20.100 2798.080 20.360 ;
      LAYER met2 ;
        RECT 2785.000 20.390 2785.140 54.000 ;
        RECT 2784.940 20.070 2785.200 20.390 ;
        RECT 2797.820 20.070 2798.080 20.390 ;
        RECT 2797.880 2.400 2798.020 20.070 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.820 2.400 2815.960 54.000 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2780.310 15.880 2780.630 15.940 ;
        RECT 2833.670 15.880 2833.990 15.940 ;
        RECT 2780.310 15.740 2833.990 15.880 ;
        RECT 2780.310 15.680 2780.630 15.740 ;
        RECT 2833.670 15.680 2833.990 15.740 ;
      LAYER via ;
        RECT 2780.340 15.680 2780.600 15.940 ;
        RECT 2833.700 15.680 2833.960 15.940 ;
      LAYER met2 ;
        RECT 2780.400 15.970 2780.540 54.000 ;
        RECT 2780.340 15.650 2780.600 15.970 ;
        RECT 2833.700 15.650 2833.960 15.970 ;
        RECT 2833.760 2.400 2833.900 15.650 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2851.150 20.300 2851.470 20.360 ;
        RECT 2798.800 20.160 2851.470 20.300 ;
        RECT 2786.290 19.620 2786.610 19.680 ;
        RECT 2798.800 19.620 2798.940 20.160 ;
        RECT 2851.150 20.100 2851.470 20.160 ;
        RECT 2786.290 19.480 2798.940 19.620 ;
        RECT 2786.290 19.420 2786.610 19.480 ;
      LAYER via ;
        RECT 2786.320 19.420 2786.580 19.680 ;
        RECT 2851.180 20.100 2851.440 20.360 ;
      LAYER met2 ;
        RECT 2786.380 19.710 2786.520 54.000 ;
        RECT 2851.180 20.070 2851.440 20.390 ;
        RECT 2786.320 19.390 2786.580 19.710 ;
        RECT 2851.240 2.400 2851.380 20.070 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2799.245 18.445 2799.415 19.975 ;
      LAYER mcon ;
        RECT 2799.245 19.805 2799.415 19.975 ;
      LAYER met1 ;
        RECT 2799.185 19.960 2799.475 20.005 ;
        RECT 2869.090 19.960 2869.410 20.020 ;
        RECT 2799.185 19.820 2869.410 19.960 ;
        RECT 2799.185 19.775 2799.475 19.820 ;
        RECT 2869.090 19.760 2869.410 19.820 ;
        RECT 2792.730 18.600 2793.050 18.660 ;
        RECT 2799.185 18.600 2799.475 18.645 ;
        RECT 2792.730 18.460 2799.475 18.600 ;
        RECT 2792.730 18.400 2793.050 18.460 ;
        RECT 2799.185 18.415 2799.475 18.460 ;
      LAYER via ;
        RECT 2869.120 19.760 2869.380 20.020 ;
        RECT 2792.760 18.400 2793.020 18.660 ;
      LAYER met2 ;
        RECT 2792.820 18.690 2792.960 54.000 ;
        RECT 2869.120 19.730 2869.380 20.050 ;
        RECT 2792.760 18.370 2793.020 18.690 ;
        RECT 2869.180 2.400 2869.320 19.730 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2798.710 18.940 2799.030 19.000 ;
        RECT 2887.030 18.940 2887.350 19.000 ;
        RECT 2798.710 18.800 2887.350 18.940 ;
        RECT 2798.710 18.740 2799.030 18.800 ;
        RECT 2887.030 18.740 2887.350 18.800 ;
      LAYER via ;
        RECT 2798.740 18.740 2799.000 19.000 ;
        RECT 2887.060 18.740 2887.320 19.000 ;
      LAYER met2 ;
        RECT 2798.800 19.030 2798.940 54.000 ;
        RECT 2798.740 18.710 2799.000 19.030 ;
        RECT 2887.060 18.710 2887.320 19.030 ;
        RECT 2887.120 2.400 2887.260 18.710 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2904.970 17.580 2905.290 17.640 ;
        RECT 2822.260 17.440 2905.290 17.580 ;
        RECT 2807.450 17.240 2807.770 17.300 ;
        RECT 2822.260 17.240 2822.400 17.440 ;
        RECT 2904.970 17.380 2905.290 17.440 ;
        RECT 2807.450 17.100 2822.400 17.240 ;
        RECT 2807.450 17.040 2807.770 17.100 ;
      LAYER via ;
        RECT 2807.480 17.040 2807.740 17.300 ;
        RECT 2905.000 17.380 2905.260 17.640 ;
      LAYER met2 ;
        RECT 2807.540 17.330 2807.680 54.000 ;
        RECT 2905.000 17.350 2905.260 17.670 ;
        RECT 2807.480 17.010 2807.740 17.330 ;
        RECT 2905.060 2.400 2905.200 17.350 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 931.185 16.745 931.355 39.355 ;
      LAYER mcon ;
        RECT 931.185 39.185 931.355 39.355 ;
      LAYER met1 ;
        RECT 931.125 39.340 931.415 39.385 ;
        RECT 2141.830 39.340 2142.150 39.400 ;
        RECT 931.125 39.200 2142.150 39.340 ;
        RECT 931.125 39.155 931.415 39.200 ;
        RECT 2141.830 39.140 2142.150 39.200 ;
        RECT 852.910 16.900 853.230 16.960 ;
        RECT 931.125 16.900 931.415 16.945 ;
        RECT 852.910 16.760 931.415 16.900 ;
        RECT 852.910 16.700 853.230 16.760 ;
        RECT 931.125 16.715 931.415 16.760 ;
      LAYER via ;
        RECT 2141.860 39.140 2142.120 39.400 ;
        RECT 852.940 16.700 853.200 16.960 ;
      LAYER met2 ;
        RECT 2141.920 39.430 2142.060 54.000 ;
        RECT 2141.860 39.110 2142.120 39.430 ;
        RECT 852.940 16.670 853.200 16.990 ;
        RECT 853.000 2.400 853.140 16.670 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 38.660 871.170 38.720 ;
        RECT 2147.350 38.660 2147.670 38.720 ;
        RECT 870.850 38.520 2147.670 38.660 ;
        RECT 870.850 38.460 871.170 38.520 ;
        RECT 2147.350 38.460 2147.670 38.520 ;
      LAYER via ;
        RECT 870.880 38.460 871.140 38.720 ;
        RECT 2147.380 38.460 2147.640 38.720 ;
      LAYER met2 ;
        RECT 2147.440 38.750 2147.580 54.000 ;
        RECT 870.880 38.430 871.140 38.750 ;
        RECT 2147.380 38.430 2147.640 38.750 ;
        RECT 870.940 2.400 871.080 38.430 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 888.790 39.000 889.110 39.060 ;
        RECT 2153.330 39.000 2153.650 39.060 ;
        RECT 888.790 38.860 2153.650 39.000 ;
        RECT 888.790 38.800 889.110 38.860 ;
        RECT 2153.330 38.800 2153.650 38.860 ;
      LAYER via ;
        RECT 888.820 38.800 889.080 39.060 ;
        RECT 2153.360 38.800 2153.620 39.060 ;
      LAYER met2 ;
        RECT 2153.420 39.090 2153.560 54.000 ;
        RECT 888.820 38.770 889.080 39.090 ;
        RECT 2153.360 38.770 2153.620 39.090 ;
        RECT 888.880 2.400 889.020 38.770 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 931.645 16.235 931.815 16.915 ;
        RECT 931.185 16.065 931.815 16.235 ;
      LAYER mcon ;
        RECT 931.645 16.745 931.815 16.915 ;
      LAYER met1 ;
        RECT 977.570 39.680 977.890 39.740 ;
        RECT 2158.850 39.680 2159.170 39.740 ;
        RECT 977.570 39.540 2159.170 39.680 ;
        RECT 977.570 39.480 977.890 39.540 ;
        RECT 2158.850 39.480 2159.170 39.540 ;
        RECT 931.585 16.900 931.875 16.945 ;
        RECT 931.585 16.760 945.600 16.900 ;
        RECT 931.585 16.715 931.875 16.760 ;
        RECT 945.460 16.560 945.600 16.760 ;
        RECT 977.570 16.560 977.890 16.620 ;
        RECT 945.460 16.420 977.890 16.560 ;
        RECT 977.570 16.360 977.890 16.420 ;
        RECT 906.730 16.220 907.050 16.280 ;
        RECT 931.125 16.220 931.415 16.265 ;
        RECT 906.730 16.080 931.415 16.220 ;
        RECT 906.730 16.020 907.050 16.080 ;
        RECT 931.125 16.035 931.415 16.080 ;
      LAYER via ;
        RECT 977.600 39.480 977.860 39.740 ;
        RECT 2158.880 39.480 2159.140 39.740 ;
        RECT 977.600 16.360 977.860 16.620 ;
        RECT 906.760 16.020 907.020 16.280 ;
      LAYER met2 ;
        RECT 2158.940 39.770 2159.080 54.000 ;
        RECT 977.600 39.450 977.860 39.770 ;
        RECT 2158.880 39.450 2159.140 39.770 ;
        RECT 977.660 16.650 977.800 39.450 ;
        RECT 977.600 16.330 977.860 16.650 ;
        RECT 906.760 15.990 907.020 16.310 ;
        RECT 906.820 2.400 906.960 15.990 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 976.265 19.125 976.435 20.655 ;
      LAYER mcon ;
        RECT 976.265 20.485 976.435 20.655 ;
      LAYER met1 ;
        RECT 1104.070 40.020 1104.390 40.080 ;
        RECT 2164.830 40.020 2165.150 40.080 ;
        RECT 1104.070 39.880 2165.150 40.020 ;
        RECT 1104.070 39.820 1104.390 39.880 ;
        RECT 2164.830 39.820 2165.150 39.880 ;
        RECT 976.205 20.640 976.495 20.685 ;
        RECT 1104.070 20.640 1104.390 20.700 ;
        RECT 976.205 20.500 1104.390 20.640 ;
        RECT 976.205 20.455 976.495 20.500 ;
        RECT 1104.070 20.440 1104.390 20.500 ;
        RECT 923.750 19.280 924.070 19.340 ;
        RECT 976.205 19.280 976.495 19.325 ;
        RECT 923.750 19.140 976.495 19.280 ;
        RECT 923.750 19.080 924.070 19.140 ;
        RECT 976.205 19.095 976.495 19.140 ;
      LAYER via ;
        RECT 1104.100 39.820 1104.360 40.080 ;
        RECT 2164.860 39.820 2165.120 40.080 ;
        RECT 1104.100 20.440 1104.360 20.700 ;
        RECT 923.780 19.080 924.040 19.340 ;
      LAYER met2 ;
        RECT 2164.920 40.110 2165.060 54.000 ;
        RECT 1104.100 39.790 1104.360 40.110 ;
        RECT 2164.860 39.790 2165.120 40.110 ;
        RECT 1104.160 20.730 1104.300 39.790 ;
        RECT 1104.100 20.410 1104.360 20.730 ;
        RECT 923.780 19.050 924.040 19.370 ;
        RECT 923.840 9.930 923.980 19.050 ;
        RECT 923.840 9.790 924.440 9.930 ;
        RECT 924.300 2.400 924.440 9.790 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 942.150 16.560 942.470 16.620 ;
        RECT 944.910 16.560 945.230 16.620 ;
        RECT 942.150 16.420 945.230 16.560 ;
        RECT 942.150 16.360 942.470 16.420 ;
        RECT 944.910 16.360 945.230 16.420 ;
      LAYER via ;
        RECT 942.180 16.360 942.440 16.620 ;
        RECT 944.940 16.360 945.200 16.620 ;
      LAYER met2 ;
        RECT 945.000 16.650 945.140 54.000 ;
        RECT 942.180 16.330 942.440 16.650 ;
        RECT 944.940 16.330 945.200 16.650 ;
        RECT 942.240 2.400 942.380 16.330 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1737.105 10.625 1738.195 10.795 ;
        RECT 1929.845 10.625 1931.395 10.795 ;
      LAYER mcon ;
        RECT 1738.025 10.625 1738.195 10.795 ;
        RECT 1931.225 10.625 1931.395 10.795 ;
      LAYER met1 ;
        RECT 960.090 10.780 960.410 10.840 ;
        RECT 1737.045 10.780 1737.335 10.825 ;
        RECT 960.090 10.640 1737.335 10.780 ;
        RECT 960.090 10.580 960.410 10.640 ;
        RECT 1737.045 10.595 1737.335 10.640 ;
        RECT 1737.965 10.780 1738.255 10.825 ;
        RECT 1929.785 10.780 1930.075 10.825 ;
        RECT 1737.965 10.640 1930.075 10.780 ;
        RECT 1737.965 10.595 1738.255 10.640 ;
        RECT 1929.785 10.595 1930.075 10.640 ;
        RECT 1931.165 10.780 1931.455 10.825 ;
        RECT 2174.490 10.780 2174.810 10.840 ;
        RECT 1931.165 10.640 2174.810 10.780 ;
        RECT 1931.165 10.595 1931.455 10.640 ;
        RECT 2174.490 10.580 2174.810 10.640 ;
      LAYER via ;
        RECT 960.120 10.580 960.380 10.840 ;
        RECT 2174.520 10.580 2174.780 10.840 ;
      LAYER met2 ;
        RECT 2177.340 49.485 2177.480 54.000 ;
        RECT 2177.270 49.115 2177.550 49.485 ;
        RECT 2174.050 48.435 2174.330 48.805 ;
        RECT 2174.120 48.010 2174.260 48.435 ;
        RECT 2174.120 47.870 2174.720 48.010 ;
        RECT 2174.580 10.870 2174.720 47.870 ;
        RECT 960.120 10.550 960.380 10.870 ;
        RECT 2174.520 10.550 2174.780 10.870 ;
        RECT 960.180 2.400 960.320 10.550 ;
        RECT 959.970 -4.800 960.530 2.400 ;
      LAYER via2 ;
        RECT 2177.270 49.160 2177.550 49.440 ;
        RECT 2174.050 48.480 2174.330 48.760 ;
      LAYER met3 ;
        RECT 2177.245 49.450 2177.575 49.465 ;
        RECT 2173.350 49.150 2177.575 49.450 ;
        RECT 2173.350 48.770 2173.650 49.150 ;
        RECT 2177.245 49.135 2177.575 49.150 ;
        RECT 2174.025 48.770 2174.355 48.785 ;
        RECT 2173.350 48.470 2174.355 48.770 ;
        RECT 2174.025 48.455 2174.355 48.470 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.500 3.130 979.640 54.000 ;
        RECT 978.120 2.990 979.640 3.130 ;
        RECT 978.120 2.400 978.260 2.990 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2078.440 38.605 2078.580 54.000 ;
        RECT 656.970 38.235 657.250 38.605 ;
        RECT 2078.370 38.235 2078.650 38.605 ;
        RECT 657.040 2.400 657.180 38.235 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 656.970 38.280 657.250 38.560 ;
        RECT 2078.370 38.280 2078.650 38.560 ;
      LAYER met3 ;
        RECT 656.945 38.570 657.275 38.585 ;
        RECT 2078.345 38.570 2078.675 38.585 ;
        RECT 656.945 38.270 2078.675 38.570 ;
        RECT 656.945 38.255 657.275 38.270 ;
        RECT 2078.345 38.255 2078.675 38.270 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1640.505 10.965 1641.135 11.135 ;
        RECT 1930.305 10.965 1930.935 11.135 ;
      LAYER mcon ;
        RECT 1640.965 10.965 1641.135 11.135 ;
        RECT 1930.765 10.965 1930.935 11.135 ;
      LAYER met1 ;
        RECT 1737.030 11.260 1737.350 11.520 ;
        RECT 995.970 11.120 996.290 11.180 ;
        RECT 1640.445 11.120 1640.735 11.165 ;
        RECT 995.970 10.980 1640.735 11.120 ;
        RECT 995.970 10.920 996.290 10.980 ;
        RECT 1640.445 10.935 1640.735 10.980 ;
        RECT 1640.905 11.120 1641.195 11.165 ;
        RECT 1737.120 11.120 1737.260 11.260 ;
        RECT 1640.905 10.980 1737.260 11.120 ;
        RECT 1738.410 11.120 1738.730 11.180 ;
        RECT 1930.245 11.120 1930.535 11.165 ;
        RECT 1738.410 10.980 1930.535 11.120 ;
        RECT 1640.905 10.935 1641.195 10.980 ;
        RECT 1738.410 10.920 1738.730 10.980 ;
        RECT 1930.245 10.935 1930.535 10.980 ;
        RECT 1930.705 11.120 1930.995 11.165 ;
        RECT 2188.750 11.120 2189.070 11.180 ;
        RECT 1930.705 10.980 2189.070 11.120 ;
        RECT 1930.705 10.935 1930.995 10.980 ;
        RECT 2188.750 10.920 2189.070 10.980 ;
      LAYER via ;
        RECT 1737.060 11.260 1737.320 11.520 ;
        RECT 996.000 10.920 996.260 11.180 ;
        RECT 1738.440 10.920 1738.700 11.180 ;
        RECT 2188.780 10.920 2189.040 11.180 ;
      LAYER met2 ;
        RECT 1737.060 11.230 1737.320 11.550 ;
        RECT 996.000 10.890 996.260 11.210 ;
        RECT 996.060 2.400 996.200 10.890 ;
        RECT 1737.120 10.610 1737.260 11.230 ;
        RECT 2188.840 11.210 2188.980 54.000 ;
        RECT 1738.440 10.890 1738.700 11.210 ;
        RECT 2188.780 10.890 2189.040 11.210 ;
        RECT 1738.500 10.610 1738.640 10.890 ;
        RECT 1737.120 10.470 1738.640 10.610 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1013.985 2.805 1014.155 48.195 ;
      LAYER mcon ;
        RECT 1013.985 48.025 1014.155 48.195 ;
      LAYER met1 ;
        RECT 1013.910 48.180 1014.230 48.240 ;
        RECT 1013.715 48.040 1014.230 48.180 ;
        RECT 1013.910 47.980 1014.230 48.040 ;
        RECT 1013.450 2.960 1013.770 3.020 ;
        RECT 1013.925 2.960 1014.215 3.005 ;
        RECT 1013.450 2.820 1014.215 2.960 ;
        RECT 1013.450 2.760 1013.770 2.820 ;
        RECT 1013.925 2.775 1014.215 2.820 ;
      LAYER via ;
        RECT 1013.940 47.980 1014.200 48.240 ;
        RECT 1013.480 2.760 1013.740 3.020 ;
      LAYER met2 ;
        RECT 1014.000 48.270 1014.140 54.000 ;
        RECT 1013.940 47.950 1014.200 48.270 ;
        RECT 1013.480 2.730 1013.740 3.050 ;
        RECT 1013.540 2.400 1013.680 2.730 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2199.420 46.085 2199.560 54.000 ;
        RECT 1031.410 45.715 1031.690 46.085 ;
        RECT 2199.350 45.715 2199.630 46.085 ;
        RECT 1031.480 2.400 1031.620 45.715 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
      LAYER via2 ;
        RECT 1031.410 45.760 1031.690 46.040 ;
        RECT 2199.350 45.760 2199.630 46.040 ;
      LAYER met3 ;
        RECT 1031.385 46.050 1031.715 46.065 ;
        RECT 2199.325 46.050 2199.655 46.065 ;
        RECT 1031.385 45.750 2199.655 46.050 ;
        RECT 1031.385 45.735 1031.715 45.750 ;
        RECT 2199.325 45.735 2199.655 45.750 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.330 44.780 1049.650 44.840 ;
        RECT 2204.850 44.780 2205.170 44.840 ;
        RECT 1049.330 44.640 2205.170 44.780 ;
        RECT 1049.330 44.580 1049.650 44.640 ;
        RECT 2204.850 44.580 2205.170 44.640 ;
      LAYER via ;
        RECT 1049.360 44.580 1049.620 44.840 ;
        RECT 2204.880 44.580 2205.140 44.840 ;
      LAYER met2 ;
        RECT 2204.940 44.870 2205.080 54.000 ;
        RECT 1049.360 44.550 1049.620 44.870 ;
        RECT 2204.880 44.550 2205.140 44.870 ;
        RECT 1049.420 2.400 1049.560 44.550 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1067.270 45.120 1067.590 45.180 ;
        RECT 2210.830 45.120 2211.150 45.180 ;
        RECT 1067.270 44.980 2211.150 45.120 ;
        RECT 1067.270 44.920 1067.590 44.980 ;
        RECT 2210.830 44.920 2211.150 44.980 ;
      LAYER via ;
        RECT 1067.300 44.920 1067.560 45.180 ;
        RECT 2210.860 44.920 2211.120 45.180 ;
      LAYER met2 ;
        RECT 2210.920 45.210 2211.060 54.000 ;
        RECT 1067.300 44.890 1067.560 45.210 ;
        RECT 2210.860 44.890 2211.120 45.210 ;
        RECT 1067.360 2.400 1067.500 44.890 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1085.210 45.460 1085.530 45.520 ;
        RECT 2214.970 45.460 2215.290 45.520 ;
        RECT 1085.210 45.320 2215.290 45.460 ;
        RECT 1085.210 45.260 1085.530 45.320 ;
        RECT 2214.970 45.260 2215.290 45.320 ;
      LAYER via ;
        RECT 1085.240 45.260 1085.500 45.520 ;
        RECT 2215.000 45.260 2215.260 45.520 ;
      LAYER met2 ;
        RECT 2215.060 45.550 2215.200 54.000 ;
        RECT 1085.240 45.230 1085.500 45.550 ;
        RECT 2215.000 45.230 2215.260 45.550 ;
        RECT 1085.300 2.400 1085.440 45.230 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1102.690 45.800 1103.010 45.860 ;
        RECT 2222.330 45.800 2222.650 45.860 ;
        RECT 1102.690 45.660 2222.650 45.800 ;
        RECT 1102.690 45.600 1103.010 45.660 ;
        RECT 2222.330 45.600 2222.650 45.660 ;
      LAYER via ;
        RECT 1102.720 45.600 1102.980 45.860 ;
        RECT 2222.360 45.600 2222.620 45.860 ;
      LAYER met2 ;
        RECT 2222.420 45.890 2222.560 54.000 ;
        RECT 1102.720 45.570 1102.980 45.890 ;
        RECT 2222.360 45.570 2222.620 45.890 ;
        RECT 1102.780 2.400 1102.920 45.570 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2227.850 46.480 2228.170 46.540 ;
        RECT 2217.820 46.340 2228.170 46.480 ;
        RECT 1120.630 46.140 1120.950 46.200 ;
        RECT 2217.820 46.140 2217.960 46.340 ;
        RECT 2227.850 46.280 2228.170 46.340 ;
        RECT 1120.630 46.000 2217.960 46.140 ;
        RECT 1120.630 45.940 1120.950 46.000 ;
      LAYER via ;
        RECT 1120.660 45.940 1120.920 46.200 ;
        RECT 2227.880 46.280 2228.140 46.540 ;
      LAYER met2 ;
        RECT 2227.940 46.570 2228.080 54.000 ;
        RECT 2227.880 46.250 2228.140 46.570 ;
        RECT 1120.660 45.910 1120.920 46.230 ;
        RECT 1120.720 2.400 1120.860 45.910 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2233.830 46.820 2234.150 46.880 ;
        RECT 2217.360 46.680 2234.150 46.820 ;
        RECT 1138.570 46.480 1138.890 46.540 ;
        RECT 2217.360 46.480 2217.500 46.680 ;
        RECT 2233.830 46.620 2234.150 46.680 ;
        RECT 1138.570 46.340 2217.500 46.480 ;
        RECT 1138.570 46.280 1138.890 46.340 ;
      LAYER via ;
        RECT 1138.600 46.280 1138.860 46.540 ;
        RECT 2233.860 46.620 2234.120 46.880 ;
      LAYER met2 ;
        RECT 2233.920 46.910 2234.060 54.000 ;
        RECT 2233.860 46.590 2234.120 46.910 ;
        RECT 1138.600 46.250 1138.860 46.570 ;
        RECT 1138.660 2.400 1138.800 46.250 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2239.350 47.160 2239.670 47.220 ;
        RECT 2216.900 47.020 2239.670 47.160 ;
        RECT 1156.510 46.820 1156.830 46.880 ;
        RECT 2216.900 46.820 2217.040 47.020 ;
        RECT 2239.350 46.960 2239.670 47.020 ;
        RECT 1156.510 46.680 2217.040 46.820 ;
        RECT 1156.510 46.620 1156.830 46.680 ;
      LAYER via ;
        RECT 1156.540 46.620 1156.800 46.880 ;
        RECT 2239.380 46.960 2239.640 47.220 ;
      LAYER met2 ;
        RECT 2239.440 47.250 2239.580 54.000 ;
        RECT 2239.380 46.930 2239.640 47.250 ;
        RECT 1156.540 46.590 1156.800 46.910 ;
        RECT 1156.600 2.400 1156.740 46.590 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.420 44.725 2084.560 54.000 ;
        RECT 674.450 44.355 674.730 44.725 ;
        RECT 2084.350 44.355 2084.630 44.725 ;
        RECT 674.520 2.400 674.660 44.355 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 674.450 44.400 674.730 44.680 ;
        RECT 2084.350 44.400 2084.630 44.680 ;
      LAYER met3 ;
        RECT 674.425 44.690 674.755 44.705 ;
        RECT 2084.325 44.690 2084.655 44.705 ;
        RECT 674.425 44.390 2084.655 44.690 ;
        RECT 674.425 44.375 674.755 44.390 ;
        RECT 2084.325 44.375 2084.655 44.390 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2243.950 47.500 2244.270 47.560 ;
        RECT 2216.440 47.360 2244.270 47.500 ;
        RECT 1173.990 47.160 1174.310 47.220 ;
        RECT 2216.440 47.160 2216.580 47.360 ;
        RECT 2243.950 47.300 2244.270 47.360 ;
        RECT 1173.990 47.020 2216.580 47.160 ;
        RECT 1173.990 46.960 1174.310 47.020 ;
      LAYER via ;
        RECT 1174.020 46.960 1174.280 47.220 ;
        RECT 2243.980 47.300 2244.240 47.560 ;
      LAYER met2 ;
        RECT 2244.040 47.590 2244.180 54.000 ;
        RECT 2243.980 47.270 2244.240 47.590 ;
        RECT 1174.020 46.930 1174.280 47.250 ;
        RECT 1174.080 2.400 1174.220 46.930 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2215.965 45.305 2216.135 47.515 ;
      LAYER mcon ;
        RECT 2215.965 47.345 2216.135 47.515 ;
      LAYER met1 ;
        RECT 1191.930 47.500 1192.250 47.560 ;
        RECT 2215.905 47.500 2216.195 47.545 ;
        RECT 1191.930 47.360 2216.195 47.500 ;
        RECT 1191.930 47.300 1192.250 47.360 ;
        RECT 2215.905 47.315 2216.195 47.360 ;
        RECT 2215.905 45.460 2216.195 45.505 ;
        RECT 2250.850 45.460 2251.170 45.520 ;
        RECT 2215.905 45.320 2251.170 45.460 ;
        RECT 2215.905 45.275 2216.195 45.320 ;
        RECT 2250.850 45.260 2251.170 45.320 ;
      LAYER via ;
        RECT 1191.960 47.300 1192.220 47.560 ;
        RECT 2250.880 45.260 2251.140 45.520 ;
      LAYER met2 ;
        RECT 1191.960 47.270 1192.220 47.590 ;
        RECT 1192.020 2.400 1192.160 47.270 ;
        RECT 2250.940 45.550 2251.080 54.000 ;
        RECT 2250.880 45.230 2251.140 45.550 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1209.870 47.840 1210.190 47.900 ;
        RECT 2256.370 47.840 2256.690 47.900 ;
        RECT 1209.870 47.700 2256.690 47.840 ;
        RECT 1209.870 47.640 1210.190 47.700 ;
        RECT 2256.370 47.640 2256.690 47.700 ;
      LAYER via ;
        RECT 1209.900 47.640 1210.160 47.900 ;
        RECT 2256.400 47.640 2256.660 47.900 ;
      LAYER met2 ;
        RECT 2256.460 47.930 2256.600 54.000 ;
        RECT 1209.900 47.610 1210.160 47.930 ;
        RECT 2256.400 47.610 2256.660 47.930 ;
        RECT 1209.960 2.400 1210.100 47.610 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 48.180 1228.130 48.240 ;
        RECT 1227.810 48.040 2257.060 48.180 ;
        RECT 1227.810 47.980 1228.130 48.040 ;
        RECT 2256.920 47.840 2257.060 48.040 ;
        RECT 2262.350 47.840 2262.670 47.900 ;
        RECT 2256.920 47.700 2262.670 47.840 ;
        RECT 2262.350 47.640 2262.670 47.700 ;
      LAYER via ;
        RECT 1227.840 47.980 1228.100 48.240 ;
        RECT 2262.380 47.640 2262.640 47.900 ;
      LAYER met2 ;
        RECT 1227.840 47.950 1228.100 48.270 ;
        RECT 1227.900 2.400 1228.040 47.950 ;
        RECT 2262.440 47.930 2262.580 54.000 ;
        RECT 2262.380 47.610 2262.640 47.930 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.750 44.440 1246.070 44.500 ;
        RECT 2268.330 44.440 2268.650 44.500 ;
        RECT 1245.750 44.300 2268.650 44.440 ;
        RECT 1245.750 44.240 1246.070 44.300 ;
        RECT 2268.330 44.240 2268.650 44.300 ;
      LAYER via ;
        RECT 1245.780 44.240 1246.040 44.500 ;
        RECT 2268.360 44.240 2268.620 44.500 ;
      LAYER met2 ;
        RECT 2268.420 44.530 2268.560 54.000 ;
        RECT 1245.780 44.210 1246.040 44.530 ;
        RECT 2268.360 44.210 2268.620 44.530 ;
        RECT 1245.840 2.400 1245.980 44.210 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1263.230 44.100 1263.550 44.160 ;
        RECT 2273.850 44.100 2274.170 44.160 ;
        RECT 1263.230 43.960 2274.170 44.100 ;
        RECT 1263.230 43.900 1263.550 43.960 ;
        RECT 2273.850 43.900 2274.170 43.960 ;
      LAYER via ;
        RECT 1263.260 43.900 1263.520 44.160 ;
        RECT 2273.880 43.900 2274.140 44.160 ;
      LAYER met2 ;
        RECT 2273.940 44.190 2274.080 54.000 ;
        RECT 1263.260 43.870 1263.520 44.190 ;
        RECT 2273.880 43.870 2274.140 44.190 ;
        RECT 1263.320 2.400 1263.460 43.870 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1281.170 43.760 1281.490 43.820 ;
        RECT 2279.830 43.760 2280.150 43.820 ;
        RECT 1281.170 43.620 2280.150 43.760 ;
        RECT 1281.170 43.560 1281.490 43.620 ;
        RECT 2279.830 43.560 2280.150 43.620 ;
      LAYER via ;
        RECT 1281.200 43.560 1281.460 43.820 ;
        RECT 2279.860 43.560 2280.120 43.820 ;
      LAYER met2 ;
        RECT 2279.920 43.850 2280.060 54.000 ;
        RECT 1281.200 43.530 1281.460 43.850 ;
        RECT 2279.860 43.530 2280.120 43.850 ;
        RECT 1281.260 2.400 1281.400 43.530 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.110 43.420 1299.430 43.480 ;
        RECT 2285.350 43.420 2285.670 43.480 ;
        RECT 1299.110 43.280 2285.670 43.420 ;
        RECT 1299.110 43.220 1299.430 43.280 ;
        RECT 2285.350 43.220 2285.670 43.280 ;
      LAYER via ;
        RECT 1299.140 43.220 1299.400 43.480 ;
        RECT 2285.380 43.220 2285.640 43.480 ;
      LAYER met2 ;
        RECT 2285.440 43.510 2285.580 54.000 ;
        RECT 1299.140 43.190 1299.400 43.510 ;
        RECT 2285.380 43.190 2285.640 43.510 ;
        RECT 1299.200 2.400 1299.340 43.190 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 43.080 1317.370 43.140 ;
        RECT 2291.330 43.080 2291.650 43.140 ;
        RECT 1317.050 42.940 2291.650 43.080 ;
        RECT 1317.050 42.880 1317.370 42.940 ;
        RECT 2291.330 42.880 2291.650 42.940 ;
      LAYER via ;
        RECT 1317.080 42.880 1317.340 43.140 ;
        RECT 2291.360 42.880 2291.620 43.140 ;
      LAYER met2 ;
        RECT 2291.420 43.170 2291.560 54.000 ;
        RECT 1317.080 42.850 1317.340 43.170 ;
        RECT 2291.360 42.850 2291.620 43.170 ;
        RECT 1317.140 2.400 1317.280 42.850 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.990 42.740 1335.310 42.800 ;
        RECT 2296.850 42.740 2297.170 42.800 ;
        RECT 1334.990 42.600 2297.170 42.740 ;
        RECT 1334.990 42.540 1335.310 42.600 ;
        RECT 2296.850 42.540 2297.170 42.600 ;
      LAYER via ;
        RECT 1335.020 42.540 1335.280 42.800 ;
        RECT 2296.880 42.540 2297.140 42.800 ;
      LAYER met2 ;
        RECT 2296.940 42.830 2297.080 54.000 ;
        RECT 1335.020 42.510 1335.280 42.830 ;
        RECT 2296.880 42.510 2297.140 42.830 ;
        RECT 1335.080 2.400 1335.220 42.510 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2088.560 45.405 2088.700 54.000 ;
        RECT 692.390 45.035 692.670 45.405 ;
        RECT 2088.490 45.035 2088.770 45.405 ;
        RECT 692.460 2.400 692.600 45.035 ;
        RECT 692.250 -4.800 692.810 2.400 ;
      LAYER via2 ;
        RECT 692.390 45.080 692.670 45.360 ;
        RECT 2088.490 45.080 2088.770 45.360 ;
      LAYER met3 ;
        RECT 692.365 45.370 692.695 45.385 ;
        RECT 2088.465 45.370 2088.795 45.385 ;
        RECT 692.365 45.070 2088.795 45.370 ;
        RECT 692.365 45.055 692.695 45.070 ;
        RECT 2088.465 45.055 2088.795 45.070 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 42.400 1352.790 42.460 ;
        RECT 2302.830 42.400 2303.150 42.460 ;
        RECT 1352.470 42.260 2303.150 42.400 ;
        RECT 1352.470 42.200 1352.790 42.260 ;
        RECT 2302.830 42.200 2303.150 42.260 ;
      LAYER via ;
        RECT 1352.500 42.200 1352.760 42.460 ;
        RECT 2302.860 42.200 2303.120 42.460 ;
      LAYER met2 ;
        RECT 2302.920 42.490 2303.060 54.000 ;
        RECT 1352.500 42.170 1352.760 42.490 ;
        RECT 2302.860 42.170 2303.120 42.490 ;
        RECT 1352.560 2.400 1352.700 42.170 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 13.840 1370.730 13.900 ;
        RECT 2305.130 13.840 2305.450 13.900 ;
        RECT 1370.410 13.700 2305.450 13.840 ;
        RECT 1370.410 13.640 1370.730 13.700 ;
        RECT 2305.130 13.640 2305.450 13.700 ;
      LAYER via ;
        RECT 1370.440 13.640 1370.700 13.900 ;
        RECT 2305.160 13.640 2305.420 13.900 ;
      LAYER met2 ;
        RECT 2305.220 13.930 2305.360 54.000 ;
        RECT 1370.440 13.610 1370.700 13.930 ;
        RECT 2305.160 13.610 2305.420 13.930 ;
        RECT 1370.500 2.400 1370.640 13.610 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1388.350 16.900 1388.670 16.960 ;
        RECT 1393.410 16.900 1393.730 16.960 ;
        RECT 1388.350 16.760 1393.730 16.900 ;
        RECT 1388.350 16.700 1388.670 16.760 ;
        RECT 1393.410 16.700 1393.730 16.760 ;
      LAYER via ;
        RECT 1388.380 16.700 1388.640 16.960 ;
        RECT 1393.440 16.700 1393.700 16.960 ;
      LAYER met2 ;
        RECT 1393.500 16.990 1393.640 54.000 ;
        RECT 1388.380 16.670 1388.640 16.990 ;
        RECT 1393.440 16.670 1393.700 16.990 ;
        RECT 1388.440 2.400 1388.580 16.670 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1640.505 9.605 1642.055 9.775 ;
      LAYER mcon ;
        RECT 1641.885 9.605 1642.055 9.775 ;
      LAYER met1 ;
        RECT 1406.290 9.760 1406.610 9.820 ;
        RECT 1640.445 9.760 1640.735 9.805 ;
        RECT 1406.290 9.620 1640.735 9.760 ;
        RECT 1406.290 9.560 1406.610 9.620 ;
        RECT 1640.445 9.575 1640.735 9.620 ;
        RECT 1641.825 9.760 1642.115 9.805 ;
        RECT 2319.390 9.760 2319.710 9.820 ;
        RECT 1641.825 9.620 2319.710 9.760 ;
        RECT 1641.825 9.575 1642.115 9.620 ;
        RECT 2319.390 9.560 2319.710 9.620 ;
      LAYER via ;
        RECT 1406.320 9.560 1406.580 9.820 ;
        RECT 2319.420 9.560 2319.680 9.820 ;
      LAYER met2 ;
        RECT 2319.480 9.850 2319.620 54.000 ;
        RECT 1406.320 9.530 1406.580 9.850 ;
        RECT 2319.420 9.530 2319.680 9.850 ;
        RECT 1406.380 2.400 1406.520 9.530 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1423.770 16.900 1424.090 16.960 ;
        RECT 1427.910 16.900 1428.230 16.960 ;
        RECT 1423.770 16.760 1428.230 16.900 ;
        RECT 1423.770 16.700 1424.090 16.760 ;
        RECT 1427.910 16.700 1428.230 16.760 ;
      LAYER via ;
        RECT 1423.800 16.700 1424.060 16.960 ;
        RECT 1427.940 16.700 1428.200 16.960 ;
      LAYER met2 ;
        RECT 1428.000 16.990 1428.140 54.000 ;
        RECT 1423.800 16.670 1424.060 16.990 ;
        RECT 1427.940 16.670 1428.200 16.990 ;
        RECT 1423.860 2.400 1424.000 16.670 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1640.045 9.265 1641.135 9.435 ;
        RECT 1737.105 9.265 1738.655 9.435 ;
        RECT 1930.765 9.265 1931.395 9.435 ;
      LAYER mcon ;
        RECT 1640.965 9.265 1641.135 9.435 ;
        RECT 1738.485 9.265 1738.655 9.435 ;
        RECT 1931.225 9.265 1931.395 9.435 ;
      LAYER met1 ;
        RECT 1441.710 9.420 1442.030 9.480 ;
        RECT 1639.985 9.420 1640.275 9.465 ;
        RECT 1441.710 9.280 1640.275 9.420 ;
        RECT 1441.710 9.220 1442.030 9.280 ;
        RECT 1639.985 9.235 1640.275 9.280 ;
        RECT 1640.905 9.420 1641.195 9.465 ;
        RECT 1737.045 9.420 1737.335 9.465 ;
        RECT 1640.905 9.280 1737.335 9.420 ;
        RECT 1640.905 9.235 1641.195 9.280 ;
        RECT 1737.045 9.235 1737.335 9.280 ;
        RECT 1738.425 9.420 1738.715 9.465 ;
        RECT 1930.705 9.420 1930.995 9.465 ;
        RECT 1738.425 9.280 1930.995 9.420 ;
        RECT 1738.425 9.235 1738.715 9.280 ;
        RECT 1930.705 9.235 1930.995 9.280 ;
        RECT 1931.165 9.420 1931.455 9.465 ;
        RECT 2326.750 9.420 2327.070 9.480 ;
        RECT 1931.165 9.280 2327.070 9.420 ;
        RECT 1931.165 9.235 1931.455 9.280 ;
        RECT 2326.750 9.220 2327.070 9.280 ;
      LAYER via ;
        RECT 1441.740 9.220 1442.000 9.480 ;
        RECT 2326.780 9.220 2327.040 9.480 ;
      LAYER met2 ;
        RECT 2326.840 9.510 2326.980 54.000 ;
        RECT 1441.740 9.190 1442.000 9.510 ;
        RECT 2326.780 9.190 2327.040 9.510 ;
        RECT 1441.800 2.400 1441.940 9.190 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1459.650 22.340 1459.970 22.400 ;
        RECT 2333.650 22.340 2333.970 22.400 ;
        RECT 1459.650 22.200 2333.970 22.340 ;
        RECT 1459.650 22.140 1459.970 22.200 ;
        RECT 2333.650 22.140 2333.970 22.200 ;
      LAYER via ;
        RECT 1459.680 22.140 1459.940 22.400 ;
        RECT 2333.680 22.140 2333.940 22.400 ;
      LAYER met2 ;
        RECT 2333.740 22.430 2333.880 54.000 ;
        RECT 1459.680 22.110 1459.940 22.430 ;
        RECT 2333.680 22.110 2333.940 22.430 ;
        RECT 1459.740 2.400 1459.880 22.110 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1477.590 17.920 1477.910 17.980 ;
        RECT 1483.110 17.920 1483.430 17.980 ;
        RECT 1477.590 17.780 1483.430 17.920 ;
        RECT 1477.590 17.720 1477.910 17.780 ;
        RECT 1483.110 17.720 1483.430 17.780 ;
      LAYER via ;
        RECT 1477.620 17.720 1477.880 17.980 ;
        RECT 1483.140 17.720 1483.400 17.980 ;
      LAYER met2 ;
        RECT 1483.200 18.010 1483.340 54.000 ;
        RECT 1477.620 17.690 1477.880 18.010 ;
        RECT 1483.140 17.690 1483.400 18.010 ;
        RECT 1477.680 2.400 1477.820 17.690 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1495.530 9.080 1495.850 9.140 ;
        RECT 1929.770 9.080 1930.090 9.140 ;
        RECT 1495.530 8.940 1930.090 9.080 ;
        RECT 1495.530 8.880 1495.850 8.940 ;
        RECT 1929.770 8.880 1930.090 8.940 ;
        RECT 1931.610 9.080 1931.930 9.140 ;
        RECT 2347.450 9.080 2347.770 9.140 ;
        RECT 1931.610 8.940 2347.770 9.080 ;
        RECT 1931.610 8.880 1931.930 8.940 ;
        RECT 2347.450 8.880 2347.770 8.940 ;
      LAYER via ;
        RECT 1495.560 8.880 1495.820 9.140 ;
        RECT 1929.800 8.880 1930.060 9.140 ;
        RECT 1931.640 8.880 1931.900 9.140 ;
        RECT 2347.480 8.880 2347.740 9.140 ;
      LAYER met2 ;
        RECT 2347.540 9.170 2347.680 54.000 ;
        RECT 1495.560 8.850 1495.820 9.170 ;
        RECT 1929.800 8.850 1930.060 9.170 ;
        RECT 1931.640 8.850 1931.900 9.170 ;
        RECT 2347.480 8.850 2347.740 9.170 ;
        RECT 1495.620 2.400 1495.760 8.850 ;
        RECT 1929.860 8.570 1930.000 8.850 ;
        RECT 1931.700 8.570 1931.840 8.850 ;
        RECT 1929.860 8.430 1931.840 8.570 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1517.610 51.920 1517.930 51.980 ;
        RECT 2354.350 51.920 2354.670 51.980 ;
        RECT 1517.610 51.780 2354.670 51.920 ;
        RECT 1517.610 51.720 1517.930 51.780 ;
        RECT 2354.350 51.720 2354.670 51.780 ;
        RECT 1513.010 17.920 1513.330 17.980 ;
        RECT 1517.610 17.920 1517.930 17.980 ;
        RECT 1513.010 17.780 1517.930 17.920 ;
        RECT 1513.010 17.720 1513.330 17.780 ;
        RECT 1517.610 17.720 1517.930 17.780 ;
      LAYER via ;
        RECT 1517.640 51.720 1517.900 51.980 ;
        RECT 2354.380 51.720 2354.640 51.980 ;
        RECT 1513.040 17.720 1513.300 17.980 ;
        RECT 1517.640 17.720 1517.900 17.980 ;
      LAYER met2 ;
        RECT 2354.440 52.010 2354.580 54.000 ;
        RECT 1517.640 51.690 1517.900 52.010 ;
        RECT 2354.380 51.690 2354.640 52.010 ;
        RECT 1517.700 18.010 1517.840 51.690 ;
        RECT 1513.040 17.690 1513.300 18.010 ;
        RECT 1517.640 17.690 1517.900 18.010 ;
        RECT 1513.100 2.400 1513.240 17.690 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2095.920 52.205 2096.060 54.000 ;
        RECT 710.330 51.835 710.610 52.205 ;
        RECT 2095.850 51.835 2096.130 52.205 ;
        RECT 710.400 2.400 710.540 51.835 ;
        RECT 710.190 -4.800 710.750 2.400 ;
      LAYER via2 ;
        RECT 710.330 51.880 710.610 52.160 ;
        RECT 2095.850 51.880 2096.130 52.160 ;
      LAYER met3 ;
        RECT 710.305 52.170 710.635 52.185 ;
        RECT 2095.825 52.170 2096.155 52.185 ;
        RECT 710.305 51.870 2096.155 52.170 ;
        RECT 710.305 51.855 710.635 51.870 ;
        RECT 2095.825 51.855 2096.155 51.870 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1531.410 52.600 1531.730 52.660 ;
        RECT 2360.330 52.600 2360.650 52.660 ;
        RECT 1531.410 52.460 2360.650 52.600 ;
        RECT 1531.410 52.400 1531.730 52.460 ;
        RECT 2360.330 52.400 2360.650 52.460 ;
      LAYER via ;
        RECT 1531.440 52.400 1531.700 52.660 ;
        RECT 2360.360 52.400 2360.620 52.660 ;
      LAYER met2 ;
        RECT 2360.420 52.690 2360.560 54.000 ;
        RECT 1531.440 52.370 1531.700 52.690 ;
        RECT 2360.360 52.370 2360.620 52.690 ;
        RECT 1531.500 17.410 1531.640 52.370 ;
        RECT 1531.040 17.270 1531.640 17.410 ;
        RECT 1531.040 2.400 1531.180 17.270 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.110 52.940 1552.430 53.000 ;
        RECT 2365.850 52.940 2366.170 53.000 ;
        RECT 1552.110 52.800 2366.170 52.940 ;
        RECT 1552.110 52.740 1552.430 52.800 ;
        RECT 2365.850 52.740 2366.170 52.800 ;
        RECT 1548.890 16.900 1549.210 16.960 ;
        RECT 1552.110 16.900 1552.430 16.960 ;
        RECT 1548.890 16.760 1552.430 16.900 ;
        RECT 1548.890 16.700 1549.210 16.760 ;
        RECT 1552.110 16.700 1552.430 16.760 ;
      LAYER via ;
        RECT 1552.140 52.740 1552.400 53.000 ;
        RECT 2365.880 52.740 2366.140 53.000 ;
        RECT 1548.920 16.700 1549.180 16.960 ;
        RECT 1552.140 16.700 1552.400 16.960 ;
      LAYER met2 ;
        RECT 2365.940 53.030 2366.080 54.000 ;
        RECT 1552.140 52.710 1552.400 53.030 ;
        RECT 2365.880 52.710 2366.140 53.030 ;
        RECT 1552.200 16.990 1552.340 52.710 ;
        RECT 1548.920 16.670 1549.180 16.990 ;
        RECT 1552.140 16.670 1552.400 16.990 ;
        RECT 1548.980 2.400 1549.120 16.670 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1572.810 52.260 1573.130 52.320 ;
        RECT 2371.830 52.260 2372.150 52.320 ;
        RECT 1572.810 52.120 2372.150 52.260 ;
        RECT 1572.810 52.060 1573.130 52.120 ;
        RECT 2371.830 52.060 2372.150 52.120 ;
        RECT 1566.830 16.900 1567.150 16.960 ;
        RECT 1572.810 16.900 1573.130 16.960 ;
        RECT 1566.830 16.760 1573.130 16.900 ;
        RECT 1566.830 16.700 1567.150 16.760 ;
        RECT 1572.810 16.700 1573.130 16.760 ;
      LAYER via ;
        RECT 1572.840 52.060 1573.100 52.320 ;
        RECT 2371.860 52.060 2372.120 52.320 ;
        RECT 1566.860 16.700 1567.120 16.960 ;
        RECT 1572.840 16.700 1573.100 16.960 ;
      LAYER met2 ;
        RECT 2371.920 52.350 2372.060 54.000 ;
        RECT 1572.840 52.030 1573.100 52.350 ;
        RECT 2371.860 52.030 2372.120 52.350 ;
        RECT 1572.900 16.990 1573.040 52.030 ;
        RECT 1566.860 16.670 1567.120 16.990 ;
        RECT 1572.840 16.670 1573.100 16.990 ;
        RECT 1566.920 2.400 1567.060 16.670 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.610 53.280 1586.930 53.340 ;
        RECT 2377.350 53.280 2377.670 53.340 ;
        RECT 1586.610 53.140 2377.670 53.280 ;
        RECT 1586.610 53.080 1586.930 53.140 ;
        RECT 2377.350 53.080 2377.670 53.140 ;
      LAYER via ;
        RECT 1586.640 53.080 1586.900 53.340 ;
        RECT 2377.380 53.080 2377.640 53.340 ;
      LAYER met2 ;
        RECT 2377.440 53.370 2377.580 54.000 ;
        RECT 1586.640 53.050 1586.900 53.370 ;
        RECT 2377.380 53.050 2377.640 53.370 ;
        RECT 1586.700 17.410 1586.840 53.050 ;
        RECT 1584.860 17.270 1586.840 17.410 ;
        RECT 1584.860 2.400 1585.000 17.270 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 53.620 1607.630 53.680 ;
        RECT 2383.330 53.620 2383.650 53.680 ;
        RECT 1607.310 53.480 2383.650 53.620 ;
        RECT 1607.310 53.420 1607.630 53.480 ;
        RECT 2383.330 53.420 2383.650 53.480 ;
        RECT 1602.250 16.900 1602.570 16.960 ;
        RECT 1607.310 16.900 1607.630 16.960 ;
        RECT 1602.250 16.760 1607.630 16.900 ;
        RECT 1602.250 16.700 1602.570 16.760 ;
        RECT 1607.310 16.700 1607.630 16.760 ;
      LAYER via ;
        RECT 1607.340 53.420 1607.600 53.680 ;
        RECT 2383.360 53.420 2383.620 53.680 ;
        RECT 1602.280 16.700 1602.540 16.960 ;
        RECT 1607.340 16.700 1607.600 16.960 ;
      LAYER met2 ;
        RECT 2383.420 53.710 2383.560 54.000 ;
        RECT 1607.340 53.390 1607.600 53.710 ;
        RECT 2383.360 53.390 2383.620 53.710 ;
        RECT 1607.400 16.990 1607.540 53.390 ;
        RECT 1602.280 16.670 1602.540 16.990 ;
        RECT 1607.340 16.670 1607.600 16.990 ;
        RECT 1602.340 2.400 1602.480 16.670 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1621.110 53.960 1621.430 54.000 ;
        RECT 2388.850 53.960 2389.170 54.000 ;
        RECT 1621.110 53.820 2389.170 53.960 ;
        RECT 1621.110 53.760 1621.430 53.820 ;
        RECT 2388.850 53.760 2389.170 53.820 ;
      LAYER via ;
        RECT 1621.140 53.760 1621.400 54.000 ;
        RECT 2388.880 53.760 2389.140 54.000 ;
      LAYER met2 ;
        RECT 1621.140 53.730 1621.400 54.000 ;
        RECT 2388.880 53.730 2389.140 54.000 ;
        RECT 1621.200 17.410 1621.340 53.730 ;
        RECT 1620.280 17.270 1621.340 17.410 ;
        RECT 1620.280 2.400 1620.420 17.270 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1638.130 15.880 1638.450 15.940 ;
        RECT 1641.810 15.880 1642.130 15.940 ;
        RECT 1638.130 15.740 1642.130 15.880 ;
        RECT 1638.130 15.680 1638.450 15.740 ;
        RECT 1641.810 15.680 1642.130 15.740 ;
      LAYER via ;
        RECT 1638.160 15.680 1638.420 15.940 ;
        RECT 1641.840 15.680 1642.100 15.940 ;
      LAYER met2 ;
        RECT 1641.900 15.970 1642.040 54.000 ;
        RECT 1638.160 15.650 1638.420 15.970 ;
        RECT 1641.840 15.650 1642.100 15.970 ;
        RECT 1638.220 2.400 1638.360 15.650 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.050 51.580 1662.370 51.640 ;
        RECT 2400.350 51.580 2400.670 51.640 ;
        RECT 1662.050 51.440 2400.670 51.580 ;
        RECT 1662.050 51.380 1662.370 51.440 ;
        RECT 2400.350 51.380 2400.670 51.440 ;
        RECT 1656.070 19.280 1656.390 19.340 ;
        RECT 1662.050 19.280 1662.370 19.340 ;
        RECT 1656.070 19.140 1662.370 19.280 ;
        RECT 1656.070 19.080 1656.390 19.140 ;
        RECT 1662.050 19.080 1662.370 19.140 ;
      LAYER via ;
        RECT 1662.080 51.380 1662.340 51.640 ;
        RECT 2400.380 51.380 2400.640 51.640 ;
        RECT 1656.100 19.080 1656.360 19.340 ;
        RECT 1662.080 19.080 1662.340 19.340 ;
      LAYER met2 ;
        RECT 2400.440 51.670 2400.580 54.000 ;
        RECT 1662.080 51.350 1662.340 51.670 ;
        RECT 2400.380 51.350 2400.640 51.670 ;
        RECT 1662.140 19.370 1662.280 51.350 ;
        RECT 1656.100 19.050 1656.360 19.370 ;
        RECT 1662.080 19.050 1662.340 19.370 ;
        RECT 1656.160 2.400 1656.300 19.050 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1673.550 16.900 1673.870 16.960 ;
        RECT 1676.310 16.900 1676.630 16.960 ;
        RECT 1673.550 16.760 1676.630 16.900 ;
        RECT 1673.550 16.700 1673.870 16.760 ;
        RECT 1676.310 16.700 1676.630 16.760 ;
      LAYER via ;
        RECT 1673.580 16.700 1673.840 16.960 ;
        RECT 1676.340 16.700 1676.600 16.960 ;
      LAYER met2 ;
        RECT 1676.400 16.990 1676.540 54.000 ;
        RECT 1673.580 16.670 1673.840 16.990 ;
        RECT 1676.340 16.670 1676.600 16.990 ;
        RECT 1673.640 2.400 1673.780 16.670 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1691.490 16.900 1691.810 16.960 ;
        RECT 1697.010 16.900 1697.330 16.960 ;
        RECT 1691.490 16.760 1697.330 16.900 ;
        RECT 1691.490 16.700 1691.810 16.760 ;
        RECT 1697.010 16.700 1697.330 16.760 ;
      LAYER via ;
        RECT 1691.520 16.700 1691.780 16.960 ;
        RECT 1697.040 16.700 1697.300 16.960 ;
      LAYER met2 ;
        RECT 1697.100 16.990 1697.240 54.000 ;
        RECT 1691.520 16.670 1691.780 16.990 ;
        RECT 1697.040 16.670 1697.300 16.990 ;
        RECT 1691.580 2.400 1691.720 16.670 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.440 52.885 2101.580 54.000 ;
        RECT 728.270 52.515 728.550 52.885 ;
        RECT 2101.370 52.515 2101.650 52.885 ;
        RECT 728.340 2.400 728.480 52.515 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 728.270 52.560 728.550 52.840 ;
        RECT 2101.370 52.560 2101.650 52.840 ;
      LAYER met3 ;
        RECT 728.245 52.850 728.575 52.865 ;
        RECT 2101.345 52.850 2101.675 52.865 ;
        RECT 728.245 52.550 2101.675 52.850 ;
        RECT 728.245 52.535 728.575 52.550 ;
        RECT 2101.345 52.535 2101.675 52.550 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1710.810 51.240 1711.130 51.300 ;
        RECT 2417.830 51.240 2418.150 51.300 ;
        RECT 1710.810 51.100 2418.150 51.240 ;
        RECT 1710.810 51.040 1711.130 51.100 ;
        RECT 2417.830 51.040 2418.150 51.100 ;
      LAYER via ;
        RECT 1710.840 51.040 1711.100 51.300 ;
        RECT 2417.860 51.040 2418.120 51.300 ;
      LAYER met2 ;
        RECT 2417.920 51.330 2418.060 54.000 ;
        RECT 1710.840 51.010 1711.100 51.330 ;
        RECT 2417.860 51.010 2418.120 51.330 ;
        RECT 1710.900 17.410 1711.040 51.010 ;
        RECT 1709.520 17.270 1711.040 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.510 50.900 1731.830 50.960 ;
        RECT 2423.350 50.900 2423.670 50.960 ;
        RECT 1731.510 50.760 2423.670 50.900 ;
        RECT 1731.510 50.700 1731.830 50.760 ;
        RECT 2423.350 50.700 2423.670 50.760 ;
        RECT 1727.370 16.900 1727.690 16.960 ;
        RECT 1731.510 16.900 1731.830 16.960 ;
        RECT 1727.370 16.760 1731.830 16.900 ;
        RECT 1727.370 16.700 1727.690 16.760 ;
        RECT 1731.510 16.700 1731.830 16.760 ;
      LAYER via ;
        RECT 1731.540 50.700 1731.800 50.960 ;
        RECT 2423.380 50.700 2423.640 50.960 ;
        RECT 1727.400 16.700 1727.660 16.960 ;
        RECT 1731.540 16.700 1731.800 16.960 ;
      LAYER met2 ;
        RECT 2423.440 50.990 2423.580 54.000 ;
        RECT 1731.540 50.670 1731.800 50.990 ;
        RECT 2423.380 50.670 2423.640 50.990 ;
        RECT 1731.600 16.990 1731.740 50.670 ;
        RECT 1727.400 16.670 1727.660 16.990 ;
        RECT 1731.540 16.670 1731.800 16.990 ;
        RECT 1727.460 2.400 1727.600 16.670 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1744.850 50.560 1745.170 50.620 ;
        RECT 2429.330 50.560 2429.650 50.620 ;
        RECT 1744.850 50.420 2429.650 50.560 ;
        RECT 1744.850 50.360 1745.170 50.420 ;
        RECT 2429.330 50.360 2429.650 50.420 ;
      LAYER via ;
        RECT 1744.880 50.360 1745.140 50.620 ;
        RECT 2429.360 50.360 2429.620 50.620 ;
      LAYER met2 ;
        RECT 2429.420 50.650 2429.560 54.000 ;
        RECT 1744.880 50.330 1745.140 50.650 ;
        RECT 2429.360 50.330 2429.620 50.650 ;
        RECT 1744.940 7.890 1745.080 50.330 ;
        RECT 1744.940 7.750 1745.540 7.890 ;
        RECT 1745.400 2.400 1745.540 7.750 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.010 50.220 1766.330 50.280 ;
        RECT 2433.470 50.220 2433.790 50.280 ;
        RECT 1766.010 50.080 2433.790 50.220 ;
        RECT 1766.010 50.020 1766.330 50.080 ;
        RECT 2433.470 50.020 2433.790 50.080 ;
        RECT 1762.790 16.900 1763.110 16.960 ;
        RECT 1766.010 16.900 1766.330 16.960 ;
        RECT 1762.790 16.760 1766.330 16.900 ;
        RECT 1762.790 16.700 1763.110 16.760 ;
        RECT 1766.010 16.700 1766.330 16.760 ;
      LAYER via ;
        RECT 1766.040 50.020 1766.300 50.280 ;
        RECT 2433.500 50.020 2433.760 50.280 ;
        RECT 1762.820 16.700 1763.080 16.960 ;
        RECT 1766.040 16.700 1766.300 16.960 ;
      LAYER met2 ;
        RECT 2433.560 50.310 2433.700 54.000 ;
        RECT 1766.040 49.990 1766.300 50.310 ;
        RECT 2433.500 49.990 2433.760 50.310 ;
        RECT 1766.100 16.990 1766.240 49.990 ;
        RECT 1762.820 16.670 1763.080 16.990 ;
        RECT 1766.040 16.670 1766.300 16.990 ;
        RECT 1762.880 2.400 1763.020 16.670 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1786.710 49.880 1787.030 49.940 ;
        RECT 2440.830 49.880 2441.150 49.940 ;
        RECT 1786.710 49.740 2441.150 49.880 ;
        RECT 1786.710 49.680 1787.030 49.740 ;
        RECT 2440.830 49.680 2441.150 49.740 ;
        RECT 1780.730 16.900 1781.050 16.960 ;
        RECT 1786.710 16.900 1787.030 16.960 ;
        RECT 1780.730 16.760 1787.030 16.900 ;
        RECT 1780.730 16.700 1781.050 16.760 ;
        RECT 1786.710 16.700 1787.030 16.760 ;
      LAYER via ;
        RECT 1786.740 49.680 1787.000 49.940 ;
        RECT 2440.860 49.680 2441.120 49.940 ;
        RECT 1780.760 16.700 1781.020 16.960 ;
        RECT 1786.740 16.700 1787.000 16.960 ;
      LAYER met2 ;
        RECT 2440.920 49.970 2441.060 54.000 ;
        RECT 1786.740 49.650 1787.000 49.970 ;
        RECT 2440.860 49.650 2441.120 49.970 ;
        RECT 1786.800 16.990 1786.940 49.650 ;
        RECT 1780.760 16.670 1781.020 16.990 ;
        RECT 1786.740 16.670 1787.000 16.990 ;
        RECT 1780.820 2.400 1780.960 16.670 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.510 49.540 1800.830 49.600 ;
        RECT 2446.350 49.540 2446.670 49.600 ;
        RECT 1800.510 49.400 2446.670 49.540 ;
        RECT 1800.510 49.340 1800.830 49.400 ;
        RECT 2446.350 49.340 2446.670 49.400 ;
      LAYER via ;
        RECT 1800.540 49.340 1800.800 49.600 ;
        RECT 2446.380 49.340 2446.640 49.600 ;
      LAYER met2 ;
        RECT 2446.440 49.630 2446.580 54.000 ;
        RECT 1800.540 49.310 1800.800 49.630 ;
        RECT 2446.380 49.310 2446.640 49.630 ;
        RECT 1800.600 17.410 1800.740 49.310 ;
        RECT 1798.760 17.270 1800.740 17.410 ;
        RECT 1798.760 2.400 1798.900 17.270 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1816.610 49.200 1816.930 49.260 ;
        RECT 2452.330 49.200 2452.650 49.260 ;
        RECT 1816.610 49.060 2452.650 49.200 ;
        RECT 1816.610 49.000 1816.930 49.060 ;
        RECT 2452.330 49.000 2452.650 49.060 ;
      LAYER via ;
        RECT 1816.640 49.000 1816.900 49.260 ;
        RECT 2452.360 49.000 2452.620 49.260 ;
      LAYER met2 ;
        RECT 2452.420 49.290 2452.560 54.000 ;
        RECT 1816.640 48.970 1816.900 49.290 ;
        RECT 2452.360 48.970 2452.620 49.290 ;
        RECT 1816.700 2.400 1816.840 48.970 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.010 48.860 1835.330 48.920 ;
        RECT 2457.850 48.860 2458.170 48.920 ;
        RECT 1835.010 48.720 2458.170 48.860 ;
        RECT 1835.010 48.660 1835.330 48.720 ;
        RECT 2457.850 48.660 2458.170 48.720 ;
      LAYER via ;
        RECT 1835.040 48.660 1835.300 48.920 ;
        RECT 2457.880 48.660 2458.140 48.920 ;
      LAYER met2 ;
        RECT 2457.940 48.950 2458.080 54.000 ;
        RECT 1835.040 48.630 1835.300 48.950 ;
        RECT 2457.880 48.630 2458.140 48.950 ;
        RECT 1835.100 3.130 1835.240 48.630 ;
        RECT 1834.640 2.990 1835.240 3.130 ;
        RECT 1834.640 2.400 1834.780 2.990 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1852.030 42.060 1852.350 42.120 ;
        RECT 2463.830 42.060 2464.150 42.120 ;
        RECT 1852.030 41.920 2464.150 42.060 ;
        RECT 1852.030 41.860 1852.350 41.920 ;
        RECT 2463.830 41.860 2464.150 41.920 ;
      LAYER via ;
        RECT 1852.060 41.860 1852.320 42.120 ;
        RECT 2463.860 41.860 2464.120 42.120 ;
      LAYER met2 ;
        RECT 2463.920 42.150 2464.060 54.000 ;
        RECT 1852.060 41.830 1852.320 42.150 ;
        RECT 2463.860 41.830 2464.120 42.150 ;
        RECT 1852.120 2.400 1852.260 41.830 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1869.970 21.660 1870.290 21.720 ;
        RECT 2464.290 21.660 2464.610 21.720 ;
        RECT 1869.970 21.520 2464.610 21.660 ;
        RECT 1869.970 21.460 1870.290 21.520 ;
        RECT 2464.290 21.460 2464.610 21.520 ;
      LAYER via ;
        RECT 1870.000 21.460 1870.260 21.720 ;
        RECT 2464.320 21.460 2464.580 21.720 ;
      LAYER met2 ;
        RECT 2464.380 21.750 2464.520 54.000 ;
        RECT 1870.000 21.430 1870.260 21.750 ;
        RECT 2464.320 21.430 2464.580 21.750 ;
        RECT 1870.060 2.400 1870.200 21.430 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 746.190 31.180 746.510 31.240 ;
        RECT 2105.950 31.180 2106.270 31.240 ;
        RECT 746.190 31.040 2106.270 31.180 ;
        RECT 746.190 30.980 746.510 31.040 ;
        RECT 2105.950 30.980 2106.270 31.040 ;
      LAYER via ;
        RECT 746.220 30.980 746.480 31.240 ;
        RECT 2105.980 30.980 2106.240 31.240 ;
      LAYER met2 ;
        RECT 2106.040 31.270 2106.180 54.000 ;
        RECT 746.220 30.950 746.480 31.270 ;
        RECT 2105.980 30.950 2106.240 31.270 ;
        RECT 746.280 2.400 746.420 30.950 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1887.910 16.560 1888.230 16.620 ;
        RECT 1890.210 16.560 1890.530 16.620 ;
        RECT 1887.910 16.420 1890.530 16.560 ;
        RECT 1887.910 16.360 1888.230 16.420 ;
        RECT 1890.210 16.360 1890.530 16.420 ;
      LAYER via ;
        RECT 1887.940 16.360 1888.200 16.620 ;
        RECT 1890.240 16.360 1890.500 16.620 ;
      LAYER met2 ;
        RECT 1890.300 16.650 1890.440 54.000 ;
        RECT 1887.940 16.330 1888.200 16.650 ;
        RECT 1890.240 16.330 1890.500 16.650 ;
        RECT 1888.000 2.400 1888.140 16.330 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1905.850 16.560 1906.170 16.620 ;
        RECT 1910.910 16.560 1911.230 16.620 ;
        RECT 1905.850 16.420 1911.230 16.560 ;
        RECT 1905.850 16.360 1906.170 16.420 ;
        RECT 1910.910 16.360 1911.230 16.420 ;
      LAYER via ;
        RECT 1905.880 16.360 1906.140 16.620 ;
        RECT 1910.940 16.360 1911.200 16.620 ;
      LAYER met2 ;
        RECT 1911.000 16.650 1911.140 54.000 ;
        RECT 1905.880 16.330 1906.140 16.650 ;
        RECT 1910.940 16.330 1911.200 16.650 ;
        RECT 1905.940 2.400 1906.080 16.330 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1924.800 17.410 1924.940 54.000 ;
        RECT 1923.420 17.270 1924.940 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1941.270 16.220 1941.590 16.280 ;
        RECT 1945.410 16.220 1945.730 16.280 ;
        RECT 1941.270 16.080 1945.730 16.220 ;
        RECT 1941.270 16.020 1941.590 16.080 ;
        RECT 1945.410 16.020 1945.730 16.080 ;
      LAYER via ;
        RECT 1941.300 16.020 1941.560 16.280 ;
        RECT 1945.440 16.020 1945.700 16.280 ;
      LAYER met2 ;
        RECT 1945.500 16.310 1945.640 54.000 ;
        RECT 1941.300 15.990 1941.560 16.310 ;
        RECT 1945.440 15.990 1945.700 16.310 ;
        RECT 1941.360 2.400 1941.500 15.990 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.300 2.400 1959.440 54.000 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1977.150 15.540 1977.470 15.600 ;
        RECT 1979.910 15.540 1980.230 15.600 ;
        RECT 1977.150 15.400 1980.230 15.540 ;
        RECT 1977.150 15.340 1977.470 15.400 ;
        RECT 1979.910 15.340 1980.230 15.400 ;
      LAYER via ;
        RECT 1977.180 15.340 1977.440 15.600 ;
        RECT 1979.940 15.340 1980.200 15.600 ;
      LAYER met2 ;
        RECT 1980.000 15.630 1980.140 54.000 ;
        RECT 1977.180 15.310 1977.440 15.630 ;
        RECT 1979.940 15.310 1980.200 15.630 ;
        RECT 1977.240 2.400 1977.380 15.310 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.090 15.540 1995.410 15.600 ;
        RECT 2000.610 15.540 2000.930 15.600 ;
        RECT 1995.090 15.400 2000.930 15.540 ;
        RECT 1995.090 15.340 1995.410 15.400 ;
        RECT 2000.610 15.340 2000.930 15.400 ;
      LAYER via ;
        RECT 1995.120 15.340 1995.380 15.600 ;
        RECT 2000.640 15.340 2000.900 15.600 ;
      LAYER met2 ;
        RECT 2000.700 15.630 2000.840 54.000 ;
        RECT 1995.120 15.310 1995.380 15.630 ;
        RECT 2000.640 15.310 2000.900 15.630 ;
        RECT 1995.180 2.400 1995.320 15.310 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2012.570 41.720 2012.890 41.780 ;
        RECT 2515.350 41.720 2515.670 41.780 ;
        RECT 2012.570 41.580 2515.670 41.720 ;
        RECT 2012.570 41.520 2012.890 41.580 ;
        RECT 2515.350 41.520 2515.670 41.580 ;
      LAYER via ;
        RECT 2012.600 41.520 2012.860 41.780 ;
        RECT 2515.380 41.520 2515.640 41.780 ;
      LAYER met2 ;
        RECT 2515.440 41.810 2515.580 54.000 ;
        RECT 2012.600 41.490 2012.860 41.810 ;
        RECT 2515.380 41.490 2515.640 41.810 ;
        RECT 2012.660 2.400 2012.800 41.490 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2030.510 17.580 2030.830 17.640 ;
        RECT 2035.110 17.580 2035.430 17.640 ;
        RECT 2030.510 17.440 2035.430 17.580 ;
        RECT 2030.510 17.380 2030.830 17.440 ;
        RECT 2035.110 17.380 2035.430 17.440 ;
      LAYER via ;
        RECT 2030.540 17.380 2030.800 17.640 ;
        RECT 2035.140 17.380 2035.400 17.640 ;
      LAYER met2 ;
        RECT 2035.200 17.670 2035.340 54.000 ;
        RECT 2030.540 17.350 2030.800 17.670 ;
        RECT 2035.140 17.350 2035.400 17.670 ;
        RECT 2030.600 2.400 2030.740 17.350 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.540 2.400 2048.680 54.000 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 814.345 16.065 814.515 16.915 ;
        RECT 855.745 15.385 855.915 16.235 ;
        RECT 903.585 15.385 903.755 17.255 ;
        RECT 910.945 15.725 911.115 17.255 ;
        RECT 965.685 15.725 965.855 17.255 ;
        RECT 1007.545 16.405 1007.715 17.255 ;
      LAYER mcon ;
        RECT 903.585 17.085 903.755 17.255 ;
        RECT 814.345 16.745 814.515 16.915 ;
        RECT 855.745 16.065 855.915 16.235 ;
        RECT 910.945 17.085 911.115 17.255 ;
        RECT 965.685 17.085 965.855 17.255 ;
        RECT 1007.545 17.085 1007.715 17.255 ;
      LAYER met1 ;
        RECT 763.670 17.580 763.990 17.640 ;
        RECT 763.670 17.440 786.900 17.580 ;
        RECT 763.670 17.380 763.990 17.440 ;
        RECT 786.760 16.900 786.900 17.440 ;
        RECT 903.525 17.240 903.815 17.285 ;
        RECT 910.885 17.240 911.175 17.285 ;
        RECT 903.525 17.100 911.175 17.240 ;
        RECT 903.525 17.055 903.815 17.100 ;
        RECT 910.885 17.055 911.175 17.100 ;
        RECT 965.625 17.240 965.915 17.285 ;
        RECT 1007.485 17.240 1007.775 17.285 ;
        RECT 1231.490 17.240 1231.810 17.300 ;
        RECT 965.625 17.100 1007.775 17.240 ;
        RECT 965.625 17.055 965.915 17.100 ;
        RECT 1007.485 17.055 1007.775 17.100 ;
        RECT 1015.380 17.100 1231.810 17.240 ;
        RECT 814.285 16.900 814.575 16.945 ;
        RECT 786.760 16.760 814.575 16.900 ;
        RECT 814.285 16.715 814.575 16.760 ;
        RECT 1007.485 16.560 1007.775 16.605 ;
        RECT 1015.380 16.560 1015.520 17.100 ;
        RECT 1231.490 17.040 1231.810 17.100 ;
        RECT 1007.485 16.420 1015.520 16.560 ;
        RECT 1007.485 16.375 1007.775 16.420 ;
        RECT 814.285 16.220 814.575 16.265 ;
        RECT 855.685 16.220 855.975 16.265 ;
        RECT 814.285 16.080 855.975 16.220 ;
        RECT 814.285 16.035 814.575 16.080 ;
        RECT 855.685 16.035 855.975 16.080 ;
        RECT 910.885 15.880 911.175 15.925 ;
        RECT 965.625 15.880 965.915 15.925 ;
        RECT 910.885 15.740 965.915 15.880 ;
        RECT 910.885 15.695 911.175 15.740 ;
        RECT 965.625 15.695 965.915 15.740 ;
        RECT 855.685 15.540 855.975 15.585 ;
        RECT 903.525 15.540 903.815 15.585 ;
        RECT 855.685 15.400 903.815 15.540 ;
        RECT 855.685 15.355 855.975 15.400 ;
        RECT 903.525 15.355 903.815 15.400 ;
      LAYER via ;
        RECT 763.700 17.380 763.960 17.640 ;
        RECT 1231.520 17.040 1231.780 17.300 ;
      LAYER met2 ;
        RECT 763.700 17.350 763.960 17.670 ;
        RECT 763.760 2.400 763.900 17.350 ;
        RECT 1231.580 17.330 1231.720 54.000 ;
        RECT 1231.520 17.010 1231.780 17.330 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2066.390 17.580 2066.710 17.640 ;
        RECT 2069.610 17.580 2069.930 17.640 ;
        RECT 2066.390 17.440 2069.930 17.580 ;
        RECT 2066.390 17.380 2066.710 17.440 ;
        RECT 2069.610 17.380 2069.930 17.440 ;
      LAYER via ;
        RECT 2066.420 17.380 2066.680 17.640 ;
        RECT 2069.640 17.380 2069.900 17.640 ;
      LAYER met2 ;
        RECT 2069.700 17.670 2069.840 54.000 ;
        RECT 2066.420 17.350 2066.680 17.670 ;
        RECT 2069.640 17.350 2069.900 17.670 ;
        RECT 2066.480 2.400 2066.620 17.350 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2084.330 17.580 2084.650 17.640 ;
        RECT 2089.850 17.580 2090.170 17.640 ;
        RECT 2084.330 17.440 2090.170 17.580 ;
        RECT 2084.330 17.380 2084.650 17.440 ;
        RECT 2089.850 17.380 2090.170 17.440 ;
      LAYER via ;
        RECT 2084.360 17.380 2084.620 17.640 ;
        RECT 2089.880 17.380 2090.140 17.640 ;
      LAYER met2 ;
        RECT 2089.940 17.670 2090.080 54.000 ;
        RECT 2084.360 17.350 2084.620 17.670 ;
        RECT 2089.880 17.350 2090.140 17.670 ;
        RECT 2084.420 2.400 2084.560 17.350 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2101.810 30.840 2102.130 30.900 ;
        RECT 2539.270 30.840 2539.590 30.900 ;
        RECT 2101.810 30.700 2539.590 30.840 ;
        RECT 2101.810 30.640 2102.130 30.700 ;
        RECT 2539.270 30.640 2539.590 30.700 ;
      LAYER via ;
        RECT 2101.840 30.640 2102.100 30.900 ;
        RECT 2539.300 30.640 2539.560 30.900 ;
      LAYER met2 ;
        RECT 2539.360 30.930 2539.500 54.000 ;
        RECT 2101.840 30.610 2102.100 30.930 ;
        RECT 2539.300 30.610 2539.560 30.930 ;
        RECT 2101.900 2.400 2102.040 30.610 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2119.750 31.180 2120.070 31.240 ;
        RECT 2547.550 31.180 2547.870 31.240 ;
        RECT 2119.750 31.040 2547.870 31.180 ;
        RECT 2119.750 30.980 2120.070 31.040 ;
        RECT 2547.550 30.980 2547.870 31.040 ;
      LAYER via ;
        RECT 2119.780 30.980 2120.040 31.240 ;
        RECT 2547.580 30.980 2547.840 31.240 ;
      LAYER met2 ;
        RECT 2547.640 31.270 2547.780 54.000 ;
        RECT 2119.780 30.950 2120.040 31.270 ;
        RECT 2547.580 30.950 2547.840 31.270 ;
        RECT 2119.840 2.400 2119.980 30.950 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2137.690 37.980 2138.010 38.040 ;
        RECT 2555.830 37.980 2556.150 38.040 ;
        RECT 2137.690 37.840 2556.150 37.980 ;
        RECT 2137.690 37.780 2138.010 37.840 ;
        RECT 2555.830 37.780 2556.150 37.840 ;
      LAYER via ;
        RECT 2137.720 37.780 2137.980 38.040 ;
        RECT 2555.860 37.780 2556.120 38.040 ;
      LAYER met2 ;
        RECT 2555.920 38.070 2556.060 54.000 ;
        RECT 2137.720 37.750 2137.980 38.070 ;
        RECT 2555.860 37.750 2556.120 38.070 ;
        RECT 2137.780 2.400 2137.920 37.750 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2155.630 38.320 2155.950 38.380 ;
        RECT 2561.350 38.320 2561.670 38.380 ;
        RECT 2155.630 38.180 2561.670 38.320 ;
        RECT 2155.630 38.120 2155.950 38.180 ;
        RECT 2561.350 38.120 2561.670 38.180 ;
      LAYER via ;
        RECT 2155.660 38.120 2155.920 38.380 ;
        RECT 2561.380 38.120 2561.640 38.380 ;
      LAYER met2 ;
        RECT 2561.440 38.410 2561.580 54.000 ;
        RECT 2155.660 38.090 2155.920 38.410 ;
        RECT 2561.380 38.090 2561.640 38.410 ;
        RECT 2155.720 2.400 2155.860 38.090 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2173.110 38.660 2173.430 38.720 ;
        RECT 2567.330 38.660 2567.650 38.720 ;
        RECT 2173.110 38.520 2567.650 38.660 ;
        RECT 2173.110 38.460 2173.430 38.520 ;
        RECT 2567.330 38.460 2567.650 38.520 ;
      LAYER via ;
        RECT 2173.140 38.460 2173.400 38.720 ;
        RECT 2567.360 38.460 2567.620 38.720 ;
      LAYER met2 ;
        RECT 2567.420 38.750 2567.560 54.000 ;
        RECT 2173.140 38.430 2173.400 38.750 ;
        RECT 2567.360 38.430 2567.620 38.750 ;
        RECT 2173.200 2.400 2173.340 38.430 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2191.050 39.000 2191.370 39.060 ;
        RECT 2572.850 39.000 2573.170 39.060 ;
        RECT 2191.050 38.860 2573.170 39.000 ;
        RECT 2191.050 38.800 2191.370 38.860 ;
        RECT 2572.850 38.800 2573.170 38.860 ;
      LAYER via ;
        RECT 2191.080 38.800 2191.340 39.060 ;
        RECT 2572.880 38.800 2573.140 39.060 ;
      LAYER met2 ;
        RECT 2572.940 39.090 2573.080 54.000 ;
        RECT 2191.080 38.770 2191.340 39.090 ;
        RECT 2572.880 38.770 2573.140 39.090 ;
        RECT 2191.140 2.400 2191.280 38.770 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2209.450 39.340 2209.770 39.400 ;
        RECT 2578.830 39.340 2579.150 39.400 ;
        RECT 2209.450 39.200 2579.150 39.340 ;
        RECT 2209.450 39.140 2209.770 39.200 ;
        RECT 2578.830 39.140 2579.150 39.200 ;
      LAYER via ;
        RECT 2209.480 39.140 2209.740 39.400 ;
        RECT 2578.860 39.140 2579.120 39.400 ;
      LAYER met2 ;
        RECT 2578.920 39.430 2579.060 54.000 ;
        RECT 2209.480 39.110 2209.740 39.430 ;
        RECT 2578.860 39.110 2579.120 39.430 ;
        RECT 2209.540 17.410 2209.680 39.110 ;
        RECT 2209.080 17.270 2209.680 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2226.930 2.960 2227.250 3.020 ;
        RECT 2228.310 2.960 2228.630 3.020 ;
        RECT 2226.930 2.820 2228.630 2.960 ;
        RECT 2226.930 2.760 2227.250 2.820 ;
        RECT 2228.310 2.760 2228.630 2.820 ;
      LAYER via ;
        RECT 2226.960 2.760 2227.220 3.020 ;
        RECT 2228.340 2.760 2228.600 3.020 ;
      LAYER met2 ;
        RECT 2228.400 3.050 2228.540 54.000 ;
        RECT 2226.960 2.730 2227.220 3.050 ;
        RECT 2228.340 2.730 2228.600 3.050 ;
        RECT 2227.020 2.400 2227.160 2.730 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.700 2.400 781.840 54.000 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2244.945 12.325 2245.115 44.795 ;
      LAYER mcon ;
        RECT 2244.945 44.625 2245.115 44.795 ;
      LAYER met1 ;
        RECT 2244.885 44.780 2245.175 44.825 ;
        RECT 2590.330 44.780 2590.650 44.840 ;
        RECT 2244.885 44.640 2590.650 44.780 ;
        RECT 2244.885 44.595 2245.175 44.640 ;
        RECT 2590.330 44.580 2590.650 44.640 ;
        RECT 2244.870 12.480 2245.190 12.540 ;
        RECT 2244.675 12.340 2245.190 12.480 ;
        RECT 2244.870 12.280 2245.190 12.340 ;
      LAYER via ;
        RECT 2590.360 44.580 2590.620 44.840 ;
        RECT 2244.900 12.280 2245.160 12.540 ;
      LAYER met2 ;
        RECT 2590.420 44.870 2590.560 54.000 ;
        RECT 2590.360 44.550 2590.620 44.870 ;
        RECT 2244.900 12.250 2245.160 12.570 ;
        RECT 2244.960 2.400 2245.100 12.250 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2262.350 45.120 2262.670 45.180 ;
        RECT 2594.930 45.120 2595.250 45.180 ;
        RECT 2262.350 44.980 2595.250 45.120 ;
        RECT 2262.350 44.920 2262.670 44.980 ;
        RECT 2594.930 44.920 2595.250 44.980 ;
      LAYER via ;
        RECT 2262.380 44.920 2262.640 45.180 ;
        RECT 2594.960 44.920 2595.220 45.180 ;
      LAYER met2 ;
        RECT 2595.020 45.210 2595.160 54.000 ;
        RECT 2262.380 44.890 2262.640 45.210 ;
        RECT 2594.960 44.890 2595.220 45.210 ;
        RECT 2262.440 2.400 2262.580 44.890 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2280.290 45.460 2280.610 45.520 ;
        RECT 2601.370 45.460 2601.690 45.520 ;
        RECT 2280.290 45.320 2601.690 45.460 ;
        RECT 2280.290 45.260 2280.610 45.320 ;
        RECT 2601.370 45.260 2601.690 45.320 ;
      LAYER via ;
        RECT 2280.320 45.260 2280.580 45.520 ;
        RECT 2601.400 45.260 2601.660 45.520 ;
      LAYER met2 ;
        RECT 2601.460 45.550 2601.600 54.000 ;
        RECT 2280.320 45.230 2280.580 45.550 ;
        RECT 2601.400 45.230 2601.660 45.550 ;
        RECT 2280.380 2.400 2280.520 45.230 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2298.690 45.800 2299.010 45.860 ;
        RECT 2607.350 45.800 2607.670 45.860 ;
        RECT 2298.690 45.660 2607.670 45.800 ;
        RECT 2298.690 45.600 2299.010 45.660 ;
        RECT 2607.350 45.600 2607.670 45.660 ;
      LAYER via ;
        RECT 2298.720 45.600 2298.980 45.860 ;
        RECT 2607.380 45.600 2607.640 45.860 ;
      LAYER met2 ;
        RECT 2607.440 45.890 2607.580 54.000 ;
        RECT 2298.720 45.570 2298.980 45.890 ;
        RECT 2607.380 45.570 2607.640 45.890 ;
        RECT 2298.780 3.130 2298.920 45.570 ;
        RECT 2298.320 2.990 2298.920 3.130 ;
        RECT 2298.320 2.400 2298.460 2.990 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2316.170 46.140 2316.490 46.200 ;
        RECT 2613.330 46.140 2613.650 46.200 ;
        RECT 2316.170 46.000 2613.650 46.140 ;
        RECT 2316.170 45.940 2316.490 46.000 ;
        RECT 2613.330 45.940 2613.650 46.000 ;
      LAYER via ;
        RECT 2316.200 45.940 2316.460 46.200 ;
        RECT 2613.360 45.940 2613.620 46.200 ;
      LAYER met2 ;
        RECT 2613.420 46.230 2613.560 54.000 ;
        RECT 2316.200 45.910 2316.460 46.230 ;
        RECT 2613.360 45.910 2613.620 46.230 ;
        RECT 2316.260 2.400 2316.400 45.910 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2334.110 14.860 2334.430 14.920 ;
        RECT 2338.710 14.860 2339.030 14.920 ;
        RECT 2334.110 14.720 2339.030 14.860 ;
        RECT 2334.110 14.660 2334.430 14.720 ;
        RECT 2338.710 14.660 2339.030 14.720 ;
      LAYER via ;
        RECT 2334.140 14.660 2334.400 14.920 ;
        RECT 2338.740 14.660 2339.000 14.920 ;
      LAYER met2 ;
        RECT 2338.800 14.950 2338.940 54.000 ;
        RECT 2334.140 14.630 2334.400 14.950 ;
        RECT 2338.740 14.630 2339.000 14.950 ;
        RECT 2334.200 2.400 2334.340 14.630 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2351.590 31.520 2351.910 31.580 ;
        RECT 2622.070 31.520 2622.390 31.580 ;
        RECT 2351.590 31.380 2622.390 31.520 ;
        RECT 2351.590 31.320 2351.910 31.380 ;
        RECT 2622.070 31.320 2622.390 31.380 ;
      LAYER via ;
        RECT 2351.620 31.320 2351.880 31.580 ;
        RECT 2622.100 31.320 2622.360 31.580 ;
      LAYER met2 ;
        RECT 2622.160 31.610 2622.300 54.000 ;
        RECT 2351.620 31.290 2351.880 31.610 ;
        RECT 2622.100 31.290 2622.360 31.610 ;
        RECT 2351.680 2.400 2351.820 31.290 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2369.530 31.860 2369.850 31.920 ;
        RECT 2629.430 31.860 2629.750 31.920 ;
        RECT 2369.530 31.720 2629.750 31.860 ;
        RECT 2369.530 31.660 2369.850 31.720 ;
        RECT 2629.430 31.660 2629.750 31.720 ;
      LAYER via ;
        RECT 2369.560 31.660 2369.820 31.920 ;
        RECT 2629.460 31.660 2629.720 31.920 ;
      LAYER met2 ;
        RECT 2629.520 31.950 2629.660 54.000 ;
        RECT 2369.560 31.630 2369.820 31.950 ;
        RECT 2629.460 31.630 2629.720 31.950 ;
        RECT 2369.620 2.400 2369.760 31.630 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2387.470 16.900 2387.790 16.960 ;
        RECT 2393.910 16.900 2394.230 16.960 ;
        RECT 2387.470 16.760 2394.230 16.900 ;
        RECT 2387.470 16.700 2387.790 16.760 ;
        RECT 2393.910 16.700 2394.230 16.760 ;
      LAYER via ;
        RECT 2387.500 16.700 2387.760 16.960 ;
        RECT 2393.940 16.700 2394.200 16.960 ;
      LAYER met2 ;
        RECT 2394.000 16.990 2394.140 54.000 ;
        RECT 2387.500 16.670 2387.760 16.990 ;
        RECT 2393.940 16.670 2394.200 16.990 ;
        RECT 2387.560 2.400 2387.700 16.670 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2407.710 51.580 2408.030 51.640 ;
        RECT 2641.850 51.580 2642.170 51.640 ;
        RECT 2407.710 51.440 2642.170 51.580 ;
        RECT 2407.710 51.380 2408.030 51.440 ;
        RECT 2641.850 51.380 2642.170 51.440 ;
        RECT 2405.410 16.900 2405.730 16.960 ;
        RECT 2407.710 16.900 2408.030 16.960 ;
        RECT 2405.410 16.760 2408.030 16.900 ;
        RECT 2405.410 16.700 2405.730 16.760 ;
        RECT 2407.710 16.700 2408.030 16.760 ;
      LAYER via ;
        RECT 2407.740 51.380 2408.000 51.640 ;
        RECT 2641.880 51.380 2642.140 51.640 ;
        RECT 2405.440 16.700 2405.700 16.960 ;
        RECT 2407.740 16.700 2408.000 16.960 ;
      LAYER met2 ;
        RECT 2641.940 51.670 2642.080 54.000 ;
        RECT 2407.740 51.350 2408.000 51.670 ;
        RECT 2641.880 51.350 2642.140 51.670 ;
        RECT 2407.800 16.990 2407.940 51.350 ;
        RECT 2405.440 16.670 2405.700 16.990 ;
        RECT 2407.740 16.670 2408.000 16.990 ;
        RECT 2405.500 2.400 2405.640 16.670 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 800.100 3.130 800.240 54.000 ;
        RECT 799.640 2.990 800.240 3.130 ;
        RECT 799.640 2.400 799.780 2.990 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 645.080 2.400 645.220 54.000 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2428.870 16.900 2429.190 16.960 ;
        RECT 2435.310 16.900 2435.630 16.960 ;
        RECT 2428.870 16.760 2435.630 16.900 ;
        RECT 2428.870 16.700 2429.190 16.760 ;
        RECT 2435.310 16.700 2435.630 16.760 ;
      LAYER via ;
        RECT 2428.900 16.700 2429.160 16.960 ;
        RECT 2435.340 16.700 2435.600 16.960 ;
      LAYER met2 ;
        RECT 2435.400 16.990 2435.540 54.000 ;
        RECT 2428.900 16.670 2429.160 16.990 ;
        RECT 2435.340 16.670 2435.600 16.990 ;
        RECT 2428.960 2.400 2429.100 16.670 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2446.810 16.900 2447.130 16.960 ;
        RECT 2449.110 16.900 2449.430 16.960 ;
        RECT 2446.810 16.760 2449.430 16.900 ;
        RECT 2446.810 16.700 2447.130 16.760 ;
        RECT 2449.110 16.700 2449.430 16.760 ;
      LAYER via ;
        RECT 2446.840 16.700 2447.100 16.960 ;
        RECT 2449.140 16.700 2449.400 16.960 ;
      LAYER met2 ;
        RECT 2449.200 16.990 2449.340 54.000 ;
        RECT 2446.840 16.670 2447.100 16.990 ;
        RECT 2449.140 16.670 2449.400 16.990 ;
        RECT 2446.900 2.400 2447.040 16.670 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2512.205 20.145 2513.295 20.315 ;
      LAYER mcon ;
        RECT 2513.125 20.145 2513.295 20.315 ;
      LAYER met1 ;
        RECT 2591.710 20.640 2592.030 20.700 ;
        RECT 2587.660 20.500 2592.030 20.640 ;
        RECT 2464.750 20.300 2465.070 20.360 ;
        RECT 2512.145 20.300 2512.435 20.345 ;
        RECT 2464.750 20.160 2512.435 20.300 ;
        RECT 2464.750 20.100 2465.070 20.160 ;
        RECT 2512.145 20.115 2512.435 20.160 ;
        RECT 2513.065 20.300 2513.355 20.345 ;
        RECT 2587.660 20.300 2587.800 20.500 ;
        RECT 2591.710 20.440 2592.030 20.500 ;
        RECT 2513.065 20.160 2587.800 20.300 ;
        RECT 2513.065 20.115 2513.355 20.160 ;
      LAYER via ;
        RECT 2464.780 20.100 2465.040 20.360 ;
        RECT 2591.740 20.440 2592.000 20.700 ;
      LAYER met2 ;
        RECT 2591.800 20.730 2591.940 54.000 ;
        RECT 2591.740 20.410 2592.000 20.730 ;
        RECT 2464.780 20.070 2465.040 20.390 ;
        RECT 2464.840 2.400 2464.980 20.070 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2483.610 2.960 2483.930 3.020 ;
        RECT 2482.690 2.820 2483.930 2.960 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
        RECT 2483.610 2.760 2483.930 2.820 ;
      LAYER via ;
        RECT 2482.720 2.760 2482.980 3.020 ;
        RECT 2483.640 2.760 2483.900 3.020 ;
      LAYER met2 ;
        RECT 2483.700 3.050 2483.840 54.000 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2483.640 2.730 2483.900 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2577.525 19.125 2577.695 20.655 ;
      LAYER mcon ;
        RECT 2577.525 20.485 2577.695 20.655 ;
      LAYER met1 ;
        RECT 2500.630 20.640 2500.950 20.700 ;
        RECT 2511.670 20.640 2511.990 20.700 ;
        RECT 2500.630 20.500 2511.990 20.640 ;
        RECT 2500.630 20.440 2500.950 20.500 ;
        RECT 2511.670 20.440 2511.990 20.500 ;
        RECT 2512.590 20.640 2512.910 20.700 ;
        RECT 2577.465 20.640 2577.755 20.685 ;
        RECT 2512.590 20.500 2577.755 20.640 ;
        RECT 2512.590 20.440 2512.910 20.500 ;
        RECT 2577.465 20.455 2577.755 20.500 ;
        RECT 2577.465 19.280 2577.755 19.325 ;
        RECT 2598.610 19.280 2598.930 19.340 ;
        RECT 2577.465 19.140 2598.930 19.280 ;
        RECT 2577.465 19.095 2577.755 19.140 ;
        RECT 2598.610 19.080 2598.930 19.140 ;
      LAYER via ;
        RECT 2500.660 20.440 2500.920 20.700 ;
        RECT 2511.700 20.440 2511.960 20.700 ;
        RECT 2512.620 20.440 2512.880 20.700 ;
        RECT 2598.640 19.080 2598.900 19.340 ;
      LAYER met2 ;
        RECT 2511.760 20.730 2512.820 20.810 ;
        RECT 2500.660 20.410 2500.920 20.730 ;
        RECT 2511.700 20.670 2512.880 20.730 ;
        RECT 2511.700 20.410 2511.960 20.670 ;
        RECT 2512.620 20.410 2512.880 20.670 ;
        RECT 2500.720 2.400 2500.860 20.410 ;
        RECT 2598.700 19.370 2598.840 54.000 ;
        RECT 2598.640 19.050 2598.900 19.370 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2518.200 2.400 2518.340 54.000 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2536.050 17.580 2536.370 17.640 ;
        RECT 2538.810 17.580 2539.130 17.640 ;
        RECT 2536.050 17.440 2539.130 17.580 ;
        RECT 2536.050 17.380 2536.370 17.440 ;
        RECT 2538.810 17.380 2539.130 17.440 ;
      LAYER via ;
        RECT 2536.080 17.380 2536.340 17.640 ;
        RECT 2538.840 17.380 2539.100 17.640 ;
      LAYER met2 ;
        RECT 2538.900 17.670 2539.040 54.000 ;
        RECT 2536.080 17.350 2536.340 17.670 ;
        RECT 2538.840 17.350 2539.100 17.670 ;
        RECT 2536.140 2.400 2536.280 17.350 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2553.990 17.240 2554.310 17.300 ;
        RECT 2604.590 17.240 2604.910 17.300 ;
        RECT 2553.990 17.100 2604.910 17.240 ;
        RECT 2553.990 17.040 2554.310 17.100 ;
        RECT 2604.590 17.040 2604.910 17.100 ;
      LAYER via ;
        RECT 2554.020 17.040 2554.280 17.300 ;
        RECT 2604.620 17.040 2604.880 17.300 ;
      LAYER met2 ;
        RECT 2604.680 17.330 2604.820 54.000 ;
        RECT 2554.020 17.010 2554.280 17.330 ;
        RECT 2604.620 17.010 2604.880 17.330 ;
        RECT 2554.080 2.400 2554.220 17.010 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2571.930 16.900 2572.250 16.960 ;
        RECT 2611.490 16.900 2611.810 16.960 ;
        RECT 2571.930 16.760 2611.810 16.900 ;
        RECT 2571.930 16.700 2572.250 16.760 ;
        RECT 2611.490 16.700 2611.810 16.760 ;
      LAYER via ;
        RECT 2571.960 16.700 2572.220 16.960 ;
        RECT 2611.520 16.700 2611.780 16.960 ;
      LAYER met2 ;
        RECT 2611.580 16.990 2611.720 54.000 ;
        RECT 2571.960 16.670 2572.220 16.990 ;
        RECT 2611.520 16.670 2611.780 16.990 ;
        RECT 2572.020 2.400 2572.160 16.670 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2589.410 20.300 2589.730 20.360 ;
        RECT 2618.390 20.300 2618.710 20.360 ;
        RECT 2589.410 20.160 2618.710 20.300 ;
        RECT 2589.410 20.100 2589.730 20.160 ;
        RECT 2618.390 20.100 2618.710 20.160 ;
      LAYER via ;
        RECT 2589.440 20.100 2589.700 20.360 ;
        RECT 2618.420 20.100 2618.680 20.360 ;
      LAYER met2 ;
        RECT 2618.480 20.390 2618.620 54.000 ;
        RECT 2589.440 20.070 2589.700 20.390 ;
        RECT 2618.420 20.070 2618.680 20.390 ;
        RECT 2589.500 2.400 2589.640 20.070 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.560 2.400 823.700 54.000 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2607.350 16.560 2607.670 16.620 ;
        RECT 2624.830 16.560 2625.150 16.620 ;
        RECT 2607.350 16.420 2625.150 16.560 ;
        RECT 2607.350 16.360 2607.670 16.420 ;
        RECT 2624.830 16.360 2625.150 16.420 ;
      LAYER via ;
        RECT 2607.380 16.360 2607.640 16.620 ;
        RECT 2624.860 16.360 2625.120 16.620 ;
      LAYER met2 ;
        RECT 2625.840 52.770 2625.980 54.000 ;
        RECT 2624.920 52.630 2625.980 52.770 ;
        RECT 2624.920 16.650 2625.060 52.630 ;
        RECT 2607.380 16.330 2607.640 16.650 ;
        RECT 2624.860 16.330 2625.120 16.650 ;
        RECT 2607.440 2.400 2607.580 16.330 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2625.290 17.580 2625.610 17.640 ;
        RECT 2631.730 17.580 2632.050 17.640 ;
        RECT 2625.290 17.440 2632.050 17.580 ;
        RECT 2625.290 17.380 2625.610 17.440 ;
        RECT 2631.730 17.380 2632.050 17.440 ;
      LAYER via ;
        RECT 2625.320 17.380 2625.580 17.640 ;
        RECT 2631.760 17.380 2632.020 17.640 ;
      LAYER met2 ;
        RECT 2631.820 53.990 2633.340 54.000 ;
        RECT 2631.820 17.670 2631.960 53.990 ;
        RECT 2625.320 17.350 2625.580 17.670 ;
        RECT 2631.760 17.350 2632.020 17.670 ;
        RECT 2625.380 2.400 2625.520 17.350 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2643.230 17.580 2643.550 17.640 ;
        RECT 2649.210 17.580 2649.530 17.640 ;
        RECT 2643.230 17.440 2649.530 17.580 ;
        RECT 2643.230 17.380 2643.550 17.440 ;
        RECT 2649.210 17.380 2649.530 17.440 ;
      LAYER via ;
        RECT 2643.260 17.380 2643.520 17.640 ;
        RECT 2649.240 17.380 2649.500 17.640 ;
      LAYER met2 ;
        RECT 2649.300 17.670 2649.440 54.000 ;
        RECT 2643.260 17.350 2643.520 17.670 ;
        RECT 2649.240 17.350 2649.500 17.670 ;
        RECT 2643.320 2.400 2643.460 17.350 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2663.100 17.410 2663.240 54.000 ;
        RECT 2661.260 17.270 2663.240 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2678.650 16.560 2678.970 16.620 ;
        RECT 2683.710 16.560 2684.030 16.620 ;
        RECT 2678.650 16.420 2684.030 16.560 ;
        RECT 2678.650 16.360 2678.970 16.420 ;
        RECT 2683.710 16.360 2684.030 16.420 ;
      LAYER via ;
        RECT 2678.680 16.360 2678.940 16.620 ;
        RECT 2683.740 16.360 2684.000 16.620 ;
      LAYER met2 ;
        RECT 2683.800 16.650 2683.940 54.000 ;
        RECT 2678.680 16.330 2678.940 16.650 ;
        RECT 2683.740 16.330 2684.000 16.650 ;
        RECT 2678.740 2.400 2678.880 16.330 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2696.590 16.900 2696.910 16.960 ;
        RECT 2728.790 16.900 2729.110 16.960 ;
        RECT 2696.590 16.760 2729.110 16.900 ;
        RECT 2696.590 16.700 2696.910 16.760 ;
        RECT 2728.790 16.700 2729.110 16.760 ;
      LAYER via ;
        RECT 2696.620 16.700 2696.880 16.960 ;
        RECT 2728.820 16.700 2729.080 16.960 ;
      LAYER met2 ;
        RECT 2728.880 16.990 2729.020 54.000 ;
        RECT 2696.620 16.670 2696.880 16.990 ;
        RECT 2728.820 16.670 2729.080 16.990 ;
        RECT 2696.680 2.400 2696.820 16.670 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2714.530 17.240 2714.850 17.300 ;
        RECT 2718.210 17.240 2718.530 17.300 ;
        RECT 2714.530 17.100 2718.530 17.240 ;
        RECT 2714.530 17.040 2714.850 17.100 ;
        RECT 2718.210 17.040 2718.530 17.100 ;
      LAYER via ;
        RECT 2714.560 17.040 2714.820 17.300 ;
        RECT 2718.240 17.040 2718.500 17.300 ;
      LAYER met2 ;
        RECT 2718.300 17.330 2718.440 54.000 ;
        RECT 2714.560 17.010 2714.820 17.330 ;
        RECT 2718.240 17.010 2718.500 17.330 ;
        RECT 2714.620 2.400 2714.760 17.010 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2732.470 16.900 2732.790 16.960 ;
        RECT 2738.450 16.900 2738.770 16.960 ;
        RECT 2732.470 16.760 2738.770 16.900 ;
        RECT 2732.470 16.700 2732.790 16.760 ;
        RECT 2738.450 16.700 2738.770 16.760 ;
      LAYER via ;
        RECT 2732.500 16.700 2732.760 16.960 ;
        RECT 2738.480 16.700 2738.740 16.960 ;
      LAYER met2 ;
        RECT 2738.540 16.990 2738.680 54.000 ;
        RECT 2732.500 16.670 2732.760 16.990 ;
        RECT 2738.480 16.670 2738.740 16.990 ;
        RECT 2732.560 2.400 2732.700 16.670 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2750.410 20.640 2750.730 20.700 ;
        RECT 2752.710 20.640 2753.030 20.700 ;
        RECT 2750.410 20.500 2753.030 20.640 ;
        RECT 2750.410 20.440 2750.730 20.500 ;
        RECT 2752.710 20.440 2753.030 20.500 ;
      LAYER via ;
        RECT 2750.440 20.440 2750.700 20.700 ;
        RECT 2752.740 20.440 2753.000 20.700 ;
      LAYER met2 ;
        RECT 2752.800 20.730 2752.940 54.000 ;
        RECT 2750.440 20.410 2750.700 20.730 ;
        RECT 2752.740 20.410 2753.000 20.730 ;
        RECT 2750.500 2.400 2750.640 20.410 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2766.970 14.180 2767.290 14.240 ;
        RECT 2766.970 14.040 2768.120 14.180 ;
        RECT 2766.970 13.980 2767.290 14.040 ;
        RECT 2767.980 13.900 2768.120 14.040 ;
        RECT 2767.890 13.640 2768.210 13.900 ;
      LAYER via ;
        RECT 2767.000 13.980 2767.260 14.240 ;
        RECT 2767.920 13.640 2768.180 13.900 ;
      LAYER met2 ;
        RECT 2767.060 14.270 2767.200 54.000 ;
        RECT 2767.000 13.950 2767.260 14.270 ;
        RECT 2767.920 13.610 2768.180 13.930 ;
        RECT 2767.980 2.400 2768.120 13.610 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 19.960 841.270 20.020 ;
        RECT 1127.990 19.960 1128.310 20.020 ;
        RECT 840.950 19.820 1128.310 19.960 ;
        RECT 840.950 19.760 841.270 19.820 ;
        RECT 1127.990 19.760 1128.310 19.820 ;
      LAYER via ;
        RECT 840.980 19.760 841.240 20.020 ;
        RECT 1128.020 19.760 1128.280 20.020 ;
      LAYER met2 ;
        RECT 1128.080 20.050 1128.220 54.000 ;
        RECT 840.980 19.730 841.240 20.050 ;
        RECT 1128.020 19.730 1128.280 20.050 ;
        RECT 841.040 2.400 841.180 19.730 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2777.090 20.640 2777.410 20.700 ;
        RECT 2785.830 20.640 2786.150 20.700 ;
        RECT 2777.090 20.500 2786.150 20.640 ;
        RECT 2777.090 20.440 2777.410 20.500 ;
        RECT 2785.830 20.440 2786.150 20.500 ;
      LAYER via ;
        RECT 2777.120 20.440 2777.380 20.700 ;
        RECT 2785.860 20.440 2786.120 20.700 ;
      LAYER met2 ;
        RECT 2777.180 20.730 2777.320 54.000 ;
        RECT 2777.120 20.410 2777.380 20.730 ;
        RECT 2785.860 20.410 2786.120 20.730 ;
        RECT 2785.920 2.400 2786.060 20.410 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2784.450 18.260 2784.770 18.320 ;
        RECT 2803.770 18.260 2804.090 18.320 ;
        RECT 2784.450 18.120 2804.090 18.260 ;
        RECT 2784.450 18.060 2784.770 18.120 ;
        RECT 2803.770 18.060 2804.090 18.120 ;
      LAYER via ;
        RECT 2784.480 18.060 2784.740 18.320 ;
        RECT 2803.800 18.060 2804.060 18.320 ;
      LAYER met2 ;
        RECT 2784.540 18.350 2784.680 54.000 ;
        RECT 2784.480 18.030 2784.740 18.350 ;
        RECT 2803.800 18.030 2804.060 18.350 ;
        RECT 2803.860 2.400 2804.000 18.030 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2815.270 17.580 2815.590 17.640 ;
        RECT 2821.710 17.580 2822.030 17.640 ;
        RECT 2815.270 17.440 2822.030 17.580 ;
        RECT 2815.270 17.380 2815.590 17.440 ;
        RECT 2821.710 17.380 2822.030 17.440 ;
      LAYER via ;
        RECT 2815.300 17.380 2815.560 17.640 ;
        RECT 2821.740 17.380 2822.000 17.640 ;
      LAYER met2 ;
        RECT 2815.360 17.670 2815.500 54.000 ;
        RECT 2815.300 17.350 2815.560 17.670 ;
        RECT 2821.740 17.350 2822.000 17.670 ;
        RECT 2821.800 2.400 2821.940 17.350 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2786.750 16.220 2787.070 16.280 ;
        RECT 2839.190 16.220 2839.510 16.280 ;
        RECT 2786.750 16.080 2839.510 16.220 ;
        RECT 2786.750 16.020 2787.070 16.080 ;
        RECT 2839.190 16.020 2839.510 16.080 ;
      LAYER via ;
        RECT 2786.780 16.020 2787.040 16.280 ;
        RECT 2839.220 16.020 2839.480 16.280 ;
      LAYER met2 ;
        RECT 2786.840 16.310 2786.980 54.000 ;
        RECT 2786.780 15.990 2787.040 16.310 ;
        RECT 2839.220 15.990 2839.480 16.310 ;
        RECT 2839.280 2.400 2839.420 15.990 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2823.165 15.045 2823.335 16.915 ;
      LAYER mcon ;
        RECT 2823.165 16.745 2823.335 16.915 ;
      LAYER met1 ;
        RECT 2823.105 16.900 2823.395 16.945 ;
        RECT 2857.130 16.900 2857.450 16.960 ;
        RECT 2823.105 16.760 2857.450 16.900 ;
        RECT 2823.105 16.715 2823.395 16.760 ;
        RECT 2857.130 16.700 2857.450 16.760 ;
        RECT 2794.110 15.200 2794.430 15.260 ;
        RECT 2823.105 15.200 2823.395 15.245 ;
        RECT 2794.110 15.060 2823.395 15.200 ;
        RECT 2794.110 15.000 2794.430 15.060 ;
        RECT 2823.105 15.015 2823.395 15.060 ;
      LAYER via ;
        RECT 2857.160 16.700 2857.420 16.960 ;
        RECT 2794.140 15.000 2794.400 15.260 ;
      LAYER met2 ;
        RECT 2794.200 15.290 2794.340 54.000 ;
        RECT 2857.160 16.670 2857.420 16.990 ;
        RECT 2794.140 14.970 2794.400 15.290 ;
        RECT 2857.220 2.400 2857.360 16.670 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2793.650 19.280 2793.970 19.340 ;
        RECT 2875.070 19.280 2875.390 19.340 ;
        RECT 2793.650 19.140 2875.390 19.280 ;
        RECT 2793.650 19.080 2793.970 19.140 ;
        RECT 2875.070 19.080 2875.390 19.140 ;
      LAYER via ;
        RECT 2793.680 19.080 2793.940 19.340 ;
        RECT 2875.100 19.080 2875.360 19.340 ;
      LAYER met2 ;
        RECT 2793.740 19.370 2793.880 54.000 ;
        RECT 2793.680 19.050 2793.940 19.370 ;
        RECT 2875.100 19.050 2875.360 19.370 ;
        RECT 2875.160 2.400 2875.300 19.050 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2801.010 18.600 2801.330 18.660 ;
        RECT 2893.010 18.600 2893.330 18.660 ;
        RECT 2801.010 18.460 2893.330 18.600 ;
        RECT 2801.010 18.400 2801.330 18.460 ;
        RECT 2893.010 18.400 2893.330 18.460 ;
      LAYER via ;
        RECT 2801.040 18.400 2801.300 18.660 ;
        RECT 2893.040 18.400 2893.300 18.660 ;
      LAYER met2 ;
        RECT 2801.100 18.690 2801.240 54.000 ;
        RECT 2801.040 18.370 2801.300 18.690 ;
        RECT 2893.040 18.370 2893.300 18.690 ;
        RECT 2893.100 2.400 2893.240 18.370 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2807.910 18.260 2808.230 18.320 ;
        RECT 2910.950 18.260 2911.270 18.320 ;
        RECT 2807.910 18.120 2911.270 18.260 ;
        RECT 2807.910 18.060 2808.230 18.120 ;
        RECT 2910.950 18.060 2911.270 18.120 ;
      LAYER via ;
        RECT 2807.940 18.060 2808.200 18.320 ;
        RECT 2910.980 18.060 2911.240 18.320 ;
      LAYER met2 ;
        RECT 2808.000 18.350 2808.140 54.000 ;
        RECT 2807.940 18.030 2808.200 18.350 ;
        RECT 2910.980 18.030 2911.240 18.350 ;
        RECT 2911.040 2.400 2911.180 18.030 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.980 2.400 859.120 54.000 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 877.380 33.730 877.520 54.000 ;
        RECT 876.920 33.590 877.520 33.730 ;
        RECT 876.920 2.400 877.060 33.590 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.770 2.960 895.090 3.020 ;
        RECT 896.610 2.960 896.930 3.020 ;
        RECT 894.770 2.820 896.930 2.960 ;
        RECT 894.770 2.760 895.090 2.820 ;
        RECT 896.610 2.760 896.930 2.820 ;
      LAYER via ;
        RECT 894.800 2.760 895.060 3.020 ;
        RECT 896.640 2.760 896.900 3.020 ;
      LAYER met2 ;
        RECT 896.700 3.050 896.840 54.000 ;
        RECT 894.800 2.730 895.060 3.050 ;
        RECT 896.640 2.730 896.900 3.050 ;
        RECT 894.860 2.400 895.000 2.730 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.800 2.400 912.940 54.000 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 931.200 3.130 931.340 54.000 ;
        RECT 930.280 2.990 931.340 3.130 ;
        RECT 930.280 2.400 930.420 2.990 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 16.900 948.450 16.960 ;
        RECT 951.810 16.900 952.130 16.960 ;
        RECT 948.130 16.760 952.130 16.900 ;
        RECT 948.130 16.700 948.450 16.760 ;
        RECT 951.810 16.700 952.130 16.760 ;
      LAYER via ;
        RECT 948.160 16.700 948.420 16.960 ;
        RECT 951.840 16.700 952.100 16.960 ;
      LAYER met2 ;
        RECT 951.900 16.990 952.040 54.000 ;
        RECT 948.160 16.670 948.420 16.990 ;
        RECT 951.840 16.670 952.100 16.990 ;
        RECT 948.220 2.400 948.360 16.670 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.070 15.540 966.390 15.600 ;
        RECT 972.510 15.540 972.830 15.600 ;
        RECT 966.070 15.400 972.830 15.540 ;
        RECT 966.070 15.340 966.390 15.400 ;
        RECT 972.510 15.340 972.830 15.400 ;
      LAYER via ;
        RECT 966.100 15.340 966.360 15.600 ;
        RECT 972.540 15.340 972.800 15.600 ;
      LAYER met2 ;
        RECT 972.600 15.630 972.740 54.000 ;
        RECT 966.100 15.310 966.360 15.630 ;
        RECT 972.540 15.310 972.800 15.630 ;
        RECT 966.160 2.400 966.300 15.310 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.100 2.400 984.240 54.000 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.560 36.450 662.700 54.000 ;
        RECT 662.560 36.310 663.160 36.450 ;
        RECT 663.020 2.400 663.160 36.310 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1736.645 11.305 1738.195 11.475 ;
      LAYER mcon ;
        RECT 1738.025 11.305 1738.195 11.475 ;
      LAYER met1 ;
        RECT 1001.950 11.460 1002.270 11.520 ;
        RECT 1736.585 11.460 1736.875 11.505 ;
        RECT 1001.950 11.320 1736.875 11.460 ;
        RECT 1001.950 11.260 1002.270 11.320 ;
        RECT 1736.585 11.275 1736.875 11.320 ;
        RECT 1737.965 11.460 1738.255 11.505 ;
        RECT 2187.830 11.460 2188.150 11.520 ;
        RECT 1737.965 11.320 2188.150 11.460 ;
        RECT 1737.965 11.275 1738.255 11.320 ;
        RECT 2187.830 11.260 2188.150 11.320 ;
      LAYER via ;
        RECT 1001.980 11.260 1002.240 11.520 ;
        RECT 2187.860 11.260 2188.120 11.520 ;
      LAYER met2 ;
        RECT 2187.920 11.550 2188.060 54.000 ;
        RECT 1001.980 11.230 1002.240 11.550 ;
        RECT 2187.860 11.230 2188.120 11.550 ;
        RECT 1002.040 2.400 1002.180 11.230 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.900 12.650 1021.040 54.000 ;
        RECT 1019.520 12.510 1021.040 12.650 ;
        RECT 1019.520 2.400 1019.660 12.510 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 20.300 1037.690 20.360 ;
        RECT 1041.510 20.300 1041.830 20.360 ;
        RECT 1037.370 20.160 1041.830 20.300 ;
        RECT 1037.370 20.100 1037.690 20.160 ;
        RECT 1041.510 20.100 1041.830 20.160 ;
      LAYER via ;
        RECT 1037.400 20.100 1037.660 20.360 ;
        RECT 1041.540 20.100 1041.800 20.360 ;
      LAYER met2 ;
        RECT 1041.600 20.390 1041.740 54.000 ;
        RECT 1037.400 20.070 1037.660 20.390 ;
        RECT 1041.540 20.070 1041.800 20.390 ;
        RECT 1037.460 2.400 1037.600 20.070 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.400 2.400 1055.540 54.000 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1073.250 11.800 1073.570 11.860 ;
        RECT 1714.490 11.800 1714.810 11.860 ;
        RECT 1073.250 11.660 1714.810 11.800 ;
        RECT 1073.250 11.600 1073.570 11.660 ;
        RECT 1714.490 11.600 1714.810 11.660 ;
        RECT 1738.410 11.800 1738.730 11.860 ;
        RECT 2209.910 11.800 2210.230 11.860 ;
        RECT 1738.410 11.660 2210.230 11.800 ;
        RECT 1738.410 11.600 1738.730 11.660 ;
        RECT 2209.910 11.600 2210.230 11.660 ;
      LAYER via ;
        RECT 1073.280 11.600 1073.540 11.860 ;
        RECT 1714.520 11.600 1714.780 11.860 ;
        RECT 1738.440 11.600 1738.700 11.860 ;
        RECT 2209.940 11.600 2210.200 11.860 ;
      LAYER met2 ;
        RECT 2211.840 44.610 2211.980 54.000 ;
        RECT 2210.000 44.470 2211.980 44.610 ;
        RECT 1073.280 11.570 1073.540 11.890 ;
        RECT 1714.510 11.715 1714.790 12.085 ;
        RECT 1738.430 11.715 1738.710 12.085 ;
        RECT 2210.000 11.890 2210.140 44.470 ;
        RECT 1714.520 11.570 1714.780 11.715 ;
        RECT 1738.440 11.570 1738.700 11.715 ;
        RECT 2209.940 11.570 2210.200 11.890 ;
        RECT 1073.340 2.400 1073.480 11.570 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 1714.510 11.760 1714.790 12.040 ;
        RECT 1738.430 11.760 1738.710 12.040 ;
      LAYER met3 ;
        RECT 1714.485 12.050 1714.815 12.065 ;
        RECT 1738.405 12.050 1738.735 12.065 ;
        RECT 1714.485 11.750 1738.735 12.050 ;
        RECT 1714.485 11.735 1714.815 11.750 ;
        RECT 1738.405 11.735 1738.735 11.750 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.730 16.900 1091.050 16.960 ;
        RECT 1096.250 16.900 1096.570 16.960 ;
        RECT 1090.730 16.760 1096.570 16.900 ;
        RECT 1090.730 16.700 1091.050 16.760 ;
        RECT 1096.250 16.700 1096.570 16.760 ;
      LAYER via ;
        RECT 1090.760 16.700 1091.020 16.960 ;
        RECT 1096.280 16.700 1096.540 16.960 ;
      LAYER met2 ;
        RECT 1096.340 16.990 1096.480 54.000 ;
        RECT 1090.760 16.670 1091.020 16.990 ;
        RECT 1096.280 16.670 1096.540 16.990 ;
        RECT 1090.820 2.400 1090.960 16.670 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.600 17.410 1110.740 54.000 ;
        RECT 1108.760 17.270 1110.740 17.410 ;
        RECT 1108.760 2.400 1108.900 17.270 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.610 20.300 1126.930 20.360 ;
        RECT 1376.390 20.300 1376.710 20.360 ;
        RECT 1126.610 20.160 1376.710 20.300 ;
        RECT 1126.610 20.100 1126.930 20.160 ;
        RECT 1376.390 20.100 1376.710 20.160 ;
      LAYER via ;
        RECT 1126.640 20.100 1126.900 20.360 ;
        RECT 1376.420 20.100 1376.680 20.360 ;
      LAYER met2 ;
        RECT 1376.480 20.390 1376.620 54.000 ;
        RECT 1126.640 20.070 1126.900 20.390 ;
        RECT 1376.420 20.070 1376.680 20.390 ;
        RECT 1126.700 2.400 1126.840 20.070 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1144.550 12.140 1144.870 12.200 ;
        RECT 2076.970 12.140 2077.290 12.200 ;
        RECT 1144.550 12.000 2077.290 12.140 ;
        RECT 1144.550 11.940 1144.870 12.000 ;
        RECT 2076.970 11.940 2077.290 12.000 ;
        RECT 2124.810 12.140 2125.130 12.200 ;
        RECT 2173.570 12.140 2173.890 12.200 ;
        RECT 2124.810 12.000 2173.890 12.140 ;
        RECT 2124.810 11.940 2125.130 12.000 ;
        RECT 2173.570 11.940 2173.890 12.000 ;
        RECT 2210.370 11.800 2210.690 11.860 ;
        RECT 2236.130 11.800 2236.450 11.860 ;
        RECT 2210.370 11.660 2236.450 11.800 ;
        RECT 2210.370 11.600 2210.690 11.660 ;
        RECT 2236.130 11.600 2236.450 11.660 ;
      LAYER via ;
        RECT 1144.580 11.940 1144.840 12.200 ;
        RECT 2077.000 11.940 2077.260 12.200 ;
        RECT 2124.840 11.940 2125.100 12.200 ;
        RECT 2173.600 11.940 2173.860 12.200 ;
        RECT 2210.400 11.600 2210.660 11.860 ;
        RECT 2236.160 11.600 2236.420 11.860 ;
      LAYER met2 ;
        RECT 2234.840 49.485 2234.980 54.000 ;
        RECT 2234.770 49.115 2235.050 49.485 ;
        RECT 2236.150 48.435 2236.430 48.805 ;
        RECT 1144.580 11.910 1144.840 12.230 ;
        RECT 2077.000 12.085 2077.260 12.230 ;
        RECT 2124.840 12.085 2125.100 12.230 ;
        RECT 2173.600 12.085 2173.860 12.230 ;
        RECT 1144.640 2.400 1144.780 11.910 ;
        RECT 2076.990 11.715 2077.270 12.085 ;
        RECT 2124.830 11.715 2125.110 12.085 ;
        RECT 2173.590 11.715 2173.870 12.085 ;
        RECT 2210.390 11.715 2210.670 12.085 ;
        RECT 2236.220 11.890 2236.360 48.435 ;
        RECT 2210.400 11.570 2210.660 11.715 ;
        RECT 2236.160 11.570 2236.420 11.890 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
      LAYER via2 ;
        RECT 2234.770 49.160 2235.050 49.440 ;
        RECT 2236.150 48.480 2236.430 48.760 ;
        RECT 2076.990 11.760 2077.270 12.040 ;
        RECT 2124.830 11.760 2125.110 12.040 ;
        RECT 2173.590 11.760 2173.870 12.040 ;
        RECT 2210.390 11.760 2210.670 12.040 ;
      LAYER met3 ;
        RECT 2234.745 49.450 2235.075 49.465 ;
        RECT 2234.745 49.150 2237.130 49.450 ;
        RECT 2234.745 49.135 2235.075 49.150 ;
        RECT 2236.125 48.770 2236.455 48.785 ;
        RECT 2236.830 48.770 2237.130 49.150 ;
        RECT 2236.125 48.470 2237.130 48.770 ;
        RECT 2236.125 48.455 2236.455 48.470 ;
        RECT 2076.965 12.050 2077.295 12.065 ;
        RECT 2124.805 12.050 2125.135 12.065 ;
        RECT 2076.965 11.750 2125.135 12.050 ;
        RECT 2076.965 11.735 2077.295 11.750 ;
        RECT 2124.805 11.735 2125.135 11.750 ;
        RECT 2173.565 12.050 2173.895 12.065 ;
        RECT 2210.365 12.050 2210.695 12.065 ;
        RECT 2173.565 11.750 2210.695 12.050 ;
        RECT 2173.565 11.735 2173.895 11.750 ;
        RECT 2210.365 11.735 2210.695 11.750 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 16.900 1162.810 16.960 ;
        RECT 1165.710 16.900 1166.030 16.960 ;
        RECT 1162.490 16.760 1166.030 16.900 ;
        RECT 1162.490 16.700 1162.810 16.760 ;
        RECT 1165.710 16.700 1166.030 16.760 ;
      LAYER via ;
        RECT 1162.520 16.700 1162.780 16.960 ;
        RECT 1165.740 16.700 1166.000 16.960 ;
      LAYER met2 ;
        RECT 1165.800 16.990 1165.940 54.000 ;
        RECT 1162.520 16.670 1162.780 16.990 ;
        RECT 1165.740 16.670 1166.000 16.990 ;
        RECT 1162.580 2.400 1162.720 16.670 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2086.260 51.525 2086.400 54.000 ;
        RECT 680.430 51.155 680.710 51.525 ;
        RECT 2086.190 51.155 2086.470 51.525 ;
        RECT 680.500 2.400 680.640 51.155 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 680.430 51.200 680.710 51.480 ;
        RECT 2086.190 51.200 2086.470 51.480 ;
      LAYER met3 ;
        RECT 680.405 51.490 680.735 51.505 ;
        RECT 2086.165 51.490 2086.495 51.505 ;
        RECT 680.405 51.190 2086.495 51.490 ;
        RECT 680.405 51.175 680.735 51.190 ;
        RECT 2086.165 51.175 2086.495 51.190 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 12.480 1180.290 12.540 ;
        RECT 1179.970 12.340 2234.060 12.480 ;
        RECT 1179.970 12.280 1180.290 12.340 ;
        RECT 2233.920 12.140 2234.060 12.340 ;
        RECT 2245.330 12.140 2245.650 12.200 ;
        RECT 2233.920 12.000 2245.650 12.140 ;
        RECT 2245.330 11.940 2245.650 12.000 ;
      LAYER via ;
        RECT 1180.000 12.280 1180.260 12.540 ;
        RECT 2245.360 11.940 2245.620 12.200 ;
      LAYER met2 ;
        RECT 2245.880 14.010 2246.020 54.000 ;
        RECT 2245.420 13.870 2246.020 14.010 ;
        RECT 1180.000 12.250 1180.260 12.570 ;
        RECT 1180.060 2.400 1180.200 12.250 ;
        RECT 2245.420 12.230 2245.560 13.870 ;
        RECT 2245.360 11.910 2245.620 12.230 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1197.910 17.580 1198.230 17.640 ;
        RECT 1200.210 17.580 1200.530 17.640 ;
        RECT 1197.910 17.440 1200.530 17.580 ;
        RECT 1197.910 17.380 1198.230 17.440 ;
        RECT 1200.210 17.380 1200.530 17.440 ;
      LAYER via ;
        RECT 1197.940 17.380 1198.200 17.640 ;
        RECT 1200.240 17.380 1200.500 17.640 ;
      LAYER met2 ;
        RECT 1200.300 17.670 1200.440 54.000 ;
        RECT 1197.940 17.350 1198.200 17.670 ;
        RECT 1200.240 17.350 1200.500 17.670 ;
        RECT 1198.000 2.400 1198.140 17.350 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1215.850 12.820 1216.170 12.880 ;
        RECT 2257.750 12.820 2258.070 12.880 ;
        RECT 1215.850 12.680 2258.070 12.820 ;
        RECT 1215.850 12.620 1216.170 12.680 ;
        RECT 2257.750 12.620 2258.070 12.680 ;
      LAYER via ;
        RECT 1215.880 12.620 1216.140 12.880 ;
        RECT 2257.780 12.620 2258.040 12.880 ;
      LAYER met2 ;
        RECT 2257.840 12.910 2257.980 54.000 ;
        RECT 1215.880 12.590 1216.140 12.910 ;
        RECT 2257.780 12.590 2258.040 12.910 ;
        RECT 1215.940 2.400 1216.080 12.590 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 19.960 1234.110 20.020 ;
        RECT 1431.590 19.960 1431.910 20.020 ;
        RECT 1233.790 19.820 1431.910 19.960 ;
        RECT 1233.790 19.760 1234.110 19.820 ;
        RECT 1431.590 19.760 1431.910 19.820 ;
      LAYER via ;
        RECT 1233.820 19.760 1234.080 20.020 ;
        RECT 1431.620 19.760 1431.880 20.020 ;
      LAYER met2 ;
        RECT 1431.680 20.050 1431.820 54.000 ;
        RECT 1233.820 19.730 1234.080 20.050 ;
        RECT 1431.620 19.730 1431.880 20.050 ;
        RECT 1233.880 2.400 1234.020 19.730 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1251.730 18.260 1252.050 18.320 ;
        RECT 1521.290 18.260 1521.610 18.320 ;
        RECT 1251.730 18.120 1521.610 18.260 ;
        RECT 1251.730 18.060 1252.050 18.120 ;
        RECT 1521.290 18.060 1521.610 18.120 ;
      LAYER via ;
        RECT 1251.760 18.060 1252.020 18.320 ;
        RECT 1521.320 18.060 1521.580 18.320 ;
      LAYER met2 ;
        RECT 1521.380 18.350 1521.520 54.000 ;
        RECT 1251.760 18.030 1252.020 18.350 ;
        RECT 1521.320 18.030 1521.580 18.350 ;
        RECT 1251.820 2.400 1251.960 18.030 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 14.520 1269.530 14.580 ;
        RECT 1462.870 14.520 1463.190 14.580 ;
        RECT 1269.210 14.380 1463.190 14.520 ;
        RECT 1269.210 14.320 1269.530 14.380 ;
        RECT 1462.870 14.320 1463.190 14.380 ;
        RECT 1462.870 8.740 1463.190 8.800 ;
        RECT 2271.090 8.740 2271.410 8.800 ;
        RECT 1462.870 8.600 2271.410 8.740 ;
        RECT 1462.870 8.540 1463.190 8.600 ;
        RECT 2271.090 8.540 2271.410 8.600 ;
      LAYER via ;
        RECT 1269.240 14.320 1269.500 14.580 ;
        RECT 1462.900 14.320 1463.160 14.580 ;
        RECT 1462.900 8.540 1463.160 8.800 ;
        RECT 2271.120 8.540 2271.380 8.800 ;
      LAYER met2 ;
        RECT 2274.860 37.130 2275.000 54.000 ;
        RECT 2271.180 36.990 2275.000 37.130 ;
        RECT 1269.240 14.290 1269.500 14.610 ;
        RECT 1462.900 14.290 1463.160 14.610 ;
        RECT 1269.300 2.400 1269.440 14.290 ;
        RECT 1462.960 8.830 1463.100 14.290 ;
        RECT 2271.180 8.830 2271.320 36.990 ;
        RECT 1462.900 8.510 1463.160 8.830 ;
        RECT 2271.120 8.510 2271.380 8.830 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.150 19.620 1287.470 19.680 ;
        RECT 1500.590 19.620 1500.910 19.680 ;
        RECT 1287.150 19.480 1500.910 19.620 ;
        RECT 1287.150 19.420 1287.470 19.480 ;
        RECT 1500.590 19.420 1500.910 19.480 ;
      LAYER via ;
        RECT 1287.180 19.420 1287.440 19.680 ;
        RECT 1500.620 19.420 1500.880 19.680 ;
      LAYER met2 ;
        RECT 1500.680 19.710 1500.820 54.000 ;
        RECT 1287.180 19.390 1287.440 19.710 ;
        RECT 1500.620 19.390 1500.880 19.710 ;
        RECT 1287.240 2.400 1287.380 19.390 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1305.090 14.180 1305.410 14.240 ;
        RECT 1555.790 14.180 1556.110 14.240 ;
        RECT 1305.090 14.040 1556.110 14.180 ;
        RECT 1305.090 13.980 1305.410 14.040 ;
        RECT 1555.790 13.980 1556.110 14.040 ;
        RECT 1555.790 8.400 1556.110 8.460 ;
        RECT 2284.890 8.400 2285.210 8.460 ;
        RECT 1555.790 8.260 2285.210 8.400 ;
        RECT 1555.790 8.200 1556.110 8.260 ;
        RECT 2284.890 8.200 2285.210 8.260 ;
      LAYER via ;
        RECT 1305.120 13.980 1305.380 14.240 ;
        RECT 1555.820 13.980 1556.080 14.240 ;
        RECT 1555.820 8.200 1556.080 8.460 ;
        RECT 2284.920 8.200 2285.180 8.460 ;
      LAYER met2 ;
        RECT 1305.120 13.950 1305.380 14.270 ;
        RECT 1555.820 13.950 1556.080 14.270 ;
        RECT 1305.180 2.400 1305.320 13.950 ;
        RECT 1555.880 8.490 1556.020 13.950 ;
        RECT 2284.980 8.490 2285.120 54.000 ;
        RECT 1555.820 8.170 1556.080 8.490 ;
        RECT 2284.920 8.170 2285.180 8.490 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1323.030 18.600 1323.350 18.660 ;
        RECT 1590.290 18.600 1590.610 18.660 ;
        RECT 1323.030 18.460 1590.610 18.600 ;
        RECT 1323.030 18.400 1323.350 18.460 ;
        RECT 1590.290 18.400 1590.610 18.460 ;
      LAYER via ;
        RECT 1323.060 18.400 1323.320 18.660 ;
        RECT 1590.320 18.400 1590.580 18.660 ;
      LAYER met2 ;
        RECT 1590.380 18.690 1590.520 54.000 ;
        RECT 1323.060 18.370 1323.320 18.690 ;
        RECT 1590.320 18.370 1590.580 18.690 ;
        RECT 1323.120 2.400 1323.260 18.370 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1461.490 40.360 1461.810 40.420 ;
        RECT 2297.770 40.360 2298.090 40.420 ;
        RECT 1461.490 40.220 2298.090 40.360 ;
        RECT 1461.490 40.160 1461.810 40.220 ;
        RECT 2297.770 40.160 2298.090 40.220 ;
        RECT 1340.510 17.920 1340.830 17.980 ;
        RECT 1461.490 17.920 1461.810 17.980 ;
        RECT 1340.510 17.780 1461.810 17.920 ;
        RECT 1340.510 17.720 1340.830 17.780 ;
        RECT 1461.490 17.720 1461.810 17.780 ;
      LAYER via ;
        RECT 1461.520 40.160 1461.780 40.420 ;
        RECT 2297.800 40.160 2298.060 40.420 ;
        RECT 1340.540 17.720 1340.800 17.980 ;
        RECT 1461.520 17.720 1461.780 17.980 ;
      LAYER met2 ;
        RECT 2297.860 40.450 2298.000 54.000 ;
        RECT 1461.520 40.130 1461.780 40.450 ;
        RECT 2297.800 40.130 2298.060 40.450 ;
        RECT 1461.580 18.010 1461.720 40.130 ;
        RECT 1340.540 17.690 1340.800 18.010 ;
        RECT 1461.520 17.690 1461.780 18.010 ;
        RECT 1340.600 2.400 1340.740 17.690 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 20.640 698.670 20.700 ;
        RECT 703.410 20.640 703.730 20.700 ;
        RECT 698.350 20.500 703.730 20.640 ;
        RECT 698.350 20.440 698.670 20.500 ;
        RECT 703.410 20.440 703.730 20.500 ;
      LAYER via ;
        RECT 698.380 20.440 698.640 20.700 ;
        RECT 703.440 20.440 703.700 20.700 ;
      LAYER met2 ;
        RECT 703.500 20.730 703.640 54.000 ;
        RECT 698.380 20.410 698.640 20.730 ;
        RECT 703.440 20.410 703.700 20.730 ;
        RECT 698.440 2.400 698.580 20.410 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2030.125 15.045 2030.295 17.595 ;
      LAYER mcon ;
        RECT 2030.125 17.425 2030.295 17.595 ;
      LAYER met1 ;
        RECT 1358.450 17.580 1358.770 17.640 ;
        RECT 2030.065 17.580 2030.355 17.625 ;
        RECT 1358.450 17.440 2030.355 17.580 ;
        RECT 1358.450 17.380 1358.770 17.440 ;
        RECT 2030.065 17.395 2030.355 17.440 ;
        RECT 2030.065 15.200 2030.355 15.245 ;
        RECT 2052.590 15.200 2052.910 15.260 ;
        RECT 2030.065 15.060 2052.910 15.200 ;
        RECT 2030.065 15.015 2030.355 15.060 ;
        RECT 2052.590 15.000 2052.910 15.060 ;
      LAYER via ;
        RECT 1358.480 17.380 1358.740 17.640 ;
        RECT 2052.620 15.000 2052.880 15.260 ;
      LAYER met2 ;
        RECT 1358.480 17.350 1358.740 17.670 ;
        RECT 1358.540 2.400 1358.680 17.350 ;
        RECT 2052.680 15.290 2052.820 54.000 ;
        RECT 2052.620 14.970 2052.880 15.290 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2098.665 14.025 2098.835 17.255 ;
      LAYER mcon ;
        RECT 2098.665 17.085 2098.835 17.255 ;
      LAYER met1 ;
        RECT 2098.605 17.240 2098.895 17.285 ;
        RECT 1387.980 17.100 2098.895 17.240 ;
        RECT 1376.390 16.900 1376.710 16.960 ;
        RECT 1387.980 16.900 1388.120 17.100 ;
        RECT 2098.605 17.055 2098.895 17.100 ;
        RECT 1376.390 16.760 1388.120 16.900 ;
        RECT 1376.390 16.700 1376.710 16.760 ;
        RECT 2098.605 14.180 2098.895 14.225 ;
        RECT 2125.270 14.180 2125.590 14.240 ;
        RECT 2098.605 14.040 2125.590 14.180 ;
        RECT 2098.605 13.995 2098.895 14.040 ;
        RECT 2125.270 13.980 2125.590 14.040 ;
      LAYER via ;
        RECT 1376.420 16.700 1376.680 16.960 ;
        RECT 2125.300 13.980 2125.560 14.240 ;
      LAYER met2 ;
        RECT 1376.420 16.670 1376.680 16.990 ;
        RECT 1376.480 2.400 1376.620 16.670 ;
        RECT 2125.360 14.270 2125.500 54.000 ;
        RECT 2125.300 13.950 2125.560 14.270 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2146.060 48.690 2146.200 54.000 ;
        RECT 2145.600 48.550 2146.200 48.690 ;
        RECT 2145.600 16.845 2145.740 48.550 ;
        RECT 1394.350 16.475 1394.630 16.845 ;
        RECT 2145.530 16.475 2145.810 16.845 ;
        RECT 1394.420 2.400 1394.560 16.475 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
      LAYER via2 ;
        RECT 1394.350 16.520 1394.630 16.800 ;
        RECT 2145.530 16.520 2145.810 16.800 ;
      LAYER met3 ;
        RECT 1394.325 16.810 1394.655 16.825 ;
        RECT 2145.505 16.810 2145.835 16.825 ;
        RECT 1394.325 16.510 2145.835 16.810 ;
        RECT 1394.325 16.495 1394.655 16.510 ;
        RECT 2145.505 16.495 2145.835 16.510 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1412.270 16.560 1412.590 16.620 ;
        RECT 1824.890 16.560 1825.210 16.620 ;
        RECT 1412.270 16.420 1825.210 16.560 ;
        RECT 1412.270 16.360 1412.590 16.420 ;
        RECT 1824.890 16.360 1825.210 16.420 ;
      LAYER via ;
        RECT 1412.300 16.360 1412.560 16.620 ;
        RECT 1824.920 16.360 1825.180 16.620 ;
      LAYER met2 ;
        RECT 1824.980 16.650 1825.120 54.000 ;
        RECT 1412.300 16.330 1412.560 16.650 ;
        RECT 1824.920 16.330 1825.180 16.650 ;
        RECT 1412.360 2.400 1412.500 16.330 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2152.500 17.525 2152.640 54.000 ;
        RECT 1429.770 17.155 1430.050 17.525 ;
        RECT 2152.430 17.155 2152.710 17.525 ;
        RECT 1429.840 2.400 1429.980 17.155 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
      LAYER via2 ;
        RECT 1429.770 17.200 1430.050 17.480 ;
        RECT 2152.430 17.200 2152.710 17.480 ;
      LAYER met3 ;
        RECT 1429.745 17.490 1430.075 17.505 ;
        RECT 2152.405 17.490 2152.735 17.505 ;
        RECT 1429.745 17.190 2152.735 17.490 ;
        RECT 1429.745 17.175 1430.075 17.190 ;
        RECT 2152.405 17.175 2152.735 17.190 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.610 51.920 1448.930 51.980 ;
        RECT 1511.170 51.920 1511.490 51.980 ;
        RECT 1448.610 51.780 1511.490 51.920 ;
        RECT 1448.610 51.720 1448.930 51.780 ;
        RECT 1511.170 51.720 1511.490 51.780 ;
      LAYER via ;
        RECT 1448.640 51.720 1448.900 51.980 ;
        RECT 1511.200 51.720 1511.460 51.980 ;
      LAYER met2 ;
        RECT 1511.260 52.010 1511.400 54.000 ;
        RECT 1448.640 51.690 1448.900 52.010 ;
        RECT 1511.200 51.690 1511.460 52.010 ;
        RECT 1448.700 16.730 1448.840 51.690 ;
        RECT 1447.780 16.590 1448.840 16.730 ;
        RECT 1447.780 2.400 1447.920 16.590 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2158.480 18.205 2158.620 54.000 ;
        RECT 1465.650 17.835 1465.930 18.205 ;
        RECT 2158.410 17.835 2158.690 18.205 ;
        RECT 1465.720 2.400 1465.860 17.835 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
      LAYER via2 ;
        RECT 1465.650 17.880 1465.930 18.160 ;
        RECT 2158.410 17.880 2158.690 18.160 ;
      LAYER met3 ;
        RECT 1465.625 18.170 1465.955 18.185 ;
        RECT 2158.385 18.170 2158.715 18.185 ;
        RECT 1465.625 17.870 2158.715 18.170 ;
        RECT 1465.625 17.855 1465.955 17.870 ;
        RECT 2158.385 17.855 2158.715 17.870 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 53.280 1490.330 53.340 ;
        RECT 1524.970 53.280 1525.290 53.340 ;
        RECT 1490.010 53.140 1525.290 53.280 ;
        RECT 1490.010 53.080 1490.330 53.140 ;
        RECT 1524.970 53.080 1525.290 53.140 ;
        RECT 1483.570 17.920 1483.890 17.980 ;
        RECT 1490.010 17.920 1490.330 17.980 ;
        RECT 1483.570 17.780 1490.330 17.920 ;
        RECT 1483.570 17.720 1483.890 17.780 ;
        RECT 1490.010 17.720 1490.330 17.780 ;
      LAYER via ;
        RECT 1490.040 53.080 1490.300 53.340 ;
        RECT 1525.000 53.080 1525.260 53.340 ;
        RECT 1483.600 17.720 1483.860 17.980 ;
        RECT 1490.040 17.720 1490.300 17.980 ;
      LAYER met2 ;
        RECT 1525.060 53.370 1525.200 54.000 ;
        RECT 1490.040 53.050 1490.300 53.370 ;
        RECT 1525.000 53.050 1525.260 53.370 ;
        RECT 1490.100 18.010 1490.240 53.050 ;
        RECT 1483.600 17.690 1483.860 18.010 ;
        RECT 1490.040 17.690 1490.300 18.010 ;
        RECT 1483.660 2.400 1483.800 17.690 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1518.145 16.745 1518.315 17.935 ;
      LAYER mcon ;
        RECT 1518.145 17.765 1518.315 17.935 ;
      LAYER met1 ;
        RECT 2169.890 18.260 2170.210 18.320 ;
        RECT 2154.340 18.120 2170.210 18.260 ;
        RECT 1518.085 17.920 1518.375 17.965 ;
        RECT 2154.340 17.920 2154.480 18.120 ;
        RECT 2169.890 18.060 2170.210 18.120 ;
        RECT 1518.085 17.780 2154.480 17.920 ;
        RECT 1518.085 17.735 1518.375 17.780 ;
        RECT 1501.510 16.900 1501.830 16.960 ;
        RECT 1518.085 16.900 1518.375 16.945 ;
        RECT 1501.510 16.760 1518.375 16.900 ;
        RECT 1501.510 16.700 1501.830 16.760 ;
        RECT 1518.085 16.715 1518.375 16.760 ;
      LAYER via ;
        RECT 2169.920 18.060 2170.180 18.320 ;
        RECT 1501.540 16.700 1501.800 16.960 ;
      LAYER met2 ;
        RECT 2169.980 18.350 2170.120 54.000 ;
        RECT 2169.920 18.030 2170.180 18.350 ;
        RECT 1501.540 16.670 1501.800 16.990 ;
        RECT 1501.600 2.400 1501.740 16.670 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1928.850 27.780 1929.170 27.840 ;
        RECT 2354.350 27.780 2354.670 27.840 ;
        RECT 1928.850 27.640 2354.670 27.780 ;
        RECT 1928.850 27.580 1929.170 27.640 ;
        RECT 2354.350 27.580 2354.670 27.640 ;
        RECT 1518.990 15.540 1519.310 15.600 ;
        RECT 1928.850 15.540 1929.170 15.600 ;
        RECT 1518.990 15.400 1929.170 15.540 ;
        RECT 1518.990 15.340 1519.310 15.400 ;
        RECT 1928.850 15.340 1929.170 15.400 ;
      LAYER via ;
        RECT 1928.880 27.580 1929.140 27.840 ;
        RECT 2354.380 27.580 2354.640 27.840 ;
        RECT 1519.020 15.340 1519.280 15.600 ;
        RECT 1928.880 15.340 1929.140 15.600 ;
      LAYER met2 ;
        RECT 2355.360 51.410 2355.500 54.000 ;
        RECT 2354.440 51.270 2355.500 51.410 ;
        RECT 2354.440 27.870 2354.580 51.270 ;
        RECT 1928.880 27.550 1929.140 27.870 ;
        RECT 2354.380 27.550 2354.640 27.870 ;
        RECT 1928.940 15.630 1929.080 27.550 ;
        RECT 1519.020 15.310 1519.280 15.630 ;
        RECT 1928.880 15.310 1929.140 15.630 ;
        RECT 1519.080 2.400 1519.220 15.310 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 716.290 37.980 716.610 38.040 ;
        RECT 720.890 37.980 721.210 38.040 ;
        RECT 716.290 37.840 721.210 37.980 ;
        RECT 716.290 37.780 716.610 37.840 ;
        RECT 720.890 37.780 721.210 37.840 ;
      LAYER via ;
        RECT 716.320 37.780 716.580 38.040 ;
        RECT 720.920 37.780 721.180 38.040 ;
      LAYER met2 ;
        RECT 720.980 38.070 721.120 54.000 ;
        RECT 716.320 37.750 716.580 38.070 ;
        RECT 720.920 37.750 721.180 38.070 ;
        RECT 716.380 2.400 716.520 37.750 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2153.865 18.105 2154.955 18.275 ;
        RECT 2154.785 17.765 2154.955 18.105 ;
        RECT 2163.065 17.595 2163.235 17.935 ;
        RECT 2163.065 17.425 2164.615 17.595 ;
      LAYER mcon ;
        RECT 2163.065 17.765 2163.235 17.935 ;
        RECT 2164.445 17.425 2164.615 17.595 ;
      LAYER met1 ;
        RECT 1536.930 18.260 1537.250 18.320 ;
        RECT 2153.805 18.260 2154.095 18.305 ;
        RECT 1536.930 18.120 2154.095 18.260 ;
        RECT 1536.930 18.060 1537.250 18.120 ;
        RECT 2153.805 18.075 2154.095 18.120 ;
        RECT 2154.725 17.920 2155.015 17.965 ;
        RECT 2163.005 17.920 2163.295 17.965 ;
        RECT 2154.725 17.780 2163.295 17.920 ;
        RECT 2154.725 17.735 2155.015 17.780 ;
        RECT 2163.005 17.735 2163.295 17.780 ;
        RECT 2164.385 17.580 2164.675 17.625 ;
        RECT 2167.130 17.580 2167.450 17.640 ;
        RECT 2164.385 17.440 2167.450 17.580 ;
        RECT 2164.385 17.395 2164.675 17.440 ;
        RECT 2167.130 17.380 2167.450 17.440 ;
      LAYER via ;
        RECT 1536.960 18.060 1537.220 18.320 ;
        RECT 2167.160 17.380 2167.420 17.640 ;
      LAYER met2 ;
        RECT 1536.960 18.030 1537.220 18.350 ;
        RECT 1537.020 2.400 1537.160 18.030 ;
        RECT 2167.220 17.670 2167.360 54.000 ;
        RECT 2167.160 17.350 2167.420 17.670 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1554.870 16.900 1555.190 16.960 ;
        RECT 1559.010 16.900 1559.330 16.960 ;
        RECT 1554.870 16.760 1559.330 16.900 ;
        RECT 1554.870 16.700 1555.190 16.760 ;
        RECT 1559.010 16.700 1559.330 16.760 ;
      LAYER via ;
        RECT 1554.900 16.700 1555.160 16.960 ;
        RECT 1559.040 16.700 1559.300 16.960 ;
      LAYER met2 ;
        RECT 1559.100 16.990 1559.240 54.000 ;
        RECT 1554.900 16.670 1555.160 16.990 ;
        RECT 1559.040 16.670 1559.300 16.990 ;
        RECT 1554.960 2.400 1555.100 16.670 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.350 18.940 1572.670 19.000 ;
        RECT 2176.790 18.940 2177.110 19.000 ;
        RECT 1572.350 18.800 2177.110 18.940 ;
        RECT 1572.350 18.740 1572.670 18.800 ;
        RECT 2176.790 18.740 2177.110 18.800 ;
      LAYER via ;
        RECT 1572.380 18.740 1572.640 19.000 ;
        RECT 2176.820 18.740 2177.080 19.000 ;
      LAYER met2 ;
        RECT 2176.880 19.030 2177.020 54.000 ;
        RECT 1572.380 18.710 1572.640 19.030 ;
        RECT 2176.820 18.710 2177.080 19.030 ;
        RECT 1572.440 9.930 1572.580 18.710 ;
        RECT 1572.440 9.790 1573.040 9.930 ;
        RECT 1572.900 2.400 1573.040 9.790 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1590.290 16.900 1590.610 16.960 ;
        RECT 1593.510 16.900 1593.830 16.960 ;
        RECT 1590.290 16.760 1593.830 16.900 ;
        RECT 1590.290 16.700 1590.610 16.760 ;
        RECT 1593.510 16.700 1593.830 16.760 ;
      LAYER via ;
        RECT 1590.320 16.700 1590.580 16.960 ;
        RECT 1593.540 16.700 1593.800 16.960 ;
      LAYER met2 ;
        RECT 1593.600 16.990 1593.740 54.000 ;
        RECT 1590.320 16.670 1590.580 16.990 ;
        RECT 1593.540 16.670 1593.800 16.990 ;
        RECT 1590.380 2.400 1590.520 16.670 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2259.665 45.985 2259.835 48.195 ;
      LAYER mcon ;
        RECT 2259.665 48.025 2259.835 48.195 ;
      LAYER met1 ;
        RECT 2259.605 48.180 2259.895 48.225 ;
        RECT 2385.170 48.180 2385.490 48.240 ;
        RECT 2259.605 48.040 2385.490 48.180 ;
        RECT 2259.605 47.995 2259.895 48.040 ;
        RECT 2385.170 47.980 2385.490 48.040 ;
        RECT 2226.470 46.140 2226.790 46.200 ;
        RECT 2259.605 46.140 2259.895 46.185 ;
        RECT 2226.470 46.000 2259.895 46.140 ;
        RECT 2226.470 45.940 2226.790 46.000 ;
        RECT 2259.605 45.955 2259.895 46.000 ;
        RECT 1608.230 18.600 1608.550 18.660 ;
        RECT 2226.470 18.600 2226.790 18.660 ;
        RECT 1608.230 18.460 2226.790 18.600 ;
        RECT 1608.230 18.400 1608.550 18.460 ;
        RECT 2226.470 18.400 2226.790 18.460 ;
      LAYER via ;
        RECT 2385.200 47.980 2385.460 48.240 ;
        RECT 2226.500 45.940 2226.760 46.200 ;
        RECT 1608.260 18.400 1608.520 18.660 ;
        RECT 2226.500 18.400 2226.760 18.660 ;
      LAYER met2 ;
        RECT 2385.260 48.270 2385.400 54.000 ;
        RECT 2385.200 47.950 2385.460 48.270 ;
        RECT 2226.500 45.910 2226.760 46.230 ;
        RECT 2226.560 18.690 2226.700 45.910 ;
        RECT 1608.260 18.370 1608.520 18.690 ;
        RECT 2226.500 18.370 2226.760 18.690 ;
        RECT 1608.320 2.400 1608.460 18.370 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1628.100 17.410 1628.240 54.000 ;
        RECT 1626.260 17.270 1628.240 17.410 ;
        RECT 1626.260 2.400 1626.400 17.270 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1644.110 19.620 1644.430 19.680 ;
        RECT 2180.470 19.620 2180.790 19.680 ;
        RECT 1644.110 19.480 2180.790 19.620 ;
        RECT 1644.110 19.420 1644.430 19.480 ;
        RECT 2180.470 19.420 2180.790 19.480 ;
      LAYER via ;
        RECT 1644.140 19.420 1644.400 19.680 ;
        RECT 2180.500 19.420 2180.760 19.680 ;
      LAYER met2 ;
        RECT 2180.560 19.710 2180.700 54.000 ;
        RECT 1644.140 19.390 1644.400 19.710 ;
        RECT 2180.500 19.390 2180.760 19.710 ;
        RECT 1644.200 2.400 1644.340 19.390 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1662.600 17.410 1662.740 54.000 ;
        RECT 1662.140 17.270 1662.740 17.410 ;
        RECT 1662.140 2.400 1662.280 17.270 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2231.070 46.480 2231.390 46.540 ;
        RECT 2408.170 46.480 2408.490 46.540 ;
        RECT 2231.070 46.340 2408.490 46.480 ;
        RECT 2231.070 46.280 2231.390 46.340 ;
        RECT 2408.170 46.280 2408.490 46.340 ;
        RECT 1679.530 19.280 1679.850 19.340 ;
        RECT 2231.070 19.280 2231.390 19.340 ;
        RECT 1679.530 19.140 2231.390 19.280 ;
        RECT 1679.530 19.080 1679.850 19.140 ;
        RECT 2231.070 19.080 2231.390 19.140 ;
      LAYER via ;
        RECT 2231.100 46.280 2231.360 46.540 ;
        RECT 2408.200 46.280 2408.460 46.540 ;
        RECT 1679.560 19.080 1679.820 19.340 ;
        RECT 2231.100 19.080 2231.360 19.340 ;
      LAYER met2 ;
        RECT 2408.260 46.570 2408.400 54.000 ;
        RECT 2231.100 46.250 2231.360 46.570 ;
        RECT 2408.200 46.250 2408.460 46.570 ;
        RECT 2231.160 19.370 2231.300 46.250 ;
        RECT 1679.560 19.050 1679.820 19.370 ;
        RECT 2231.100 19.050 2231.360 19.370 ;
        RECT 1679.620 2.400 1679.760 19.050 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.470 16.900 1697.790 16.960 ;
        RECT 1703.910 16.900 1704.230 16.960 ;
        RECT 1697.470 16.760 1704.230 16.900 ;
        RECT 1697.470 16.700 1697.790 16.760 ;
        RECT 1703.910 16.700 1704.230 16.760 ;
      LAYER via ;
        RECT 1697.500 16.700 1697.760 16.960 ;
        RECT 1703.940 16.700 1704.200 16.960 ;
      LAYER met2 ;
        RECT 1704.000 16.990 1704.140 54.000 ;
        RECT 1697.500 16.670 1697.760 16.990 ;
        RECT 1703.940 16.670 1704.200 16.990 ;
        RECT 1697.560 2.400 1697.700 16.670 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 734.230 52.260 734.550 52.320 ;
        RECT 1566.370 52.260 1566.690 52.320 ;
        RECT 734.230 52.120 1566.690 52.260 ;
        RECT 734.230 52.060 734.550 52.120 ;
        RECT 1566.370 52.060 1566.690 52.120 ;
      LAYER via ;
        RECT 734.260 52.060 734.520 52.320 ;
        RECT 1566.400 52.060 1566.660 52.320 ;
      LAYER met2 ;
        RECT 1566.460 52.350 1566.600 54.000 ;
        RECT 734.260 52.030 734.520 52.350 ;
        RECT 1566.400 52.030 1566.660 52.350 ;
        RECT 734.320 2.400 734.460 52.030 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2255.910 47.500 2256.230 47.560 ;
        RECT 2419.670 47.500 2419.990 47.560 ;
        RECT 2255.910 47.360 2419.990 47.500 ;
        RECT 2255.910 47.300 2256.230 47.360 ;
        RECT 2419.670 47.300 2419.990 47.360 ;
        RECT 1715.410 19.960 1715.730 20.020 ;
        RECT 2255.910 19.960 2256.230 20.020 ;
        RECT 1715.410 19.820 2256.230 19.960 ;
        RECT 1715.410 19.760 1715.730 19.820 ;
        RECT 2255.910 19.760 2256.230 19.820 ;
      LAYER via ;
        RECT 2255.940 47.300 2256.200 47.560 ;
        RECT 2419.700 47.300 2419.960 47.560 ;
        RECT 1715.440 19.760 1715.700 20.020 ;
        RECT 2255.940 19.760 2256.200 20.020 ;
      LAYER met2 ;
        RECT 2419.760 47.590 2419.900 54.000 ;
        RECT 2255.940 47.270 2256.200 47.590 ;
        RECT 2419.700 47.270 2419.960 47.590 ;
        RECT 2256.000 20.050 2256.140 47.270 ;
        RECT 1715.440 19.730 1715.700 20.050 ;
        RECT 2255.940 19.730 2256.200 20.050 ;
        RECT 1715.500 2.400 1715.640 19.730 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2098.205 14.025 2098.375 15.215 ;
        RECT 2107.405 15.045 2107.575 17.595 ;
        RECT 2113.385 17.425 2118.615 17.595 ;
      LAYER mcon ;
        RECT 2107.405 17.425 2107.575 17.595 ;
        RECT 2118.445 17.425 2118.615 17.595 ;
        RECT 2098.205 15.045 2098.375 15.215 ;
      LAYER met1 ;
        RECT 2107.345 17.580 2107.635 17.625 ;
        RECT 2113.325 17.580 2113.615 17.625 ;
        RECT 2107.345 17.440 2113.615 17.580 ;
        RECT 2107.345 17.395 2107.635 17.440 ;
        RECT 2113.325 17.395 2113.615 17.440 ;
        RECT 2118.385 17.580 2118.675 17.625 ;
        RECT 2132.170 17.580 2132.490 17.640 ;
        RECT 2118.385 17.440 2132.490 17.580 ;
        RECT 2118.385 17.395 2118.675 17.440 ;
        RECT 2132.170 17.380 2132.490 17.440 ;
        RECT 2098.145 15.200 2098.435 15.245 ;
        RECT 2107.345 15.200 2107.635 15.245 ;
        RECT 2098.145 15.060 2107.635 15.200 ;
        RECT 2098.145 15.015 2098.435 15.060 ;
        RECT 2107.345 15.015 2107.635 15.060 ;
        RECT 1733.350 14.180 1733.670 14.240 ;
        RECT 2098.145 14.180 2098.435 14.225 ;
        RECT 1733.350 14.040 2098.435 14.180 ;
        RECT 1733.350 13.980 1733.670 14.040 ;
        RECT 2098.145 13.995 2098.435 14.040 ;
      LAYER via ;
        RECT 2132.200 17.380 2132.460 17.640 ;
        RECT 1733.380 13.980 1733.640 14.240 ;
      LAYER met2 ;
        RECT 2132.260 17.670 2132.400 54.000 ;
        RECT 2132.200 17.350 2132.460 17.670 ;
        RECT 1733.380 13.950 1733.640 14.270 ;
        RECT 1733.440 2.400 1733.580 13.950 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2208.145 18.785 2208.315 20.315 ;
      LAYER mcon ;
        RECT 2208.145 20.145 2208.315 20.315 ;
      LAYER met1 ;
        RECT 2263.270 47.840 2263.590 47.900 ;
        RECT 2431.170 47.840 2431.490 47.900 ;
        RECT 2263.270 47.700 2431.490 47.840 ;
        RECT 2263.270 47.640 2263.590 47.700 ;
        RECT 2431.170 47.640 2431.490 47.700 ;
        RECT 1751.290 20.300 1751.610 20.360 ;
        RECT 2208.085 20.300 2208.375 20.345 ;
        RECT 1751.290 20.160 2208.375 20.300 ;
        RECT 1751.290 20.100 1751.610 20.160 ;
        RECT 2208.085 20.115 2208.375 20.160 ;
        RECT 2208.085 18.940 2208.375 18.985 ;
        RECT 2263.270 18.940 2263.590 19.000 ;
        RECT 2208.085 18.800 2263.590 18.940 ;
        RECT 2208.085 18.755 2208.375 18.800 ;
        RECT 2263.270 18.740 2263.590 18.800 ;
      LAYER via ;
        RECT 2263.300 47.640 2263.560 47.900 ;
        RECT 2431.200 47.640 2431.460 47.900 ;
        RECT 1751.320 20.100 1751.580 20.360 ;
        RECT 2263.300 18.740 2263.560 19.000 ;
      LAYER met2 ;
        RECT 2431.260 47.930 2431.400 54.000 ;
        RECT 2263.300 47.610 2263.560 47.930 ;
        RECT 2431.200 47.610 2431.460 47.930 ;
        RECT 1751.320 20.070 1751.580 20.390 ;
        RECT 1751.380 2.400 1751.520 20.070 ;
        RECT 2263.360 19.030 2263.500 47.610 ;
        RECT 2263.300 18.710 2263.560 19.030 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.770 16.900 1769.090 16.960 ;
        RECT 1772.910 16.900 1773.230 16.960 ;
        RECT 1768.770 16.760 1773.230 16.900 ;
        RECT 1768.770 16.700 1769.090 16.760 ;
        RECT 1772.910 16.700 1773.230 16.760 ;
      LAYER via ;
        RECT 1768.800 16.700 1769.060 16.960 ;
        RECT 1772.940 16.700 1773.200 16.960 ;
      LAYER met2 ;
        RECT 1773.000 16.990 1773.140 54.000 ;
        RECT 1768.800 16.670 1769.060 16.990 ;
        RECT 1772.940 16.670 1773.200 16.990 ;
        RECT 1768.860 2.400 1769.000 16.670 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1801.045 16.065 1801.215 16.915 ;
      LAYER mcon ;
        RECT 1801.045 16.745 1801.215 16.915 ;
      LAYER met1 ;
        RECT 2263.730 46.820 2264.050 46.880 ;
        RECT 2442.670 46.820 2442.990 46.880 ;
        RECT 2263.730 46.680 2442.990 46.820 ;
        RECT 2263.730 46.620 2264.050 46.680 ;
        RECT 2442.670 46.620 2442.990 46.680 ;
        RECT 1800.985 16.900 1801.275 16.945 ;
        RECT 2263.730 16.900 2264.050 16.960 ;
        RECT 1800.985 16.760 2264.050 16.900 ;
        RECT 1800.985 16.715 1801.275 16.760 ;
        RECT 2263.730 16.700 2264.050 16.760 ;
        RECT 1786.710 16.220 1787.030 16.280 ;
        RECT 1800.985 16.220 1801.275 16.265 ;
        RECT 1786.710 16.080 1801.275 16.220 ;
        RECT 1786.710 16.020 1787.030 16.080 ;
        RECT 1800.985 16.035 1801.275 16.080 ;
      LAYER via ;
        RECT 2263.760 46.620 2264.020 46.880 ;
        RECT 2442.700 46.620 2442.960 46.880 ;
        RECT 2263.760 16.700 2264.020 16.960 ;
        RECT 1786.740 16.020 1787.000 16.280 ;
      LAYER met2 ;
        RECT 2442.760 46.910 2442.900 54.000 ;
        RECT 2263.760 46.590 2264.020 46.910 ;
        RECT 2442.700 46.590 2442.960 46.910 ;
        RECT 2263.820 16.990 2263.960 46.590 ;
        RECT 2263.760 16.670 2264.020 16.990 ;
        RECT 1786.740 15.990 1787.000 16.310 ;
        RECT 1786.800 2.400 1786.940 15.990 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1804.650 20.640 1804.970 20.700 ;
        RECT 1807.410 20.640 1807.730 20.700 ;
        RECT 1804.650 20.500 1807.730 20.640 ;
        RECT 1804.650 20.440 1804.970 20.500 ;
        RECT 1807.410 20.440 1807.730 20.500 ;
      LAYER via ;
        RECT 1804.680 20.440 1804.940 20.700 ;
        RECT 1807.440 20.440 1807.700 20.700 ;
      LAYER met2 ;
        RECT 1807.500 20.730 1807.640 54.000 ;
        RECT 1804.680 20.410 1804.940 20.730 ;
        RECT 1807.440 20.410 1807.700 20.730 ;
        RECT 1804.740 2.400 1804.880 20.410 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1822.590 20.640 1822.910 20.700 ;
        RECT 2307.890 20.640 2308.210 20.700 ;
        RECT 1822.590 20.500 2308.210 20.640 ;
        RECT 1822.590 20.440 1822.910 20.500 ;
        RECT 2307.890 20.440 2308.210 20.500 ;
      LAYER via ;
        RECT 1822.620 20.440 1822.880 20.700 ;
        RECT 2307.920 20.440 2308.180 20.700 ;
      LAYER met2 ;
        RECT 2307.980 20.730 2308.120 54.000 ;
        RECT 1822.620 20.410 1822.880 20.730 ;
        RECT 2307.920 20.410 2308.180 20.730 ;
        RECT 1822.680 2.400 1822.820 20.410 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1842.000 3.130 1842.140 54.000 ;
        RECT 1840.160 2.990 1842.140 3.130 ;
        RECT 1840.160 2.400 1840.300 2.990 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2292.710 47.160 2293.030 47.220 ;
        RECT 2465.670 47.160 2465.990 47.220 ;
        RECT 2292.710 47.020 2465.990 47.160 ;
        RECT 2292.710 46.960 2293.030 47.020 ;
        RECT 2465.670 46.960 2465.990 47.020 ;
        RECT 1858.010 15.880 1858.330 15.940 ;
        RECT 2292.710 15.880 2293.030 15.940 ;
        RECT 1858.010 15.740 2293.030 15.880 ;
        RECT 1858.010 15.680 1858.330 15.740 ;
        RECT 2292.710 15.680 2293.030 15.740 ;
      LAYER via ;
        RECT 2292.740 46.960 2293.000 47.220 ;
        RECT 2465.700 46.960 2465.960 47.220 ;
        RECT 1858.040 15.680 1858.300 15.940 ;
        RECT 2292.740 15.680 2293.000 15.940 ;
      LAYER met2 ;
        RECT 2465.760 47.250 2465.900 54.000 ;
        RECT 2292.740 46.930 2293.000 47.250 ;
        RECT 2465.700 46.930 2465.960 47.250 ;
        RECT 2292.800 15.970 2292.940 46.930 ;
        RECT 1858.040 15.650 1858.300 15.970 ;
        RECT 2292.740 15.650 2293.000 15.970 ;
        RECT 1858.100 2.400 1858.240 15.650 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1876.040 2.400 1876.180 54.000 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 753.090 45.120 753.410 45.180 ;
        RECT 870.850 45.120 871.170 45.180 ;
        RECT 753.090 44.980 871.170 45.120 ;
        RECT 753.090 44.920 753.410 44.980 ;
        RECT 870.850 44.920 871.170 44.980 ;
      LAYER via ;
        RECT 753.120 44.920 753.380 45.180 ;
        RECT 870.880 44.920 871.140 45.180 ;
      LAYER met2 ;
        RECT 870.940 45.210 871.080 54.000 ;
        RECT 753.120 44.890 753.380 45.210 ;
        RECT 870.880 44.890 871.140 45.210 ;
        RECT 753.180 14.010 753.320 44.890 ;
        RECT 752.260 13.870 753.320 14.010 ;
        RECT 752.260 2.400 752.400 13.870 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1916.965 15.045 1917.135 16.575 ;
      LAYER mcon ;
        RECT 1916.965 16.405 1917.135 16.575 ;
      LAYER met1 ;
        RECT 2359.410 32.540 2359.730 32.600 ;
        RECT 2478.090 32.540 2478.410 32.600 ;
        RECT 2359.410 32.400 2478.410 32.540 ;
        RECT 2359.410 32.340 2359.730 32.400 ;
        RECT 2478.090 32.340 2478.410 32.400 ;
        RECT 1916.905 16.560 1917.195 16.605 ;
        RECT 2359.410 16.560 2359.730 16.620 ;
        RECT 1916.905 16.420 2359.730 16.560 ;
        RECT 1916.905 16.375 1917.195 16.420 ;
        RECT 2359.410 16.360 2359.730 16.420 ;
        RECT 1893.890 15.200 1894.210 15.260 ;
        RECT 1916.905 15.200 1917.195 15.245 ;
        RECT 1893.890 15.060 1917.195 15.200 ;
        RECT 1893.890 15.000 1894.210 15.060 ;
        RECT 1916.905 15.015 1917.195 15.060 ;
      LAYER via ;
        RECT 2359.440 32.340 2359.700 32.600 ;
        RECT 2478.120 32.340 2478.380 32.600 ;
        RECT 2359.440 16.360 2359.700 16.620 ;
        RECT 1893.920 15.000 1894.180 15.260 ;
      LAYER met2 ;
        RECT 2478.180 32.630 2478.320 54.000 ;
        RECT 2359.440 32.310 2359.700 32.630 ;
        RECT 2478.120 32.310 2478.380 32.630 ;
        RECT 2359.500 16.650 2359.640 32.310 ;
        RECT 2359.440 16.330 2359.700 16.650 ;
        RECT 1893.920 14.970 1894.180 15.290 ;
        RECT 1893.980 2.400 1894.120 14.970 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1916.430 20.980 1916.750 21.040 ;
        RECT 1917.810 20.980 1918.130 21.040 ;
        RECT 1916.430 20.840 1918.130 20.980 ;
        RECT 1916.430 20.780 1916.750 20.840 ;
        RECT 1917.810 20.780 1918.130 20.840 ;
        RECT 1911.830 16.560 1912.150 16.620 ;
        RECT 1916.430 16.560 1916.750 16.620 ;
        RECT 1911.830 16.420 1916.750 16.560 ;
        RECT 1911.830 16.360 1912.150 16.420 ;
        RECT 1916.430 16.360 1916.750 16.420 ;
      LAYER via ;
        RECT 1916.460 20.780 1916.720 21.040 ;
        RECT 1917.840 20.780 1918.100 21.040 ;
        RECT 1911.860 16.360 1912.120 16.620 ;
        RECT 1916.460 16.360 1916.720 16.620 ;
      LAYER met2 ;
        RECT 1917.900 21.070 1918.040 54.000 ;
        RECT 1916.460 20.750 1916.720 21.070 ;
        RECT 1917.840 20.750 1918.100 21.070 ;
        RECT 1916.520 16.650 1916.660 20.750 ;
        RECT 1911.860 16.330 1912.120 16.650 ;
        RECT 1916.460 16.330 1916.720 16.650 ;
        RECT 1911.920 2.400 1912.060 16.330 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1952.845 15.045 1953.015 16.235 ;
      LAYER mcon ;
        RECT 1952.845 16.065 1953.015 16.235 ;
      LAYER met1 ;
        RECT 2380.570 33.220 2380.890 33.280 ;
        RECT 2484.530 33.220 2484.850 33.280 ;
        RECT 2380.570 33.080 2484.850 33.220 ;
        RECT 2380.570 33.020 2380.890 33.080 ;
        RECT 2484.530 33.020 2484.850 33.080 ;
        RECT 1952.785 16.220 1953.075 16.265 ;
        RECT 2380.570 16.220 2380.890 16.280 ;
        RECT 1952.785 16.080 2380.890 16.220 ;
        RECT 1952.785 16.035 1953.075 16.080 ;
        RECT 2380.570 16.020 2380.890 16.080 ;
        RECT 1929.310 15.200 1929.630 15.260 ;
        RECT 1952.785 15.200 1953.075 15.245 ;
        RECT 1929.310 15.060 1953.075 15.200 ;
        RECT 1929.310 15.000 1929.630 15.060 ;
        RECT 1952.785 15.015 1953.075 15.060 ;
      LAYER via ;
        RECT 2380.600 33.020 2380.860 33.280 ;
        RECT 2484.560 33.020 2484.820 33.280 ;
        RECT 2380.600 16.020 2380.860 16.280 ;
        RECT 1929.340 15.000 1929.600 15.260 ;
      LAYER met2 ;
        RECT 2485.540 36.450 2485.680 54.000 ;
        RECT 2484.620 36.310 2485.680 36.450 ;
        RECT 2484.620 33.310 2484.760 36.310 ;
        RECT 2380.600 32.990 2380.860 33.310 ;
        RECT 2484.560 32.990 2484.820 33.310 ;
        RECT 2380.660 16.310 2380.800 32.990 ;
        RECT 2380.600 15.990 2380.860 16.310 ;
        RECT 1929.340 14.970 1929.600 15.290 ;
        RECT 1929.400 2.400 1929.540 14.970 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1947.250 16.220 1947.570 16.280 ;
        RECT 1952.310 16.220 1952.630 16.280 ;
        RECT 1947.250 16.080 1952.630 16.220 ;
        RECT 1947.250 16.020 1947.570 16.080 ;
        RECT 1952.310 16.020 1952.630 16.080 ;
      LAYER via ;
        RECT 1947.280 16.020 1947.540 16.280 ;
        RECT 1952.340 16.020 1952.600 16.280 ;
      LAYER met2 ;
        RECT 1952.400 16.310 1952.540 54.000 ;
        RECT 1947.280 15.990 1947.540 16.310 ;
        RECT 1952.340 15.990 1952.600 16.310 ;
        RECT 1947.340 2.400 1947.480 15.990 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1965.190 14.860 1965.510 14.920 ;
        RECT 2321.230 14.860 2321.550 14.920 ;
        RECT 1965.190 14.720 2321.550 14.860 ;
        RECT 1965.190 14.660 1965.510 14.720 ;
        RECT 2321.230 14.660 2321.550 14.720 ;
      LAYER via ;
        RECT 1965.220 14.660 1965.480 14.920 ;
        RECT 2321.260 14.660 2321.520 14.920 ;
      LAYER met2 ;
        RECT 2321.320 14.950 2321.460 54.000 ;
        RECT 1965.220 14.630 1965.480 14.950 ;
        RECT 2321.260 14.630 2321.520 14.950 ;
        RECT 1965.280 2.400 1965.420 14.630 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1983.130 15.540 1983.450 15.600 ;
        RECT 1986.810 15.540 1987.130 15.600 ;
        RECT 1983.130 15.400 1987.130 15.540 ;
        RECT 1983.130 15.340 1983.450 15.400 ;
        RECT 1986.810 15.340 1987.130 15.400 ;
      LAYER via ;
        RECT 1983.160 15.340 1983.420 15.600 ;
        RECT 1986.840 15.340 1987.100 15.600 ;
      LAYER met2 ;
        RECT 1986.900 15.630 1987.040 54.000 ;
        RECT 1983.160 15.310 1983.420 15.630 ;
        RECT 1986.840 15.310 1987.100 15.630 ;
        RECT 1983.220 2.400 1983.360 15.310 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2018.090 48.520 2018.410 48.580 ;
        RECT 2511.670 48.520 2511.990 48.580 ;
        RECT 2018.090 48.380 2511.990 48.520 ;
        RECT 2018.090 48.320 2018.410 48.380 ;
        RECT 2511.670 48.320 2511.990 48.380 ;
        RECT 2001.070 15.540 2001.390 15.600 ;
        RECT 2018.090 15.540 2018.410 15.600 ;
        RECT 2001.070 15.400 2018.410 15.540 ;
        RECT 2001.070 15.340 2001.390 15.400 ;
        RECT 2018.090 15.340 2018.410 15.400 ;
      LAYER via ;
        RECT 2018.120 48.320 2018.380 48.580 ;
        RECT 2511.700 48.320 2511.960 48.580 ;
        RECT 2001.100 15.340 2001.360 15.600 ;
        RECT 2018.120 15.340 2018.380 15.600 ;
      LAYER met2 ;
        RECT 2511.760 48.610 2511.900 54.000 ;
        RECT 2018.120 48.290 2018.380 48.610 ;
        RECT 2511.700 48.290 2511.960 48.610 ;
        RECT 2018.180 15.630 2018.320 48.290 ;
        RECT 2001.100 15.310 2001.360 15.630 ;
        RECT 2018.120 15.310 2018.380 15.630 ;
        RECT 2001.160 2.400 2001.300 15.310 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2387.930 32.200 2388.250 32.260 ;
        RECT 2512.590 32.200 2512.910 32.260 ;
        RECT 2387.930 32.060 2512.910 32.200 ;
        RECT 2387.930 32.000 2388.250 32.060 ;
        RECT 2512.590 32.000 2512.910 32.060 ;
        RECT 2018.550 15.540 2018.870 15.600 ;
        RECT 2387.930 15.540 2388.250 15.600 ;
        RECT 2018.550 15.400 2388.250 15.540 ;
        RECT 2018.550 15.340 2018.870 15.400 ;
        RECT 2387.930 15.340 2388.250 15.400 ;
      LAYER via ;
        RECT 2387.960 32.000 2388.220 32.260 ;
        RECT 2512.620 32.000 2512.880 32.260 ;
        RECT 2018.580 15.340 2018.840 15.600 ;
        RECT 2387.960 15.340 2388.220 15.600 ;
      LAYER met2 ;
        RECT 2512.680 32.290 2512.820 54.000 ;
        RECT 2387.960 31.970 2388.220 32.290 ;
        RECT 2512.620 31.970 2512.880 32.290 ;
        RECT 2388.020 15.630 2388.160 31.970 ;
        RECT 2018.580 15.310 2018.840 15.630 ;
        RECT 2387.960 15.310 2388.220 15.630 ;
        RECT 2018.640 2.400 2018.780 15.310 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2036.490 17.580 2036.810 17.640 ;
        RECT 2042.010 17.580 2042.330 17.640 ;
        RECT 2036.490 17.440 2042.330 17.580 ;
        RECT 2036.490 17.380 2036.810 17.440 ;
        RECT 2042.010 17.380 2042.330 17.440 ;
      LAYER via ;
        RECT 2036.520 17.380 2036.780 17.640 ;
        RECT 2042.040 17.380 2042.300 17.640 ;
      LAYER met2 ;
        RECT 2042.100 17.670 2042.240 54.000 ;
        RECT 2036.520 17.350 2036.780 17.670 ;
        RECT 2042.040 17.350 2042.300 17.670 ;
        RECT 2036.580 2.400 2036.720 17.350 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2397.590 52.940 2397.910 53.000 ;
        RECT 2528.690 52.940 2529.010 53.000 ;
        RECT 2397.590 52.800 2529.010 52.940 ;
        RECT 2397.590 52.740 2397.910 52.800 ;
        RECT 2528.690 52.740 2529.010 52.800 ;
        RECT 2054.430 14.520 2054.750 14.580 ;
        RECT 2397.590 14.520 2397.910 14.580 ;
        RECT 2054.430 14.380 2397.910 14.520 ;
        RECT 2054.430 14.320 2054.750 14.380 ;
        RECT 2397.590 14.320 2397.910 14.380 ;
      LAYER via ;
        RECT 2397.620 52.740 2397.880 53.000 ;
        RECT 2528.720 52.740 2528.980 53.000 ;
        RECT 2054.460 14.320 2054.720 14.580 ;
        RECT 2397.620 14.320 2397.880 14.580 ;
      LAYER met2 ;
        RECT 2528.780 53.030 2528.920 54.000 ;
        RECT 2397.620 52.710 2397.880 53.030 ;
        RECT 2528.720 52.710 2528.980 53.030 ;
        RECT 2397.680 14.610 2397.820 52.710 ;
        RECT 2054.460 14.290 2054.720 14.610 ;
        RECT 2397.620 14.290 2397.880 14.610 ;
        RECT 2054.520 2.400 2054.660 14.290 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 769.650 44.780 769.970 44.840 ;
        RECT 1024.490 44.780 1024.810 44.840 ;
        RECT 769.650 44.640 1024.810 44.780 ;
        RECT 769.650 44.580 769.970 44.640 ;
        RECT 1024.490 44.580 1024.810 44.640 ;
      LAYER via ;
        RECT 769.680 44.580 769.940 44.840 ;
        RECT 1024.520 44.580 1024.780 44.840 ;
      LAYER met2 ;
        RECT 1024.580 44.870 1024.720 54.000 ;
        RECT 769.680 44.550 769.940 44.870 ;
        RECT 1024.520 44.550 1024.780 44.870 ;
        RECT 769.740 2.400 769.880 44.550 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2090.385 15.045 2090.555 17.595 ;
      LAYER mcon ;
        RECT 2090.385 17.425 2090.555 17.595 ;
      LAYER met1 ;
        RECT 2196.570 17.920 2196.890 17.980 ;
        RECT 2164.000 17.780 2196.890 17.920 ;
        RECT 2090.325 17.580 2090.615 17.625 ;
        RECT 2106.870 17.580 2107.190 17.640 ;
        RECT 2090.325 17.440 2107.190 17.580 ;
        RECT 2090.325 17.395 2090.615 17.440 ;
        RECT 2106.870 17.380 2107.190 17.440 ;
        RECT 2132.630 17.580 2132.950 17.640 ;
        RECT 2164.000 17.580 2164.140 17.780 ;
        RECT 2196.570 17.720 2196.890 17.780 ;
        RECT 2132.630 17.440 2164.140 17.580 ;
        RECT 2132.630 17.380 2132.950 17.440 ;
        RECT 2072.370 15.200 2072.690 15.260 ;
        RECT 2090.325 15.200 2090.615 15.245 ;
        RECT 2072.370 15.060 2090.615 15.200 ;
        RECT 2072.370 15.000 2072.690 15.060 ;
        RECT 2090.325 15.015 2090.615 15.060 ;
      LAYER via ;
        RECT 2106.900 17.380 2107.160 17.640 ;
        RECT 2132.660 17.380 2132.920 17.640 ;
        RECT 2196.600 17.720 2196.860 17.980 ;
        RECT 2072.400 15.000 2072.660 15.260 ;
      LAYER met2 ;
        RECT 2106.890 18.515 2107.170 18.885 ;
        RECT 2132.650 18.515 2132.930 18.885 ;
        RECT 2106.960 17.670 2107.100 18.515 ;
        RECT 2132.720 17.670 2132.860 18.515 ;
        RECT 2196.660 18.010 2196.800 54.000 ;
        RECT 2196.600 17.690 2196.860 18.010 ;
        RECT 2106.900 17.350 2107.160 17.670 ;
        RECT 2132.660 17.350 2132.920 17.670 ;
        RECT 2072.400 14.970 2072.660 15.290 ;
        RECT 2072.460 2.400 2072.600 14.970 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
      LAYER via2 ;
        RECT 2106.890 18.560 2107.170 18.840 ;
        RECT 2132.650 18.560 2132.930 18.840 ;
      LAYER met3 ;
        RECT 2106.865 18.850 2107.195 18.865 ;
        RECT 2132.625 18.850 2132.955 18.865 ;
        RECT 2106.865 18.550 2132.955 18.850 ;
        RECT 2106.865 18.535 2107.195 18.550 ;
        RECT 2132.625 18.535 2132.955 18.550 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 20.980 2090.630 21.040 ;
        RECT 2104.110 20.980 2104.430 21.040 ;
        RECT 2090.310 20.840 2104.430 20.980 ;
        RECT 2090.310 20.780 2090.630 20.840 ;
        RECT 2104.110 20.780 2104.430 20.840 ;
      LAYER via ;
        RECT 2090.340 20.780 2090.600 21.040 ;
        RECT 2104.140 20.780 2104.400 21.040 ;
      LAYER met2 ;
        RECT 2104.200 21.070 2104.340 54.000 ;
        RECT 2090.340 20.750 2090.600 21.070 ;
        RECT 2104.140 20.750 2104.400 21.070 ;
        RECT 2090.400 16.730 2090.540 20.750 ;
        RECT 2089.940 16.590 2090.540 16.730 ;
        RECT 2089.940 2.400 2090.080 16.590 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2403.570 32.880 2403.890 32.940 ;
        RECT 2546.630 32.880 2546.950 32.940 ;
        RECT 2403.570 32.740 2546.950 32.880 ;
        RECT 2403.570 32.680 2403.890 32.740 ;
        RECT 2546.630 32.680 2546.950 32.740 ;
        RECT 2107.790 15.200 2108.110 15.260 ;
        RECT 2403.570 15.200 2403.890 15.260 ;
        RECT 2107.790 15.060 2403.890 15.200 ;
        RECT 2107.790 15.000 2108.110 15.060 ;
        RECT 2403.570 15.000 2403.890 15.060 ;
      LAYER via ;
        RECT 2403.600 32.680 2403.860 32.940 ;
        RECT 2546.660 32.680 2546.920 32.940 ;
        RECT 2107.820 15.000 2108.080 15.260 ;
        RECT 2403.600 15.000 2403.860 15.260 ;
      LAYER met2 ;
        RECT 2546.720 32.970 2546.860 54.000 ;
        RECT 2403.600 32.650 2403.860 32.970 ;
        RECT 2546.660 32.650 2546.920 32.970 ;
        RECT 2403.660 15.290 2403.800 32.650 ;
        RECT 2107.820 14.970 2108.080 15.290 ;
        RECT 2403.600 14.970 2403.860 15.290 ;
        RECT 2107.880 2.400 2108.020 14.970 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2425.190 53.280 2425.510 53.340 ;
        RECT 2551.690 53.280 2552.010 53.340 ;
        RECT 2425.190 53.140 2552.010 53.280 ;
        RECT 2425.190 53.080 2425.510 53.140 ;
        RECT 2551.690 53.080 2552.010 53.140 ;
        RECT 2125.730 14.180 2126.050 14.240 ;
        RECT 2425.190 14.180 2425.510 14.240 ;
        RECT 2125.730 14.040 2425.510 14.180 ;
        RECT 2125.730 13.980 2126.050 14.040 ;
        RECT 2425.190 13.980 2425.510 14.040 ;
      LAYER via ;
        RECT 2425.220 53.080 2425.480 53.340 ;
        RECT 2551.720 53.080 2551.980 53.340 ;
        RECT 2125.760 13.980 2126.020 14.240 ;
        RECT 2425.220 13.980 2425.480 14.240 ;
      LAYER met2 ;
        RECT 2551.780 53.370 2551.920 54.000 ;
        RECT 2425.220 53.050 2425.480 53.370 ;
        RECT 2551.720 53.050 2551.980 53.370 ;
        RECT 2425.280 14.270 2425.420 53.050 ;
        RECT 2125.760 13.950 2126.020 14.270 ;
        RECT 2425.220 13.950 2425.480 14.270 ;
        RECT 2125.820 2.400 2125.960 13.950 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2144.680 48.690 2144.820 54.000 ;
        RECT 2144.680 48.550 2145.280 48.690 ;
        RECT 2145.140 16.050 2145.280 48.550 ;
        RECT 2145.140 15.910 2145.740 16.050 ;
        RECT 2145.600 3.130 2145.740 15.910 ;
        RECT 2143.760 2.990 2145.740 3.130 ;
        RECT 2143.760 2.400 2143.900 2.990 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2366.845 17.085 2367.935 17.255 ;
      LAYER mcon ;
        RECT 2367.765 17.085 2367.935 17.255 ;
      LAYER met1 ;
        RECT 2161.610 17.240 2161.930 17.300 ;
        RECT 2366.785 17.240 2367.075 17.285 ;
        RECT 2161.610 17.100 2367.075 17.240 ;
        RECT 2161.610 17.040 2161.930 17.100 ;
        RECT 2366.785 17.055 2367.075 17.100 ;
        RECT 2367.705 17.240 2367.995 17.285 ;
        RECT 2549.390 17.240 2549.710 17.300 ;
        RECT 2367.705 17.100 2549.710 17.240 ;
        RECT 2367.705 17.055 2367.995 17.100 ;
        RECT 2549.390 17.040 2549.710 17.100 ;
      LAYER via ;
        RECT 2161.640 17.040 2161.900 17.300 ;
        RECT 2549.420 17.040 2549.680 17.300 ;
      LAYER met2 ;
        RECT 2549.480 17.330 2549.620 54.000 ;
        RECT 2161.640 17.010 2161.900 17.330 ;
        RECT 2549.420 17.010 2549.680 17.330 ;
        RECT 2161.700 2.400 2161.840 17.010 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2415.145 17.425 2416.695 17.595 ;
        RECT 2505.765 16.745 2505.935 17.595 ;
      LAYER mcon ;
        RECT 2416.525 17.425 2416.695 17.595 ;
        RECT 2505.765 17.425 2505.935 17.595 ;
      LAYER met1 ;
        RECT 2179.090 17.580 2179.410 17.640 ;
        RECT 2415.085 17.580 2415.375 17.625 ;
        RECT 2179.090 17.440 2415.375 17.580 ;
        RECT 2179.090 17.380 2179.410 17.440 ;
        RECT 2415.085 17.395 2415.375 17.440 ;
        RECT 2416.465 17.580 2416.755 17.625 ;
        RECT 2505.705 17.580 2505.995 17.625 ;
        RECT 2416.465 17.440 2505.995 17.580 ;
        RECT 2416.465 17.395 2416.755 17.440 ;
        RECT 2505.705 17.395 2505.995 17.440 ;
        RECT 2505.705 16.900 2505.995 16.945 ;
        RECT 2556.290 16.900 2556.610 16.960 ;
        RECT 2505.705 16.760 2556.610 16.900 ;
        RECT 2505.705 16.715 2505.995 16.760 ;
        RECT 2556.290 16.700 2556.610 16.760 ;
      LAYER via ;
        RECT 2179.120 17.380 2179.380 17.640 ;
        RECT 2556.320 16.700 2556.580 16.960 ;
      LAYER met2 ;
        RECT 2179.120 17.350 2179.380 17.670 ;
        RECT 2179.180 2.400 2179.320 17.350 ;
        RECT 2556.380 16.990 2556.520 54.000 ;
        RECT 2556.320 16.670 2556.580 16.990 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2197.030 19.620 2197.350 19.680 ;
        RECT 2217.730 19.620 2218.050 19.680 ;
        RECT 2197.030 19.480 2218.050 19.620 ;
        RECT 2197.030 19.420 2197.350 19.480 ;
        RECT 2217.730 19.420 2218.050 19.480 ;
      LAYER via ;
        RECT 2197.060 19.420 2197.320 19.680 ;
        RECT 2217.760 19.420 2218.020 19.680 ;
      LAYER met2 ;
        RECT 2219.200 53.450 2219.340 54.000 ;
        RECT 2217.820 53.310 2219.340 53.450 ;
        RECT 2217.820 19.710 2217.960 53.310 ;
        RECT 2197.060 19.390 2197.320 19.710 ;
        RECT 2217.760 19.390 2218.020 19.710 ;
        RECT 2197.120 2.400 2197.260 19.390 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2319.005 17.765 2319.635 17.935 ;
        RECT 2416.065 17.765 2417.155 17.935 ;
      LAYER mcon ;
        RECT 2319.465 17.765 2319.635 17.935 ;
        RECT 2416.985 17.765 2417.155 17.935 ;
      LAYER met1 ;
        RECT 2214.970 18.260 2215.290 18.320 ;
        RECT 2214.970 18.120 2259.820 18.260 ;
        RECT 2214.970 18.060 2215.290 18.120 ;
        RECT 2259.680 17.920 2259.820 18.120 ;
        RECT 2318.945 17.920 2319.235 17.965 ;
        RECT 2259.680 17.780 2319.235 17.920 ;
        RECT 2318.945 17.735 2319.235 17.780 ;
        RECT 2319.405 17.920 2319.695 17.965 ;
        RECT 2366.770 17.920 2367.090 17.980 ;
        RECT 2319.405 17.780 2367.090 17.920 ;
        RECT 2319.405 17.735 2319.695 17.780 ;
        RECT 2366.770 17.720 2367.090 17.780 ;
        RECT 2367.230 17.920 2367.550 17.980 ;
        RECT 2416.005 17.920 2416.295 17.965 ;
        RECT 2367.230 17.780 2416.295 17.920 ;
        RECT 2367.230 17.720 2367.550 17.780 ;
        RECT 2416.005 17.735 2416.295 17.780 ;
        RECT 2416.925 17.920 2417.215 17.965 ;
        RECT 2581.130 17.920 2581.450 17.980 ;
        RECT 2416.925 17.780 2581.450 17.920 ;
        RECT 2416.925 17.735 2417.215 17.780 ;
        RECT 2581.130 17.720 2581.450 17.780 ;
      LAYER via ;
        RECT 2215.000 18.060 2215.260 18.320 ;
        RECT 2366.800 17.720 2367.060 17.980 ;
        RECT 2367.260 17.720 2367.520 17.980 ;
        RECT 2581.160 17.720 2581.420 17.980 ;
      LAYER met2 ;
        RECT 2215.000 18.030 2215.260 18.350 ;
        RECT 2215.060 2.400 2215.200 18.030 ;
        RECT 2581.220 18.010 2581.360 54.000 ;
        RECT 2366.800 17.690 2367.060 18.010 ;
        RECT 2367.260 17.690 2367.520 18.010 ;
        RECT 2581.160 17.690 2581.420 18.010 ;
        RECT 2366.860 17.410 2367.000 17.690 ;
        RECT 2367.320 17.410 2367.460 17.690 ;
        RECT 2366.860 17.270 2367.460 17.410 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2232.910 17.920 2233.230 17.980 ;
        RECT 2238.890 17.920 2239.210 17.980 ;
        RECT 2232.910 17.780 2239.210 17.920 ;
        RECT 2232.910 17.720 2233.230 17.780 ;
        RECT 2238.890 17.720 2239.210 17.780 ;
      LAYER via ;
        RECT 2232.940 17.720 2233.200 17.980 ;
        RECT 2238.920 17.720 2239.180 17.980 ;
      LAYER met2 ;
        RECT 2238.980 18.010 2239.120 54.000 ;
        RECT 2232.940 17.690 2233.200 18.010 ;
        RECT 2238.920 17.690 2239.180 18.010 ;
        RECT 2233.000 2.400 2233.140 17.690 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1020.425 16.745 1020.595 20.315 ;
      LAYER mcon ;
        RECT 1020.425 20.145 1020.595 20.315 ;
      LAYER met1 ;
        RECT 787.590 20.300 787.910 20.360 ;
        RECT 1020.365 20.300 1020.655 20.345 ;
        RECT 787.590 20.160 1020.655 20.300 ;
        RECT 787.590 20.100 787.910 20.160 ;
        RECT 1020.365 20.115 1020.655 20.160 ;
        RECT 1020.365 16.900 1020.655 16.945 ;
        RECT 1072.790 16.900 1073.110 16.960 ;
        RECT 1020.365 16.760 1073.110 16.900 ;
        RECT 1020.365 16.715 1020.655 16.760 ;
        RECT 1072.790 16.700 1073.110 16.760 ;
      LAYER via ;
        RECT 787.620 20.100 787.880 20.360 ;
        RECT 1072.820 16.700 1073.080 16.960 ;
      LAYER met2 ;
        RECT 787.620 20.070 787.880 20.390 ;
        RECT 787.680 2.400 787.820 20.070 ;
        RECT 1072.880 16.990 1073.020 54.000 ;
        RECT 1072.820 16.670 1073.080 16.990 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2269.785 10.285 2269.955 19.295 ;
        RECT 2317.625 18.105 2317.795 19.975 ;
        RECT 2318.545 18.105 2318.715 19.975 ;
        RECT 2366.385 18.105 2366.555 19.975 ;
        RECT 2415.605 18.105 2416.695 18.275 ;
        RECT 2463.445 16.405 2463.615 18.275 ;
        RECT 2511.285 16.405 2511.455 18.275 ;
        RECT 2511.745 18.105 2513.295 18.275 ;
      LAYER mcon ;
        RECT 2317.625 19.805 2317.795 19.975 ;
        RECT 2269.785 19.125 2269.955 19.295 ;
        RECT 2318.545 19.805 2318.715 19.975 ;
        RECT 2366.385 19.805 2366.555 19.975 ;
        RECT 2416.525 18.105 2416.695 18.275 ;
        RECT 2463.445 18.105 2463.615 18.275 ;
        RECT 2511.285 18.105 2511.455 18.275 ;
        RECT 2513.125 18.105 2513.295 18.275 ;
      LAYER met1 ;
        RECT 2317.565 19.960 2317.855 20.005 ;
        RECT 2270.260 19.820 2317.855 19.960 ;
        RECT 2269.725 19.280 2270.015 19.325 ;
        RECT 2270.260 19.280 2270.400 19.820 ;
        RECT 2317.565 19.775 2317.855 19.820 ;
        RECT 2318.485 19.960 2318.775 20.005 ;
        RECT 2366.325 19.960 2366.615 20.005 ;
        RECT 2318.485 19.820 2366.615 19.960 ;
        RECT 2318.485 19.775 2318.775 19.820 ;
        RECT 2366.325 19.775 2366.615 19.820 ;
        RECT 2269.725 19.140 2270.400 19.280 ;
        RECT 2269.725 19.095 2270.015 19.140 ;
        RECT 2317.565 18.260 2317.855 18.305 ;
        RECT 2318.485 18.260 2318.775 18.305 ;
        RECT 2317.565 18.120 2318.775 18.260 ;
        RECT 2317.565 18.075 2317.855 18.120 ;
        RECT 2318.485 18.075 2318.775 18.120 ;
        RECT 2366.325 18.260 2366.615 18.305 ;
        RECT 2415.545 18.260 2415.835 18.305 ;
        RECT 2366.325 18.120 2415.835 18.260 ;
        RECT 2366.325 18.075 2366.615 18.120 ;
        RECT 2415.545 18.075 2415.835 18.120 ;
        RECT 2416.465 18.260 2416.755 18.305 ;
        RECT 2463.385 18.260 2463.675 18.305 ;
        RECT 2416.465 18.120 2463.675 18.260 ;
        RECT 2416.465 18.075 2416.755 18.120 ;
        RECT 2463.385 18.075 2463.675 18.120 ;
        RECT 2511.225 18.260 2511.515 18.305 ;
        RECT 2511.685 18.260 2511.975 18.305 ;
        RECT 2511.225 18.120 2511.975 18.260 ;
        RECT 2511.225 18.075 2511.515 18.120 ;
        RECT 2511.685 18.075 2511.975 18.120 ;
        RECT 2513.065 18.260 2513.355 18.305 ;
        RECT 2590.790 18.260 2591.110 18.320 ;
        RECT 2513.065 18.120 2591.110 18.260 ;
        RECT 2513.065 18.075 2513.355 18.120 ;
        RECT 2590.790 18.060 2591.110 18.120 ;
        RECT 2463.385 16.560 2463.675 16.605 ;
        RECT 2511.225 16.560 2511.515 16.605 ;
        RECT 2463.385 16.420 2511.515 16.560 ;
        RECT 2463.385 16.375 2463.675 16.420 ;
        RECT 2511.225 16.375 2511.515 16.420 ;
        RECT 2250.850 10.440 2251.170 10.500 ;
        RECT 2269.725 10.440 2270.015 10.485 ;
        RECT 2250.850 10.300 2270.015 10.440 ;
        RECT 2250.850 10.240 2251.170 10.300 ;
        RECT 2269.725 10.255 2270.015 10.300 ;
      LAYER via ;
        RECT 2590.820 18.060 2591.080 18.320 ;
        RECT 2250.880 10.240 2251.140 10.500 ;
      LAYER met2 ;
        RECT 2590.880 18.350 2591.020 54.000 ;
        RECT 2590.820 18.030 2591.080 18.350 ;
        RECT 2250.880 10.210 2251.140 10.530 ;
        RECT 2250.940 2.400 2251.080 10.210 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2268.330 16.900 2268.650 16.960 ;
        RECT 2287.190 16.900 2287.510 16.960 ;
        RECT 2268.330 16.760 2287.510 16.900 ;
        RECT 2268.330 16.700 2268.650 16.760 ;
        RECT 2287.190 16.700 2287.510 16.760 ;
      LAYER via ;
        RECT 2268.360 16.700 2268.620 16.960 ;
        RECT 2287.220 16.700 2287.480 16.960 ;
      LAYER met2 ;
        RECT 2287.280 16.990 2287.420 54.000 ;
        RECT 2268.360 16.670 2268.620 16.990 ;
        RECT 2287.220 16.670 2287.480 16.990 ;
        RECT 2268.420 2.400 2268.560 16.670 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2415.145 18.445 2416.235 18.615 ;
      LAYER mcon ;
        RECT 2416.065 18.445 2416.235 18.615 ;
      LAYER met1 ;
        RECT 2286.270 18.600 2286.590 18.660 ;
        RECT 2415.085 18.600 2415.375 18.645 ;
        RECT 2286.270 18.460 2415.375 18.600 ;
        RECT 2286.270 18.400 2286.590 18.460 ;
        RECT 2415.085 18.415 2415.375 18.460 ;
        RECT 2416.005 18.600 2416.295 18.645 ;
        RECT 2602.750 18.600 2603.070 18.660 ;
        RECT 2416.005 18.460 2512.360 18.600 ;
        RECT 2416.005 18.415 2416.295 18.460 ;
        RECT 2512.220 18.260 2512.360 18.460 ;
        RECT 2512.680 18.460 2603.070 18.600 ;
        RECT 2512.680 18.260 2512.820 18.460 ;
        RECT 2602.750 18.400 2603.070 18.460 ;
        RECT 2512.220 18.120 2512.820 18.260 ;
      LAYER via ;
        RECT 2286.300 18.400 2286.560 18.660 ;
        RECT 2602.780 18.400 2603.040 18.660 ;
      LAYER met2 ;
        RECT 2602.840 18.690 2602.980 54.000 ;
        RECT 2286.300 18.370 2286.560 18.690 ;
        RECT 2602.780 18.370 2603.040 18.690 ;
        RECT 2286.360 2.400 2286.500 18.370 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2415.145 19.125 2416.235 19.295 ;
      LAYER mcon ;
        RECT 2416.065 19.125 2416.235 19.295 ;
      LAYER met1 ;
        RECT 2304.210 19.280 2304.530 19.340 ;
        RECT 2415.085 19.280 2415.375 19.325 ;
        RECT 2304.210 19.140 2415.375 19.280 ;
        RECT 2304.210 19.080 2304.530 19.140 ;
        RECT 2415.085 19.095 2415.375 19.140 ;
        RECT 2416.005 19.280 2416.295 19.325 ;
        RECT 2570.090 19.280 2570.410 19.340 ;
        RECT 2416.005 19.140 2570.410 19.280 ;
        RECT 2416.005 19.095 2416.295 19.140 ;
        RECT 2570.090 19.080 2570.410 19.140 ;
      LAYER via ;
        RECT 2304.240 19.080 2304.500 19.340 ;
        RECT 2570.120 19.080 2570.380 19.340 ;
      LAYER met2 ;
        RECT 2570.180 19.370 2570.320 54.000 ;
        RECT 2304.240 19.050 2304.500 19.370 ;
        RECT 2570.120 19.050 2570.380 19.370 ;
        RECT 2304.300 2.400 2304.440 19.050 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2415.605 18.785 2416.695 18.955 ;
        RECT 2512.205 18.785 2513.295 18.955 ;
      LAYER mcon ;
        RECT 2416.525 18.785 2416.695 18.955 ;
        RECT 2513.125 18.785 2513.295 18.955 ;
      LAYER met1 ;
        RECT 2322.150 18.940 2322.470 19.000 ;
        RECT 2415.545 18.940 2415.835 18.985 ;
        RECT 2322.150 18.800 2415.835 18.940 ;
        RECT 2322.150 18.740 2322.470 18.800 ;
        RECT 2415.545 18.755 2415.835 18.800 ;
        RECT 2416.465 18.940 2416.755 18.985 ;
        RECT 2512.145 18.940 2512.435 18.985 ;
        RECT 2416.465 18.800 2512.435 18.940 ;
        RECT 2416.465 18.755 2416.755 18.800 ;
        RECT 2512.145 18.755 2512.435 18.800 ;
        RECT 2513.065 18.940 2513.355 18.985 ;
        RECT 2616.090 18.940 2616.410 19.000 ;
        RECT 2513.065 18.800 2616.410 18.940 ;
        RECT 2513.065 18.755 2513.355 18.800 ;
        RECT 2616.090 18.740 2616.410 18.800 ;
      LAYER via ;
        RECT 2322.180 18.740 2322.440 19.000 ;
        RECT 2616.120 18.740 2616.380 19.000 ;
      LAYER met2 ;
        RECT 2616.180 19.030 2616.320 54.000 ;
        RECT 2322.180 18.710 2322.440 19.030 ;
        RECT 2616.120 18.710 2616.380 19.030 ;
        RECT 2322.240 2.400 2322.380 18.710 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2339.630 16.900 2339.950 16.960 ;
        RECT 2345.150 16.900 2345.470 16.960 ;
        RECT 2339.630 16.760 2345.470 16.900 ;
        RECT 2339.630 16.700 2339.950 16.760 ;
        RECT 2345.150 16.700 2345.470 16.760 ;
      LAYER via ;
        RECT 2339.660 16.700 2339.920 16.960 ;
        RECT 2345.180 16.700 2345.440 16.960 ;
      LAYER met2 ;
        RECT 2345.240 16.990 2345.380 54.000 ;
        RECT 2339.660 16.670 2339.920 16.990 ;
        RECT 2345.180 16.670 2345.440 16.990 ;
        RECT 2339.720 2.400 2339.860 16.670 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2511.745 19.465 2513.295 19.635 ;
      LAYER mcon ;
        RECT 2513.125 19.465 2513.295 19.635 ;
      LAYER met1 ;
        RECT 2357.570 19.620 2357.890 19.680 ;
        RECT 2511.685 19.620 2511.975 19.665 ;
        RECT 2357.570 19.480 2511.975 19.620 ;
        RECT 2357.570 19.420 2357.890 19.480 ;
        RECT 2511.685 19.435 2511.975 19.480 ;
        RECT 2513.065 19.620 2513.355 19.665 ;
        RECT 2623.450 19.620 2623.770 19.680 ;
        RECT 2513.065 19.480 2623.770 19.620 ;
        RECT 2513.065 19.435 2513.355 19.480 ;
        RECT 2623.450 19.420 2623.770 19.480 ;
      LAYER via ;
        RECT 2357.600 19.420 2357.860 19.680 ;
        RECT 2623.480 19.420 2623.740 19.680 ;
      LAYER met2 ;
        RECT 2623.540 19.710 2623.680 54.000 ;
        RECT 2357.600 19.390 2357.860 19.710 ;
        RECT 2623.480 19.390 2623.740 19.710 ;
        RECT 2357.660 2.400 2357.800 19.390 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2375.510 16.900 2375.830 16.960 ;
        RECT 2380.110 16.900 2380.430 16.960 ;
        RECT 2375.510 16.760 2380.430 16.900 ;
        RECT 2375.510 16.700 2375.830 16.760 ;
        RECT 2380.110 16.700 2380.430 16.760 ;
      LAYER via ;
        RECT 2375.540 16.700 2375.800 16.960 ;
        RECT 2380.140 16.700 2380.400 16.960 ;
      LAYER met2 ;
        RECT 2380.200 16.990 2380.340 54.000 ;
        RECT 2375.540 16.670 2375.800 16.990 ;
        RECT 2380.140 16.670 2380.400 16.990 ;
        RECT 2375.600 2.400 2375.740 16.670 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2512.665 19.805 2513.755 19.975 ;
      LAYER mcon ;
        RECT 2513.585 19.805 2513.755 19.975 ;
      LAYER met1 ;
        RECT 2393.450 19.960 2393.770 20.020 ;
        RECT 2512.605 19.960 2512.895 20.005 ;
        RECT 2393.450 19.820 2512.895 19.960 ;
        RECT 2393.450 19.760 2393.770 19.820 ;
        RECT 2512.605 19.775 2512.895 19.820 ;
        RECT 2513.525 19.960 2513.815 20.005 ;
        RECT 2636.790 19.960 2637.110 20.020 ;
        RECT 2513.525 19.820 2637.110 19.960 ;
        RECT 2513.525 19.775 2513.815 19.820 ;
        RECT 2636.790 19.760 2637.110 19.820 ;
      LAYER via ;
        RECT 2393.480 19.760 2393.740 20.020 ;
        RECT 2636.820 19.760 2637.080 20.020 ;
      LAYER met2 ;
        RECT 2636.880 20.050 2637.020 54.000 ;
        RECT 2393.480 19.730 2393.740 20.050 ;
        RECT 2636.820 19.730 2637.080 20.050 ;
        RECT 2393.540 2.400 2393.680 19.730 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2411.390 16.900 2411.710 16.960 ;
        RECT 2414.610 16.900 2414.930 16.960 ;
        RECT 2411.390 16.760 2414.930 16.900 ;
        RECT 2411.390 16.700 2411.710 16.760 ;
        RECT 2414.610 16.700 2414.930 16.760 ;
      LAYER via ;
        RECT 2411.420 16.700 2411.680 16.960 ;
        RECT 2414.640 16.700 2414.900 16.960 ;
      LAYER met2 ;
        RECT 2414.700 16.990 2414.840 54.000 ;
        RECT 2411.420 16.670 2411.680 16.990 ;
        RECT 2414.640 16.670 2414.900 16.990 ;
        RECT 2411.480 2.400 2411.620 16.670 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 51.580 807.230 51.640 ;
        RECT 1651.470 51.580 1651.790 51.640 ;
        RECT 806.910 51.440 1651.790 51.580 ;
        RECT 806.910 51.380 807.230 51.440 ;
        RECT 1651.470 51.380 1651.790 51.440 ;
        RECT 805.530 2.960 805.850 3.020 ;
        RECT 806.910 2.960 807.230 3.020 ;
        RECT 805.530 2.820 807.230 2.960 ;
        RECT 805.530 2.760 805.850 2.820 ;
        RECT 806.910 2.760 807.230 2.820 ;
      LAYER via ;
        RECT 806.940 51.380 807.200 51.640 ;
        RECT 1651.500 51.380 1651.760 51.640 ;
        RECT 805.560 2.760 805.820 3.020 ;
        RECT 806.940 2.760 807.200 3.020 ;
      LAYER met2 ;
        RECT 1651.560 51.670 1651.700 54.000 ;
        RECT 806.940 51.350 807.200 51.670 ;
        RECT 1651.500 51.350 1651.760 51.670 ;
        RECT 807.000 3.050 807.140 51.350 ;
        RECT 805.560 2.730 805.820 3.050 ;
        RECT 806.940 2.730 807.200 3.050 ;
        RECT 805.620 2.400 805.760 2.730 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2818.490 17.920 2818.810 17.980 ;
        RECT 2916.930 17.920 2917.250 17.980 ;
        RECT 2818.490 17.780 2917.250 17.920 ;
        RECT 2818.490 17.720 2818.810 17.780 ;
        RECT 2916.930 17.720 2917.250 17.780 ;
      LAYER via ;
        RECT 2818.520 17.720 2818.780 17.980 ;
        RECT 2916.960 17.720 2917.220 17.980 ;
      LAYER met2 ;
        RECT 2818.580 18.010 2818.720 54.000 ;
        RECT 2818.520 17.690 2818.780 18.010 ;
        RECT 2916.960 17.690 2917.220 18.010 ;
        RECT 2917.020 2.400 2917.160 17.690 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.610 1128.020 45.930 1128.080 ;
        RECT 45.610 1127.880 54.000 1128.020 ;
        RECT 45.610 1127.820 45.930 1127.880 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 45.610 17.240 45.930 17.300 ;
        RECT 2.830 17.100 45.930 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 45.610 17.040 45.930 17.100 ;
      LAYER via ;
        RECT 45.640 1127.820 45.900 1128.080 ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 45.640 17.040 45.900 17.300 ;
      LAYER met2 ;
        RECT 45.640 1127.790 45.900 1128.110 ;
        RECT 45.700 17.330 45.840 1127.790 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 45.640 17.010 45.900 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 52.050 51.580 52.370 51.640 ;
        RECT 600.370 51.580 600.690 51.640 ;
        RECT 52.050 51.440 600.690 51.580 ;
        RECT 52.050 51.380 52.370 51.440 ;
        RECT 600.370 51.380 600.690 51.440 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 52.050 17.580 52.370 17.640 ;
        RECT 8.350 17.440 52.370 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 52.050 17.380 52.370 17.440 ;
      LAYER via ;
        RECT 52.080 51.380 52.340 51.640 ;
        RECT 600.400 51.380 600.660 51.640 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 52.080 17.380 52.340 17.640 ;
      LAYER met2 ;
        RECT 600.460 51.670 600.600 54.000 ;
        RECT 52.080 51.350 52.340 51.670 ;
        RECT 600.400 51.350 600.660 51.670 ;
        RECT 52.140 17.670 52.280 51.350 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 52.080 17.350 52.340 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 51.590 141.340 51.910 141.400 ;
        RECT 51.590 141.200 54.000 141.340 ;
        RECT 51.590 141.140 51.910 141.200 ;
        RECT 14.330 18.600 14.650 18.660 ;
        RECT 51.590 18.600 51.910 18.660 ;
        RECT 14.330 18.460 51.910 18.600 ;
        RECT 14.330 18.400 14.650 18.460 ;
        RECT 51.590 18.400 51.910 18.460 ;
      LAYER via ;
        RECT 51.620 141.140 51.880 141.400 ;
        RECT 14.360 18.400 14.620 18.660 ;
        RECT 51.620 18.400 51.880 18.660 ;
      LAYER met2 ;
        RECT 51.620 141.110 51.880 141.430 ;
        RECT 51.680 18.690 51.820 141.110 ;
        RECT 14.360 18.370 14.620 18.690 ;
        RECT 51.620 18.370 51.880 18.690 ;
        RECT 14.420 2.400 14.560 18.370 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 16.900 38.570 16.960 ;
        RECT 58.490 16.900 58.810 16.960 ;
        RECT 38.250 16.760 58.810 16.900 ;
        RECT 38.250 16.700 38.570 16.760 ;
        RECT 58.490 16.700 58.810 16.760 ;
      LAYER via ;
        RECT 38.280 16.700 38.540 16.960 ;
        RECT 58.520 16.700 58.780 16.960 ;
      LAYER met2 ;
        RECT 58.580 16.990 58.720 54.000 ;
        RECT 38.280 16.670 38.540 16.990 ;
        RECT 58.520 16.670 58.780 16.990 ;
        RECT 38.340 2.400 38.480 16.670 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.200 17.410 241.340 54.000 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 16.900 258.450 16.960 ;
        RECT 261.810 16.900 262.130 16.960 ;
        RECT 258.130 16.760 262.130 16.900 ;
        RECT 258.130 16.700 258.450 16.760 ;
        RECT 261.810 16.700 262.130 16.760 ;
      LAYER via ;
        RECT 258.160 16.700 258.420 16.960 ;
        RECT 261.840 16.700 262.100 16.960 ;
      LAYER met2 ;
        RECT 261.900 16.990 262.040 54.000 ;
        RECT 258.160 16.670 258.420 16.990 ;
        RECT 261.840 16.670 262.100 16.990 ;
        RECT 258.220 2.400 258.360 16.670 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 15.540 276.390 15.600 ;
        RECT 282.510 15.540 282.830 15.600 ;
        RECT 276.070 15.400 282.830 15.540 ;
        RECT 276.070 15.340 276.390 15.400 ;
        RECT 282.510 15.340 282.830 15.400 ;
      LAYER via ;
        RECT 276.100 15.340 276.360 15.600 ;
        RECT 282.540 15.340 282.800 15.600 ;
      LAYER met2 ;
        RECT 282.600 15.630 282.740 54.000 ;
        RECT 276.100 15.310 276.360 15.630 ;
        RECT 282.540 15.310 282.800 15.630 ;
        RECT 276.160 2.400 276.300 15.310 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 16.560 294.330 16.620 ;
        RECT 296.310 16.560 296.630 16.620 ;
        RECT 294.010 16.420 296.630 16.560 ;
        RECT 294.010 16.360 294.330 16.420 ;
        RECT 296.310 16.360 296.630 16.420 ;
      LAYER via ;
        RECT 294.040 16.360 294.300 16.620 ;
        RECT 296.340 16.360 296.600 16.620 ;
      LAYER met2 ;
        RECT 296.400 16.650 296.540 54.000 ;
        RECT 294.040 16.330 294.300 16.650 ;
        RECT 296.340 16.330 296.600 16.650 ;
        RECT 294.100 2.400 294.240 16.330 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 14.860 312.270 14.920 ;
        RECT 317.010 14.860 317.330 14.920 ;
        RECT 311.950 14.720 317.330 14.860 ;
        RECT 311.950 14.660 312.270 14.720 ;
        RECT 317.010 14.660 317.330 14.720 ;
      LAYER via ;
        RECT 311.980 14.660 312.240 14.920 ;
        RECT 317.040 14.660 317.300 14.920 ;
      LAYER met2 ;
        RECT 317.100 14.950 317.240 54.000 ;
        RECT 311.980 14.630 312.240 14.950 ;
        RECT 317.040 14.630 317.300 14.950 ;
        RECT 312.040 2.400 312.180 14.630 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 329.965 48.365 330.135 54.000 ;
      LAYER met1 ;
        RECT 329.890 48.520 330.210 48.580 ;
        RECT 329.695 48.380 330.210 48.520 ;
        RECT 329.890 48.320 330.210 48.380 ;
        RECT 329.430 2.960 329.750 3.020 ;
        RECT 329.890 2.960 330.210 3.020 ;
        RECT 329.430 2.820 330.210 2.960 ;
        RECT 329.430 2.760 329.750 2.820 ;
        RECT 329.890 2.760 330.210 2.820 ;
      LAYER via ;
        RECT 329.920 48.320 330.180 48.580 ;
        RECT 329.460 2.760 329.720 3.020 ;
        RECT 329.920 2.760 330.180 3.020 ;
      LAYER met2 ;
        RECT 329.920 48.290 330.180 48.610 ;
        RECT 329.980 48.010 330.120 48.290 ;
        RECT 329.520 47.870 330.120 48.010 ;
        RECT 329.520 3.050 329.660 47.870 ;
        RECT 329.460 2.730 329.720 3.050 ;
        RECT 329.920 2.730 330.180 3.050 ;
        RECT 329.980 2.400 330.120 2.730 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 25.740 347.690 25.800 ;
        RECT 848.770 25.740 849.090 25.800 ;
        RECT 347.370 25.600 849.090 25.740 ;
        RECT 347.370 25.540 347.690 25.600 ;
        RECT 848.770 25.540 849.090 25.600 ;
      LAYER via ;
        RECT 347.400 25.540 347.660 25.800 ;
        RECT 848.800 25.540 849.060 25.800 ;
      LAYER met2 ;
        RECT 848.860 25.830 849.000 54.000 ;
        RECT 347.400 25.510 347.660 25.830 ;
        RECT 848.800 25.510 849.060 25.830 ;
        RECT 347.460 2.400 347.600 25.510 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 25.400 365.630 25.460 ;
        RECT 862.570 25.400 862.890 25.460 ;
        RECT 365.310 25.260 862.890 25.400 ;
        RECT 365.310 25.200 365.630 25.260 ;
        RECT 862.570 25.200 862.890 25.260 ;
      LAYER via ;
        RECT 365.340 25.200 365.600 25.460 ;
        RECT 862.600 25.200 862.860 25.460 ;
      LAYER met2 ;
        RECT 862.660 25.490 862.800 54.000 ;
        RECT 365.340 25.170 365.600 25.490 ;
        RECT 862.600 25.170 862.860 25.490 ;
        RECT 365.400 2.400 365.540 25.170 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 26.080 383.570 26.140 ;
        RECT 876.370 26.080 876.690 26.140 ;
        RECT 383.250 25.940 876.690 26.080 ;
        RECT 383.250 25.880 383.570 25.940 ;
        RECT 876.370 25.880 876.690 25.940 ;
      LAYER via ;
        RECT 383.280 25.880 383.540 26.140 ;
        RECT 876.400 25.880 876.660 26.140 ;
      LAYER met2 ;
        RECT 876.460 26.170 876.600 54.000 ;
        RECT 383.280 25.850 383.540 26.170 ;
        RECT 876.400 25.850 876.660 26.170 ;
        RECT 383.340 2.400 383.480 25.850 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 26.420 401.510 26.480 ;
        RECT 890.170 26.420 890.490 26.480 ;
        RECT 401.190 26.280 890.490 26.420 ;
        RECT 401.190 26.220 401.510 26.280 ;
        RECT 890.170 26.220 890.490 26.280 ;
      LAYER via ;
        RECT 401.220 26.220 401.480 26.480 ;
        RECT 890.200 26.220 890.460 26.480 ;
      LAYER met2 ;
        RECT 890.260 26.510 890.400 54.000 ;
        RECT 401.220 26.190 401.480 26.510 ;
        RECT 890.200 26.190 890.460 26.510 ;
        RECT 401.280 2.400 401.420 26.190 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 641.860 24.325 642.000 54.000 ;
        RECT 62.190 23.955 62.470 24.325 ;
        RECT 641.790 23.955 642.070 24.325 ;
        RECT 62.260 2.400 62.400 23.955 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 62.190 24.000 62.470 24.280 ;
        RECT 641.790 24.000 642.070 24.280 ;
      LAYER met3 ;
        RECT 62.165 24.290 62.495 24.305 ;
        RECT 641.765 24.290 642.095 24.305 ;
        RECT 62.165 23.990 642.095 24.290 ;
        RECT 62.165 23.975 62.495 23.990 ;
        RECT 641.765 23.975 642.095 23.990 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 897.145 48.365 897.315 54.000 ;
      LAYER met1 ;
        RECT 897.070 48.520 897.390 48.580 ;
        RECT 896.875 48.380 897.390 48.520 ;
        RECT 897.070 48.320 897.390 48.380 ;
        RECT 419.130 26.760 419.450 26.820 ;
        RECT 897.070 26.760 897.390 26.820 ;
        RECT 419.130 26.620 897.390 26.760 ;
        RECT 419.130 26.560 419.450 26.620 ;
        RECT 897.070 26.560 897.390 26.620 ;
      LAYER via ;
        RECT 897.100 48.320 897.360 48.580 ;
        RECT 419.160 26.560 419.420 26.820 ;
        RECT 897.100 26.560 897.360 26.820 ;
      LAYER met2 ;
        RECT 897.100 48.290 897.360 48.610 ;
        RECT 897.160 26.850 897.300 48.290 ;
        RECT 419.160 26.530 419.420 26.850 ;
        RECT 897.100 26.530 897.360 26.850 ;
        RECT 419.220 2.400 419.360 26.530 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 910.945 48.365 911.115 54.000 ;
      LAYER met1 ;
        RECT 910.870 48.520 911.190 48.580 ;
        RECT 910.675 48.380 911.190 48.520 ;
        RECT 910.870 48.320 911.190 48.380 ;
        RECT 436.610 27.100 436.930 27.160 ;
        RECT 910.870 27.100 911.190 27.160 ;
        RECT 436.610 26.960 911.190 27.100 ;
        RECT 436.610 26.900 436.930 26.960 ;
        RECT 910.870 26.900 911.190 26.960 ;
      LAYER via ;
        RECT 910.900 48.320 911.160 48.580 ;
        RECT 436.640 26.900 436.900 27.160 ;
        RECT 910.900 26.900 911.160 27.160 ;
      LAYER met2 ;
        RECT 910.900 48.290 911.160 48.610 ;
        RECT 910.960 27.190 911.100 48.290 ;
        RECT 436.640 26.870 436.900 27.190 ;
        RECT 910.900 26.870 911.160 27.190 ;
        RECT 436.700 2.400 436.840 26.870 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 27.440 454.870 27.500 ;
        RECT 923.750 27.440 924.070 27.500 ;
        RECT 454.550 27.300 924.070 27.440 ;
        RECT 454.550 27.240 454.870 27.300 ;
        RECT 923.750 27.240 924.070 27.300 ;
      LAYER via ;
        RECT 454.580 27.240 454.840 27.500 ;
        RECT 923.780 27.240 924.040 27.500 ;
      LAYER met2 ;
        RECT 922.920 48.805 923.060 54.000 ;
        RECT 922.850 48.435 923.130 48.805 ;
        RECT 923.770 48.435 924.050 48.805 ;
        RECT 923.840 27.530 923.980 48.435 ;
        RECT 454.580 27.210 454.840 27.530 ;
        RECT 923.780 27.210 924.040 27.530 ;
        RECT 454.640 2.400 454.780 27.210 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 922.850 48.480 923.130 48.760 ;
        RECT 923.770 48.480 924.050 48.760 ;
      LAYER met3 ;
        RECT 922.825 48.770 923.155 48.785 ;
        RECT 923.745 48.770 924.075 48.785 ;
        RECT 922.825 48.470 924.075 48.770 ;
        RECT 922.825 48.455 923.155 48.470 ;
        RECT 923.745 48.455 924.075 48.470 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 23.700 472.810 23.760 ;
        RECT 938.470 23.700 938.790 23.760 ;
        RECT 472.490 23.560 938.790 23.700 ;
        RECT 472.490 23.500 472.810 23.560 ;
        RECT 938.470 23.500 938.790 23.560 ;
      LAYER via ;
        RECT 472.520 23.500 472.780 23.760 ;
        RECT 938.500 23.500 938.760 23.760 ;
      LAYER met2 ;
        RECT 938.560 23.790 938.700 54.000 ;
        RECT 472.520 23.470 472.780 23.790 ;
        RECT 938.500 23.470 938.760 23.790 ;
        RECT 472.580 2.400 472.720 23.470 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 23.360 490.750 23.420 ;
        RECT 952.270 23.360 952.590 23.420 ;
        RECT 490.430 23.220 952.590 23.360 ;
        RECT 490.430 23.160 490.750 23.220 ;
        RECT 952.270 23.160 952.590 23.220 ;
      LAYER via ;
        RECT 490.460 23.160 490.720 23.420 ;
        RECT 952.300 23.160 952.560 23.420 ;
      LAYER met2 ;
        RECT 952.360 23.450 952.500 54.000 ;
        RECT 490.460 23.130 490.720 23.450 ;
        RECT 952.300 23.130 952.560 23.450 ;
        RECT 490.520 2.400 490.660 23.130 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 23.020 508.230 23.080 ;
        RECT 966.070 23.020 966.390 23.080 ;
        RECT 507.910 22.880 966.390 23.020 ;
        RECT 507.910 22.820 508.230 22.880 ;
        RECT 966.070 22.820 966.390 22.880 ;
      LAYER via ;
        RECT 507.940 22.820 508.200 23.080 ;
        RECT 966.100 22.820 966.360 23.080 ;
      LAYER met2 ;
        RECT 966.160 23.110 966.300 54.000 ;
        RECT 507.940 22.790 508.200 23.110 ;
        RECT 966.100 22.790 966.360 23.110 ;
        RECT 508.000 2.400 508.140 22.790 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 22.340 526.170 22.400 ;
        RECT 979.870 22.340 980.190 22.400 ;
        RECT 525.850 22.200 980.190 22.340 ;
        RECT 525.850 22.140 526.170 22.200 ;
        RECT 979.870 22.140 980.190 22.200 ;
      LAYER via ;
        RECT 525.880 22.140 526.140 22.400 ;
        RECT 979.900 22.140 980.160 22.400 ;
      LAYER met2 ;
        RECT 979.960 22.430 980.100 54.000 ;
        RECT 525.880 22.110 526.140 22.430 ;
        RECT 979.900 22.110 980.160 22.430 ;
        RECT 525.940 2.400 526.080 22.110 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 22.680 544.110 22.740 ;
        RECT 993.670 22.680 993.990 22.740 ;
        RECT 543.790 22.540 993.990 22.680 ;
        RECT 543.790 22.480 544.110 22.540 ;
        RECT 993.670 22.480 993.990 22.540 ;
      LAYER via ;
        RECT 543.820 22.480 544.080 22.740 ;
        RECT 993.700 22.480 993.960 22.740 ;
      LAYER met2 ;
        RECT 993.760 22.770 993.900 54.000 ;
        RECT 543.820 22.450 544.080 22.770 ;
        RECT 993.700 22.450 993.960 22.770 ;
        RECT 543.880 2.400 544.020 22.450 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 22.000 562.050 22.060 ;
        RECT 1007.010 22.000 1007.330 22.060 ;
        RECT 561.730 21.860 1007.330 22.000 ;
        RECT 561.730 21.800 562.050 21.860 ;
        RECT 1007.010 21.800 1007.330 21.860 ;
      LAYER via ;
        RECT 561.760 21.800 562.020 22.060 ;
        RECT 1007.040 21.800 1007.300 22.060 ;
      LAYER met2 ;
        RECT 1007.560 24.890 1007.700 54.000 ;
        RECT 1007.100 24.750 1007.700 24.890 ;
        RECT 1007.100 22.090 1007.240 24.750 ;
        RECT 561.760 21.770 562.020 22.090 ;
        RECT 1007.040 21.770 1007.300 22.090 ;
        RECT 561.820 2.400 561.960 21.770 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 21.320 579.990 21.380 ;
        RECT 1015.290 21.320 1015.610 21.380 ;
        RECT 579.670 21.180 1015.610 21.320 ;
        RECT 579.670 21.120 579.990 21.180 ;
        RECT 1015.290 21.120 1015.610 21.180 ;
      LAYER via ;
        RECT 579.700 21.120 579.960 21.380 ;
        RECT 1015.320 21.120 1015.580 21.380 ;
      LAYER met2 ;
        RECT 1015.380 21.410 1015.520 54.000 ;
        RECT 579.700 21.090 579.960 21.410 ;
        RECT 1015.320 21.090 1015.580 21.410 ;
        RECT 579.760 2.400 579.900 21.090 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 24.380 86.410 24.440 ;
        RECT 656.030 24.380 656.350 24.440 ;
        RECT 86.090 24.240 656.350 24.380 ;
        RECT 86.090 24.180 86.410 24.240 ;
        RECT 656.030 24.180 656.350 24.240 ;
      LAYER via ;
        RECT 86.120 24.180 86.380 24.440 ;
        RECT 656.060 24.180 656.320 24.440 ;
      LAYER met2 ;
        RECT 656.120 24.470 656.260 54.000 ;
        RECT 86.120 24.150 86.380 24.470 ;
        RECT 656.060 24.150 656.320 24.470 ;
        RECT 86.180 2.400 86.320 24.150 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1028.630 48.520 1028.950 48.580 ;
        RECT 1030.010 48.520 1030.330 48.580 ;
        RECT 1028.630 48.380 1030.330 48.520 ;
        RECT 1028.630 48.320 1028.950 48.380 ;
        RECT 1030.010 48.320 1030.330 48.380 ;
        RECT 597.150 21.660 597.470 21.720 ;
        RECT 614.630 21.660 614.950 21.720 ;
        RECT 597.150 21.520 614.950 21.660 ;
        RECT 597.150 21.460 597.470 21.520 ;
        RECT 614.630 21.460 614.950 21.520 ;
        RECT 628.430 21.660 628.750 21.720 ;
        RECT 1030.010 21.660 1030.330 21.720 ;
        RECT 628.430 21.520 1030.330 21.660 ;
        RECT 628.430 21.460 628.750 21.520 ;
        RECT 1030.010 21.460 1030.330 21.520 ;
      LAYER via ;
        RECT 1028.660 48.320 1028.920 48.580 ;
        RECT 1030.040 48.320 1030.300 48.580 ;
        RECT 597.180 21.460 597.440 21.720 ;
        RECT 614.660 21.460 614.920 21.720 ;
        RECT 628.460 21.460 628.720 21.720 ;
        RECT 1030.040 21.460 1030.300 21.720 ;
      LAYER met2 ;
        RECT 1028.720 48.610 1028.860 54.000 ;
        RECT 1028.660 48.290 1028.920 48.610 ;
        RECT 1030.040 48.290 1030.300 48.610 ;
        RECT 1030.100 21.750 1030.240 48.290 ;
        RECT 597.180 21.430 597.440 21.750 ;
        RECT 614.660 21.605 614.920 21.750 ;
        RECT 628.460 21.605 628.720 21.750 ;
        RECT 597.240 2.400 597.380 21.430 ;
        RECT 614.650 21.235 614.930 21.605 ;
        RECT 628.450 21.235 628.730 21.605 ;
        RECT 1030.040 21.430 1030.300 21.750 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 614.650 21.280 614.930 21.560 ;
        RECT 628.450 21.280 628.730 21.560 ;
      LAYER met3 ;
        RECT 614.625 21.570 614.955 21.585 ;
        RECT 628.425 21.570 628.755 21.585 ;
        RECT 614.625 21.270 628.755 21.570 ;
        RECT 614.625 21.255 614.955 21.270 ;
        RECT 628.425 21.255 628.755 21.270 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 628.045 20.825 628.215 21.675 ;
      LAYER mcon ;
        RECT 628.045 21.505 628.215 21.675 ;
      LAYER met1 ;
        RECT 1042.430 48.520 1042.750 48.580 ;
        RECT 1044.270 48.520 1044.590 48.580 ;
        RECT 1042.430 48.380 1044.590 48.520 ;
        RECT 1042.430 48.320 1042.750 48.380 ;
        RECT 1044.270 48.320 1044.590 48.380 ;
        RECT 615.090 21.660 615.410 21.720 ;
        RECT 627.985 21.660 628.275 21.705 ;
        RECT 615.090 21.520 628.275 21.660 ;
        RECT 615.090 21.460 615.410 21.520 ;
        RECT 627.985 21.475 628.275 21.520 ;
        RECT 627.985 20.980 628.275 21.025 ;
        RECT 1044.270 20.980 1044.590 21.040 ;
        RECT 627.985 20.840 1044.590 20.980 ;
        RECT 627.985 20.795 628.275 20.840 ;
        RECT 1044.270 20.780 1044.590 20.840 ;
      LAYER via ;
        RECT 1042.460 48.320 1042.720 48.580 ;
        RECT 1044.300 48.320 1044.560 48.580 ;
        RECT 615.120 21.460 615.380 21.720 ;
        RECT 1044.300 20.780 1044.560 21.040 ;
      LAYER met2 ;
        RECT 1042.520 48.610 1042.660 54.000 ;
        RECT 1042.460 48.290 1042.720 48.610 ;
        RECT 1044.300 48.290 1044.560 48.610 ;
        RECT 615.120 21.430 615.380 21.750 ;
        RECT 615.180 2.400 615.320 21.430 ;
        RECT 1044.360 21.070 1044.500 48.290 ;
        RECT 1044.300 20.750 1044.560 21.070 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 24.040 109.870 24.100 ;
        RECT 676.730 24.040 677.050 24.100 ;
        RECT 109.550 23.900 677.050 24.040 ;
        RECT 109.550 23.840 109.870 23.900 ;
        RECT 676.730 23.840 677.050 23.900 ;
      LAYER via ;
        RECT 109.580 23.840 109.840 24.100 ;
        RECT 676.760 23.840 677.020 24.100 ;
      LAYER met2 ;
        RECT 676.820 24.130 676.960 54.000 ;
        RECT 109.580 23.810 109.840 24.130 ;
        RECT 676.760 23.810 677.020 24.130 ;
        RECT 109.640 2.400 109.780 23.810 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 24.720 133.790 24.780 ;
        RECT 690.530 24.720 690.850 24.780 ;
        RECT 133.470 24.580 690.850 24.720 ;
        RECT 133.470 24.520 133.790 24.580 ;
        RECT 690.530 24.520 690.850 24.580 ;
      LAYER via ;
        RECT 133.500 24.520 133.760 24.780 ;
        RECT 690.560 24.520 690.820 24.780 ;
      LAYER met2 ;
        RECT 690.620 24.810 690.760 54.000 ;
        RECT 133.500 24.490 133.760 24.810 ;
        RECT 690.560 24.490 690.820 24.810 ;
        RECT 133.560 2.400 133.700 24.490 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 25.060 151.730 25.120 ;
        RECT 704.330 25.060 704.650 25.120 ;
        RECT 151.410 24.920 704.650 25.060 ;
        RECT 151.410 24.860 151.730 24.920 ;
        RECT 704.330 24.860 704.650 24.920 ;
      LAYER via ;
        RECT 151.440 24.860 151.700 25.120 ;
        RECT 704.360 24.860 704.620 25.120 ;
      LAYER met2 ;
        RECT 704.420 25.150 704.560 54.000 ;
        RECT 151.440 24.830 151.700 25.150 ;
        RECT 704.360 24.830 704.620 25.150 ;
        RECT 151.500 2.400 151.640 24.830 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 31.520 169.670 31.580 ;
        RECT 717.670 31.520 717.990 31.580 ;
        RECT 169.350 31.380 717.990 31.520 ;
        RECT 169.350 31.320 169.670 31.380 ;
        RECT 717.670 31.320 717.990 31.380 ;
      LAYER via ;
        RECT 169.380 31.320 169.640 31.580 ;
        RECT 717.700 31.320 717.960 31.580 ;
      LAYER met2 ;
        RECT 717.760 31.610 717.900 54.000 ;
        RECT 169.380 31.290 169.640 31.610 ;
        RECT 717.700 31.290 717.960 31.610 ;
        RECT 169.440 2.400 169.580 31.290 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 31.860 187.150 31.920 ;
        RECT 731.470 31.860 731.790 31.920 ;
        RECT 186.830 31.720 731.790 31.860 ;
        RECT 186.830 31.660 187.150 31.720 ;
        RECT 731.470 31.660 731.790 31.720 ;
      LAYER via ;
        RECT 186.860 31.660 187.120 31.920 ;
        RECT 731.500 31.660 731.760 31.920 ;
      LAYER met2 ;
        RECT 731.560 31.950 731.700 54.000 ;
        RECT 186.860 31.630 187.120 31.950 ;
        RECT 731.500 31.630 731.760 31.950 ;
        RECT 186.920 2.400 187.060 31.630 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 32.200 205.090 32.260 ;
        RECT 745.730 32.200 746.050 32.260 ;
        RECT 204.770 32.060 746.050 32.200 ;
        RECT 204.770 32.000 205.090 32.060 ;
        RECT 745.730 32.000 746.050 32.060 ;
      LAYER via ;
        RECT 204.800 32.000 205.060 32.260 ;
        RECT 745.760 32.000 746.020 32.260 ;
      LAYER met2 ;
        RECT 745.820 32.290 745.960 54.000 ;
        RECT 204.800 31.970 205.060 32.290 ;
        RECT 745.760 31.970 746.020 32.290 ;
        RECT 204.860 2.400 205.000 31.970 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 32.540 223.030 32.600 ;
        RECT 759.070 32.540 759.390 32.600 ;
        RECT 222.710 32.400 759.390 32.540 ;
        RECT 222.710 32.340 223.030 32.400 ;
        RECT 759.070 32.340 759.390 32.400 ;
      LAYER via ;
        RECT 222.740 32.340 223.000 32.600 ;
        RECT 759.100 32.340 759.360 32.600 ;
      LAYER met2 ;
        RECT 759.160 32.630 759.300 54.000 ;
        RECT 222.740 32.310 223.000 32.630 ;
        RECT 759.100 32.310 759.360 32.630 ;
        RECT 222.800 2.400 222.940 32.310 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 30.840 20.630 30.900 ;
        RECT 608.190 30.840 608.510 30.900 ;
        RECT 20.310 30.700 608.510 30.840 ;
        RECT 20.310 30.640 20.630 30.700 ;
        RECT 608.190 30.640 608.510 30.700 ;
      LAYER via ;
        RECT 20.340 30.640 20.600 30.900 ;
        RECT 608.220 30.640 608.480 30.900 ;
      LAYER met2 ;
        RECT 608.280 30.930 608.420 54.000 ;
        RECT 20.340 30.610 20.600 30.930 ;
        RECT 608.220 30.610 608.480 30.930 ;
        RECT 20.400 2.400 20.540 30.610 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 31.180 44.550 31.240 ;
        RECT 628.430 31.180 628.750 31.240 ;
        RECT 44.230 31.040 628.750 31.180 ;
        RECT 44.230 30.980 44.550 31.040 ;
        RECT 628.430 30.980 628.750 31.040 ;
      LAYER via ;
        RECT 44.260 30.980 44.520 31.240 ;
        RECT 628.460 30.980 628.720 31.240 ;
      LAYER met2 ;
        RECT 628.520 31.270 628.660 54.000 ;
        RECT 44.260 30.950 44.520 31.270 ;
        RECT 628.460 30.950 628.720 31.270 ;
        RECT 44.320 2.400 44.460 30.950 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 32.880 246.950 32.940 ;
        RECT 772.870 32.880 773.190 32.940 ;
        RECT 246.630 32.740 773.190 32.880 ;
        RECT 246.630 32.680 246.950 32.740 ;
        RECT 772.870 32.680 773.190 32.740 ;
      LAYER via ;
        RECT 246.660 32.680 246.920 32.940 ;
        RECT 772.900 32.680 773.160 32.940 ;
      LAYER met2 ;
        RECT 772.960 32.970 773.100 54.000 ;
        RECT 246.660 32.650 246.920 32.970 ;
        RECT 772.900 32.650 773.160 32.970 ;
        RECT 246.720 2.400 246.860 32.650 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 16.900 264.430 16.960 ;
        RECT 268.710 16.900 269.030 16.960 ;
        RECT 264.110 16.760 269.030 16.900 ;
        RECT 264.110 16.700 264.430 16.760 ;
        RECT 268.710 16.700 269.030 16.760 ;
      LAYER via ;
        RECT 264.140 16.700 264.400 16.960 ;
        RECT 268.740 16.700 269.000 16.960 ;
      LAYER met2 ;
        RECT 268.800 16.990 268.940 54.000 ;
        RECT 264.140 16.670 264.400 16.990 ;
        RECT 268.740 16.670 269.000 16.990 ;
        RECT 264.200 2.400 264.340 16.670 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 33.220 282.370 33.280 ;
        RECT 800.470 33.220 800.790 33.280 ;
        RECT 282.050 33.080 800.790 33.220 ;
        RECT 282.050 33.020 282.370 33.080 ;
        RECT 800.470 33.020 800.790 33.080 ;
      LAYER via ;
        RECT 282.080 33.020 282.340 33.280 ;
        RECT 800.500 33.020 800.760 33.280 ;
      LAYER met2 ;
        RECT 800.560 33.310 800.700 54.000 ;
        RECT 282.080 32.990 282.340 33.310 ;
        RECT 800.500 32.990 800.760 33.310 ;
        RECT 282.140 2.400 282.280 32.990 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 16.560 300.310 16.620 ;
        RECT 303.210 16.560 303.530 16.620 ;
        RECT 299.990 16.420 303.530 16.560 ;
        RECT 299.990 16.360 300.310 16.420 ;
        RECT 303.210 16.360 303.530 16.420 ;
      LAYER via ;
        RECT 300.020 16.360 300.280 16.620 ;
        RECT 303.240 16.360 303.500 16.620 ;
      LAYER met2 ;
        RECT 303.300 16.650 303.440 54.000 ;
        RECT 300.020 16.330 300.280 16.650 ;
        RECT 303.240 16.330 303.500 16.650 ;
        RECT 300.080 2.400 300.220 16.330 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 33.560 318.250 33.620 ;
        RECT 828.530 33.560 828.850 33.620 ;
        RECT 317.930 33.420 828.850 33.560 ;
        RECT 317.930 33.360 318.250 33.420 ;
        RECT 828.530 33.360 828.850 33.420 ;
      LAYER via ;
        RECT 317.960 33.360 318.220 33.620 ;
        RECT 828.560 33.360 828.820 33.620 ;
      LAYER met2 ;
        RECT 828.620 33.650 828.760 54.000 ;
        RECT 317.960 33.330 318.220 33.650 ;
        RECT 828.560 33.330 828.820 33.650 ;
        RECT 318.020 2.400 318.160 33.330 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 335.945 48.365 336.115 54.000 ;
      LAYER met1 ;
        RECT 335.870 48.520 336.190 48.580 ;
        RECT 335.675 48.380 336.190 48.520 ;
        RECT 335.870 48.320 336.190 48.380 ;
      LAYER via ;
        RECT 335.900 48.320 336.160 48.580 ;
      LAYER met2 ;
        RECT 335.900 48.290 336.160 48.610 ;
        RECT 335.960 2.400 336.100 48.290 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 353.350 33.900 353.670 33.960 ;
        RECT 856.130 33.900 856.450 33.960 ;
        RECT 353.350 33.760 856.450 33.900 ;
        RECT 353.350 33.700 353.670 33.760 ;
        RECT 856.130 33.700 856.450 33.760 ;
      LAYER via ;
        RECT 353.380 33.700 353.640 33.960 ;
        RECT 856.160 33.700 856.420 33.960 ;
      LAYER met2 ;
        RECT 856.220 33.990 856.360 54.000 ;
        RECT 353.380 33.670 353.640 33.990 ;
        RECT 856.160 33.670 856.420 33.990 ;
        RECT 353.440 2.400 353.580 33.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.300 17.410 372.440 54.000 ;
        RECT 371.380 17.270 372.440 17.410 ;
        RECT 371.380 2.400 371.520 17.270 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 34.240 389.550 34.300 ;
        RECT 876.830 34.240 877.150 34.300 ;
        RECT 389.230 34.100 877.150 34.240 ;
        RECT 389.230 34.040 389.550 34.100 ;
        RECT 876.830 34.040 877.150 34.100 ;
      LAYER via ;
        RECT 389.260 34.040 389.520 34.300 ;
        RECT 876.860 34.040 877.120 34.300 ;
      LAYER met2 ;
        RECT 876.920 34.330 877.060 54.000 ;
        RECT 389.260 34.010 389.520 34.330 ;
        RECT 876.860 34.010 877.120 34.330 ;
        RECT 389.320 2.400 389.460 34.010 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 15.880 407.490 15.940 ;
        RECT 413.610 15.880 413.930 15.940 ;
        RECT 407.170 15.740 413.930 15.880 ;
        RECT 407.170 15.680 407.490 15.740 ;
        RECT 413.610 15.680 413.930 15.740 ;
      LAYER via ;
        RECT 407.200 15.680 407.460 15.940 ;
        RECT 413.640 15.680 413.900 15.940 ;
      LAYER met2 ;
        RECT 413.700 15.970 413.840 54.000 ;
        RECT 407.200 15.650 407.460 15.970 ;
        RECT 413.640 15.650 413.900 15.970 ;
        RECT 407.260 2.400 407.400 15.650 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.700 17.410 68.840 54.000 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.650 15.540 424.970 15.600 ;
        RECT 427.410 15.540 427.730 15.600 ;
        RECT 424.650 15.400 427.730 15.540 ;
        RECT 424.650 15.340 424.970 15.400 ;
        RECT 427.410 15.340 427.730 15.400 ;
      LAYER via ;
        RECT 424.680 15.340 424.940 15.600 ;
        RECT 427.440 15.340 427.700 15.600 ;
      LAYER met2 ;
        RECT 427.500 15.630 427.640 54.000 ;
        RECT 424.680 15.310 424.940 15.630 ;
        RECT 427.440 15.310 427.700 15.630 ;
        RECT 424.740 2.400 424.880 15.310 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 442.590 15.540 442.910 15.600 ;
        RECT 448.110 15.540 448.430 15.600 ;
        RECT 442.590 15.400 448.430 15.540 ;
        RECT 442.590 15.340 442.910 15.400 ;
        RECT 448.110 15.340 448.430 15.400 ;
      LAYER via ;
        RECT 442.620 15.340 442.880 15.600 ;
        RECT 448.140 15.340 448.400 15.600 ;
      LAYER met2 ;
        RECT 448.200 15.630 448.340 54.000 ;
        RECT 442.620 15.310 442.880 15.630 ;
        RECT 448.140 15.310 448.400 15.630 ;
        RECT 442.680 2.400 442.820 15.310 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.000 17.410 462.140 54.000 ;
        RECT 460.620 17.270 462.140 17.410 ;
        RECT 460.620 2.400 460.760 17.270 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 478.470 14.520 478.790 14.580 ;
        RECT 482.610 14.520 482.930 14.580 ;
        RECT 478.470 14.380 482.930 14.520 ;
        RECT 478.470 14.320 478.790 14.380 ;
        RECT 482.610 14.320 482.930 14.380 ;
      LAYER via ;
        RECT 478.500 14.320 478.760 14.580 ;
        RECT 482.640 14.320 482.900 14.580 ;
      LAYER met2 ;
        RECT 482.700 14.610 482.840 54.000 ;
        RECT 478.500 14.290 478.760 14.610 ;
        RECT 482.640 14.290 482.900 14.610 ;
        RECT 478.560 2.400 478.700 14.290 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.040 17.410 496.180 54.000 ;
        RECT 496.040 17.270 496.640 17.410 ;
        RECT 496.500 2.400 496.640 17.270 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 14.520 514.210 14.580 ;
        RECT 517.110 14.520 517.430 14.580 ;
        RECT 513.890 14.380 517.430 14.520 ;
        RECT 513.890 14.320 514.210 14.380 ;
        RECT 517.110 14.320 517.430 14.380 ;
      LAYER via ;
        RECT 513.920 14.320 514.180 14.580 ;
        RECT 517.140 14.320 517.400 14.580 ;
      LAYER met2 ;
        RECT 517.200 14.610 517.340 54.000 ;
        RECT 513.920 14.290 514.180 14.610 ;
        RECT 517.140 14.290 517.400 14.610 ;
        RECT 513.980 2.400 514.120 14.290 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 531.830 14.520 532.150 14.580 ;
        RECT 537.810 14.520 538.130 14.580 ;
        RECT 531.830 14.380 538.130 14.520 ;
        RECT 531.830 14.320 532.150 14.380 ;
        RECT 537.810 14.320 538.130 14.380 ;
      LAYER via ;
        RECT 531.860 14.320 532.120 14.580 ;
        RECT 537.840 14.320 538.100 14.580 ;
      LAYER met2 ;
        RECT 537.900 14.610 538.040 54.000 ;
        RECT 531.860 14.290 532.120 14.610 ;
        RECT 537.840 14.290 538.100 14.610 ;
        RECT 531.920 2.400 532.060 14.290 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.700 16.730 551.840 54.000 ;
        RECT 549.860 16.590 551.840 16.730 ;
        RECT 549.860 2.400 550.000 16.590 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 17.920 568.030 17.980 ;
        RECT 572.310 17.920 572.630 17.980 ;
        RECT 567.710 17.780 572.630 17.920 ;
        RECT 567.710 17.720 568.030 17.780 ;
        RECT 572.310 17.720 572.630 17.780 ;
      LAYER via ;
        RECT 567.740 17.720 568.000 17.980 ;
        RECT 572.340 17.720 572.600 17.980 ;
      LAYER met2 ;
        RECT 572.400 18.010 572.540 54.000 ;
        RECT 567.740 17.690 568.000 18.010 ;
        RECT 572.340 17.690 572.600 18.010 ;
        RECT 567.800 2.400 567.940 17.690 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.740 2.400 585.880 54.000 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 44.780 91.930 44.840 ;
        RECT 662.930 44.780 663.250 44.840 ;
        RECT 91.610 44.640 663.250 44.780 ;
        RECT 91.610 44.580 91.930 44.640 ;
        RECT 662.930 44.580 663.250 44.640 ;
      LAYER via ;
        RECT 91.640 44.580 91.900 44.840 ;
        RECT 662.960 44.580 663.220 44.840 ;
      LAYER met2 ;
        RECT 663.020 44.870 663.160 54.000 ;
        RECT 91.640 44.550 91.900 44.870 ;
        RECT 662.960 44.550 663.220 44.870 ;
        RECT 91.700 2.400 91.840 44.550 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 18.600 603.450 18.660 ;
        RECT 606.810 18.600 607.130 18.660 ;
        RECT 603.130 18.460 607.130 18.600 ;
        RECT 603.130 18.400 603.450 18.460 ;
        RECT 606.810 18.400 607.130 18.460 ;
      LAYER via ;
        RECT 603.160 18.400 603.420 18.660 ;
        RECT 606.840 18.400 607.100 18.660 ;
      LAYER met2 ;
        RECT 606.900 18.690 607.040 54.000 ;
        RECT 603.160 18.370 603.420 18.690 ;
        RECT 606.840 18.370 607.100 18.690 ;
        RECT 603.220 2.400 603.360 18.370 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 18.600 621.390 18.660 ;
        RECT 627.050 18.600 627.370 18.660 ;
        RECT 621.070 18.460 627.370 18.600 ;
        RECT 621.070 18.400 621.390 18.460 ;
        RECT 627.050 18.400 627.370 18.460 ;
      LAYER via ;
        RECT 621.100 18.400 621.360 18.660 ;
        RECT 627.080 18.400 627.340 18.660 ;
      LAYER met2 ;
        RECT 627.140 18.690 627.280 54.000 ;
        RECT 621.100 18.370 621.360 18.690 ;
        RECT 627.080 18.370 627.340 18.690 ;
        RECT 621.160 2.400 621.300 18.370 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 677.190 17.580 677.510 17.640 ;
        RECT 649.680 17.440 677.510 17.580 ;
        RECT 115.530 17.240 115.850 17.300 ;
        RECT 649.680 17.240 649.820 17.440 ;
        RECT 677.190 17.380 677.510 17.440 ;
        RECT 115.530 17.100 649.820 17.240 ;
        RECT 115.530 17.040 115.850 17.100 ;
      LAYER via ;
        RECT 115.560 17.040 115.820 17.300 ;
        RECT 677.220 17.380 677.480 17.640 ;
      LAYER met2 ;
        RECT 677.280 17.670 677.420 54.000 ;
        RECT 677.220 17.350 677.480 17.670 ;
        RECT 115.560 17.010 115.820 17.330 ;
        RECT 115.620 2.400 115.760 17.010 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 665.765 18.105 665.935 19.295 ;
      LAYER mcon ;
        RECT 665.765 19.125 665.935 19.295 ;
      LAYER met1 ;
        RECT 665.705 19.280 665.995 19.325 ;
        RECT 665.705 19.140 693.520 19.280 ;
        RECT 665.705 19.095 665.995 19.140 ;
        RECT 693.380 18.940 693.520 19.140 ;
        RECT 696.970 18.940 697.290 19.000 ;
        RECT 693.380 18.800 697.290 18.940 ;
        RECT 696.970 18.740 697.290 18.800 ;
        RECT 139.450 18.260 139.770 18.320 ;
        RECT 665.705 18.260 665.995 18.305 ;
        RECT 139.450 18.120 665.995 18.260 ;
        RECT 139.450 18.060 139.770 18.120 ;
        RECT 665.705 18.075 665.995 18.120 ;
      LAYER via ;
        RECT 697.000 18.740 697.260 19.000 ;
        RECT 139.480 18.060 139.740 18.320 ;
      LAYER met2 ;
        RECT 697.060 19.030 697.200 54.000 ;
        RECT 697.000 18.710 697.260 19.030 ;
        RECT 139.480 18.030 139.740 18.350 ;
        RECT 139.540 2.400 139.680 18.030 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 157.390 37.980 157.710 38.040 ;
        RECT 711.230 37.980 711.550 38.040 ;
        RECT 157.390 37.840 711.550 37.980 ;
        RECT 157.390 37.780 157.710 37.840 ;
        RECT 711.230 37.780 711.550 37.840 ;
      LAYER via ;
        RECT 157.420 37.780 157.680 38.040 ;
        RECT 711.260 37.780 711.520 38.040 ;
      LAYER met2 ;
        RECT 711.320 38.070 711.460 54.000 ;
        RECT 157.420 37.750 157.680 38.070 ;
        RECT 711.260 37.750 711.520 38.070 ;
        RECT 157.480 2.400 157.620 37.750 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 692.905 17.425 693.075 18.955 ;
      LAYER mcon ;
        RECT 692.905 18.785 693.075 18.955 ;
      LAYER met1 ;
        RECT 174.870 18.940 175.190 19.000 ;
        RECT 692.845 18.940 693.135 18.985 ;
        RECT 174.870 18.800 693.135 18.940 ;
        RECT 174.870 18.740 175.190 18.800 ;
        RECT 692.845 18.755 693.135 18.800 ;
        RECT 692.845 17.580 693.135 17.625 ;
        RECT 725.030 17.580 725.350 17.640 ;
        RECT 692.845 17.440 725.350 17.580 ;
        RECT 692.845 17.395 693.135 17.440 ;
        RECT 725.030 17.380 725.350 17.440 ;
      LAYER via ;
        RECT 174.900 18.740 175.160 19.000 ;
        RECT 725.060 17.380 725.320 17.640 ;
      LAYER met2 ;
        RECT 174.900 18.710 175.160 19.030 ;
        RECT 174.960 2.400 175.100 18.710 ;
        RECT 725.120 17.670 725.260 54.000 ;
        RECT 725.060 17.350 725.320 17.670 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.900 2.400 193.040 54.000 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 210.750 19.620 211.070 19.680 ;
        RECT 745.270 19.620 745.590 19.680 ;
        RECT 210.750 19.480 745.590 19.620 ;
        RECT 210.750 19.420 211.070 19.480 ;
        RECT 745.270 19.420 745.590 19.480 ;
      LAYER via ;
        RECT 210.780 19.420 211.040 19.680 ;
        RECT 745.300 19.420 745.560 19.680 ;
      LAYER met2 ;
        RECT 745.360 19.710 745.500 54.000 ;
        RECT 210.780 19.390 211.040 19.710 ;
        RECT 745.300 19.390 745.560 19.710 ;
        RECT 210.840 2.400 210.980 19.390 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 228.690 16.900 229.010 16.960 ;
        RECT 234.210 16.900 234.530 16.960 ;
        RECT 228.690 16.760 234.530 16.900 ;
        RECT 228.690 16.700 229.010 16.760 ;
        RECT 234.210 16.700 234.530 16.760 ;
      LAYER via ;
        RECT 228.720 16.700 228.980 16.960 ;
        RECT 234.240 16.700 234.500 16.960 ;
      LAYER met2 ;
        RECT 234.300 16.990 234.440 54.000 ;
        RECT 228.720 16.670 228.980 16.990 ;
        RECT 234.240 16.670 234.500 16.990 ;
        RECT 228.780 2.400 228.920 16.670 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 18.260 50.530 18.320 ;
        RECT 127.490 18.260 127.810 18.320 ;
        RECT 50.210 18.120 127.810 18.260 ;
        RECT 50.210 18.060 50.530 18.120 ;
        RECT 127.490 18.060 127.810 18.120 ;
      LAYER via ;
        RECT 50.240 18.060 50.500 18.320 ;
        RECT 127.520 18.060 127.780 18.320 ;
      LAYER met2 ;
        RECT 127.580 18.350 127.720 54.000 ;
        RECT 50.240 18.030 50.500 18.350 ;
        RECT 127.520 18.030 127.780 18.350 ;
        RECT 50.300 2.400 50.440 18.030 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 300.525 16.065 300.695 20.655 ;
      LAYER mcon ;
        RECT 300.525 20.485 300.695 20.655 ;
      LAYER met1 ;
        RECT 300.465 20.640 300.755 20.685 ;
        RECT 300.465 20.500 698.120 20.640 ;
        RECT 300.465 20.455 300.755 20.500 ;
        RECT 697.980 20.300 698.120 20.500 ;
        RECT 762.290 20.300 762.610 20.360 ;
        RECT 697.980 20.160 762.610 20.300 ;
        RECT 762.290 20.100 762.610 20.160 ;
        RECT 252.610 16.560 252.930 16.620 ;
        RECT 252.610 16.420 293.780 16.560 ;
        RECT 252.610 16.360 252.930 16.420 ;
        RECT 293.640 16.220 293.780 16.420 ;
        RECT 300.465 16.220 300.755 16.265 ;
        RECT 293.640 16.080 300.755 16.220 ;
        RECT 300.465 16.035 300.755 16.080 ;
      LAYER via ;
        RECT 762.320 20.100 762.580 20.360 ;
        RECT 252.640 16.360 252.900 16.620 ;
      LAYER met2 ;
        RECT 762.380 20.390 762.520 54.000 ;
        RECT 762.320 20.070 762.580 20.390 ;
        RECT 252.640 16.330 252.900 16.650 ;
        RECT 252.700 2.400 252.840 16.330 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 16.900 270.410 16.960 ;
        RECT 782.990 16.900 783.310 16.960 ;
        RECT 270.090 16.760 783.310 16.900 ;
        RECT 270.090 16.700 270.410 16.760 ;
        RECT 782.990 16.700 783.310 16.760 ;
      LAYER via ;
        RECT 270.120 16.700 270.380 16.960 ;
        RECT 783.020 16.700 783.280 16.960 ;
      LAYER met2 ;
        RECT 783.080 16.990 783.220 54.000 ;
        RECT 270.120 16.670 270.380 16.990 ;
        RECT 783.020 16.670 783.280 16.990 ;
        RECT 270.180 2.400 270.320 16.670 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 20.640 288.350 20.700 ;
        RECT 299.990 20.640 300.310 20.700 ;
        RECT 288.030 20.500 300.310 20.640 ;
        RECT 288.030 20.440 288.350 20.500 ;
        RECT 299.990 20.440 300.310 20.500 ;
      LAYER via ;
        RECT 288.060 20.440 288.320 20.700 ;
        RECT 300.020 20.440 300.280 20.700 ;
      LAYER met2 ;
        RECT 300.080 20.730 300.220 54.000 ;
        RECT 288.060 20.410 288.320 20.730 ;
        RECT 300.020 20.410 300.280 20.730 ;
        RECT 288.120 2.400 288.260 20.410 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 16.560 306.290 16.620 ;
        RECT 796.790 16.560 797.110 16.620 ;
        RECT 305.970 16.420 797.110 16.560 ;
        RECT 305.970 16.360 306.290 16.420 ;
        RECT 796.790 16.360 797.110 16.420 ;
      LAYER via ;
        RECT 306.000 16.360 306.260 16.620 ;
        RECT 796.820 16.360 797.080 16.620 ;
      LAYER met2 ;
        RECT 796.880 16.650 797.020 54.000 ;
        RECT 306.000 16.330 306.260 16.650 ;
        RECT 796.820 16.330 797.080 16.650 ;
        RECT 306.060 2.400 306.200 16.330 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 19.280 324.230 19.340 ;
        RECT 334.490 19.280 334.810 19.340 ;
        RECT 323.910 19.140 334.810 19.280 ;
        RECT 323.910 19.080 324.230 19.140 ;
        RECT 334.490 19.080 334.810 19.140 ;
      LAYER via ;
        RECT 323.940 19.080 324.200 19.340 ;
        RECT 334.520 19.080 334.780 19.340 ;
      LAYER met2 ;
        RECT 334.580 19.370 334.720 54.000 ;
        RECT 323.940 19.050 324.200 19.370 ;
        RECT 334.520 19.050 334.780 19.370 ;
        RECT 324.000 2.400 324.140 19.050 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 16.220 341.710 16.280 ;
        RECT 810.590 16.220 810.910 16.280 ;
        RECT 341.390 16.080 810.910 16.220 ;
        RECT 341.390 16.020 341.710 16.080 ;
        RECT 810.590 16.020 810.910 16.080 ;
      LAYER via ;
        RECT 341.420 16.020 341.680 16.280 ;
        RECT 810.620 16.020 810.880 16.280 ;
      LAYER met2 ;
        RECT 810.680 16.310 810.820 54.000 ;
        RECT 341.420 15.990 341.680 16.310 ;
        RECT 810.620 15.990 810.880 16.310 ;
        RECT 341.480 2.400 341.620 15.990 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 14.860 359.650 14.920 ;
        RECT 375.890 14.860 376.210 14.920 ;
        RECT 359.330 14.720 376.210 14.860 ;
        RECT 359.330 14.660 359.650 14.720 ;
        RECT 375.890 14.660 376.210 14.720 ;
      LAYER via ;
        RECT 359.360 14.660 359.620 14.920 ;
        RECT 375.920 14.660 376.180 14.920 ;
      LAYER met2 ;
        RECT 375.980 14.950 376.120 54.000 ;
        RECT 359.360 14.630 359.620 14.950 ;
        RECT 375.920 14.630 376.180 14.950 ;
        RECT 359.420 2.400 359.560 14.630 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.030 15.880 817.350 15.940 ;
        RECT 414.160 15.740 817.350 15.880 ;
        RECT 414.160 15.540 414.300 15.740 ;
        RECT 817.030 15.680 817.350 15.740 ;
        RECT 411.400 15.400 414.300 15.540 ;
        RECT 377.270 15.200 377.590 15.260 ;
        RECT 411.400 15.200 411.540 15.400 ;
        RECT 377.270 15.060 411.540 15.200 ;
        RECT 377.270 15.000 377.590 15.060 ;
      LAYER via ;
        RECT 817.060 15.680 817.320 15.940 ;
        RECT 377.300 15.000 377.560 15.260 ;
      LAYER met2 ;
        RECT 817.580 38.490 817.720 54.000 ;
        RECT 817.120 38.350 817.720 38.490 ;
        RECT 817.120 15.970 817.260 38.350 ;
        RECT 817.060 15.650 817.320 15.970 ;
        RECT 377.300 14.970 377.560 15.290 ;
        RECT 377.360 2.400 377.500 14.970 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 15.540 395.530 15.600 ;
        RECT 410.390 15.540 410.710 15.600 ;
        RECT 395.210 15.400 410.710 15.540 ;
        RECT 395.210 15.340 395.530 15.400 ;
        RECT 410.390 15.340 410.710 15.400 ;
      LAYER via ;
        RECT 395.240 15.340 395.500 15.600 ;
        RECT 410.420 15.340 410.680 15.600 ;
      LAYER met2 ;
        RECT 410.480 15.630 410.620 54.000 ;
        RECT 395.240 15.310 395.500 15.630 ;
        RECT 410.420 15.310 410.680 15.630 ;
        RECT 395.300 2.400 395.440 15.310 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 824.390 15.540 824.710 15.600 ;
        RECT 448.660 15.400 824.710 15.540 ;
        RECT 413.150 15.200 413.470 15.260 ;
        RECT 448.660 15.200 448.800 15.400 ;
        RECT 824.390 15.340 824.710 15.400 ;
        RECT 413.150 15.060 448.800 15.200 ;
        RECT 413.150 15.000 413.470 15.060 ;
      LAYER via ;
        RECT 413.180 15.000 413.440 15.260 ;
        RECT 824.420 15.340 824.680 15.600 ;
      LAYER met2 ;
        RECT 824.480 15.630 824.620 54.000 ;
        RECT 824.420 15.310 824.680 15.630 ;
        RECT 413.180 14.970 413.440 15.290 ;
        RECT 413.240 2.400 413.380 14.970 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 74.130 18.600 74.450 18.660 ;
        RECT 141.290 18.600 141.610 18.660 ;
        RECT 74.130 18.460 141.610 18.600 ;
        RECT 74.130 18.400 74.450 18.460 ;
        RECT 141.290 18.400 141.610 18.460 ;
      LAYER via ;
        RECT 74.160 18.400 74.420 18.660 ;
        RECT 141.320 18.400 141.580 18.660 ;
      LAYER met2 ;
        RECT 141.380 18.690 141.520 54.000 ;
        RECT 74.160 18.370 74.420 18.690 ;
        RECT 141.320 18.370 141.580 18.690 ;
        RECT 74.220 2.400 74.360 18.370 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 831.290 15.200 831.610 15.260 ;
        RECT 449.120 15.060 831.610 15.200 ;
        RECT 430.630 14.860 430.950 14.920 ;
        RECT 449.120 14.860 449.260 15.060 ;
        RECT 831.290 15.000 831.610 15.060 ;
        RECT 430.630 14.720 449.260 14.860 ;
        RECT 430.630 14.660 430.950 14.720 ;
      LAYER via ;
        RECT 430.660 14.660 430.920 14.920 ;
        RECT 831.320 15.000 831.580 15.260 ;
      LAYER met2 ;
        RECT 831.380 15.290 831.520 54.000 ;
        RECT 831.320 14.970 831.580 15.290 ;
        RECT 430.660 14.630 430.920 14.950 ;
        RECT 430.720 2.400 430.860 14.630 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 14.180 448.890 14.240 ;
        RECT 477.090 14.180 477.410 14.240 ;
        RECT 448.570 14.040 477.410 14.180 ;
        RECT 448.570 13.980 448.890 14.040 ;
        RECT 477.090 13.980 477.410 14.040 ;
      LAYER via ;
        RECT 448.600 13.980 448.860 14.240 ;
        RECT 477.120 13.980 477.380 14.240 ;
      LAYER met2 ;
        RECT 479.480 15.370 479.620 54.000 ;
        RECT 478.100 15.230 479.620 15.370 ;
        RECT 448.600 13.950 448.860 14.270 ;
        RECT 477.120 14.010 477.380 14.270 ;
        RECT 478.100 14.010 478.240 15.230 ;
        RECT 477.120 13.950 478.240 14.010 ;
        RECT 448.660 2.400 448.800 13.950 ;
        RECT 477.180 13.870 478.240 13.950 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 14.860 466.830 14.920 ;
        RECT 845.550 14.860 845.870 14.920 ;
        RECT 466.510 14.720 845.870 14.860 ;
        RECT 466.510 14.660 466.830 14.720 ;
        RECT 845.550 14.660 845.870 14.720 ;
      LAYER via ;
        RECT 466.540 14.660 466.800 14.920 ;
        RECT 845.580 14.660 845.840 14.920 ;
      LAYER met2 ;
        RECT 845.640 14.950 845.780 54.000 ;
        RECT 466.540 14.630 466.800 14.950 ;
        RECT 845.580 14.630 845.840 14.950 ;
        RECT 466.600 2.400 466.740 14.630 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 14.520 484.770 14.580 ;
        RECT 513.430 14.520 513.750 14.580 ;
        RECT 484.450 14.380 513.750 14.520 ;
        RECT 484.450 14.320 484.770 14.380 ;
        RECT 513.430 14.320 513.750 14.380 ;
      LAYER via ;
        RECT 484.480 14.320 484.740 14.580 ;
        RECT 513.460 14.320 513.720 14.580 ;
      LAYER met2 ;
        RECT 513.980 15.370 514.120 54.000 ;
        RECT 513.520 15.230 514.120 15.370 ;
        RECT 513.520 14.610 513.660 15.230 ;
        RECT 484.480 14.290 484.740 14.610 ;
        RECT 513.460 14.290 513.720 14.610 ;
        RECT 484.540 2.400 484.680 14.290 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 554.905 14.025 556.455 14.195 ;
      LAYER mcon ;
        RECT 556.285 14.025 556.455 14.195 ;
      LAYER met1 ;
        RECT 845.090 14.520 845.410 14.580 ;
        RECT 559.060 14.380 845.410 14.520 ;
        RECT 502.390 14.180 502.710 14.240 ;
        RECT 554.845 14.180 555.135 14.225 ;
        RECT 502.390 14.040 555.135 14.180 ;
        RECT 502.390 13.980 502.710 14.040 ;
        RECT 554.845 13.995 555.135 14.040 ;
        RECT 556.225 14.180 556.515 14.225 ;
        RECT 559.060 14.180 559.200 14.380 ;
        RECT 845.090 14.320 845.410 14.380 ;
        RECT 556.225 14.040 559.200 14.180 ;
        RECT 556.225 13.995 556.515 14.040 ;
      LAYER via ;
        RECT 502.420 13.980 502.680 14.240 ;
        RECT 845.120 14.320 845.380 14.580 ;
      LAYER met2 ;
        RECT 845.180 14.610 845.320 54.000 ;
        RECT 845.120 14.290 845.380 14.610 ;
        RECT 502.420 13.950 502.680 14.270 ;
        RECT 502.480 2.400 502.620 13.950 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 14.520 520.190 14.580 ;
        RECT 527.690 14.520 528.010 14.580 ;
        RECT 519.870 14.380 528.010 14.520 ;
        RECT 519.870 14.320 520.190 14.380 ;
        RECT 527.690 14.320 528.010 14.380 ;
      LAYER via ;
        RECT 519.900 14.320 520.160 14.580 ;
        RECT 527.720 14.320 527.980 14.580 ;
      LAYER met2 ;
        RECT 527.780 14.610 527.920 54.000 ;
        RECT 519.900 14.290 520.160 14.610 ;
        RECT 527.720 14.290 527.980 14.610 ;
        RECT 519.960 2.400 520.100 14.290 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 538.270 14.520 538.590 14.580 ;
        RECT 538.270 14.380 555.520 14.520 ;
        RECT 538.270 14.320 538.590 14.380 ;
        RECT 555.380 13.840 555.520 14.380 ;
        RECT 857.970 14.180 858.290 14.240 ;
        RECT 559.520 14.040 858.290 14.180 ;
        RECT 559.520 13.840 559.660 14.040 ;
        RECT 857.970 13.980 858.290 14.040 ;
        RECT 555.380 13.700 559.660 13.840 ;
      LAYER via ;
        RECT 538.300 14.320 538.560 14.580 ;
        RECT 858.000 13.980 858.260 14.240 ;
      LAYER met2 ;
        RECT 538.300 14.290 538.560 14.610 ;
        RECT 538.360 14.010 538.500 14.290 ;
        RECT 858.060 14.270 858.200 54.000 ;
        RECT 537.900 13.870 538.500 14.010 ;
        RECT 858.000 13.950 858.260 14.270 ;
        RECT 537.900 2.400 538.040 13.870 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 14.520 556.070 14.580 ;
        RECT 558.510 14.520 558.830 14.580 ;
        RECT 555.750 14.380 558.830 14.520 ;
        RECT 555.750 14.320 556.070 14.380 ;
        RECT 558.510 14.320 558.830 14.380 ;
      LAYER via ;
        RECT 555.780 14.320 556.040 14.580 ;
        RECT 558.540 14.320 558.800 14.580 ;
      LAYER met2 ;
        RECT 558.600 14.610 558.740 54.000 ;
        RECT 555.780 14.290 556.040 14.610 ;
        RECT 558.540 14.290 558.800 14.610 ;
        RECT 555.840 2.400 555.980 14.290 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 17.920 574.010 17.980 ;
        RECT 579.210 17.920 579.530 17.980 ;
        RECT 573.690 17.780 579.530 17.920 ;
        RECT 573.690 17.720 574.010 17.780 ;
        RECT 579.210 17.720 579.530 17.780 ;
      LAYER via ;
        RECT 573.720 17.720 573.980 17.980 ;
        RECT 579.240 17.720 579.500 17.980 ;
      LAYER met2 ;
        RECT 579.300 18.010 579.440 54.000 ;
        RECT 573.720 17.690 573.980 18.010 ;
        RECT 579.240 17.690 579.500 18.010 ;
        RECT 573.780 2.400 573.920 17.690 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 17.920 591.490 17.980 ;
        RECT 865.790 17.920 866.110 17.980 ;
        RECT 591.170 17.780 866.110 17.920 ;
        RECT 591.170 17.720 591.490 17.780 ;
        RECT 865.790 17.720 866.110 17.780 ;
      LAYER via ;
        RECT 591.200 17.720 591.460 17.980 ;
        RECT 865.820 17.720 866.080 17.980 ;
      LAYER met2 ;
        RECT 865.880 18.010 866.020 54.000 ;
        RECT 591.200 17.690 591.460 18.010 ;
        RECT 865.820 17.690 866.080 18.010 ;
        RECT 591.260 2.400 591.400 17.690 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 20.300 97.910 20.360 ;
        RECT 230.990 20.300 231.310 20.360 ;
        RECT 97.590 20.160 231.310 20.300 ;
        RECT 97.590 20.100 97.910 20.160 ;
        RECT 230.990 20.100 231.310 20.160 ;
      LAYER via ;
        RECT 97.620 20.100 97.880 20.360 ;
        RECT 231.020 20.100 231.280 20.360 ;
      LAYER met2 ;
        RECT 231.080 20.390 231.220 54.000 ;
        RECT 97.620 20.070 97.880 20.390 ;
        RECT 231.020 20.070 231.280 20.390 ;
        RECT 97.680 2.400 97.820 20.070 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 18.600 609.430 18.660 ;
        RECT 613.710 18.600 614.030 18.660 ;
        RECT 609.110 18.460 614.030 18.600 ;
        RECT 609.110 18.400 609.430 18.460 ;
        RECT 613.710 18.400 614.030 18.460 ;
      LAYER via ;
        RECT 609.140 18.400 609.400 18.660 ;
        RECT 613.740 18.400 614.000 18.660 ;
      LAYER met2 ;
        RECT 613.800 18.690 613.940 54.000 ;
        RECT 609.140 18.370 609.400 18.690 ;
        RECT 613.740 18.370 614.000 18.690 ;
        RECT 609.200 2.400 609.340 18.370 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.600 18.090 627.740 54.000 ;
        RECT 627.140 17.950 627.740 18.090 ;
        RECT 627.140 2.400 627.280 17.950 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 666.150 18.260 666.470 18.320 ;
        RECT 683.170 18.260 683.490 18.320 ;
        RECT 666.150 18.120 683.490 18.260 ;
        RECT 666.150 18.060 666.470 18.120 ;
        RECT 683.170 18.060 683.490 18.120 ;
        RECT 121.510 17.580 121.830 17.640 ;
        RECT 649.130 17.580 649.450 17.640 ;
        RECT 121.510 17.440 649.450 17.580 ;
        RECT 121.510 17.380 121.830 17.440 ;
        RECT 649.130 17.380 649.450 17.440 ;
      LAYER via ;
        RECT 666.180 18.060 666.440 18.320 ;
        RECT 683.200 18.060 683.460 18.320 ;
        RECT 121.540 17.380 121.800 17.640 ;
        RECT 649.160 17.380 649.420 17.640 ;
      LAYER met2 ;
        RECT 683.260 18.350 683.400 54.000 ;
        RECT 666.180 18.205 666.440 18.350 ;
        RECT 649.150 17.835 649.430 18.205 ;
        RECT 666.170 17.835 666.450 18.205 ;
        RECT 683.200 18.030 683.460 18.350 ;
        RECT 649.220 17.670 649.360 17.835 ;
        RECT 121.540 17.350 121.800 17.670 ;
        RECT 649.160 17.350 649.420 17.670 ;
        RECT 121.600 2.400 121.740 17.350 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 649.150 17.880 649.430 18.160 ;
        RECT 666.170 17.880 666.450 18.160 ;
      LAYER met3 ;
        RECT 649.125 18.170 649.455 18.185 ;
        RECT 666.145 18.170 666.475 18.185 ;
        RECT 649.125 17.870 666.475 18.170 ;
        RECT 649.125 17.855 649.455 17.870 ;
        RECT 666.145 17.855 666.475 17.870 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 179.545 18.445 179.715 20.655 ;
        RECT 276.145 14.705 276.315 18.615 ;
        RECT 311.565 14.705 311.735 18.615 ;
        RECT 372.745 15.045 372.915 18.615 ;
        RECT 420.585 14.705 420.755 18.615 ;
        RECT 469.345 14.365 469.515 18.615 ;
        RECT 517.185 13.685 517.355 18.615 ;
        RECT 565.945 18.445 566.115 20.995 ;
        RECT 627.585 18.445 627.755 20.995 ;
        RECT 650.125 17.085 650.295 18.615 ;
      LAYER mcon ;
        RECT 565.945 20.825 566.115 20.995 ;
        RECT 179.545 20.485 179.715 20.655 ;
        RECT 276.145 18.445 276.315 18.615 ;
        RECT 311.565 18.445 311.735 18.615 ;
        RECT 372.745 18.445 372.915 18.615 ;
        RECT 420.585 18.445 420.755 18.615 ;
        RECT 469.345 18.445 469.515 18.615 ;
        RECT 517.185 18.445 517.355 18.615 ;
        RECT 627.585 20.825 627.755 20.995 ;
        RECT 650.125 18.445 650.295 18.615 ;
      LAYER met1 ;
        RECT 565.885 20.980 566.175 21.025 ;
        RECT 627.525 20.980 627.815 21.025 ;
        RECT 565.885 20.840 627.815 20.980 ;
        RECT 565.885 20.795 566.175 20.840 ;
        RECT 627.525 20.795 627.815 20.840 ;
        RECT 179.485 20.640 179.775 20.685 ;
        RECT 227.310 20.640 227.630 20.700 ;
        RECT 179.485 20.500 227.630 20.640 ;
        RECT 179.485 20.455 179.775 20.500 ;
        RECT 227.310 20.440 227.630 20.500 ;
        RECT 145.430 18.600 145.750 18.660 ;
        RECT 179.485 18.600 179.775 18.645 ;
        RECT 145.430 18.460 179.775 18.600 ;
        RECT 145.430 18.400 145.750 18.460 ;
        RECT 179.485 18.415 179.775 18.460 ;
        RECT 227.310 18.600 227.630 18.660 ;
        RECT 276.085 18.600 276.375 18.645 ;
        RECT 227.310 18.460 276.375 18.600 ;
        RECT 227.310 18.400 227.630 18.460 ;
        RECT 276.085 18.415 276.375 18.460 ;
        RECT 311.505 18.600 311.795 18.645 ;
        RECT 372.685 18.600 372.975 18.645 ;
        RECT 311.505 18.460 372.975 18.600 ;
        RECT 311.505 18.415 311.795 18.460 ;
        RECT 372.685 18.415 372.975 18.460 ;
        RECT 420.525 18.600 420.815 18.645 ;
        RECT 469.285 18.600 469.575 18.645 ;
        RECT 420.525 18.460 469.575 18.600 ;
        RECT 420.525 18.415 420.815 18.460 ;
        RECT 469.285 18.415 469.575 18.460 ;
        RECT 517.125 18.600 517.415 18.645 ;
        RECT 565.885 18.600 566.175 18.645 ;
        RECT 517.125 18.460 566.175 18.600 ;
        RECT 517.125 18.415 517.415 18.460 ;
        RECT 565.885 18.415 566.175 18.460 ;
        RECT 627.525 18.600 627.815 18.645 ;
        RECT 650.065 18.600 650.355 18.645 ;
        RECT 627.525 18.460 650.355 18.600 ;
        RECT 627.525 18.415 627.815 18.460 ;
        RECT 650.065 18.415 650.355 18.460 ;
        RECT 650.065 17.240 650.355 17.285 ;
        RECT 703.870 17.240 704.190 17.300 ;
        RECT 650.065 17.100 704.190 17.240 ;
        RECT 650.065 17.055 650.355 17.100 ;
        RECT 703.870 17.040 704.190 17.100 ;
        RECT 372.685 15.200 372.975 15.245 ;
        RECT 372.685 15.060 376.580 15.200 ;
        RECT 372.685 15.015 372.975 15.060 ;
        RECT 276.085 14.860 276.375 14.905 ;
        RECT 311.505 14.860 311.795 14.905 ;
        RECT 276.085 14.720 311.795 14.860 ;
        RECT 376.440 14.860 376.580 15.060 ;
        RECT 420.525 14.860 420.815 14.905 ;
        RECT 376.440 14.720 420.815 14.860 ;
        RECT 276.085 14.675 276.375 14.720 ;
        RECT 311.505 14.675 311.795 14.720 ;
        RECT 420.525 14.675 420.815 14.720 ;
        RECT 469.285 14.520 469.575 14.565 ;
        RECT 469.285 14.380 478.240 14.520 ;
        RECT 469.285 14.335 469.575 14.380 ;
        RECT 478.100 13.840 478.240 14.380 ;
        RECT 479.940 14.040 502.160 14.180 ;
        RECT 479.940 13.840 480.080 14.040 ;
        RECT 478.100 13.700 480.080 13.840 ;
        RECT 502.020 13.840 502.160 14.040 ;
        RECT 517.125 13.840 517.415 13.885 ;
        RECT 502.020 13.700 517.415 13.840 ;
        RECT 517.125 13.655 517.415 13.700 ;
      LAYER via ;
        RECT 227.340 20.440 227.600 20.700 ;
        RECT 145.460 18.400 145.720 18.660 ;
        RECT 227.340 18.400 227.600 18.660 ;
        RECT 703.900 17.040 704.160 17.300 ;
      LAYER met2 ;
        RECT 227.340 20.410 227.600 20.730 ;
        RECT 227.400 18.690 227.540 20.410 ;
        RECT 145.460 18.370 145.720 18.690 ;
        RECT 227.340 18.370 227.600 18.690 ;
        RECT 145.520 2.400 145.660 18.370 ;
        RECT 703.960 17.330 704.100 54.000 ;
        RECT 703.900 17.010 704.160 17.330 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 228.305 16.745 228.475 20.655 ;
      LAYER mcon ;
        RECT 228.305 20.485 228.475 20.655 ;
      LAYER met1 ;
        RECT 228.245 20.640 228.535 20.685 ;
        RECT 251.690 20.640 252.010 20.700 ;
        RECT 228.245 20.500 252.010 20.640 ;
        RECT 228.245 20.455 228.535 20.500 ;
        RECT 251.690 20.440 252.010 20.500 ;
        RECT 163.370 16.900 163.690 16.960 ;
        RECT 228.245 16.900 228.535 16.945 ;
        RECT 163.370 16.760 228.535 16.900 ;
        RECT 163.370 16.700 163.690 16.760 ;
        RECT 228.245 16.715 228.535 16.760 ;
      LAYER via ;
        RECT 251.720 20.440 251.980 20.700 ;
        RECT 163.400 16.700 163.660 16.960 ;
      LAYER met2 ;
        RECT 251.780 20.730 251.920 54.000 ;
        RECT 251.720 20.410 251.980 20.730 ;
        RECT 163.400 16.670 163.660 16.990 ;
        RECT 163.460 2.400 163.600 16.670 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 276.145 19.125 276.775 19.295 ;
        RECT 276.605 14.365 276.775 19.125 ;
        RECT 335.025 14.365 335.195 19.295 ;
        RECT 372.745 19.125 373.375 19.295 ;
        RECT 373.205 14.365 373.375 19.125 ;
        RECT 420.125 19.125 420.755 19.295 ;
        RECT 469.345 19.125 469.515 20.995 ;
        RECT 517.185 19.125 517.355 20.995 ;
        RECT 420.125 14.365 420.295 19.125 ;
        RECT 650.585 18.445 650.755 19.295 ;
      LAYER mcon ;
        RECT 469.345 20.825 469.515 20.995 ;
        RECT 335.025 19.125 335.195 19.295 ;
        RECT 420.585 19.125 420.755 19.295 ;
        RECT 517.185 20.825 517.355 20.995 ;
        RECT 650.585 19.125 650.755 19.295 ;
      LAYER met1 ;
        RECT 469.285 20.980 469.575 21.025 ;
        RECT 517.125 20.980 517.415 21.025 ;
        RECT 469.285 20.840 517.415 20.980 ;
        RECT 469.285 20.795 469.575 20.840 ;
        RECT 517.125 20.795 517.415 20.840 ;
        RECT 180.850 19.280 181.170 19.340 ;
        RECT 276.085 19.280 276.375 19.325 ;
        RECT 180.850 19.140 276.375 19.280 ;
        RECT 180.850 19.080 181.170 19.140 ;
        RECT 276.085 19.095 276.375 19.140 ;
        RECT 334.965 19.280 335.255 19.325 ;
        RECT 372.685 19.280 372.975 19.325 ;
        RECT 334.965 19.140 372.975 19.280 ;
        RECT 334.965 19.095 335.255 19.140 ;
        RECT 372.685 19.095 372.975 19.140 ;
        RECT 420.525 19.280 420.815 19.325 ;
        RECT 469.285 19.280 469.575 19.325 ;
        RECT 420.525 19.140 469.575 19.280 ;
        RECT 420.525 19.095 420.815 19.140 ;
        RECT 469.285 19.095 469.575 19.140 ;
        RECT 517.125 19.280 517.415 19.325 ;
        RECT 565.870 19.280 566.190 19.340 ;
        RECT 517.125 19.140 566.190 19.280 ;
        RECT 517.125 19.095 517.415 19.140 ;
        RECT 565.870 19.080 566.190 19.140 ;
        RECT 593.470 19.280 593.790 19.340 ;
        RECT 650.525 19.280 650.815 19.325 ;
        RECT 593.470 19.140 650.815 19.280 ;
        RECT 593.470 19.080 593.790 19.140 ;
        RECT 650.525 19.095 650.815 19.140 ;
        RECT 650.525 18.600 650.815 18.645 ;
        RECT 724.570 18.600 724.890 18.660 ;
        RECT 650.525 18.460 724.890 18.600 ;
        RECT 650.525 18.415 650.815 18.460 ;
        RECT 724.570 18.400 724.890 18.460 ;
        RECT 276.545 14.520 276.835 14.565 ;
        RECT 334.965 14.520 335.255 14.565 ;
        RECT 276.545 14.380 335.255 14.520 ;
        RECT 276.545 14.335 276.835 14.380 ;
        RECT 334.965 14.335 335.255 14.380 ;
        RECT 373.145 14.520 373.435 14.565 ;
        RECT 420.065 14.520 420.355 14.565 ;
        RECT 373.145 14.380 420.355 14.520 ;
        RECT 373.145 14.335 373.435 14.380 ;
        RECT 420.065 14.335 420.355 14.380 ;
      LAYER via ;
        RECT 180.880 19.080 181.140 19.340 ;
        RECT 565.900 19.080 566.160 19.340 ;
        RECT 593.500 19.080 593.760 19.340 ;
        RECT 724.600 18.400 724.860 18.660 ;
      LAYER met2 ;
        RECT 180.880 19.050 181.140 19.370 ;
        RECT 565.890 19.195 566.170 19.565 ;
        RECT 593.490 19.195 593.770 19.565 ;
        RECT 565.900 19.050 566.160 19.195 ;
        RECT 593.500 19.050 593.760 19.195 ;
        RECT 180.940 2.400 181.080 19.050 ;
        RECT 724.660 18.690 724.800 54.000 ;
        RECT 724.600 18.370 724.860 18.690 ;
        RECT 180.730 -4.800 181.290 2.400 ;
      LAYER via2 ;
        RECT 565.890 19.240 566.170 19.520 ;
        RECT 593.490 19.240 593.770 19.520 ;
      LAYER met3 ;
        RECT 565.865 19.530 566.195 19.545 ;
        RECT 593.465 19.530 593.795 19.545 ;
        RECT 565.865 19.230 593.795 19.530 ;
        RECT 565.865 19.215 566.195 19.230 ;
        RECT 593.465 19.215 593.795 19.230 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 15.540 199.110 15.600 ;
        RECT 265.490 15.540 265.810 15.600 ;
        RECT 198.790 15.400 265.810 15.540 ;
        RECT 198.790 15.340 199.110 15.400 ;
        RECT 265.490 15.340 265.810 15.400 ;
      LAYER via ;
        RECT 198.820 15.340 199.080 15.600 ;
        RECT 265.520 15.340 265.780 15.600 ;
      LAYER met2 ;
        RECT 265.580 15.630 265.720 54.000 ;
        RECT 198.820 15.310 199.080 15.630 ;
        RECT 265.520 15.310 265.780 15.630 ;
        RECT 198.880 2.400 199.020 15.310 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 19.960 217.050 20.020 ;
        RECT 752.170 19.960 752.490 20.020 ;
        RECT 216.730 19.820 752.490 19.960 ;
        RECT 216.730 19.760 217.050 19.820 ;
        RECT 752.170 19.760 752.490 19.820 ;
      LAYER via ;
        RECT 216.760 19.760 217.020 20.020 ;
        RECT 752.200 19.760 752.460 20.020 ;
      LAYER met2 ;
        RECT 752.260 20.050 752.400 54.000 ;
        RECT 216.760 19.730 217.020 20.050 ;
        RECT 752.200 19.730 752.460 20.050 ;
        RECT 216.820 2.400 216.960 19.730 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 697.505 18.785 697.675 20.315 ;
      LAYER mcon ;
        RECT 697.505 20.145 697.675 20.315 ;
      LAYER met1 ;
        RECT 234.670 20.300 234.990 20.360 ;
        RECT 697.445 20.300 697.735 20.345 ;
        RECT 234.670 20.160 697.735 20.300 ;
        RECT 234.670 20.100 234.990 20.160 ;
        RECT 697.445 20.115 697.735 20.160 ;
        RECT 697.445 18.940 697.735 18.985 ;
        RECT 765.970 18.940 766.290 19.000 ;
        RECT 697.445 18.800 766.290 18.940 ;
        RECT 697.445 18.755 697.735 18.800 ;
        RECT 765.970 18.740 766.290 18.800 ;
      LAYER via ;
        RECT 234.700 20.100 234.960 20.360 ;
        RECT 766.000 18.740 766.260 19.000 ;
      LAYER met2 ;
        RECT 234.700 20.070 234.960 20.390 ;
        RECT 234.760 2.400 234.900 20.070 ;
        RECT 766.060 19.030 766.200 54.000 ;
        RECT 766.000 18.710 766.260 19.030 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 18.940 56.510 19.000 ;
        RECT 155.090 18.940 155.410 19.000 ;
        RECT 56.190 18.800 155.410 18.940 ;
        RECT 56.190 18.740 56.510 18.800 ;
        RECT 155.090 18.740 155.410 18.800 ;
      LAYER via ;
        RECT 56.220 18.740 56.480 19.000 ;
        RECT 155.120 18.740 155.380 19.000 ;
      LAYER met2 ;
        RECT 155.180 19.030 155.320 54.000 ;
        RECT 56.220 18.710 56.480 19.030 ;
        RECT 155.120 18.710 155.380 19.030 ;
        RECT 56.280 2.400 56.420 18.710 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 251.765 15.045 251.935 16.575 ;
      LAYER mcon ;
        RECT 251.765 16.405 251.935 16.575 ;
      LAYER met1 ;
        RECT 80.110 16.560 80.430 16.620 ;
        RECT 251.705 16.560 251.995 16.605 ;
        RECT 80.110 16.420 251.995 16.560 ;
        RECT 80.110 16.360 80.430 16.420 ;
        RECT 251.705 16.375 251.995 16.420 ;
        RECT 251.705 15.200 251.995 15.245 ;
        RECT 286.190 15.200 286.510 15.260 ;
        RECT 251.705 15.060 286.510 15.200 ;
        RECT 251.705 15.015 251.995 15.060 ;
        RECT 286.190 15.000 286.510 15.060 ;
      LAYER via ;
        RECT 80.140 16.360 80.400 16.620 ;
        RECT 286.220 15.000 286.480 15.260 ;
      LAYER met2 ;
        RECT 80.140 16.330 80.400 16.650 ;
        RECT 80.200 2.400 80.340 16.330 ;
        RECT 286.280 15.290 286.420 54.000 ;
        RECT 286.220 14.970 286.480 15.290 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 289.945 15.385 290.115 16.235 ;
      LAYER mcon ;
        RECT 289.945 16.065 290.115 16.235 ;
      LAYER met1 ;
        RECT 103.570 16.220 103.890 16.280 ;
        RECT 289.885 16.220 290.175 16.265 ;
        RECT 103.570 16.080 290.175 16.220 ;
        RECT 103.570 16.020 103.890 16.080 ;
        RECT 289.885 16.035 290.175 16.080 ;
        RECT 289.885 15.540 290.175 15.585 ;
        RECT 306.890 15.540 307.210 15.600 ;
        RECT 289.885 15.400 307.210 15.540 ;
        RECT 289.885 15.355 290.175 15.400 ;
        RECT 306.890 15.340 307.210 15.400 ;
      LAYER via ;
        RECT 103.600 16.020 103.860 16.280 ;
        RECT 306.920 15.340 307.180 15.600 ;
      LAYER met2 ;
        RECT 103.600 15.990 103.860 16.310 ;
        RECT 103.660 2.400 103.800 15.990 ;
        RECT 306.980 15.630 307.120 54.000 ;
        RECT 306.920 15.310 307.180 15.630 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 691.080 16.845 691.220 54.000 ;
        RECT 127.510 16.475 127.790 16.845 ;
        RECT 691.010 16.475 691.290 16.845 ;
        RECT 127.580 2.400 127.720 16.475 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 127.510 16.520 127.790 16.800 ;
        RECT 691.010 16.520 691.290 16.800 ;
      LAYER met3 ;
        RECT 127.485 16.810 127.815 16.825 ;
        RECT 690.985 16.810 691.315 16.825 ;
        RECT 127.485 16.510 691.315 16.810 ;
        RECT 127.485 16.495 127.815 16.510 ;
        RECT 690.985 16.495 691.315 16.510 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 15.880 26.610 15.940 ;
        RECT 340.470 15.880 340.790 15.940 ;
        RECT 26.290 15.740 340.790 15.880 ;
        RECT 26.290 15.680 26.610 15.740 ;
        RECT 340.470 15.680 340.790 15.740 ;
      LAYER via ;
        RECT 26.320 15.680 26.580 15.940 ;
        RECT 340.500 15.680 340.760 15.940 ;
      LAYER met2 ;
        RECT 340.560 15.970 340.700 54.000 ;
        RECT 26.320 15.650 26.580 15.970 ;
        RECT 340.500 15.650 340.760 15.970 ;
        RECT 26.380 2.400 26.520 15.650 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 17.920 32.590 17.980 ;
        RECT 567.250 17.920 567.570 17.980 ;
        RECT 32.270 17.780 567.570 17.920 ;
        RECT 32.270 17.720 32.590 17.780 ;
        RECT 567.250 17.720 567.570 17.780 ;
        RECT 580.130 17.920 580.450 17.980 ;
        RECT 589.790 17.920 590.110 17.980 ;
        RECT 580.130 17.780 590.110 17.920 ;
        RECT 580.130 17.720 580.450 17.780 ;
        RECT 589.790 17.720 590.110 17.780 ;
      LAYER via ;
        RECT 32.300 17.720 32.560 17.980 ;
        RECT 567.280 17.720 567.540 17.980 ;
        RECT 580.160 17.720 580.420 17.980 ;
        RECT 589.820 17.720 590.080 17.980 ;
      LAYER met2 ;
        RECT 32.300 17.690 32.560 18.010 ;
        RECT 567.270 17.835 567.550 18.205 ;
        RECT 580.150 17.835 580.430 18.205 ;
        RECT 589.880 18.010 590.020 54.000 ;
        RECT 567.280 17.690 567.540 17.835 ;
        RECT 580.160 17.690 580.420 17.835 ;
        RECT 589.820 17.690 590.080 18.010 ;
        RECT 32.360 2.400 32.500 17.690 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 567.270 17.880 567.550 18.160 ;
        RECT 580.150 17.880 580.430 18.160 ;
      LAYER met3 ;
        RECT 567.245 18.170 567.575 18.185 ;
        RECT 580.125 18.170 580.455 18.185 ;
        RECT 567.245 17.870 580.455 18.170 ;
        RECT 567.245 17.855 567.575 17.870 ;
        RECT 580.125 17.855 580.455 17.870 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 3466.000 187.020 3529.000 ;
        RECT 364.020 3466.000 367.020 3529.000 ;
        RECT 544.020 3466.000 547.020 3529.000 ;
        RECT 724.020 3466.000 727.020 3529.000 ;
        RECT 904.020 3466.000 907.020 3529.000 ;
        RECT 1084.020 3466.000 1087.020 3529.000 ;
        RECT 1264.020 3466.000 1267.020 3529.000 ;
        RECT 1444.020 3466.000 1447.020 3529.000 ;
        RECT 1624.020 3466.000 1627.020 3529.000 ;
        RECT 1804.020 3466.000 1807.020 3529.000 ;
        RECT 1984.020 3466.000 1987.020 3529.000 ;
        RECT 2164.020 3466.000 2167.020 3529.000 ;
        RECT 2344.020 3466.000 2347.020 3529.000 ;
        RECT 2524.020 3466.000 2527.020 3529.000 ;
        RECT 2704.020 3466.000 2707.020 3529.000 ;
        RECT 184.020 -9.320 187.020 54.000 ;
        RECT 364.020 -9.320 367.020 54.000 ;
        RECT 544.020 -9.320 547.020 54.000 ;
        RECT 724.020 -9.320 727.020 54.000 ;
        RECT 904.020 -9.320 907.020 54.000 ;
        RECT 1084.020 -9.320 1087.020 54.000 ;
        RECT 1264.020 -9.320 1267.020 54.000 ;
        RECT 1444.020 -9.320 1447.020 54.000 ;
        RECT 1624.020 -9.320 1627.020 54.000 ;
        RECT 1804.020 -9.320 1807.020 54.000 ;
        RECT 1984.020 -9.320 1987.020 54.000 ;
        RECT 2164.020 -9.320 2167.020 54.000 ;
        RECT 2344.020 -9.320 2347.020 54.000 ;
        RECT 2524.020 -9.320 2527.020 54.000 ;
        RECT 2704.020 -9.320 2707.020 54.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 54.000 3432.380 ;
        RECT 2866.000 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 54.000 3252.380 ;
        RECT 2866.000 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 54.000 3072.380 ;
        RECT 2866.000 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 54.000 2892.380 ;
        RECT 2866.000 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 54.000 2712.380 ;
        RECT 2866.000 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 54.000 2532.380 ;
        RECT 2866.000 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 54.000 2352.380 ;
        RECT 2866.000 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 54.000 2172.380 ;
        RECT 2866.000 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 54.000 1992.380 ;
        RECT 2866.000 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 54.000 1812.380 ;
        RECT 2866.000 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 54.000 1632.380 ;
        RECT 2866.000 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 54.000 1452.380 ;
        RECT 2866.000 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 54.000 1272.380 ;
        RECT 2866.000 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 54.000 1092.380 ;
        RECT 2866.000 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 54.000 912.380 ;
        RECT 2866.000 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 54.000 732.380 ;
        RECT 2866.000 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 54.000 552.380 ;
        RECT 2866.000 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 54.000 372.380 ;
        RECT 2866.000 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 54.000 192.380 ;
        RECT 2866.000 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 3466.000 97.020 3529.000 ;
        RECT 274.020 3466.000 277.020 3529.000 ;
        RECT 454.020 3466.000 457.020 3529.000 ;
        RECT 634.020 3466.000 637.020 3529.000 ;
        RECT 814.020 3466.000 817.020 3529.000 ;
        RECT 994.020 3466.000 997.020 3529.000 ;
        RECT 1174.020 3466.000 1177.020 3529.000 ;
        RECT 1354.020 3466.000 1357.020 3529.000 ;
        RECT 1534.020 3466.000 1537.020 3529.000 ;
        RECT 1714.020 3466.000 1717.020 3529.000 ;
        RECT 1894.020 3466.000 1897.020 3529.000 ;
        RECT 2074.020 3466.000 2077.020 3529.000 ;
        RECT 2254.020 3466.000 2257.020 3529.000 ;
        RECT 2434.020 3466.000 2437.020 3529.000 ;
        RECT 2614.020 3466.000 2617.020 3529.000 ;
        RECT 2794.020 3466.000 2797.020 3529.000 ;
        RECT 94.020 -9.320 97.020 54.000 ;
        RECT 274.020 -9.320 277.020 54.000 ;
        RECT 454.020 -9.320 457.020 54.000 ;
        RECT 634.020 -9.320 637.020 54.000 ;
        RECT 814.020 -9.320 817.020 54.000 ;
        RECT 994.020 -9.320 997.020 54.000 ;
        RECT 1174.020 -9.320 1177.020 54.000 ;
        RECT 1354.020 -9.320 1357.020 54.000 ;
        RECT 1534.020 -9.320 1537.020 54.000 ;
        RECT 1714.020 -9.320 1717.020 54.000 ;
        RECT 1894.020 -9.320 1897.020 54.000 ;
        RECT 2074.020 -9.320 2077.020 54.000 ;
        RECT 2254.020 -9.320 2257.020 54.000 ;
        RECT 2434.020 -9.320 2437.020 54.000 ;
        RECT 2614.020 -9.320 2617.020 54.000 ;
        RECT 2794.020 -9.320 2797.020 54.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 54.000 3342.380 ;
        RECT 2866.000 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 54.000 3162.380 ;
        RECT 2866.000 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 54.000 2982.380 ;
        RECT 2866.000 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 54.000 2802.380 ;
        RECT 2866.000 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 54.000 2622.380 ;
        RECT 2866.000 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 54.000 2442.380 ;
        RECT 2866.000 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 54.000 2262.380 ;
        RECT 2866.000 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 54.000 2082.380 ;
        RECT 2866.000 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 54.000 1902.380 ;
        RECT 2866.000 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 54.000 1722.380 ;
        RECT 2866.000 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 54.000 1542.380 ;
        RECT 2866.000 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 54.000 1362.380 ;
        RECT 2866.000 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 54.000 1182.380 ;
        RECT 2866.000 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 54.000 1002.380 ;
        RECT 2866.000 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 54.000 822.380 ;
        RECT 2866.000 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 54.000 642.380 ;
        RECT 2866.000 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 54.000 462.380 ;
        RECT 2866.000 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 54.000 282.380 ;
        RECT 2866.000 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 54.000 102.380 ;
        RECT 2866.000 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 54.000 2633.765 2866.000 3415.555 ;
        RECT 54.000 2524.795 1593.750 2633.765 ;
      LAYER li1 ;
        RECT 1593.750 2524.795 2870.710 2633.765 ;
      LAYER li1 ;
        RECT 54.000 1087.745 2866.000 2524.795 ;
      LAYER li1 ;
        RECT 51.520 646.935 501.255 1087.745 ;
      LAYER li1 ;
        RECT 501.255 646.935 2866.000 1087.745 ;
        RECT 54.000 486.405 2866.000 646.935 ;
      LAYER li1 ;
        RECT 51.520 167.995 454.480 486.405 ;
      LAYER li1 ;
        RECT 454.480 167.995 2866.000 486.405 ;
        RECT 54.000 54.000 2866.000 167.995 ;
      LAYER met1 ;
        RECT 54.000 2666.860 2866.000 3463.880 ;
        RECT 2871.850 2666.860 2872.170 2666.920 ;
        RECT 54.000 2666.720 2872.170 2666.860 ;
        RECT 54.000 2639.420 2866.000 2666.720 ;
        RECT 2871.850 2666.660 2872.170 2666.720 ;
        RECT 54.000 2524.640 1591.060 2639.420 ;
      LAYER met1 ;
        RECT 1591.060 2524.640 2873.860 2639.420 ;
      LAYER met1 ;
        RECT 54.000 2494.140 2866.000 2524.640 ;
        RECT 2870.470 2494.140 2870.790 2494.200 ;
        RECT 54.000 2494.000 2870.790 2494.140 ;
        RECT 54.000 1087.900 2866.000 2494.000 ;
        RECT 2870.470 2493.940 2870.790 2494.000 ;
      LAYER met1 ;
        RECT 51.520 646.780 501.330 1087.900 ;
      LAYER met1 ;
        RECT 501.330 646.780 2866.000 1087.900 ;
        RECT 54.000 486.560 2866.000 646.780 ;
      LAYER met1 ;
        RECT 51.520 167.840 454.480 486.560 ;
      LAYER met1 ;
        RECT 454.480 167.840 2866.000 486.560 ;
        RECT 54.000 54.000 2866.000 167.840 ;
      LAYER via ;
        RECT 2871.880 2666.660 2872.140 2666.920 ;
        RECT 2870.500 2493.940 2870.760 2494.200 ;
      LAYER met2 ;
        RECT 54.840 2644.930 2866.000 3466.000 ;
        RECT 2871.880 2666.630 2872.140 2666.950 ;
        RECT 54.840 2643.570 2866.100 2644.930 ;
        RECT 2868.500 2643.570 2868.780 2644.560 ;
        RECT 2871.940 2644.250 2872.080 2666.630 ;
        RECT 2873.560 2644.250 2873.840 2644.560 ;
        RECT 2871.940 2644.110 2873.840 2644.250 ;
        RECT 54.840 2643.430 2868.780 2643.570 ;
        RECT 54.840 2640.560 2866.000 2643.430 ;
        RECT 2868.500 2640.560 2868.780 2643.430 ;
        RECT 2873.560 2640.560 2873.840 2644.110 ;
        RECT 54.840 2640.280 2863.540 2640.560 ;
      LAYER met2 ;
        RECT 2863.540 2640.280 2868.220 2640.560 ;
        RECT 2869.060 2640.280 2873.280 2640.560 ;
      LAYER met2 ;
        RECT 54.840 2518.280 1591.090 2640.280 ;
      LAYER met2 ;
        RECT 1591.090 2518.280 2873.830 2640.280 ;
      LAYER met2 ;
        RECT 54.840 2518.000 2863.540 2518.280 ;
      LAYER met2 ;
        RECT 2863.540 2518.000 2868.220 2518.280 ;
        RECT 2869.060 2518.000 2873.280 2518.280 ;
      LAYER met2 ;
        RECT 54.840 2514.370 2866.000 2518.000 ;
        RECT 2868.500 2514.370 2868.780 2518.000 ;
        RECT 2873.560 2514.370 2873.840 2518.000 ;
        RECT 54.840 2514.230 2868.780 2514.370 ;
        RECT 54.840 54.000 2866.000 2514.230 ;
        RECT 2868.500 2514.000 2868.780 2514.230 ;
        RECT 2870.560 2514.230 2873.840 2514.370 ;
        RECT 2870.560 2494.230 2870.700 2514.230 ;
        RECT 2873.560 2514.000 2873.840 2514.230 ;
        RECT 2870.500 2493.910 2870.760 2494.230 ;
      LAYER met3 ;
        RECT 54.000 1095.645 2830.165 3416.145 ;
      LAYER met3 ;
        RECT 50.000 1094.780 501.600 1095.645 ;
      LAYER met3 ;
        RECT 501.600 1094.780 2830.165 1095.645 ;
      LAYER met3 ;
        RECT 50.000 1090.060 502.000 1094.780 ;
      LAYER met3 ;
        RECT 502.000 1090.060 2830.165 1094.780 ;
      LAYER met3 ;
        RECT 50.000 1088.660 501.600 1090.060 ;
      LAYER met3 ;
        RECT 501.600 1088.660 2830.165 1090.060 ;
      LAYER met3 ;
        RECT 50.000 1083.940 502.000 1088.660 ;
      LAYER met3 ;
        RECT 502.000 1083.940 2830.165 1088.660 ;
      LAYER met3 ;
        RECT 50.000 1082.540 501.600 1083.940 ;
      LAYER met3 ;
        RECT 501.600 1082.540 2830.165 1083.940 ;
      LAYER met3 ;
        RECT 50.000 1077.820 502.000 1082.540 ;
      LAYER met3 ;
        RECT 502.000 1077.820 2830.165 1082.540 ;
      LAYER met3 ;
        RECT 50.000 1076.420 501.600 1077.820 ;
      LAYER met3 ;
        RECT 501.600 1076.420 2830.165 1077.820 ;
      LAYER met3 ;
        RECT 50.000 1071.700 502.000 1076.420 ;
      LAYER met3 ;
        RECT 502.000 1071.700 2830.165 1076.420 ;
      LAYER met3 ;
        RECT 50.000 1070.300 501.600 1071.700 ;
      LAYER met3 ;
        RECT 501.600 1070.300 2830.165 1071.700 ;
      LAYER met3 ;
        RECT 50.000 1065.580 502.000 1070.300 ;
      LAYER met3 ;
        RECT 502.000 1065.580 2830.165 1070.300 ;
      LAYER met3 ;
        RECT 50.000 1064.180 501.600 1065.580 ;
      LAYER met3 ;
        RECT 501.600 1064.180 2830.165 1065.580 ;
      LAYER met3 ;
        RECT 50.000 1059.460 502.000 1064.180 ;
      LAYER met3 ;
        RECT 502.000 1059.460 2830.165 1064.180 ;
      LAYER met3 ;
        RECT 50.000 1058.060 501.600 1059.460 ;
      LAYER met3 ;
        RECT 501.600 1058.060 2830.165 1059.460 ;
      LAYER met3 ;
        RECT 50.000 1053.340 502.000 1058.060 ;
      LAYER met3 ;
        RECT 502.000 1053.340 2830.165 1058.060 ;
      LAYER met3 ;
        RECT 50.000 1051.940 501.600 1053.340 ;
      LAYER met3 ;
        RECT 501.600 1051.940 2830.165 1053.340 ;
      LAYER met3 ;
        RECT 50.000 1047.220 502.000 1051.940 ;
      LAYER met3 ;
        RECT 502.000 1047.220 2830.165 1051.940 ;
      LAYER met3 ;
        RECT 50.000 1045.820 501.600 1047.220 ;
      LAYER met3 ;
        RECT 501.600 1045.820 2830.165 1047.220 ;
      LAYER met3 ;
        RECT 50.000 1041.100 502.000 1045.820 ;
      LAYER met3 ;
        RECT 502.000 1041.100 2830.165 1045.820 ;
      LAYER met3 ;
        RECT 50.000 1039.700 501.600 1041.100 ;
      LAYER met3 ;
        RECT 501.600 1039.700 2830.165 1041.100 ;
      LAYER met3 ;
        RECT 50.000 1034.980 502.000 1039.700 ;
      LAYER met3 ;
        RECT 502.000 1034.980 2830.165 1039.700 ;
      LAYER met3 ;
        RECT 50.000 1033.580 501.600 1034.980 ;
      LAYER met3 ;
        RECT 501.600 1033.580 2830.165 1034.980 ;
      LAYER met3 ;
        RECT 50.000 1028.860 502.000 1033.580 ;
      LAYER met3 ;
        RECT 502.000 1028.860 2830.165 1033.580 ;
      LAYER met3 ;
        RECT 50.000 1027.460 501.600 1028.860 ;
      LAYER met3 ;
        RECT 501.600 1027.460 2830.165 1028.860 ;
      LAYER met3 ;
        RECT 50.000 1022.740 502.000 1027.460 ;
      LAYER met3 ;
        RECT 502.000 1022.740 2830.165 1027.460 ;
      LAYER met3 ;
        RECT 50.000 1021.340 501.600 1022.740 ;
      LAYER met3 ;
        RECT 501.600 1021.340 2830.165 1022.740 ;
      LAYER met3 ;
        RECT 50.000 1016.620 502.000 1021.340 ;
      LAYER met3 ;
        RECT 502.000 1016.620 2830.165 1021.340 ;
      LAYER met3 ;
        RECT 50.000 1015.220 501.600 1016.620 ;
      LAYER met3 ;
        RECT 501.600 1015.220 2830.165 1016.620 ;
      LAYER met3 ;
        RECT 50.000 1010.500 502.000 1015.220 ;
      LAYER met3 ;
        RECT 502.000 1010.500 2830.165 1015.220 ;
      LAYER met3 ;
        RECT 50.000 1009.100 501.600 1010.500 ;
      LAYER met3 ;
        RECT 501.600 1009.100 2830.165 1010.500 ;
      LAYER met3 ;
        RECT 50.000 1004.380 502.000 1009.100 ;
      LAYER met3 ;
        RECT 502.000 1004.380 2830.165 1009.100 ;
      LAYER met3 ;
        RECT 50.000 1002.980 501.600 1004.380 ;
      LAYER met3 ;
        RECT 501.600 1002.980 2830.165 1004.380 ;
      LAYER met3 ;
        RECT 50.000 998.260 502.000 1002.980 ;
      LAYER met3 ;
        RECT 502.000 998.260 2830.165 1002.980 ;
      LAYER met3 ;
        RECT 50.000 996.860 501.600 998.260 ;
      LAYER met3 ;
        RECT 501.600 996.860 2830.165 998.260 ;
      LAYER met3 ;
        RECT 50.000 992.140 502.000 996.860 ;
      LAYER met3 ;
        RECT 502.000 992.140 2830.165 996.860 ;
      LAYER met3 ;
        RECT 50.000 990.740 501.600 992.140 ;
      LAYER met3 ;
        RECT 501.600 990.740 2830.165 992.140 ;
      LAYER met3 ;
        RECT 50.000 986.700 502.000 990.740 ;
      LAYER met3 ;
        RECT 502.000 986.700 2830.165 990.740 ;
      LAYER met3 ;
        RECT 50.000 985.300 501.600 986.700 ;
      LAYER met3 ;
        RECT 501.600 985.300 2830.165 986.700 ;
      LAYER met3 ;
        RECT 50.000 980.580 502.000 985.300 ;
      LAYER met3 ;
        RECT 502.000 980.580 2830.165 985.300 ;
      LAYER met3 ;
        RECT 50.000 979.180 501.600 980.580 ;
      LAYER met3 ;
        RECT 501.600 979.180 2830.165 980.580 ;
      LAYER met3 ;
        RECT 50.000 974.460 502.000 979.180 ;
      LAYER met3 ;
        RECT 502.000 974.460 2830.165 979.180 ;
      LAYER met3 ;
        RECT 50.000 973.060 501.600 974.460 ;
      LAYER met3 ;
        RECT 501.600 973.060 2830.165 974.460 ;
      LAYER met3 ;
        RECT 50.000 968.340 502.000 973.060 ;
      LAYER met3 ;
        RECT 502.000 968.340 2830.165 973.060 ;
      LAYER met3 ;
        RECT 50.000 966.940 501.600 968.340 ;
      LAYER met3 ;
        RECT 501.600 966.940 2830.165 968.340 ;
      LAYER met3 ;
        RECT 50.000 962.220 502.000 966.940 ;
      LAYER met3 ;
        RECT 502.000 962.220 2830.165 966.940 ;
      LAYER met3 ;
        RECT 50.000 960.820 501.600 962.220 ;
      LAYER met3 ;
        RECT 501.600 960.820 2830.165 962.220 ;
      LAYER met3 ;
        RECT 50.000 956.100 502.000 960.820 ;
      LAYER met3 ;
        RECT 502.000 956.100 2830.165 960.820 ;
      LAYER met3 ;
        RECT 50.000 954.700 501.600 956.100 ;
      LAYER met3 ;
        RECT 501.600 954.700 2830.165 956.100 ;
      LAYER met3 ;
        RECT 50.000 949.980 502.000 954.700 ;
      LAYER met3 ;
        RECT 502.000 949.980 2830.165 954.700 ;
      LAYER met3 ;
        RECT 50.000 948.580 501.600 949.980 ;
      LAYER met3 ;
        RECT 501.600 948.580 2830.165 949.980 ;
      LAYER met3 ;
        RECT 50.000 943.860 502.000 948.580 ;
      LAYER met3 ;
        RECT 502.000 943.860 2830.165 948.580 ;
      LAYER met3 ;
        RECT 50.000 942.460 501.600 943.860 ;
      LAYER met3 ;
        RECT 501.600 942.460 2830.165 943.860 ;
      LAYER met3 ;
        RECT 50.000 937.740 502.000 942.460 ;
      LAYER met3 ;
        RECT 502.000 937.740 2830.165 942.460 ;
      LAYER met3 ;
        RECT 50.000 936.340 501.600 937.740 ;
      LAYER met3 ;
        RECT 501.600 936.340 2830.165 937.740 ;
      LAYER met3 ;
        RECT 50.000 931.620 502.000 936.340 ;
      LAYER met3 ;
        RECT 502.000 931.620 2830.165 936.340 ;
      LAYER met3 ;
        RECT 50.000 930.220 501.600 931.620 ;
      LAYER met3 ;
        RECT 501.600 930.220 2830.165 931.620 ;
      LAYER met3 ;
        RECT 50.000 925.500 502.000 930.220 ;
      LAYER met3 ;
        RECT 502.000 925.500 2830.165 930.220 ;
      LAYER met3 ;
        RECT 50.000 924.100 501.600 925.500 ;
      LAYER met3 ;
        RECT 501.600 924.100 2830.165 925.500 ;
      LAYER met3 ;
        RECT 50.000 919.380 502.000 924.100 ;
      LAYER met3 ;
        RECT 502.000 919.380 2830.165 924.100 ;
      LAYER met3 ;
        RECT 50.000 917.980 501.600 919.380 ;
      LAYER met3 ;
        RECT 501.600 917.980 2830.165 919.380 ;
      LAYER met3 ;
        RECT 50.000 913.260 502.000 917.980 ;
      LAYER met3 ;
        RECT 502.000 913.260 2830.165 917.980 ;
      LAYER met3 ;
        RECT 50.000 911.860 501.600 913.260 ;
      LAYER met3 ;
        RECT 501.600 911.860 2830.165 913.260 ;
      LAYER met3 ;
        RECT 50.000 907.140 502.000 911.860 ;
      LAYER met3 ;
        RECT 502.000 907.140 2830.165 911.860 ;
      LAYER met3 ;
        RECT 50.000 905.740 501.600 907.140 ;
      LAYER met3 ;
        RECT 501.600 905.740 2830.165 907.140 ;
      LAYER met3 ;
        RECT 50.000 901.020 502.000 905.740 ;
      LAYER met3 ;
        RECT 502.000 901.020 2830.165 905.740 ;
      LAYER met3 ;
        RECT 50.000 899.620 501.600 901.020 ;
      LAYER met3 ;
        RECT 501.600 899.620 2830.165 901.020 ;
      LAYER met3 ;
        RECT 50.000 894.900 502.000 899.620 ;
      LAYER met3 ;
        RECT 502.000 894.900 2830.165 899.620 ;
      LAYER met3 ;
        RECT 50.000 893.500 501.600 894.900 ;
      LAYER met3 ;
        RECT 501.600 893.500 2830.165 894.900 ;
      LAYER met3 ;
        RECT 50.000 888.780 502.000 893.500 ;
      LAYER met3 ;
        RECT 502.000 888.780 2830.165 893.500 ;
      LAYER met3 ;
        RECT 50.000 887.380 501.600 888.780 ;
      LAYER met3 ;
        RECT 501.600 887.380 2830.165 888.780 ;
      LAYER met3 ;
        RECT 50.000 882.660 502.000 887.380 ;
      LAYER met3 ;
        RECT 502.000 882.660 2830.165 887.380 ;
      LAYER met3 ;
        RECT 50.000 881.260 501.600 882.660 ;
      LAYER met3 ;
        RECT 501.600 881.260 2830.165 882.660 ;
      LAYER met3 ;
        RECT 50.000 876.540 502.000 881.260 ;
      LAYER met3 ;
        RECT 502.000 876.540 2830.165 881.260 ;
      LAYER met3 ;
        RECT 50.000 875.140 501.600 876.540 ;
      LAYER met3 ;
        RECT 501.600 875.140 2830.165 876.540 ;
      LAYER met3 ;
        RECT 50.000 871.100 502.000 875.140 ;
      LAYER met3 ;
        RECT 502.000 871.100 2830.165 875.140 ;
      LAYER met3 ;
        RECT 50.000 869.700 501.600 871.100 ;
      LAYER met3 ;
        RECT 501.600 869.700 2830.165 871.100 ;
      LAYER met3 ;
        RECT 50.000 868.380 502.000 869.700 ;
        RECT 50.400 866.980 502.000 868.380 ;
        RECT 50.000 864.980 502.000 866.980 ;
      LAYER met3 ;
        RECT 502.000 864.980 2830.165 869.700 ;
      LAYER met3 ;
        RECT 50.000 863.580 501.600 864.980 ;
      LAYER met3 ;
        RECT 501.600 863.580 2830.165 864.980 ;
      LAYER met3 ;
        RECT 50.000 858.860 502.000 863.580 ;
      LAYER met3 ;
        RECT 502.000 858.860 2830.165 863.580 ;
      LAYER met3 ;
        RECT 50.000 857.460 501.600 858.860 ;
      LAYER met3 ;
        RECT 501.600 857.460 2830.165 858.860 ;
      LAYER met3 ;
        RECT 50.000 852.740 502.000 857.460 ;
      LAYER met3 ;
        RECT 502.000 852.740 2830.165 857.460 ;
      LAYER met3 ;
        RECT 50.000 851.340 501.600 852.740 ;
      LAYER met3 ;
        RECT 501.600 851.340 2830.165 852.740 ;
      LAYER met3 ;
        RECT 50.000 846.620 502.000 851.340 ;
      LAYER met3 ;
        RECT 502.000 846.620 2830.165 851.340 ;
      LAYER met3 ;
        RECT 50.000 845.220 501.600 846.620 ;
      LAYER met3 ;
        RECT 501.600 845.220 2830.165 846.620 ;
      LAYER met3 ;
        RECT 50.000 840.500 502.000 845.220 ;
      LAYER met3 ;
        RECT 502.000 840.500 2830.165 845.220 ;
      LAYER met3 ;
        RECT 50.000 839.100 501.600 840.500 ;
      LAYER met3 ;
        RECT 501.600 839.100 2830.165 840.500 ;
      LAYER met3 ;
        RECT 50.000 834.380 502.000 839.100 ;
      LAYER met3 ;
        RECT 502.000 834.380 2830.165 839.100 ;
      LAYER met3 ;
        RECT 50.000 832.980 501.600 834.380 ;
      LAYER met3 ;
        RECT 501.600 832.980 2830.165 834.380 ;
      LAYER met3 ;
        RECT 50.000 828.260 502.000 832.980 ;
      LAYER met3 ;
        RECT 502.000 828.260 2830.165 832.980 ;
      LAYER met3 ;
        RECT 50.000 826.860 501.600 828.260 ;
      LAYER met3 ;
        RECT 501.600 826.860 2830.165 828.260 ;
      LAYER met3 ;
        RECT 50.000 822.140 502.000 826.860 ;
      LAYER met3 ;
        RECT 502.000 822.140 2830.165 826.860 ;
      LAYER met3 ;
        RECT 50.000 820.740 501.600 822.140 ;
      LAYER met3 ;
        RECT 501.600 820.740 2830.165 822.140 ;
      LAYER met3 ;
        RECT 50.000 816.020 502.000 820.740 ;
      LAYER met3 ;
        RECT 502.000 816.020 2830.165 820.740 ;
      LAYER met3 ;
        RECT 50.000 814.620 501.600 816.020 ;
      LAYER met3 ;
        RECT 501.600 814.620 2830.165 816.020 ;
      LAYER met3 ;
        RECT 50.000 809.900 502.000 814.620 ;
      LAYER met3 ;
        RECT 502.000 809.900 2830.165 814.620 ;
      LAYER met3 ;
        RECT 50.000 808.500 501.600 809.900 ;
      LAYER met3 ;
        RECT 501.600 808.500 2830.165 809.900 ;
      LAYER met3 ;
        RECT 50.000 803.780 502.000 808.500 ;
      LAYER met3 ;
        RECT 502.000 803.780 2830.165 808.500 ;
      LAYER met3 ;
        RECT 50.000 802.380 501.600 803.780 ;
      LAYER met3 ;
        RECT 501.600 802.380 2830.165 803.780 ;
      LAYER met3 ;
        RECT 50.000 797.660 502.000 802.380 ;
      LAYER met3 ;
        RECT 502.000 797.660 2830.165 802.380 ;
      LAYER met3 ;
        RECT 50.000 796.260 501.600 797.660 ;
      LAYER met3 ;
        RECT 501.600 796.260 2830.165 797.660 ;
      LAYER met3 ;
        RECT 50.000 791.540 502.000 796.260 ;
      LAYER met3 ;
        RECT 502.000 791.540 2830.165 796.260 ;
      LAYER met3 ;
        RECT 50.000 790.140 501.600 791.540 ;
      LAYER met3 ;
        RECT 501.600 790.140 2830.165 791.540 ;
      LAYER met3 ;
        RECT 50.000 785.420 502.000 790.140 ;
      LAYER met3 ;
        RECT 502.000 785.420 2830.165 790.140 ;
      LAYER met3 ;
        RECT 50.000 784.020 501.600 785.420 ;
      LAYER met3 ;
        RECT 501.600 784.020 2830.165 785.420 ;
      LAYER met3 ;
        RECT 50.000 779.300 502.000 784.020 ;
      LAYER met3 ;
        RECT 502.000 779.300 2830.165 784.020 ;
      LAYER met3 ;
        RECT 50.000 777.900 501.600 779.300 ;
      LAYER met3 ;
        RECT 501.600 777.900 2830.165 779.300 ;
      LAYER met3 ;
        RECT 50.000 773.180 502.000 777.900 ;
      LAYER met3 ;
        RECT 502.000 773.180 2830.165 777.900 ;
      LAYER met3 ;
        RECT 50.000 771.780 501.600 773.180 ;
      LAYER met3 ;
        RECT 501.600 771.780 2830.165 773.180 ;
      LAYER met3 ;
        RECT 50.000 767.060 502.000 771.780 ;
      LAYER met3 ;
        RECT 502.000 767.060 2830.165 771.780 ;
      LAYER met3 ;
        RECT 50.000 765.660 501.600 767.060 ;
      LAYER met3 ;
        RECT 501.600 765.660 2830.165 767.060 ;
      LAYER met3 ;
        RECT 50.000 760.940 502.000 765.660 ;
      LAYER met3 ;
        RECT 502.000 760.940 2830.165 765.660 ;
      LAYER met3 ;
        RECT 50.000 759.540 501.600 760.940 ;
      LAYER met3 ;
        RECT 501.600 759.540 2830.165 760.940 ;
      LAYER met3 ;
        RECT 50.000 755.500 502.000 759.540 ;
      LAYER met3 ;
        RECT 502.000 755.500 2830.165 759.540 ;
      LAYER met3 ;
        RECT 50.000 754.100 501.600 755.500 ;
      LAYER met3 ;
        RECT 501.600 754.100 2830.165 755.500 ;
      LAYER met3 ;
        RECT 50.000 749.380 502.000 754.100 ;
      LAYER met3 ;
        RECT 502.000 749.380 2830.165 754.100 ;
      LAYER met3 ;
        RECT 50.000 747.980 501.600 749.380 ;
      LAYER met3 ;
        RECT 501.600 747.980 2830.165 749.380 ;
      LAYER met3 ;
        RECT 50.000 743.260 502.000 747.980 ;
      LAYER met3 ;
        RECT 502.000 743.260 2830.165 747.980 ;
      LAYER met3 ;
        RECT 50.000 741.860 501.600 743.260 ;
      LAYER met3 ;
        RECT 501.600 741.860 2830.165 743.260 ;
      LAYER met3 ;
        RECT 50.000 737.140 502.000 741.860 ;
      LAYER met3 ;
        RECT 502.000 737.140 2830.165 741.860 ;
      LAYER met3 ;
        RECT 50.000 735.740 501.600 737.140 ;
      LAYER met3 ;
        RECT 501.600 735.740 2830.165 737.140 ;
      LAYER met3 ;
        RECT 50.000 731.020 502.000 735.740 ;
      LAYER met3 ;
        RECT 502.000 731.020 2830.165 735.740 ;
      LAYER met3 ;
        RECT 50.000 729.620 501.600 731.020 ;
      LAYER met3 ;
        RECT 501.600 729.620 2830.165 731.020 ;
      LAYER met3 ;
        RECT 50.000 724.900 502.000 729.620 ;
      LAYER met3 ;
        RECT 502.000 724.900 2830.165 729.620 ;
      LAYER met3 ;
        RECT 50.000 723.500 501.600 724.900 ;
      LAYER met3 ;
        RECT 501.600 723.500 2830.165 724.900 ;
      LAYER met3 ;
        RECT 50.000 718.780 502.000 723.500 ;
      LAYER met3 ;
        RECT 502.000 718.780 2830.165 723.500 ;
      LAYER met3 ;
        RECT 50.000 717.380 501.600 718.780 ;
      LAYER met3 ;
        RECT 501.600 717.380 2830.165 718.780 ;
      LAYER met3 ;
        RECT 50.000 712.660 502.000 717.380 ;
      LAYER met3 ;
        RECT 502.000 712.660 2830.165 717.380 ;
      LAYER met3 ;
        RECT 50.000 711.260 501.600 712.660 ;
      LAYER met3 ;
        RECT 501.600 711.260 2830.165 712.660 ;
      LAYER met3 ;
        RECT 50.000 706.540 502.000 711.260 ;
      LAYER met3 ;
        RECT 502.000 706.540 2830.165 711.260 ;
      LAYER met3 ;
        RECT 50.000 705.140 501.600 706.540 ;
      LAYER met3 ;
        RECT 501.600 705.140 2830.165 706.540 ;
      LAYER met3 ;
        RECT 50.000 700.420 502.000 705.140 ;
      LAYER met3 ;
        RECT 502.000 700.420 2830.165 705.140 ;
      LAYER met3 ;
        RECT 50.000 699.020 501.600 700.420 ;
      LAYER met3 ;
        RECT 501.600 699.020 2830.165 700.420 ;
      LAYER met3 ;
        RECT 50.000 694.300 502.000 699.020 ;
      LAYER met3 ;
        RECT 502.000 694.300 2830.165 699.020 ;
      LAYER met3 ;
        RECT 50.000 692.900 501.600 694.300 ;
      LAYER met3 ;
        RECT 501.600 692.900 2830.165 694.300 ;
      LAYER met3 ;
        RECT 50.000 688.180 502.000 692.900 ;
      LAYER met3 ;
        RECT 502.000 688.180 2830.165 692.900 ;
      LAYER met3 ;
        RECT 50.000 686.780 501.600 688.180 ;
      LAYER met3 ;
        RECT 501.600 686.780 2830.165 688.180 ;
      LAYER met3 ;
        RECT 50.000 682.060 502.000 686.780 ;
      LAYER met3 ;
        RECT 502.000 682.060 2830.165 686.780 ;
      LAYER met3 ;
        RECT 50.000 680.660 501.600 682.060 ;
      LAYER met3 ;
        RECT 501.600 680.660 2830.165 682.060 ;
      LAYER met3 ;
        RECT 50.000 675.940 502.000 680.660 ;
      LAYER met3 ;
        RECT 502.000 675.940 2830.165 680.660 ;
      LAYER met3 ;
        RECT 50.000 674.540 501.600 675.940 ;
      LAYER met3 ;
        RECT 501.600 674.540 2830.165 675.940 ;
      LAYER met3 ;
        RECT 50.000 669.820 502.000 674.540 ;
      LAYER met3 ;
        RECT 502.000 669.820 2830.165 674.540 ;
      LAYER met3 ;
        RECT 50.000 668.420 501.600 669.820 ;
      LAYER met3 ;
        RECT 501.600 668.420 2830.165 669.820 ;
      LAYER met3 ;
        RECT 50.000 663.700 502.000 668.420 ;
      LAYER met3 ;
        RECT 502.000 663.700 2830.165 668.420 ;
      LAYER met3 ;
        RECT 50.000 662.300 501.600 663.700 ;
      LAYER met3 ;
        RECT 501.600 662.300 2830.165 663.700 ;
      LAYER met3 ;
        RECT 50.000 657.580 502.000 662.300 ;
      LAYER met3 ;
        RECT 502.000 657.580 2830.165 662.300 ;
      LAYER met3 ;
        RECT 50.000 656.180 501.600 657.580 ;
      LAYER met3 ;
        RECT 501.600 656.180 2830.165 657.580 ;
      LAYER met3 ;
        RECT 50.000 651.460 502.000 656.180 ;
      LAYER met3 ;
        RECT 502.000 651.460 2830.165 656.180 ;
      LAYER met3 ;
        RECT 50.000 650.060 501.600 651.460 ;
      LAYER met3 ;
        RECT 501.600 650.060 2830.165 651.460 ;
      LAYER met3 ;
        RECT 50.000 645.340 502.000 650.060 ;
      LAYER met3 ;
        RECT 502.000 645.340 2830.165 650.060 ;
      LAYER met3 ;
        RECT 50.000 643.940 501.600 645.340 ;
      LAYER met3 ;
        RECT 501.600 643.940 2830.165 645.340 ;
      LAYER met3 ;
        RECT 50.000 639.900 502.000 643.940 ;
      LAYER met3 ;
        RECT 502.000 639.900 2830.165 643.940 ;
      LAYER met3 ;
        RECT 50.000 639.035 501.600 639.900 ;
      LAYER met3 ;
        RECT 501.600 639.035 2830.165 639.900 ;
        RECT 54.000 494.985 2830.165 639.035 ;
      LAYER met3 ;
        RECT 50.000 494.120 455.600 494.985 ;
      LAYER met3 ;
        RECT 455.600 494.120 2830.165 494.985 ;
      LAYER met3 ;
        RECT 50.000 490.760 456.000 494.120 ;
      LAYER met3 ;
        RECT 456.000 490.760 2830.165 494.120 ;
      LAYER met3 ;
        RECT 50.000 489.360 455.600 490.760 ;
      LAYER met3 ;
        RECT 455.600 489.360 2830.165 490.760 ;
      LAYER met3 ;
        RECT 50.000 486.680 456.000 489.360 ;
      LAYER met3 ;
        RECT 456.000 486.680 2830.165 489.360 ;
      LAYER met3 ;
        RECT 50.000 485.280 455.600 486.680 ;
      LAYER met3 ;
        RECT 455.600 485.280 2830.165 486.680 ;
      LAYER met3 ;
        RECT 50.000 481.920 456.000 485.280 ;
      LAYER met3 ;
        RECT 456.000 481.920 2830.165 485.280 ;
      LAYER met3 ;
        RECT 50.000 480.520 455.600 481.920 ;
      LAYER met3 ;
        RECT 455.600 480.520 2830.165 481.920 ;
      LAYER met3 ;
        RECT 50.000 477.840 456.000 480.520 ;
      LAYER met3 ;
        RECT 456.000 477.840 2830.165 480.520 ;
      LAYER met3 ;
        RECT 50.000 476.440 455.600 477.840 ;
      LAYER met3 ;
        RECT 455.600 476.440 2830.165 477.840 ;
      LAYER met3 ;
        RECT 50.000 473.080 456.000 476.440 ;
      LAYER met3 ;
        RECT 456.000 473.080 2830.165 476.440 ;
      LAYER met3 ;
        RECT 50.000 471.680 455.600 473.080 ;
      LAYER met3 ;
        RECT 455.600 471.680 2830.165 473.080 ;
      LAYER met3 ;
        RECT 50.000 468.320 456.000 471.680 ;
      LAYER met3 ;
        RECT 456.000 468.320 2830.165 471.680 ;
      LAYER met3 ;
        RECT 50.000 466.920 455.600 468.320 ;
      LAYER met3 ;
        RECT 455.600 466.920 2830.165 468.320 ;
      LAYER met3 ;
        RECT 50.000 464.240 456.000 466.920 ;
      LAYER met3 ;
        RECT 456.000 464.240 2830.165 466.920 ;
      LAYER met3 ;
        RECT 50.000 462.840 455.600 464.240 ;
      LAYER met3 ;
        RECT 455.600 462.840 2830.165 464.240 ;
      LAYER met3 ;
        RECT 50.000 459.480 456.000 462.840 ;
      LAYER met3 ;
        RECT 456.000 459.480 2830.165 462.840 ;
      LAYER met3 ;
        RECT 50.000 458.080 455.600 459.480 ;
      LAYER met3 ;
        RECT 455.600 458.080 2830.165 459.480 ;
      LAYER met3 ;
        RECT 50.000 455.400 456.000 458.080 ;
      LAYER met3 ;
        RECT 456.000 455.400 2830.165 458.080 ;
      LAYER met3 ;
        RECT 50.000 454.000 455.600 455.400 ;
      LAYER met3 ;
        RECT 455.600 454.000 2830.165 455.400 ;
      LAYER met3 ;
        RECT 50.000 450.640 456.000 454.000 ;
      LAYER met3 ;
        RECT 456.000 450.640 2830.165 454.000 ;
      LAYER met3 ;
        RECT 50.000 449.240 455.600 450.640 ;
      LAYER met3 ;
        RECT 455.600 449.240 2830.165 450.640 ;
      LAYER met3 ;
        RECT 50.000 446.560 456.000 449.240 ;
      LAYER met3 ;
        RECT 456.000 446.560 2830.165 449.240 ;
      LAYER met3 ;
        RECT 50.000 445.160 455.600 446.560 ;
      LAYER met3 ;
        RECT 455.600 445.160 2830.165 446.560 ;
      LAYER met3 ;
        RECT 50.000 441.800 456.000 445.160 ;
      LAYER met3 ;
        RECT 456.000 441.800 2830.165 445.160 ;
      LAYER met3 ;
        RECT 50.000 440.400 455.600 441.800 ;
      LAYER met3 ;
        RECT 455.600 440.400 2830.165 441.800 ;
      LAYER met3 ;
        RECT 50.000 437.040 456.000 440.400 ;
      LAYER met3 ;
        RECT 456.000 437.040 2830.165 440.400 ;
      LAYER met3 ;
        RECT 50.000 435.640 455.600 437.040 ;
      LAYER met3 ;
        RECT 455.600 435.640 2830.165 437.040 ;
      LAYER met3 ;
        RECT 50.000 432.960 456.000 435.640 ;
      LAYER met3 ;
        RECT 456.000 432.960 2830.165 435.640 ;
      LAYER met3 ;
        RECT 50.000 431.560 455.600 432.960 ;
      LAYER met3 ;
        RECT 455.600 431.560 2830.165 432.960 ;
      LAYER met3 ;
        RECT 50.000 428.200 456.000 431.560 ;
      LAYER met3 ;
        RECT 456.000 428.200 2830.165 431.560 ;
      LAYER met3 ;
        RECT 50.000 426.800 455.600 428.200 ;
      LAYER met3 ;
        RECT 455.600 426.800 2830.165 428.200 ;
      LAYER met3 ;
        RECT 50.000 424.120 456.000 426.800 ;
      LAYER met3 ;
        RECT 456.000 424.120 2830.165 426.800 ;
      LAYER met3 ;
        RECT 50.000 422.720 455.600 424.120 ;
      LAYER met3 ;
        RECT 455.600 422.720 2830.165 424.120 ;
      LAYER met3 ;
        RECT 50.000 419.360 456.000 422.720 ;
      LAYER met3 ;
        RECT 456.000 419.360 2830.165 422.720 ;
      LAYER met3 ;
        RECT 50.000 417.960 455.600 419.360 ;
      LAYER met3 ;
        RECT 455.600 417.960 2830.165 419.360 ;
      LAYER met3 ;
        RECT 50.000 415.280 456.000 417.960 ;
      LAYER met3 ;
        RECT 456.000 415.280 2830.165 417.960 ;
      LAYER met3 ;
        RECT 50.000 413.880 455.600 415.280 ;
      LAYER met3 ;
        RECT 455.600 413.880 2830.165 415.280 ;
      LAYER met3 ;
        RECT 50.000 410.520 456.000 413.880 ;
      LAYER met3 ;
        RECT 456.000 410.520 2830.165 413.880 ;
      LAYER met3 ;
        RECT 50.000 409.120 455.600 410.520 ;
      LAYER met3 ;
        RECT 455.600 409.120 2830.165 410.520 ;
      LAYER met3 ;
        RECT 50.000 405.760 456.000 409.120 ;
      LAYER met3 ;
        RECT 456.000 405.760 2830.165 409.120 ;
      LAYER met3 ;
        RECT 50.000 404.360 455.600 405.760 ;
      LAYER met3 ;
        RECT 455.600 404.360 2830.165 405.760 ;
      LAYER met3 ;
        RECT 50.000 401.680 456.000 404.360 ;
      LAYER met3 ;
        RECT 456.000 401.680 2830.165 404.360 ;
      LAYER met3 ;
        RECT 50.000 400.280 455.600 401.680 ;
      LAYER met3 ;
        RECT 455.600 400.280 2830.165 401.680 ;
      LAYER met3 ;
        RECT 50.000 396.920 456.000 400.280 ;
      LAYER met3 ;
        RECT 456.000 396.920 2830.165 400.280 ;
      LAYER met3 ;
        RECT 50.000 395.520 455.600 396.920 ;
      LAYER met3 ;
        RECT 455.600 395.520 2830.165 396.920 ;
      LAYER met3 ;
        RECT 50.000 392.840 456.000 395.520 ;
      LAYER met3 ;
        RECT 456.000 392.840 2830.165 395.520 ;
      LAYER met3 ;
        RECT 50.000 391.440 455.600 392.840 ;
      LAYER met3 ;
        RECT 455.600 391.440 2830.165 392.840 ;
      LAYER met3 ;
        RECT 50.000 388.080 456.000 391.440 ;
      LAYER met3 ;
        RECT 456.000 388.080 2830.165 391.440 ;
      LAYER met3 ;
        RECT 50.000 386.680 455.600 388.080 ;
      LAYER met3 ;
        RECT 455.600 386.680 2830.165 388.080 ;
      LAYER met3 ;
        RECT 50.000 383.320 456.000 386.680 ;
      LAYER met3 ;
        RECT 456.000 383.320 2830.165 386.680 ;
      LAYER met3 ;
        RECT 50.000 381.920 455.600 383.320 ;
      LAYER met3 ;
        RECT 455.600 381.920 2830.165 383.320 ;
      LAYER met3 ;
        RECT 50.000 379.240 456.000 381.920 ;
      LAYER met3 ;
        RECT 456.000 379.240 2830.165 381.920 ;
      LAYER met3 ;
        RECT 50.000 377.840 455.600 379.240 ;
      LAYER met3 ;
        RECT 455.600 377.840 2830.165 379.240 ;
      LAYER met3 ;
        RECT 50.000 374.480 456.000 377.840 ;
      LAYER met3 ;
        RECT 456.000 374.480 2830.165 377.840 ;
      LAYER met3 ;
        RECT 50.000 373.080 455.600 374.480 ;
      LAYER met3 ;
        RECT 455.600 373.080 2830.165 374.480 ;
      LAYER met3 ;
        RECT 50.000 370.400 456.000 373.080 ;
      LAYER met3 ;
        RECT 456.000 370.400 2830.165 373.080 ;
      LAYER met3 ;
        RECT 50.000 369.000 455.600 370.400 ;
      LAYER met3 ;
        RECT 455.600 369.000 2830.165 370.400 ;
      LAYER met3 ;
        RECT 50.000 365.640 456.000 369.000 ;
      LAYER met3 ;
        RECT 456.000 365.640 2830.165 369.000 ;
      LAYER met3 ;
        RECT 50.000 364.240 455.600 365.640 ;
      LAYER met3 ;
        RECT 455.600 364.240 2830.165 365.640 ;
      LAYER met3 ;
        RECT 50.000 361.560 456.000 364.240 ;
      LAYER met3 ;
        RECT 456.000 361.560 2830.165 364.240 ;
      LAYER met3 ;
        RECT 50.000 360.160 455.600 361.560 ;
      LAYER met3 ;
        RECT 455.600 360.160 2830.165 361.560 ;
      LAYER met3 ;
        RECT 50.000 356.800 456.000 360.160 ;
      LAYER met3 ;
        RECT 456.000 356.800 2830.165 360.160 ;
      LAYER met3 ;
        RECT 50.000 355.400 455.600 356.800 ;
      LAYER met3 ;
        RECT 455.600 355.400 2830.165 356.800 ;
      LAYER met3 ;
        RECT 50.000 352.040 456.000 355.400 ;
      LAYER met3 ;
        RECT 456.000 352.040 2830.165 355.400 ;
      LAYER met3 ;
        RECT 50.000 350.640 455.600 352.040 ;
      LAYER met3 ;
        RECT 455.600 350.640 2830.165 352.040 ;
      LAYER met3 ;
        RECT 50.000 347.960 456.000 350.640 ;
      LAYER met3 ;
        RECT 456.000 347.960 2830.165 350.640 ;
      LAYER met3 ;
        RECT 50.000 346.560 455.600 347.960 ;
      LAYER met3 ;
        RECT 455.600 346.560 2830.165 347.960 ;
      LAYER met3 ;
        RECT 50.000 343.200 456.000 346.560 ;
      LAYER met3 ;
        RECT 456.000 343.200 2830.165 346.560 ;
      LAYER met3 ;
        RECT 50.000 341.800 455.600 343.200 ;
      LAYER met3 ;
        RECT 455.600 341.800 2830.165 343.200 ;
      LAYER met3 ;
        RECT 50.000 339.120 456.000 341.800 ;
      LAYER met3 ;
        RECT 456.000 339.120 2830.165 341.800 ;
      LAYER met3 ;
        RECT 50.000 337.720 455.600 339.120 ;
      LAYER met3 ;
        RECT 455.600 337.720 2830.165 339.120 ;
      LAYER met3 ;
        RECT 50.000 334.360 456.000 337.720 ;
      LAYER met3 ;
        RECT 456.000 334.360 2830.165 337.720 ;
      LAYER met3 ;
        RECT 50.000 332.960 455.600 334.360 ;
      LAYER met3 ;
        RECT 455.600 332.960 2830.165 334.360 ;
      LAYER met3 ;
        RECT 50.000 330.280 456.000 332.960 ;
      LAYER met3 ;
        RECT 456.000 330.280 2830.165 332.960 ;
      LAYER met3 ;
        RECT 50.000 328.880 455.600 330.280 ;
      LAYER met3 ;
        RECT 455.600 328.880 2830.165 330.280 ;
      LAYER met3 ;
        RECT 50.000 328.240 456.000 328.880 ;
        RECT 50.400 326.840 456.000 328.240 ;
        RECT 50.000 325.520 456.000 326.840 ;
      LAYER met3 ;
        RECT 456.000 325.520 2830.165 328.880 ;
      LAYER met3 ;
        RECT 50.000 324.120 455.600 325.520 ;
      LAYER met3 ;
        RECT 455.600 324.120 2830.165 325.520 ;
      LAYER met3 ;
        RECT 50.000 320.760 456.000 324.120 ;
      LAYER met3 ;
        RECT 456.000 320.760 2830.165 324.120 ;
      LAYER met3 ;
        RECT 50.000 319.360 455.600 320.760 ;
      LAYER met3 ;
        RECT 455.600 319.360 2830.165 320.760 ;
      LAYER met3 ;
        RECT 50.000 316.680 456.000 319.360 ;
      LAYER met3 ;
        RECT 456.000 316.680 2830.165 319.360 ;
      LAYER met3 ;
        RECT 50.000 315.280 455.600 316.680 ;
      LAYER met3 ;
        RECT 455.600 315.280 2830.165 316.680 ;
      LAYER met3 ;
        RECT 50.000 311.920 456.000 315.280 ;
      LAYER met3 ;
        RECT 456.000 311.920 2830.165 315.280 ;
      LAYER met3 ;
        RECT 50.000 310.520 455.600 311.920 ;
      LAYER met3 ;
        RECT 455.600 310.520 2830.165 311.920 ;
      LAYER met3 ;
        RECT 50.000 307.840 456.000 310.520 ;
      LAYER met3 ;
        RECT 456.000 307.840 2830.165 310.520 ;
      LAYER met3 ;
        RECT 50.000 306.440 455.600 307.840 ;
      LAYER met3 ;
        RECT 455.600 306.440 2830.165 307.840 ;
      LAYER met3 ;
        RECT 50.000 303.080 456.000 306.440 ;
      LAYER met3 ;
        RECT 456.000 303.080 2830.165 306.440 ;
      LAYER met3 ;
        RECT 50.000 301.680 455.600 303.080 ;
      LAYER met3 ;
        RECT 455.600 301.680 2830.165 303.080 ;
      LAYER met3 ;
        RECT 50.000 298.320 456.000 301.680 ;
      LAYER met3 ;
        RECT 456.000 298.320 2830.165 301.680 ;
      LAYER met3 ;
        RECT 50.000 296.920 455.600 298.320 ;
      LAYER met3 ;
        RECT 455.600 296.920 2830.165 298.320 ;
      LAYER met3 ;
        RECT 50.000 294.240 456.000 296.920 ;
      LAYER met3 ;
        RECT 456.000 294.240 2830.165 296.920 ;
      LAYER met3 ;
        RECT 50.000 292.840 455.600 294.240 ;
      LAYER met3 ;
        RECT 455.600 292.840 2830.165 294.240 ;
      LAYER met3 ;
        RECT 50.000 289.480 456.000 292.840 ;
      LAYER met3 ;
        RECT 456.000 289.480 2830.165 292.840 ;
      LAYER met3 ;
        RECT 50.000 288.080 455.600 289.480 ;
      LAYER met3 ;
        RECT 455.600 288.080 2830.165 289.480 ;
      LAYER met3 ;
        RECT 50.000 285.400 456.000 288.080 ;
      LAYER met3 ;
        RECT 456.000 285.400 2830.165 288.080 ;
      LAYER met3 ;
        RECT 50.000 284.000 455.600 285.400 ;
      LAYER met3 ;
        RECT 455.600 284.000 2830.165 285.400 ;
      LAYER met3 ;
        RECT 50.000 280.640 456.000 284.000 ;
      LAYER met3 ;
        RECT 456.000 280.640 2830.165 284.000 ;
      LAYER met3 ;
        RECT 50.000 279.240 455.600 280.640 ;
      LAYER met3 ;
        RECT 455.600 279.240 2830.165 280.640 ;
      LAYER met3 ;
        RECT 50.000 276.560 456.000 279.240 ;
      LAYER met3 ;
        RECT 456.000 276.560 2830.165 279.240 ;
      LAYER met3 ;
        RECT 50.000 275.160 455.600 276.560 ;
      LAYER met3 ;
        RECT 455.600 275.160 2830.165 276.560 ;
      LAYER met3 ;
        RECT 50.000 271.800 456.000 275.160 ;
      LAYER met3 ;
        RECT 456.000 271.800 2830.165 275.160 ;
      LAYER met3 ;
        RECT 50.000 270.400 455.600 271.800 ;
      LAYER met3 ;
        RECT 455.600 270.400 2830.165 271.800 ;
      LAYER met3 ;
        RECT 50.000 267.040 456.000 270.400 ;
      LAYER met3 ;
        RECT 456.000 267.040 2830.165 270.400 ;
      LAYER met3 ;
        RECT 50.000 265.640 455.600 267.040 ;
      LAYER met3 ;
        RECT 455.600 265.640 2830.165 267.040 ;
      LAYER met3 ;
        RECT 50.000 262.960 456.000 265.640 ;
      LAYER met3 ;
        RECT 456.000 262.960 2830.165 265.640 ;
      LAYER met3 ;
        RECT 50.000 261.560 455.600 262.960 ;
      LAYER met3 ;
        RECT 455.600 261.560 2830.165 262.960 ;
      LAYER met3 ;
        RECT 50.000 258.200 456.000 261.560 ;
      LAYER met3 ;
        RECT 456.000 258.200 2830.165 261.560 ;
      LAYER met3 ;
        RECT 50.000 256.800 455.600 258.200 ;
      LAYER met3 ;
        RECT 455.600 256.800 2830.165 258.200 ;
      LAYER met3 ;
        RECT 50.000 254.120 456.000 256.800 ;
      LAYER met3 ;
        RECT 456.000 254.120 2830.165 256.800 ;
      LAYER met3 ;
        RECT 50.000 252.720 455.600 254.120 ;
      LAYER met3 ;
        RECT 455.600 252.720 2830.165 254.120 ;
      LAYER met3 ;
        RECT 50.000 249.360 456.000 252.720 ;
      LAYER met3 ;
        RECT 456.000 249.360 2830.165 252.720 ;
      LAYER met3 ;
        RECT 50.000 247.960 455.600 249.360 ;
      LAYER met3 ;
        RECT 455.600 247.960 2830.165 249.360 ;
      LAYER met3 ;
        RECT 50.000 245.280 456.000 247.960 ;
      LAYER met3 ;
        RECT 456.000 245.280 2830.165 247.960 ;
      LAYER met3 ;
        RECT 50.000 243.880 455.600 245.280 ;
      LAYER met3 ;
        RECT 455.600 243.880 2830.165 245.280 ;
      LAYER met3 ;
        RECT 50.000 240.520 456.000 243.880 ;
      LAYER met3 ;
        RECT 456.000 240.520 2830.165 243.880 ;
      LAYER met3 ;
        RECT 50.000 239.120 455.600 240.520 ;
      LAYER met3 ;
        RECT 455.600 239.120 2830.165 240.520 ;
      LAYER met3 ;
        RECT 50.000 235.760 456.000 239.120 ;
      LAYER met3 ;
        RECT 456.000 235.760 2830.165 239.120 ;
      LAYER met3 ;
        RECT 50.000 234.360 455.600 235.760 ;
      LAYER met3 ;
        RECT 455.600 234.360 2830.165 235.760 ;
      LAYER met3 ;
        RECT 50.000 231.680 456.000 234.360 ;
      LAYER met3 ;
        RECT 456.000 231.680 2830.165 234.360 ;
      LAYER met3 ;
        RECT 50.000 230.280 455.600 231.680 ;
      LAYER met3 ;
        RECT 455.600 230.280 2830.165 231.680 ;
      LAYER met3 ;
        RECT 50.000 226.920 456.000 230.280 ;
      LAYER met3 ;
        RECT 456.000 226.920 2830.165 230.280 ;
      LAYER met3 ;
        RECT 50.000 225.520 455.600 226.920 ;
      LAYER met3 ;
        RECT 455.600 225.520 2830.165 226.920 ;
      LAYER met3 ;
        RECT 50.000 222.840 456.000 225.520 ;
      LAYER met3 ;
        RECT 456.000 222.840 2830.165 225.520 ;
      LAYER met3 ;
        RECT 50.000 221.440 455.600 222.840 ;
      LAYER met3 ;
        RECT 455.600 221.440 2830.165 222.840 ;
      LAYER met3 ;
        RECT 50.000 218.080 456.000 221.440 ;
      LAYER met3 ;
        RECT 456.000 218.080 2830.165 221.440 ;
      LAYER met3 ;
        RECT 50.000 216.680 455.600 218.080 ;
      LAYER met3 ;
        RECT 455.600 216.680 2830.165 218.080 ;
      LAYER met3 ;
        RECT 50.000 213.320 456.000 216.680 ;
      LAYER met3 ;
        RECT 456.000 213.320 2830.165 216.680 ;
      LAYER met3 ;
        RECT 50.000 211.920 455.600 213.320 ;
      LAYER met3 ;
        RECT 455.600 211.920 2830.165 213.320 ;
      LAYER met3 ;
        RECT 50.000 209.240 456.000 211.920 ;
      LAYER met3 ;
        RECT 456.000 209.240 2830.165 211.920 ;
      LAYER met3 ;
        RECT 50.000 207.840 455.600 209.240 ;
      LAYER met3 ;
        RECT 455.600 207.840 2830.165 209.240 ;
      LAYER met3 ;
        RECT 50.000 204.480 456.000 207.840 ;
      LAYER met3 ;
        RECT 456.000 204.480 2830.165 207.840 ;
      LAYER met3 ;
        RECT 50.000 203.080 455.600 204.480 ;
      LAYER met3 ;
        RECT 455.600 203.080 2830.165 204.480 ;
      LAYER met3 ;
        RECT 50.000 200.400 456.000 203.080 ;
      LAYER met3 ;
        RECT 456.000 200.400 2830.165 203.080 ;
      LAYER met3 ;
        RECT 50.000 199.000 455.600 200.400 ;
      LAYER met3 ;
        RECT 455.600 199.000 2830.165 200.400 ;
      LAYER met3 ;
        RECT 50.000 195.640 456.000 199.000 ;
      LAYER met3 ;
        RECT 456.000 195.640 2830.165 199.000 ;
      LAYER met3 ;
        RECT 50.000 194.240 455.600 195.640 ;
      LAYER met3 ;
        RECT 455.600 194.240 2830.165 195.640 ;
      LAYER met3 ;
        RECT 50.000 191.560 456.000 194.240 ;
      LAYER met3 ;
        RECT 456.000 191.560 2830.165 194.240 ;
      LAYER met3 ;
        RECT 50.000 190.160 455.600 191.560 ;
      LAYER met3 ;
        RECT 455.600 190.160 2830.165 191.560 ;
      LAYER met3 ;
        RECT 50.000 186.800 456.000 190.160 ;
      LAYER met3 ;
        RECT 456.000 186.800 2830.165 190.160 ;
      LAYER met3 ;
        RECT 50.000 185.400 455.600 186.800 ;
      LAYER met3 ;
        RECT 455.600 185.400 2830.165 186.800 ;
      LAYER met3 ;
        RECT 50.000 182.040 456.000 185.400 ;
      LAYER met3 ;
        RECT 456.000 182.040 2830.165 185.400 ;
      LAYER met3 ;
        RECT 50.000 180.640 455.600 182.040 ;
      LAYER met3 ;
        RECT 455.600 180.640 2830.165 182.040 ;
      LAYER met3 ;
        RECT 50.000 177.960 456.000 180.640 ;
      LAYER met3 ;
        RECT 456.000 177.960 2830.165 180.640 ;
      LAYER met3 ;
        RECT 50.000 176.560 455.600 177.960 ;
      LAYER met3 ;
        RECT 455.600 176.560 2830.165 177.960 ;
      LAYER met3 ;
        RECT 50.000 173.200 456.000 176.560 ;
      LAYER met3 ;
        RECT 456.000 173.200 2830.165 176.560 ;
      LAYER met3 ;
        RECT 50.000 171.800 455.600 173.200 ;
      LAYER met3 ;
        RECT 455.600 171.800 2830.165 173.200 ;
      LAYER met3 ;
        RECT 50.000 169.120 456.000 171.800 ;
      LAYER met3 ;
        RECT 456.000 169.120 2830.165 171.800 ;
      LAYER met3 ;
        RECT 50.000 167.720 455.600 169.120 ;
      LAYER met3 ;
        RECT 455.600 167.720 2830.165 169.120 ;
      LAYER met3 ;
        RECT 50.000 164.360 456.000 167.720 ;
      LAYER met3 ;
        RECT 456.000 164.360 2830.165 167.720 ;
      LAYER met3 ;
        RECT 50.000 162.960 455.600 164.360 ;
      LAYER met3 ;
        RECT 455.600 162.960 2830.165 164.360 ;
      LAYER met3 ;
        RECT 50.000 160.280 456.000 162.960 ;
      LAYER met3 ;
        RECT 456.000 160.280 2830.165 162.960 ;
      LAYER met3 ;
        RECT 50.000 159.415 455.600 160.280 ;
      LAYER met3 ;
        RECT 455.600 159.415 2830.165 160.280 ;
        RECT 54.000 57.975 2830.165 159.415 ;
      LAYER met4 ;
        RECT 67.040 54.000 2797.020 3466.000 ;
      LAYER met5 ;
        RECT 54.000 99.370 2866.000 3432.390 ;
  END
END user_project_wrapper
END LIBRARY

