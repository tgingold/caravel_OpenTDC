magic
tech sky130A
magscale 1 2
timestamp 1607276359
<< locali >>
rect 28457 42687 28491 42857
rect 28457 42551 28491 42653
rect 37565 42551 37599 42721
rect 16497 41667 16531 41769
rect 62773 40919 62807 41021
rect 29101 40443 29135 40613
rect 41061 38743 41095 38981
rect 43361 38743 43395 38981
rect 15117 38403 15151 38505
rect 30573 38199 30607 38505
rect 23489 37655 23523 37893
rect 56977 37655 57011 37961
rect 61209 36771 61243 36873
rect 16405 36023 16439 36125
rect 45569 36023 45603 36125
rect 51825 36091 51859 36193
rect 40325 35479 40359 35649
rect 57161 35479 57195 35649
rect 63693 35479 63727 35785
rect 79149 35479 79183 35717
rect 79609 35615 79643 35785
rect 32873 34935 32907 35173
rect 65533 35003 65567 35105
rect 79609 34527 79643 34629
rect 29377 33643 29411 33949
rect 30573 33439 30607 34017
rect 56609 33915 56643 34153
rect 13461 32827 13495 32929
rect 57989 32487 58023 32589
rect 57977 32453 58023 32487
rect 72433 32147 72467 32453
rect 86877 31603 86911 31773
rect 9597 31195 9631 31433
rect 37289 31127 37323 31433
rect 46857 31127 46891 31433
rect 46889 31093 46891 31127
rect 48145 31229 48329 31263
rect 48145 31127 48179 31229
rect 48237 31059 48271 31093
rect 48421 31059 48455 31161
rect 48237 31025 48455 31059
rect 17693 30107 17727 30277
rect 59277 27659 59311 31569
rect 59553 27931 59587 31297
rect 87337 30855 87371 31161
rect 96537 30991 96571 31161
rect 99331 30957 99389 30991
rect 23213 27319 23247 27489
rect 28365 24123 28399 24293
rect 15117 21879 15151 21981
rect 15301 19703 15335 19873
rect 19533 18071 19567 18173
rect 26157 13311 26191 13481
rect 16037 12087 16071 12189
rect 18245 11135 18279 11305
<< viali >>
rect 6101 43877 6135 43911
rect 6285 43877 6319 43911
rect 4629 43809 4663 43843
rect 5181 43809 5215 43843
rect 5365 43809 5399 43843
rect 18889 43809 18923 43843
rect 24225 43809 24259 43843
rect 24777 43809 24811 43843
rect 24961 43809 24995 43843
rect 38485 43809 38519 43843
rect 39037 43809 39071 43843
rect 39221 43809 39255 43843
rect 47317 43809 47351 43843
rect 48513 43809 48547 43843
rect 49709 43809 49743 43843
rect 49893 43809 49927 43843
rect 61945 43809 61979 43843
rect 62037 43809 62071 43843
rect 69673 43809 69707 43843
rect 69949 43809 69983 43843
rect 4537 43741 4571 43775
rect 24041 43741 24075 43775
rect 25329 43741 25363 43775
rect 38301 43741 38335 43775
rect 48605 43741 48639 43775
rect 5549 43673 5583 43707
rect 18981 43673 19015 43707
rect 39405 43673 39439 43707
rect 61761 43673 61795 43707
rect 62589 43673 62623 43707
rect 6009 43605 6043 43639
rect 23857 43605 23891 43639
rect 25605 43605 25639 43639
rect 37841 43605 37875 43639
rect 38025 43605 38059 43639
rect 47409 43605 47443 43639
rect 49985 43605 50019 43639
rect 62221 43605 62255 43639
rect 69765 43605 69799 43639
rect 19441 43401 19475 43435
rect 36829 43401 36863 43435
rect 37013 43401 37047 43435
rect 49433 43401 49467 43435
rect 70501 43401 70535 43435
rect 50629 43333 50663 43367
rect 66269 43333 66303 43367
rect 3709 43265 3743 43299
rect 24961 43265 24995 43299
rect 32597 43265 32631 43299
rect 37197 43265 37231 43299
rect 46765 43265 46799 43299
rect 59277 43265 59311 43299
rect 3985 43197 4019 43231
rect 6837 43197 6871 43231
rect 9880 43197 9914 43231
rect 10149 43197 10183 43231
rect 18061 43197 18095 43231
rect 18337 43197 18371 43231
rect 23673 43197 23707 43231
rect 23857 43197 23891 43231
rect 24409 43197 24443 43231
rect 24593 43197 24627 43231
rect 26709 43197 26743 43231
rect 26985 43197 27019 43231
rect 32321 43197 32355 43231
rect 37381 43197 37415 43231
rect 37841 43197 37875 43231
rect 37933 43197 37967 43231
rect 40509 43197 40543 43231
rect 42349 43197 42383 43231
rect 42625 43197 42659 43231
rect 46489 43197 46523 43231
rect 48329 43197 48363 43231
rect 49065 43197 49099 43231
rect 49249 43197 49283 43231
rect 50537 43197 50571 43231
rect 55781 43197 55815 43231
rect 56057 43197 56091 43231
rect 56241 43197 56275 43231
rect 59553 43197 59587 43231
rect 66177 43197 66211 43231
rect 66545 43197 66579 43231
rect 66913 43197 66947 43231
rect 69121 43197 69155 43231
rect 69397 43197 69431 43231
rect 5549 43129 5583 43163
rect 11529 43129 11563 43163
rect 28365 43129 28399 43163
rect 33977 43129 34011 43163
rect 38485 43129 38519 43163
rect 42165 43129 42199 43163
rect 49157 43129 49191 43163
rect 55229 43129 55263 43163
rect 67189 43129 67223 43163
rect 5273 43061 5307 43095
rect 6929 43061 6963 43095
rect 11713 43061 11747 43095
rect 19809 43061 19843 43095
rect 23489 43061 23523 43095
rect 25237 43061 25271 43095
rect 26525 43061 26559 43095
rect 34161 43061 34195 43095
rect 40693 43061 40727 43095
rect 43729 43061 43763 43095
rect 47869 43061 47903 43095
rect 49893 43061 49927 43095
rect 60841 43061 60875 43095
rect 61117 43061 61151 43095
rect 67373 43061 67407 43095
rect 69029 43061 69063 43095
rect 6653 42857 6687 42891
rect 28457 42857 28491 42891
rect 40417 42857 40451 42891
rect 49433 42857 49467 42891
rect 50813 42857 50847 42891
rect 57345 42857 57379 42891
rect 6469 42789 6503 42823
rect 4813 42721 4847 42755
rect 5089 42721 5123 42755
rect 10425 42721 10459 42755
rect 12081 42721 12115 42755
rect 12909 42721 12943 42755
rect 15393 42721 15427 42755
rect 15669 42721 15703 42755
rect 16221 42721 16255 42755
rect 16405 42721 16439 42755
rect 23949 42721 23983 42755
rect 24501 42721 24535 42755
rect 24685 42721 24719 42755
rect 29009 42721 29043 42755
rect 32965 42721 32999 42755
rect 34345 42721 34379 42755
rect 35173 42721 35207 42755
rect 37473 42721 37507 42755
rect 37565 42721 37599 42755
rect 43361 42721 43395 42755
rect 45293 42721 45327 42755
rect 45385 42721 45419 42755
rect 47501 42721 47535 42755
rect 47685 42721 47719 42755
rect 48053 42721 48087 42755
rect 48973 42721 49007 42755
rect 49249 42721 49283 42755
rect 50537 42721 50571 42755
rect 50721 42721 50755 42755
rect 57437 42721 57471 42755
rect 57805 42721 57839 42755
rect 58081 42721 58115 42755
rect 60289 42721 60323 42755
rect 61577 42721 61611 42755
rect 69029 42721 69063 42755
rect 69213 42721 69247 42755
rect 69305 42721 69339 42755
rect 71421 42721 71455 42755
rect 10701 42653 10735 42687
rect 12265 42653 12299 42687
rect 15117 42653 15151 42687
rect 15485 42653 15519 42687
rect 16773 42653 16807 42687
rect 17049 42653 17083 42687
rect 17693 42653 17727 42687
rect 17969 42653 18003 42687
rect 19349 42653 19383 42687
rect 23673 42653 23707 42687
rect 23857 42653 23891 42687
rect 25053 42653 25087 42687
rect 28457 42653 28491 42687
rect 28733 42653 28767 42687
rect 30389 42653 30423 42687
rect 32689 42653 32723 42687
rect 34529 42653 34563 42687
rect 25329 42585 25363 42619
rect 39037 42653 39071 42687
rect 39313 42653 39347 42687
rect 43453 42653 43487 42687
rect 45845 42653 45879 42687
rect 54769 42653 54803 42687
rect 55045 42653 55079 42687
rect 56517 42653 56551 42687
rect 61301 42653 61335 42687
rect 63141 42653 63175 42687
rect 65809 42653 65843 42687
rect 66085 42653 66119 42687
rect 69857 42653 69891 42687
rect 49065 42585 49099 42619
rect 67649 42585 67683 42619
rect 13001 42517 13035 42551
rect 19441 42517 19475 42551
rect 23305 42517 23339 42551
rect 23397 42517 23431 42551
rect 28457 42517 28491 42551
rect 28549 42517 28583 42551
rect 35265 42517 35299 42551
rect 37289 42517 37323 42551
rect 37565 42517 37599 42551
rect 37841 42517 37875 42551
rect 38945 42517 38979 42551
rect 45109 42517 45143 42551
rect 46029 42517 46063 42551
rect 56149 42517 56183 42551
rect 58541 42517 58575 42551
rect 60381 42517 60415 42551
rect 62681 42517 62715 42551
rect 67189 42517 67223 42551
rect 69489 42517 69523 42551
rect 71513 42517 71547 42551
rect 2421 42313 2455 42347
rect 4445 42313 4479 42347
rect 23121 42313 23155 42347
rect 23305 42313 23339 42347
rect 63049 42313 63083 42347
rect 69305 42313 69339 42347
rect 10793 42245 10827 42279
rect 22937 42245 22971 42279
rect 29469 42245 29503 42279
rect 29653 42245 29687 42279
rect 44097 42245 44131 42279
rect 59369 42245 59403 42279
rect 2605 42177 2639 42211
rect 15761 42177 15795 42211
rect 17233 42177 17267 42211
rect 17509 42177 17543 42211
rect 18797 42177 18831 42211
rect 19441 42177 19475 42211
rect 23673 42177 23707 42211
rect 24961 42177 24995 42211
rect 29837 42177 29871 42211
rect 36277 42177 36311 42211
rect 44741 42177 44775 42211
rect 45293 42177 45327 42211
rect 48053 42177 48087 42211
rect 51733 42177 51767 42211
rect 53481 42177 53515 42211
rect 60565 42177 60599 42211
rect 61945 42177 61979 42211
rect 65809 42177 65843 42211
rect 66361 42177 66395 42211
rect 70777 42177 70811 42211
rect 70869 42177 70903 42211
rect 2881 42109 2915 42143
rect 5273 42109 5307 42143
rect 9689 42109 9723 42143
rect 9858 42109 9892 42143
rect 10425 42109 10459 42143
rect 10600 42109 10634 42143
rect 12441 42109 12475 42143
rect 16405 42109 16439 42143
rect 16589 42109 16623 42143
rect 16957 42109 16991 42143
rect 17049 42109 17083 42143
rect 18705 42109 18739 42143
rect 19073 42109 19107 42143
rect 19257 42109 19291 42143
rect 20085 42109 20119 42143
rect 23857 42109 23891 42143
rect 24409 42109 24443 42143
rect 24593 42109 24627 42143
rect 25973 42109 26007 42143
rect 26157 42109 26191 42143
rect 26617 42109 26651 42143
rect 26709 42109 26743 42143
rect 27445 42109 27479 42143
rect 27629 42109 27663 42143
rect 30021 42109 30055 42143
rect 30481 42109 30515 42143
rect 30573 42109 30607 42143
rect 31309 42109 31343 42143
rect 31493 42109 31527 42143
rect 34897 42109 34931 42143
rect 36461 42109 36495 42143
rect 36645 42109 36679 42143
rect 37105 42109 37139 42143
rect 37197 42109 37231 42143
rect 44649 42109 44683 42143
rect 45017 42109 45051 42143
rect 45109 42109 45143 42143
rect 46121 42109 46155 42143
rect 48697 42109 48731 42143
rect 48789 42109 48823 42143
rect 49065 42109 49099 42143
rect 49249 42109 49283 42143
rect 52009 42109 52043 42143
rect 54953 42109 54987 42143
rect 55965 42109 55999 42143
rect 56241 42109 56275 42143
rect 59737 42109 59771 42143
rect 60105 42109 60139 42143
rect 61485 42109 61519 42143
rect 61670 42109 61704 42143
rect 62957 42109 62991 42143
rect 63509 42109 63543 42143
rect 66637 42109 66671 42143
rect 66821 42109 66855 42143
rect 69489 42109 69523 42143
rect 69765 42109 69799 42143
rect 71145 42109 71179 42143
rect 15945 42041 15979 42075
rect 18061 42041 18095 42075
rect 20177 42041 20211 42075
rect 25605 42041 25639 42075
rect 25789 42041 25823 42075
rect 27261 42041 27295 42075
rect 31125 42041 31159 42075
rect 36093 42041 36127 42075
rect 37749 42041 37783 42075
rect 46213 42041 46247 42075
rect 49433 42041 49467 42075
rect 55045 42041 55079 42075
rect 66913 42041 66947 42075
rect 3985 41973 4019 42007
rect 5365 41973 5399 42007
rect 9505 41973 9539 42007
rect 11253 41973 11287 42007
rect 12541 41973 12575 42007
rect 15577 41973 15611 42007
rect 17601 41973 17635 42007
rect 17785 41973 17819 42007
rect 19625 41973 19659 42007
rect 25237 41973 25271 42007
rect 34989 41973 35023 42007
rect 38025 41973 38059 42007
rect 43821 41973 43855 42007
rect 53113 41973 53147 42007
rect 56057 41973 56091 42007
rect 59645 41973 59679 42007
rect 60841 41973 60875 42007
rect 72249 41973 72283 42007
rect 5273 41769 5307 41803
rect 10885 41769 10919 41803
rect 11253 41769 11287 41803
rect 16497 41769 16531 41803
rect 16589 41769 16623 41803
rect 17969 41769 18003 41803
rect 18337 41769 18371 41803
rect 44557 41769 44591 41803
rect 49065 41769 49099 41803
rect 51733 41769 51767 41803
rect 54217 41769 54251 41803
rect 59185 41769 59219 41803
rect 59921 41769 59955 41803
rect 63877 41769 63911 41803
rect 9413 41701 9447 41735
rect 36921 41701 36955 41735
rect 43361 41701 43395 41735
rect 59369 41701 59403 41735
rect 60197 41701 60231 41735
rect 4261 41633 4295 41667
rect 4353 41633 4387 41667
rect 4813 41633 4847 41667
rect 4997 41633 5031 41667
rect 7297 41633 7331 41667
rect 8033 41633 8067 41667
rect 8217 41633 8251 41667
rect 8585 41633 8619 41667
rect 8769 41633 8803 41667
rect 9689 41633 9723 41667
rect 9873 41633 9907 41667
rect 10425 41633 10459 41667
rect 10609 41633 10643 41667
rect 14013 41633 14047 41667
rect 16497 41633 16531 41667
rect 16773 41633 16807 41667
rect 16957 41633 16991 41667
rect 17509 41633 17543 41667
rect 17693 41633 17727 41667
rect 24041 41633 24075 41667
rect 24501 41633 24535 41667
rect 24593 41633 24627 41667
rect 25421 41633 25455 41667
rect 26249 41633 26283 41667
rect 29837 41633 29871 41667
rect 30849 41633 30883 41667
rect 35449 41633 35483 41667
rect 35633 41633 35667 41667
rect 36185 41633 36219 41667
rect 36369 41633 36403 41667
rect 37933 41633 37967 41667
rect 38393 41633 38427 41667
rect 38485 41633 38519 41667
rect 43545 41633 43579 41667
rect 43913 41633 43947 41667
rect 45017 41633 45051 41667
rect 48973 41633 49007 41667
rect 49249 41633 49283 41667
rect 51641 41633 51675 41667
rect 53113 41633 53147 41667
rect 54401 41633 54435 41667
rect 54585 41633 54619 41667
rect 59001 41633 59035 41667
rect 60749 41633 60783 41667
rect 61025 41633 61059 41667
rect 61209 41633 61243 41667
rect 62037 41633 62071 41667
rect 63601 41633 63635 41667
rect 63785 41633 63819 41667
rect 65809 41633 65843 41667
rect 66177 41633 66211 41667
rect 67005 41633 67039 41667
rect 68477 41633 68511 41667
rect 68661 41633 68695 41667
rect 69029 41633 69063 41667
rect 69857 41633 69891 41667
rect 70041 41633 70075 41667
rect 71421 41633 71455 41667
rect 7573 41565 7607 41599
rect 23857 41565 23891 41599
rect 25145 41565 25179 41599
rect 29929 41565 29963 41599
rect 37289 41565 37323 41599
rect 37749 41565 37783 41599
rect 39313 41565 39347 41599
rect 44741 41565 44775 41599
rect 54033 41565 54067 41599
rect 54953 41565 54987 41599
rect 61853 41565 61887 41599
rect 62405 41565 62439 41599
rect 67097 41565 67131 41599
rect 70317 41565 70351 41599
rect 77953 41565 77987 41599
rect 78229 41565 78263 41599
rect 5641 41497 5675 41531
rect 7481 41497 7515 41531
rect 8953 41497 8987 41531
rect 23673 41497 23707 41531
rect 26065 41497 26099 41531
rect 30941 41497 30975 41531
rect 36645 41497 36679 41531
rect 38853 41497 38887 41531
rect 55045 41497 55079 41531
rect 62175 41497 62209 41531
rect 62313 41497 62347 41531
rect 9137 41429 9171 41463
rect 11345 41429 11379 41463
rect 11529 41429 11563 41463
rect 13829 41429 13863 41463
rect 14197 41429 14231 41463
rect 18521 41429 18555 41463
rect 23581 41429 23615 41463
rect 25513 41429 25547 41463
rect 37473 41429 37507 41463
rect 46121 41429 46155 41463
rect 53205 41429 53239 41463
rect 54723 41429 54757 41463
rect 54861 41429 54895 41463
rect 55505 41429 55539 41463
rect 62681 41429 62715 41463
rect 65993 41429 66027 41463
rect 71605 41429 71639 41463
rect 77861 41429 77895 41463
rect 79517 41429 79551 41463
rect 10241 41225 10275 41259
rect 10793 41225 10827 41259
rect 18245 41225 18279 41259
rect 19349 41225 19383 41259
rect 23765 41225 23799 41259
rect 29837 41225 29871 41259
rect 31677 41225 31711 41259
rect 44925 41225 44959 41259
rect 52009 41225 52043 41259
rect 63877 41225 63911 41259
rect 68109 41225 68143 41259
rect 68707 41225 68741 41259
rect 68845 41225 68879 41259
rect 10425 41157 10459 41191
rect 27261 41157 27295 41191
rect 27537 41157 27571 41191
rect 38393 41157 38427 41191
rect 60841 41157 60875 41191
rect 63049 41157 63083 41191
rect 71237 41157 71271 41191
rect 3157 41089 3191 41123
rect 9597 41089 9631 41123
rect 12449 41089 12483 41123
rect 25697 41089 25731 41123
rect 30113 41089 30147 41123
rect 35909 41089 35943 41123
rect 37197 41089 37231 41123
rect 38264 41089 38298 41123
rect 38485 41089 38519 41123
rect 68937 41089 68971 41123
rect 70409 41089 70443 41123
rect 71145 41089 71179 41123
rect 72433 41089 72467 41123
rect 78321 41089 78355 41123
rect 3433 41021 3467 41055
rect 3525 41021 3559 41055
rect 3893 41021 3927 41055
rect 3985 41021 4019 41055
rect 5457 41021 5491 41055
rect 9505 41021 9539 41055
rect 9873 41021 9907 41055
rect 10057 41021 10091 41055
rect 12725 41021 12759 41055
rect 18061 41021 18095 41055
rect 18429 41021 18463 41055
rect 19165 41021 19199 41055
rect 19533 41021 19567 41055
rect 23949 41021 23983 41055
rect 24133 41021 24167 41055
rect 24593 41021 24627 41055
rect 24685 41021 24719 41055
rect 26341 41021 26375 41055
rect 27445 41021 27479 41055
rect 30205 41021 30239 41055
rect 30665 41021 30699 41055
rect 30757 41021 30791 41055
rect 36093 41021 36127 41055
rect 36553 41021 36587 41055
rect 36645 41021 36679 41055
rect 38117 41021 38151 41055
rect 43177 41021 43211 41055
rect 44833 41021 44867 41055
rect 52561 41021 52595 41055
rect 52653 41021 52687 41055
rect 52929 41021 52963 41055
rect 53113 41021 53147 41055
rect 54125 41021 54159 41055
rect 54493 41021 54527 41055
rect 55505 41021 55539 41055
rect 60749 41021 60783 41055
rect 61025 41021 61059 41055
rect 61761 41021 61795 41055
rect 62773 41021 62807 41055
rect 62957 41021 62991 41055
rect 63233 41021 63267 41055
rect 64705 41021 64739 41055
rect 68569 41021 68603 41055
rect 70685 41021 70719 41055
rect 72157 41021 72191 41055
rect 77125 41021 77159 41055
rect 77677 41021 77711 41055
rect 77953 41021 77987 41055
rect 79793 41021 79827 41055
rect 4537 40953 4571 40987
rect 4997 40953 5031 40987
rect 5181 40953 5215 40987
rect 8861 40953 8895 40987
rect 31309 40953 31343 40987
rect 38853 40953 38887 40987
rect 44649 40953 44683 40987
rect 53941 40953 53975 40987
rect 55321 40953 55355 40987
rect 55873 40953 55907 40987
rect 69305 40953 69339 40987
rect 70593 40953 70627 40987
rect 71973 40953 72007 40987
rect 4813 40885 4847 40919
rect 5549 40885 5583 40919
rect 10517 40885 10551 40919
rect 14013 40885 14047 40919
rect 14289 40885 14323 40919
rect 25145 40885 25179 40919
rect 25513 40885 25547 40919
rect 26157 40885 26191 40919
rect 31493 40885 31527 40919
rect 37473 40885 37507 40919
rect 43269 40885 43303 40919
rect 44465 40885 44499 40919
rect 53297 40885 53331 40919
rect 55965 40885 55999 40919
rect 61577 40885 61611 40919
rect 61853 40885 61887 40919
rect 62773 40885 62807 40919
rect 63417 40885 63451 40919
rect 64337 40885 64371 40919
rect 64521 40885 64555 40919
rect 68385 40885 68419 40919
rect 71789 40885 71823 40919
rect 76941 40885 76975 40919
rect 77217 40885 77251 40919
rect 79885 40885 79919 40919
rect 12725 40681 12759 40715
rect 13737 40681 13771 40715
rect 36185 40681 36219 40715
rect 38945 40681 38979 40715
rect 72525 40681 72559 40715
rect 78689 40681 78723 40715
rect 27352 40613 27386 40647
rect 29101 40613 29135 40647
rect 34621 40613 34655 40647
rect 38301 40613 38335 40647
rect 41061 40613 41095 40647
rect 43729 40613 43763 40647
rect 44833 40613 44867 40647
rect 45385 40613 45419 40647
rect 57069 40613 57103 40647
rect 60749 40613 60783 40647
rect 63877 40613 63911 40647
rect 64613 40613 64647 40647
rect 69581 40613 69615 40647
rect 70225 40613 70259 40647
rect 77033 40613 77067 40647
rect 4813 40545 4847 40579
rect 6653 40545 6687 40579
rect 10885 40545 10919 40579
rect 13369 40545 13403 40579
rect 16957 40545 16991 40579
rect 24041 40545 24075 40579
rect 24501 40545 24535 40579
rect 24593 40545 24627 40579
rect 27500 40545 27534 40579
rect 5089 40477 5123 40511
rect 11161 40477 11195 40511
rect 12541 40477 12575 40511
rect 16681 40477 16715 40511
rect 23857 40477 23891 40511
rect 25145 40477 25179 40511
rect 27721 40477 27755 40511
rect 28089 40477 28123 40511
rect 29193 40545 29227 40579
rect 29377 40545 29411 40579
rect 29561 40545 29595 40579
rect 30021 40545 30055 40579
rect 30113 40545 30147 40579
rect 34989 40545 35023 40579
rect 35173 40545 35207 40579
rect 35633 40545 35667 40579
rect 35725 40545 35759 40579
rect 36461 40545 36495 40579
rect 43637 40545 43671 40579
rect 45017 40545 45051 40579
rect 52009 40545 52043 40579
rect 52285 40545 52319 40579
rect 53021 40545 53055 40579
rect 53205 40545 53239 40579
rect 55321 40545 55355 40579
rect 55873 40545 55907 40579
rect 56149 40545 56183 40579
rect 57161 40545 57195 40579
rect 60657 40545 60691 40579
rect 61669 40545 61703 40579
rect 62313 40545 62347 40579
rect 62405 40545 62439 40579
rect 62647 40545 62681 40579
rect 62865 40545 62899 40579
rect 63969 40545 64003 40579
rect 64429 40545 64463 40579
rect 66729 40545 66763 40579
rect 68477 40545 68511 40579
rect 69765 40545 69799 40579
rect 71421 40545 71455 40579
rect 72617 40545 72651 40579
rect 77585 40545 77619 40579
rect 77861 40545 77895 40579
rect 78045 40545 78079 40579
rect 78137 40545 78171 40579
rect 78873 40545 78907 40579
rect 83197 40545 83231 40579
rect 83381 40545 83415 40579
rect 30665 40477 30699 40511
rect 38669 40477 38703 40511
rect 41429 40477 41463 40511
rect 41521 40477 41555 40511
rect 52101 40477 52135 40511
rect 55689 40477 55723 40511
rect 63693 40477 63727 40511
rect 72893 40477 72927 40511
rect 79149 40477 79183 40511
rect 83657 40477 83691 40511
rect 25421 40409 25455 40443
rect 29101 40409 29135 40443
rect 30941 40409 30975 40443
rect 66545 40409 66579 40443
rect 6193 40341 6227 40375
rect 13461 40341 13495 40375
rect 18245 40341 18279 40375
rect 18429 40341 18463 40375
rect 23765 40341 23799 40375
rect 25605 40341 25639 40375
rect 27629 40341 27663 40375
rect 28273 40341 28307 40375
rect 31125 40341 31159 40375
rect 34805 40341 34839 40375
rect 36645 40341 36679 40375
rect 38439 40341 38473 40375
rect 38577 40341 38611 40375
rect 41199 40341 41233 40375
rect 41337 40341 41371 40375
rect 53297 40341 53331 40375
rect 56885 40341 56919 40375
rect 57345 40341 57379 40375
rect 57805 40341 57839 40375
rect 63049 40341 63083 40375
rect 68661 40341 68695 40375
rect 69397 40341 69431 40375
rect 69857 40341 69891 40375
rect 71513 40341 71547 40375
rect 73997 40341 74031 40375
rect 80253 40341 80287 40375
rect 84761 40341 84795 40375
rect 4445 40137 4479 40171
rect 6929 40137 6963 40171
rect 11161 40137 11195 40171
rect 35725 40137 35759 40171
rect 37197 40137 37231 40171
rect 39405 40137 39439 40171
rect 43867 40137 43901 40171
rect 52653 40137 52687 40171
rect 61577 40137 61611 40171
rect 78413 40137 78447 40171
rect 83933 40137 83967 40171
rect 4721 40069 4755 40103
rect 11529 40069 11563 40103
rect 11713 40069 11747 40103
rect 17785 40069 17819 40103
rect 19625 40069 19659 40103
rect 23213 40069 23247 40103
rect 25421 40069 25455 40103
rect 25789 40069 25823 40103
rect 27629 40069 27663 40103
rect 32873 40069 32907 40103
rect 35817 40069 35851 40103
rect 37933 40069 37967 40103
rect 44005 40069 44039 40103
rect 71605 40069 71639 40103
rect 3157 40001 3191 40035
rect 9965 40001 9999 40035
rect 17693 40001 17727 40035
rect 18797 40001 18831 40035
rect 19441 40001 19475 40035
rect 23673 40001 23707 40035
rect 25237 40001 25271 40035
rect 32137 40001 32171 40035
rect 32744 40001 32778 40035
rect 32965 40001 32999 40035
rect 36001 40001 36035 40035
rect 37749 40001 37783 40035
rect 42717 40001 42751 40035
rect 44097 40001 44131 40035
rect 48973 40001 49007 40035
rect 60197 40001 60231 40035
rect 61945 40001 61979 40035
rect 63969 40001 64003 40035
rect 65533 40001 65567 40035
rect 67281 40001 67315 40035
rect 69213 40001 69247 40035
rect 69949 40001 69983 40035
rect 70501 40001 70535 40035
rect 70777 40001 70811 40035
rect 74917 40001 74951 40035
rect 2881 39933 2915 39967
rect 5733 39933 5767 39967
rect 7105 39933 7139 39967
rect 10149 39933 10183 39967
rect 10701 39933 10735 39967
rect 10885 39933 10919 39967
rect 13093 39933 13127 39967
rect 18705 39933 18739 39967
rect 19073 39933 19107 39967
rect 19257 39933 19291 39967
rect 23857 39933 23891 39967
rect 24317 39933 24351 39967
rect 24409 39933 24443 39967
rect 25513 39933 25547 39967
rect 25881 39933 25915 39967
rect 26065 39933 26099 39967
rect 26525 39933 26559 39967
rect 26617 39933 26651 39967
rect 30573 39933 30607 39967
rect 30665 39933 30699 39967
rect 31033 39933 31067 39967
rect 31125 39933 31159 39967
rect 32597 39933 32631 39967
rect 33333 39933 33367 39967
rect 36139 39933 36173 39967
rect 36645 39933 36679 39967
rect 36737 39933 36771 39967
rect 37473 39933 37507 39967
rect 38209 39933 38243 39967
rect 38393 39933 38427 39967
rect 38853 39933 38887 39967
rect 38945 39933 38979 39967
rect 39681 39933 39715 39967
rect 41153 39933 41187 39967
rect 41337 39933 41371 39967
rect 41521 39933 41555 39967
rect 41705 39933 41739 39967
rect 42165 39933 42199 39967
rect 42257 39933 42291 39967
rect 43269 39933 43303 39967
rect 43453 39933 43487 39967
rect 47593 39933 47627 39967
rect 47685 39933 47719 39967
rect 48053 39933 48087 39967
rect 48145 39933 48179 39967
rect 49157 39933 49191 39967
rect 52377 39933 52411 39967
rect 52561 39933 52595 39967
rect 53757 39933 53791 39967
rect 54033 39933 54067 39967
rect 55505 39933 55539 39967
rect 60473 39933 60507 39967
rect 63693 39933 63727 39967
rect 67465 39933 67499 39967
rect 67557 39933 67591 39967
rect 70041 39933 70075 39967
rect 70409 39933 70443 39967
rect 71421 39933 71455 39967
rect 72893 39933 72927 39967
rect 74181 39933 74215 39967
rect 74365 39933 74399 39967
rect 74457 39933 74491 39967
rect 75837 39933 75871 39967
rect 76113 39933 76147 39967
rect 77033 39933 77067 39967
rect 78229 39933 78263 39967
rect 78597 39933 78631 39967
rect 79977 39933 80011 39967
rect 83841 39933 83875 39967
rect 85589 39933 85623 39967
rect 86049 39933 86083 39967
rect 23397 39865 23431 39899
rect 24961 39865 24995 39899
rect 27445 39865 27479 39899
rect 31677 39865 31711 39899
rect 33517 39865 33551 39899
rect 43729 39865 43763 39899
rect 47225 39865 47259 39899
rect 69397 39865 69431 39899
rect 76849 39865 76883 39899
rect 77401 39865 77435 39899
rect 85405 39865 85439 39899
rect 85957 39865 85991 39899
rect 5825 39797 5859 39831
rect 7205 39797 7239 39831
rect 9781 39797 9815 39831
rect 13277 39797 13311 39831
rect 13461 39797 13495 39831
rect 18153 39797 18187 39831
rect 27077 39797 27111 39831
rect 31861 39797 31895 39831
rect 38025 39797 38059 39831
rect 39957 39797 39991 39831
rect 43085 39797 43119 39831
rect 44373 39797 44407 39831
rect 48605 39797 48639 39831
rect 55137 39797 55171 39831
rect 65073 39797 65107 39831
rect 70961 39797 70995 39831
rect 73077 39797 73111 39831
rect 73905 39797 73939 39831
rect 75929 39797 75963 39831
rect 76665 39797 76699 39831
rect 80069 39797 80103 39831
rect 5641 39593 5675 39627
rect 34805 39593 34839 39627
rect 36829 39593 36863 39627
rect 79609 39593 79643 39627
rect 80805 39593 80839 39627
rect 86049 39593 86083 39627
rect 11989 39525 12023 39559
rect 13001 39525 13035 39559
rect 18981 39525 19015 39559
rect 26525 39525 26559 39559
rect 36461 39525 36495 39559
rect 42349 39525 42383 39559
rect 44649 39525 44683 39559
rect 52193 39525 52227 39559
rect 53113 39525 53147 39559
rect 55321 39525 55355 39559
rect 55505 39525 55539 39559
rect 61669 39525 61703 39559
rect 68477 39525 68511 39559
rect 83565 39525 83599 39559
rect 83749 39525 83783 39559
rect 85589 39525 85623 39559
rect 4629 39457 4663 39491
rect 5181 39457 5215 39491
rect 5365 39457 5399 39491
rect 10885 39457 10919 39491
rect 11437 39457 11471 39491
rect 11621 39457 11655 39491
rect 12909 39457 12943 39491
rect 16405 39457 16439 39491
rect 18889 39457 18923 39491
rect 23443 39457 23477 39491
rect 23581 39457 23615 39491
rect 23949 39457 23983 39491
rect 24041 39457 24075 39491
rect 24869 39457 24903 39491
rect 25053 39457 25087 39491
rect 29837 39457 29871 39491
rect 30297 39457 30331 39491
rect 30389 39457 30423 39491
rect 31401 39457 31435 39491
rect 35173 39457 35207 39491
rect 35357 39457 35391 39491
rect 35817 39457 35851 39491
rect 35909 39457 35943 39491
rect 41245 39457 41279 39491
rect 41705 39457 41739 39491
rect 41797 39457 41831 39491
rect 43545 39457 43579 39491
rect 44097 39457 44131 39491
rect 44281 39457 44315 39491
rect 44925 39457 44959 39491
rect 45109 39457 45143 39491
rect 48973 39457 49007 39491
rect 50721 39457 50755 39491
rect 52101 39457 52135 39491
rect 53297 39457 53331 39491
rect 53665 39457 53699 39491
rect 54769 39457 54803 39491
rect 54861 39457 54895 39491
rect 56425 39457 56459 39491
rect 61853 39457 61887 39491
rect 62221 39457 62255 39491
rect 63049 39457 63083 39491
rect 63233 39457 63267 39491
rect 64453 39457 64487 39491
rect 66729 39457 66763 39491
rect 67649 39457 67683 39491
rect 67925 39457 67959 39491
rect 68661 39457 68695 39491
rect 71421 39457 71455 39491
rect 75837 39457 75871 39491
rect 77217 39457 77251 39491
rect 78045 39457 78079 39491
rect 79149 39457 79183 39491
rect 79425 39457 79459 39491
rect 80713 39457 80747 39491
rect 84393 39457 84427 39491
rect 84761 39457 84795 39491
rect 84945 39457 84979 39491
rect 85773 39457 85807 39491
rect 85957 39457 85991 39491
rect 4445 39389 4479 39423
rect 10517 39389 10551 39423
rect 10701 39389 10735 39423
rect 12725 39389 12759 39423
rect 16681 39389 16715 39423
rect 23029 39389 23063 39423
rect 26893 39389 26927 39423
rect 27261 39389 27295 39423
rect 29745 39389 29779 39423
rect 31217 39389 31251 39423
rect 36645 39389 36679 39423
rect 41153 39389 41187 39423
rect 42809 39389 42843 39423
rect 43361 39389 43395 39423
rect 49249 39389 49283 39423
rect 56149 39389 56183 39423
rect 68937 39389 68971 39423
rect 71513 39389 71547 39423
rect 77364 39389 77398 39423
rect 77585 39389 77619 39423
rect 77953 39389 77987 39423
rect 79241 39389 79275 39423
rect 84301 39389 84335 39423
rect 6009 39321 6043 39355
rect 40877 39321 40911 39355
rect 64521 39321 64555 39355
rect 66545 39321 66579 39355
rect 76021 39321 76055 39355
rect 77493 39321 77527 39355
rect 4261 39253 4295 39287
rect 17969 39253 18003 39287
rect 18245 39253 18279 39287
rect 23213 39253 23247 39287
rect 24501 39253 24535 39287
rect 26663 39253 26697 39287
rect 26801 39253 26835 39287
rect 30849 39253 30883 39287
rect 34989 39253 35023 39287
rect 42533 39253 42567 39287
rect 42901 39253 42935 39287
rect 43085 39253 43119 39287
rect 50353 39253 50387 39287
rect 54585 39253 54619 39287
rect 55965 39253 55999 39287
rect 57529 39253 57563 39287
rect 63325 39253 63359 39287
rect 63785 39253 63819 39287
rect 67741 39253 67775 39287
rect 70041 39253 70075 39287
rect 76757 39253 76791 39287
rect 77125 39253 77159 39287
rect 83381 39253 83415 39287
rect 11713 39049 11747 39083
rect 15485 39049 15519 39083
rect 18153 39049 18187 39083
rect 29745 39049 29779 39083
rect 38209 39049 38243 39083
rect 54217 39049 54251 39083
rect 69029 39049 69063 39083
rect 70961 39049 70995 39083
rect 72617 39049 72651 39083
rect 75193 39049 75227 39083
rect 77217 39049 77251 39083
rect 83473 39049 83507 39083
rect 85497 39049 85531 39083
rect 15853 38981 15887 39015
rect 26019 38981 26053 39015
rect 26157 38981 26191 39015
rect 41061 38981 41095 39015
rect 19717 38913 19751 38947
rect 26249 38913 26283 38947
rect 37749 38913 37783 38947
rect 2697 38845 2731 38879
rect 2973 38845 3007 38879
rect 5273 38845 5307 38879
rect 5733 38845 5767 38879
rect 10793 38845 10827 38879
rect 10977 38845 11011 38879
rect 11345 38845 11379 38879
rect 11529 38845 11563 38879
rect 14427 38845 14461 38879
rect 14565 38845 14599 38879
rect 15025 38845 15059 38879
rect 15209 38845 15243 38879
rect 16589 38845 16623 38879
rect 16957 38845 16991 38879
rect 18061 38845 18095 38879
rect 19441 38845 19475 38879
rect 23673 38845 23707 38879
rect 23857 38845 23891 38879
rect 24409 38845 24443 38879
rect 24593 38845 24627 38879
rect 25237 38845 25271 38879
rect 25881 38845 25915 38879
rect 29653 38845 29687 38879
rect 36461 38845 36495 38879
rect 36645 38845 36679 38879
rect 37105 38845 37139 38879
rect 37197 38845 37231 38879
rect 10333 38777 10367 38811
rect 11805 38777 11839 38811
rect 14105 38777 14139 38811
rect 23489 38777 23523 38811
rect 24961 38777 24995 38811
rect 26617 38777 26651 38811
rect 43361 38981 43395 39015
rect 43545 38981 43579 39015
rect 43867 38981 43901 39015
rect 44005 38981 44039 39015
rect 44373 38981 44407 39015
rect 48881 38981 48915 39015
rect 49065 38981 49099 39015
rect 76849 38981 76883 39015
rect 80069 38981 80103 39015
rect 80989 38981 81023 39015
rect 42717 38913 42751 38947
rect 43085 38913 43119 38947
rect 41429 38845 41463 38879
rect 41521 38845 41555 38879
rect 41705 38845 41739 38879
rect 42165 38845 42199 38879
rect 42257 38845 42291 38879
rect 44097 38913 44131 38947
rect 47409 38913 47443 38947
rect 63785 38913 63819 38947
rect 64705 38913 64739 38947
rect 72341 38913 72375 38947
rect 74917 38913 74951 38947
rect 77677 38913 77711 38947
rect 79940 38913 79974 38947
rect 80158 38913 80192 38947
rect 83749 38913 83783 38947
rect 84117 38913 84151 38947
rect 43729 38845 43763 38879
rect 47501 38845 47535 38879
rect 47961 38845 47995 38879
rect 48053 38845 48087 38879
rect 52653 38845 52687 38879
rect 52837 38845 52871 38879
rect 53297 38845 53331 38879
rect 53389 38845 53423 38879
rect 55689 38845 55723 38879
rect 55781 38845 55815 38879
rect 56057 38845 56091 38879
rect 63233 38845 63267 38879
rect 63417 38845 63451 38879
rect 64613 38845 64647 38879
rect 68569 38845 68603 38879
rect 69673 38845 69707 38879
rect 70777 38845 70811 38879
rect 72249 38845 72283 38879
rect 75377 38845 75411 38879
rect 75653 38845 75687 38879
rect 77769 38845 77803 38879
rect 78137 38845 78171 38879
rect 78321 38845 78355 38879
rect 80805 38845 80839 38879
rect 83662 38845 83696 38879
rect 83933 38845 83967 38879
rect 84485 38845 84519 38879
rect 85405 38845 85439 38879
rect 86509 38845 86543 38879
rect 86785 38845 86819 38879
rect 54309 38777 54343 38811
rect 69489 38777 69523 38811
rect 79793 38777 79827 38811
rect 80621 38777 80655 38811
rect 4261 38709 4295 38743
rect 4445 38709 4479 38743
rect 5273 38709 5307 38743
rect 16773 38709 16807 38743
rect 20821 38709 20855 38743
rect 21189 38709 21223 38743
rect 25421 38709 25455 38743
rect 38025 38709 38059 38743
rect 41061 38709 41095 38743
rect 41153 38709 41187 38743
rect 43269 38709 43303 38743
rect 43361 38709 43395 38743
rect 47225 38709 47259 38743
rect 48513 38709 48547 38743
rect 53849 38709 53883 38743
rect 68753 38709 68787 38743
rect 69857 38709 69891 38743
rect 76941 38709 76975 38743
rect 80437 38709 80471 38743
rect 86417 38709 86451 38743
rect 87889 38709 87923 38743
rect 9965 38505 9999 38539
rect 13093 38505 13127 38539
rect 14933 38505 14967 38539
rect 15117 38505 15151 38539
rect 16497 38505 16531 38539
rect 16865 38505 16899 38539
rect 25421 38505 25455 38539
rect 29653 38505 29687 38539
rect 30573 38505 30607 38539
rect 53297 38505 53331 38539
rect 63785 38505 63819 38539
rect 69213 38505 69247 38539
rect 74641 38505 74675 38539
rect 84025 38505 84059 38539
rect 7481 38437 7515 38471
rect 10885 38437 10919 38471
rect 23581 38437 23615 38471
rect 24961 38437 24995 38471
rect 4353 38369 4387 38403
rect 6101 38369 6135 38403
rect 7297 38369 7331 38403
rect 8033 38369 8067 38403
rect 8217 38369 8251 38403
rect 8585 38369 8619 38403
rect 8769 38369 8803 38403
rect 9781 38369 9815 38403
rect 11529 38369 11563 38403
rect 11897 38369 11931 38403
rect 12081 38369 12115 38403
rect 12909 38369 12943 38403
rect 14749 38369 14783 38403
rect 15117 38369 15151 38403
rect 15485 38369 15519 38403
rect 15577 38369 15611 38403
rect 16037 38369 16071 38403
rect 16221 38369 16255 38403
rect 19717 38369 19751 38403
rect 23673 38369 23707 38403
rect 23857 38369 23891 38403
rect 24407 38369 24441 38403
rect 24593 38369 24627 38403
rect 4629 38301 4663 38335
rect 7573 38301 7607 38335
rect 11621 38301 11655 38335
rect 12265 38301 12299 38335
rect 25237 38301 25271 38335
rect 27905 38301 27939 38335
rect 28089 38301 28123 38335
rect 28365 38301 28399 38335
rect 12357 38233 12391 38267
rect 75561 38437 75595 38471
rect 77033 38437 77067 38471
rect 78597 38437 78631 38471
rect 86417 38437 86451 38471
rect 30665 38369 30699 38403
rect 33241 38369 33275 38403
rect 36553 38369 36587 38403
rect 37749 38369 37783 38403
rect 37933 38369 37967 38403
rect 38393 38369 38427 38403
rect 38485 38369 38519 38403
rect 39221 38369 39255 38403
rect 40877 38369 40911 38403
rect 47593 38369 47627 38403
rect 51917 38369 51951 38403
rect 52377 38369 52411 38403
rect 52469 38369 52503 38403
rect 60933 38369 60967 38403
rect 64153 38369 64187 38403
rect 64521 38369 64555 38403
rect 69397 38369 69431 38403
rect 70133 38369 70167 38403
rect 71421 38369 71455 38403
rect 74549 38369 74583 38403
rect 75745 38369 75779 38403
rect 76205 38369 76239 38403
rect 76757 38369 76791 38403
rect 78781 38369 78815 38403
rect 83565 38369 83599 38403
rect 83657 38369 83691 38403
rect 83841 38369 83875 38403
rect 85865 38369 85899 38403
rect 85957 38369 85991 38403
rect 36645 38301 36679 38335
rect 39037 38301 39071 38335
rect 41245 38301 41279 38335
rect 41613 38301 41647 38335
rect 51825 38301 51859 38335
rect 60657 38301 60691 38335
rect 63969 38301 64003 38335
rect 64429 38301 64463 38335
rect 65073 38301 65107 38335
rect 70317 38301 70351 38335
rect 76113 38301 76147 38335
rect 77401 38301 77435 38335
rect 77677 38301 77711 38335
rect 40693 38233 40727 38267
rect 69673 38233 69707 38267
rect 76389 38233 76423 38267
rect 77309 38233 77343 38267
rect 5733 38165 5767 38199
rect 19809 38165 19843 38199
rect 30573 38165 30607 38199
rect 30757 38165 30791 38199
rect 33057 38165 33091 38199
rect 39497 38165 39531 38199
rect 41015 38165 41049 38199
rect 41153 38165 41187 38199
rect 46305 38165 46339 38199
rect 47685 38165 47719 38199
rect 52929 38165 52963 38199
rect 53389 38165 53423 38199
rect 62221 38165 62255 38199
rect 64889 38165 64923 38199
rect 71605 38165 71639 38199
rect 76573 38165 76607 38199
rect 77171 38165 77205 38199
rect 78413 38165 78447 38199
rect 78873 38165 78907 38199
rect 83381 38165 83415 38199
rect 85681 38165 85715 38199
rect 3985 37961 4019 37995
rect 6101 37961 6135 37995
rect 14197 37961 14231 37995
rect 14473 37961 14507 37995
rect 20545 37961 20579 37995
rect 54861 37961 54895 37995
rect 56977 37961 57011 37995
rect 61853 37961 61887 37995
rect 65165 37961 65199 37995
rect 69121 37961 69155 37995
rect 72065 37961 72099 37995
rect 83841 37961 83875 37995
rect 86877 37961 86911 37995
rect 20821 37893 20855 37927
rect 23489 37893 23523 37927
rect 30665 37893 30699 37927
rect 31907 37893 31941 37927
rect 32045 37893 32079 37927
rect 35357 37893 35391 37927
rect 45845 37893 45879 37927
rect 47593 37893 47627 37927
rect 2605 37825 2639 37859
rect 17049 37825 17083 37859
rect 2881 37757 2915 37791
rect 5273 37757 5307 37791
rect 5733 37757 5767 37791
rect 6929 37757 6963 37791
rect 7389 37757 7423 37791
rect 10609 37757 10643 37791
rect 10793 37757 10827 37791
rect 11161 37757 11195 37791
rect 11345 37757 11379 37791
rect 14013 37757 14047 37791
rect 15761 37757 15795 37791
rect 15945 37757 15979 37791
rect 16405 37757 16439 37791
rect 16497 37757 16531 37791
rect 18981 37757 19015 37791
rect 19257 37757 19291 37791
rect 4445 37689 4479 37723
rect 10149 37689 10183 37723
rect 27077 37825 27111 37859
rect 29561 37825 29595 37859
rect 32137 37825 32171 37859
rect 35541 37825 35575 37859
rect 35817 37825 35851 37859
rect 38117 37825 38151 37859
rect 46121 37825 46155 37859
rect 54033 37825 54067 37859
rect 25973 37757 26007 37791
rect 26065 37757 26099 37791
rect 26525 37757 26559 37791
rect 26709 37757 26743 37791
rect 29292 37757 29326 37791
rect 32505 37757 32539 37791
rect 37197 37757 37231 37791
rect 38025 37757 38059 37791
rect 41981 37757 42015 37791
rect 42073 37757 42107 37791
rect 42441 37757 42475 37791
rect 42533 37757 42567 37791
rect 46397 37757 46431 37791
rect 46581 37757 46615 37791
rect 47133 37757 47167 37791
rect 47317 37757 47351 37791
rect 48605 37757 48639 37791
rect 52285 37757 52319 37791
rect 52561 37757 52595 37791
rect 53941 37757 53975 37791
rect 54769 37757 54803 37791
rect 31769 37689 31803 37723
rect 41705 37689 41739 37723
rect 43085 37689 43119 37723
rect 57345 37893 57379 37927
rect 57529 37893 57563 37927
rect 65717 37893 65751 37927
rect 57713 37825 57747 37859
rect 59001 37825 59035 37859
rect 60565 37825 60599 37859
rect 64061 37825 64095 37859
rect 64521 37825 64555 37859
rect 75745 37825 75779 37859
rect 78045 37825 78079 37859
rect 85865 37825 85899 37859
rect 57897 37757 57931 37791
rect 58449 37757 58483 37791
rect 58633 37757 58667 37791
rect 60289 37757 60323 37791
rect 64245 37757 64279 37791
rect 64613 37757 64647 37791
rect 65625 37757 65659 37791
rect 69305 37757 69339 37791
rect 69581 37757 69615 37791
rect 71973 37757 72007 37791
rect 75653 37757 75687 37791
rect 75929 37757 75963 37791
rect 76665 37757 76699 37791
rect 76941 37757 76975 37791
rect 82737 37757 82771 37791
rect 83749 37757 83783 37791
rect 84025 37757 84059 37791
rect 85405 37757 85439 37791
rect 85589 37757 85623 37791
rect 86049 37757 86083 37791
rect 86785 37757 86819 37791
rect 63601 37689 63635 37723
rect 64981 37689 65015 37723
rect 71789 37689 71823 37723
rect 4537 37621 4571 37655
rect 5273 37621 5307 37655
rect 6929 37621 6963 37655
rect 15577 37621 15611 37655
rect 17233 37621 17267 37655
rect 23489 37621 23523 37655
rect 25513 37621 25547 37655
rect 25697 37621 25731 37655
rect 31033 37621 31067 37655
rect 31585 37621 31619 37655
rect 41521 37621 41555 37655
rect 43361 37621 43395 37655
rect 48697 37621 48731 37655
rect 52101 37621 52135 37655
rect 56977 37621 57011 37655
rect 57069 37621 57103 37655
rect 70685 37621 70719 37655
rect 71605 37621 71639 37655
rect 76573 37621 76607 37655
rect 82829 37621 82863 37655
rect 6745 37417 6779 37451
rect 10057 37417 10091 37451
rect 11069 37417 11103 37451
rect 16497 37417 16531 37451
rect 19901 37417 19935 37451
rect 21097 37417 21131 37451
rect 26065 37417 26099 37451
rect 54309 37417 54343 37451
rect 57253 37417 57287 37451
rect 57437 37417 57471 37451
rect 57713 37417 57747 37451
rect 61853 37417 61887 37451
rect 63049 37417 63083 37451
rect 67189 37417 67223 37451
rect 67373 37417 67407 37451
rect 84485 37417 84519 37451
rect 15025 37349 15059 37383
rect 18797 37349 18831 37383
rect 27813 37349 27847 37383
rect 29837 37349 29871 37383
rect 36829 37349 36863 37383
rect 40233 37349 40267 37383
rect 41981 37349 42015 37383
rect 47961 37349 47995 37383
rect 49709 37349 49743 37383
rect 51549 37349 51583 37383
rect 69489 37349 69523 37383
rect 71145 37349 71179 37383
rect 77769 37349 77803 37383
rect 4997 37281 5031 37315
rect 5273 37281 5307 37315
rect 9873 37281 9907 37315
rect 11437 37281 11471 37315
rect 11621 37281 11655 37315
rect 11989 37281 12023 37315
rect 12173 37281 12207 37315
rect 15301 37281 15335 37315
rect 15485 37281 15519 37315
rect 16037 37281 16071 37315
rect 16221 37281 16255 37315
rect 16865 37281 16899 37315
rect 17693 37281 17727 37315
rect 18245 37281 18279 37315
rect 18429 37281 18463 37315
rect 19809 37281 19843 37315
rect 20913 37281 20947 37315
rect 21281 37281 21315 37315
rect 25237 37281 25271 37315
rect 26249 37281 26283 37315
rect 26709 37281 26743 37315
rect 27261 37281 27295 37315
rect 27445 37281 27479 37315
rect 29653 37281 29687 37315
rect 29984 37281 30018 37315
rect 30176 37281 30210 37315
rect 31677 37281 31711 37315
rect 31769 37281 31803 37315
rect 34989 37281 35023 37315
rect 35173 37281 35207 37315
rect 40049 37281 40083 37315
rect 40417 37281 40451 37315
rect 40601 37281 40635 37315
rect 41061 37281 41095 37315
rect 41153 37281 41187 37315
rect 46305 37281 46339 37315
rect 46581 37281 46615 37315
rect 48053 37281 48087 37315
rect 49893 37281 49927 37315
rect 50169 37281 50203 37315
rect 51641 37281 51675 37315
rect 53021 37281 53055 37315
rect 53113 37281 53147 37315
rect 53389 37281 53423 37315
rect 53481 37281 53515 37315
rect 54585 37281 54619 37315
rect 54815 37281 54849 37315
rect 54924 37281 54958 37315
rect 55321 37281 55355 37315
rect 57989 37281 58023 37315
rect 58541 37281 58575 37315
rect 58725 37281 58759 37315
rect 61761 37281 61795 37315
rect 62589 37281 62623 37315
rect 63233 37281 63267 37315
rect 63417 37281 63451 37315
rect 63785 37281 63819 37315
rect 63969 37281 64003 37315
rect 66269 37281 66303 37315
rect 66453 37281 66487 37315
rect 66821 37281 66855 37315
rect 70041 37281 70075 37315
rect 70179 37281 70213 37315
rect 70317 37281 70351 37315
rect 71697 37281 71731 37315
rect 71973 37281 72007 37315
rect 75285 37281 75319 37315
rect 77217 37281 77251 37315
rect 77350 37281 77384 37315
rect 78597 37281 78631 37315
rect 81541 37281 81575 37315
rect 81633 37281 81667 37315
rect 83381 37281 83415 37315
rect 86141 37281 86175 37315
rect 86233 37281 86267 37315
rect 86693 37281 86727 37315
rect 17509 37213 17543 37247
rect 26525 37213 26559 37247
rect 35449 37213 35483 37247
rect 57805 37213 57839 37247
rect 59093 37213 59127 37247
rect 66729 37213 66763 37247
rect 77033 37213 77067 37247
rect 83105 37213 83139 37247
rect 25053 37145 25087 37179
rect 25421 37145 25455 37179
rect 30113 37145 30147 37179
rect 71513 37145 71547 37179
rect 75469 37145 75503 37179
rect 82921 37145 82955 37179
rect 85957 37145 85991 37179
rect 6377 37077 6411 37111
rect 17325 37077 17359 37111
rect 30481 37077 30515 37111
rect 31493 37077 31527 37111
rect 34713 37077 34747 37111
rect 41613 37077 41647 37111
rect 46029 37077 46063 37111
rect 52469 37077 52503 37111
rect 54723 37077 54757 37111
rect 66085 37077 66119 37111
rect 78689 37077 78723 37111
rect 10977 36873 11011 36907
rect 18337 36873 18371 36907
rect 41521 36873 41555 36907
rect 44649 36873 44683 36907
rect 51825 36873 51859 36907
rect 53113 36873 53147 36907
rect 61209 36873 61243 36907
rect 71145 36873 71179 36907
rect 82921 36873 82955 36907
rect 83289 36873 83323 36907
rect 86969 36873 87003 36907
rect 18797 36805 18831 36839
rect 34437 36805 34471 36839
rect 34529 36805 34563 36839
rect 36001 36805 36035 36839
rect 41153 36805 41187 36839
rect 44465 36805 44499 36839
rect 47225 36805 47259 36839
rect 71513 36805 71547 36839
rect 72893 36805 72927 36839
rect 18061 36737 18095 36771
rect 19441 36737 19475 36771
rect 34897 36737 34931 36771
rect 41024 36737 41058 36771
rect 41245 36737 41279 36771
rect 45569 36737 45603 36771
rect 45753 36737 45787 36771
rect 48881 36737 48915 36771
rect 53757 36737 53791 36771
rect 54125 36737 54159 36771
rect 61209 36737 61243 36771
rect 65073 36737 65107 36771
rect 66637 36737 66671 36771
rect 71384 36737 71418 36771
rect 71605 36737 71639 36771
rect 84301 36737 84335 36771
rect 85957 36737 85991 36771
rect 87153 36737 87187 36771
rect 87429 36737 87463 36771
rect 5273 36669 5307 36703
rect 5641 36669 5675 36703
rect 10793 36669 10827 36703
rect 15117 36669 15151 36703
rect 15301 36669 15335 36703
rect 15853 36669 15887 36703
rect 16037 36669 16071 36703
rect 18153 36669 18187 36703
rect 19717 36669 19751 36703
rect 19809 36669 19843 36703
rect 20177 36669 20211 36703
rect 20269 36669 20303 36703
rect 21741 36669 21775 36703
rect 25467 36669 25501 36703
rect 25605 36669 25639 36703
rect 26065 36669 26099 36703
rect 26249 36669 26283 36703
rect 26801 36669 26835 36703
rect 35081 36669 35115 36703
rect 35633 36669 35667 36703
rect 35817 36669 35851 36703
rect 42441 36669 42475 36703
rect 44189 36669 44223 36703
rect 44336 36669 44370 36703
rect 44528 36669 44562 36703
rect 46121 36669 46155 36703
rect 46305 36669 46339 36703
rect 46857 36669 46891 36703
rect 47041 36669 47075 36703
rect 48697 36669 48731 36703
rect 48973 36669 49007 36703
rect 49157 36669 49191 36703
rect 49617 36669 49651 36703
rect 49709 36669 49743 36703
rect 50721 36669 50755 36703
rect 51733 36669 51767 36703
rect 53665 36669 53699 36703
rect 54033 36669 54067 36703
rect 61301 36669 61335 36703
rect 61393 36669 61427 36703
rect 61577 36669 61611 36703
rect 63049 36669 63083 36703
rect 63509 36669 63543 36703
rect 63693 36669 63727 36703
rect 64061 36669 64095 36703
rect 64245 36669 64279 36703
rect 65533 36669 65567 36703
rect 65717 36669 65751 36703
rect 66085 36669 66119 36703
rect 66177 36669 66211 36703
rect 66453 36669 66487 36703
rect 68661 36669 68695 36703
rect 68937 36669 68971 36703
rect 69765 36669 69799 36703
rect 69949 36669 69983 36703
rect 72065 36669 72099 36703
rect 72801 36669 72835 36703
rect 76941 36669 76975 36703
rect 77309 36669 77343 36703
rect 77861 36669 77895 36703
rect 78229 36669 78263 36703
rect 82185 36669 82219 36703
rect 82277 36669 82311 36703
rect 83841 36669 83875 36703
rect 83933 36669 83967 36703
rect 84209 36669 84243 36703
rect 85589 36669 85623 36703
rect 86049 36669 86083 36703
rect 26617 36601 26651 36635
rect 40877 36601 40911 36635
rect 50537 36601 50571 36635
rect 68753 36601 68787 36635
rect 69857 36601 69891 36635
rect 70409 36601 70443 36635
rect 71237 36601 71271 36635
rect 71973 36601 72007 36635
rect 85405 36601 85439 36635
rect 5181 36533 5215 36567
rect 14933 36533 14967 36567
rect 16313 36533 16347 36567
rect 20729 36533 20763 36567
rect 21833 36533 21867 36567
rect 25237 36533 25271 36567
rect 42533 36533 42567 36567
rect 50169 36533 50203 36567
rect 61761 36533 61795 36567
rect 64429 36533 64463 36567
rect 77217 36533 77251 36567
rect 77401 36533 77435 36567
rect 83013 36533 83047 36567
rect 88533 36533 88567 36567
rect 4997 36329 5031 36363
rect 15485 36329 15519 36363
rect 17233 36329 17267 36363
rect 25421 36329 25455 36363
rect 26617 36329 26651 36363
rect 35817 36329 35851 36363
rect 41705 36329 41739 36363
rect 42257 36329 42291 36363
rect 44557 36329 44591 36363
rect 45109 36329 45143 36363
rect 51641 36329 51675 36363
rect 73629 36329 73663 36363
rect 77217 36329 77251 36363
rect 78689 36329 78723 36363
rect 84209 36329 84243 36363
rect 86969 36329 87003 36363
rect 10609 36261 10643 36295
rect 11345 36261 11379 36295
rect 33793 36261 33827 36295
rect 52101 36261 52135 36295
rect 69949 36261 69983 36295
rect 79793 36261 79827 36295
rect 83933 36261 83967 36295
rect 85405 36261 85439 36295
rect 85957 36261 85991 36295
rect 5181 36193 5215 36227
rect 5365 36193 5399 36227
rect 6469 36193 6503 36227
rect 10793 36193 10827 36227
rect 15301 36193 15335 36227
rect 16497 36193 16531 36227
rect 16589 36193 16623 36227
rect 25145 36193 25179 36227
rect 25237 36193 25271 36227
rect 26157 36193 26191 36227
rect 27169 36193 27203 36227
rect 27537 36193 27571 36227
rect 30113 36193 30147 36227
rect 32413 36193 32447 36227
rect 34161 36193 34195 36227
rect 34345 36193 34379 36227
rect 34805 36193 34839 36227
rect 35357 36193 35391 36227
rect 35541 36193 35575 36227
rect 39497 36193 39531 36227
rect 40693 36193 40727 36227
rect 41153 36193 41187 36227
rect 41245 36193 41279 36227
rect 42073 36193 42107 36227
rect 43545 36193 43579 36227
rect 43637 36193 43671 36227
rect 44005 36193 44039 36227
rect 44097 36193 44131 36227
rect 46029 36193 46063 36227
rect 46673 36193 46707 36227
rect 47041 36193 47075 36227
rect 47225 36193 47259 36227
rect 49525 36193 49559 36227
rect 49893 36193 49927 36227
rect 50077 36193 50111 36227
rect 50537 36193 50571 36227
rect 50629 36193 50663 36227
rect 51825 36193 51859 36227
rect 51917 36193 51951 36227
rect 52248 36193 52282 36227
rect 57345 36193 57379 36227
rect 57529 36193 57563 36227
rect 57897 36193 57931 36227
rect 58081 36193 58115 36227
rect 62681 36193 62715 36227
rect 65809 36193 65843 36227
rect 66085 36193 66119 36227
rect 70133 36193 70167 36227
rect 70501 36193 70535 36227
rect 72157 36193 72191 36227
rect 72249 36193 72283 36227
rect 77309 36193 77343 36227
rect 79977 36193 80011 36227
rect 82829 36193 82863 36227
rect 83197 36193 83231 36227
rect 84117 36193 84151 36227
rect 85589 36193 85623 36227
rect 86785 36193 86819 36227
rect 11069 36125 11103 36159
rect 16405 36125 16439 36159
rect 21005 36125 21039 36159
rect 21281 36125 21315 36159
rect 27077 36125 27111 36159
rect 27445 36125 27479 36159
rect 31953 36125 31987 36159
rect 32137 36125 32171 36159
rect 34621 36125 34655 36159
rect 40509 36125 40543 36159
rect 43177 36125 43211 36159
rect 44925 36125 44959 36159
rect 45569 36125 45603 36159
rect 45845 36125 45879 36159
rect 46765 36125 46799 36159
rect 51365 36125 51399 36159
rect 6653 36057 6687 36091
rect 22753 36057 22787 36091
rect 29929 36057 29963 36091
rect 52469 36125 52503 36159
rect 56885 36125 56919 36159
rect 62405 36125 62439 36159
rect 65901 36125 65935 36159
rect 66269 36125 66303 36159
rect 70593 36125 70627 36159
rect 72525 36125 72559 36159
rect 77585 36125 77619 36159
rect 45661 36057 45695 36091
rect 50997 36057 51031 36091
rect 51825 36057 51859 36091
rect 52377 36057 52411 36091
rect 56517 36057 56551 36091
rect 83013 36057 83047 36091
rect 83749 36057 83783 36091
rect 16405 35989 16439 36023
rect 16773 35989 16807 36023
rect 22569 35989 22603 36023
rect 26249 35989 26283 36023
rect 34529 35989 34563 36023
rect 39589 35989 39623 36023
rect 39865 35989 39899 36023
rect 40325 35989 40359 36023
rect 45569 35989 45603 36023
rect 49709 35989 49743 36023
rect 52745 35989 52779 36023
rect 56701 35989 56735 36023
rect 62221 35989 62255 36023
rect 63969 35989 64003 36023
rect 80069 35989 80103 36023
rect 16037 35785 16071 35819
rect 27169 35785 27203 35819
rect 31033 35785 31067 35819
rect 34437 35785 34471 35819
rect 39681 35785 39715 35819
rect 51089 35785 51123 35819
rect 52377 35785 52411 35819
rect 54861 35785 54895 35819
rect 55045 35785 55079 35819
rect 63693 35785 63727 35819
rect 79425 35785 79459 35819
rect 79609 35785 79643 35819
rect 80069 35785 80103 35819
rect 80437 35785 80471 35819
rect 86049 35785 86083 35819
rect 86969 35785 87003 35819
rect 21741 35717 21775 35751
rect 32689 35717 32723 35751
rect 33057 35717 33091 35751
rect 33241 35717 33275 35751
rect 42993 35717 43027 35751
rect 52009 35717 52043 35751
rect 56793 35717 56827 35751
rect 56977 35717 57011 35751
rect 3893 35649 3927 35683
rect 20637 35649 20671 35683
rect 30573 35649 30607 35683
rect 30849 35649 30883 35683
rect 35633 35649 35667 35683
rect 35817 35649 35851 35683
rect 39497 35649 39531 35683
rect 40325 35649 40359 35683
rect 41797 35649 41831 35683
rect 42864 35649 42898 35683
rect 43085 35649 43119 35683
rect 50721 35649 50755 35683
rect 51880 35649 51914 35683
rect 52101 35649 52135 35683
rect 57161 35649 57195 35683
rect 3617 35581 3651 35615
rect 6837 35581 6871 35615
rect 7389 35581 7423 35615
rect 10885 35581 10919 35615
rect 11161 35581 11195 35615
rect 11345 35581 11379 35615
rect 13369 35581 13403 35615
rect 13645 35581 13679 35615
rect 15761 35581 15795 35615
rect 15853 35581 15887 35615
rect 20361 35581 20395 35615
rect 25421 35581 25455 35615
rect 25605 35581 25639 35615
rect 25789 35581 25823 35615
rect 26249 35581 26283 35615
rect 26341 35581 26375 35615
rect 29285 35581 29319 35615
rect 29469 35581 29503 35615
rect 29929 35581 29963 35615
rect 30021 35581 30055 35615
rect 31493 35581 31527 35615
rect 31631 35581 31665 35615
rect 32137 35581 32171 35615
rect 32229 35581 32263 35615
rect 35541 35581 35575 35615
rect 35909 35581 35943 35615
rect 38209 35581 38243 35615
rect 38393 35581 38427 35615
rect 38853 35581 38887 35615
rect 38945 35581 38979 35615
rect 39865 35581 39899 35615
rect 5365 35513 5399 35547
rect 10333 35513 10367 35547
rect 15025 35513 15059 35547
rect 26893 35513 26927 35547
rect 34897 35513 34931 35547
rect 40647 35581 40681 35615
rect 40785 35581 40819 35615
rect 41153 35581 41187 35615
rect 41245 35581 41279 35615
rect 42073 35581 42107 35615
rect 49433 35581 49467 35615
rect 49617 35581 49651 35615
rect 50077 35581 50111 35615
rect 50169 35581 50203 35615
rect 53297 35581 53331 35615
rect 55689 35581 55723 35615
rect 55873 35581 55907 35615
rect 56241 35581 56275 35615
rect 56425 35581 56459 35615
rect 56609 35581 56643 35615
rect 42717 35513 42751 35547
rect 50905 35513 50939 35547
rect 51733 35513 51767 35547
rect 55229 35513 55263 35547
rect 57345 35581 57379 35615
rect 57529 35581 57563 35615
rect 58081 35581 58115 35615
rect 58265 35581 58299 35615
rect 58633 35513 58667 35547
rect 4997 35445 5031 35479
rect 6929 35445 6963 35479
rect 10241 35445 10275 35479
rect 11529 35445 11563 35479
rect 13277 35445 13311 35479
rect 22109 35445 22143 35479
rect 28825 35445 28859 35479
rect 29009 35445 29043 35479
rect 31125 35445 31159 35479
rect 31309 35445 31343 35479
rect 34621 35445 34655 35479
rect 37841 35445 37875 35479
rect 38025 35445 38059 35479
rect 40141 35445 40175 35479
rect 40325 35445 40359 35479
rect 42257 35445 42291 35479
rect 43361 35445 43395 35479
rect 49065 35445 49099 35479
rect 49249 35445 49283 35479
rect 53389 35445 53423 35479
rect 57161 35445 57195 35479
rect 69765 35717 69799 35751
rect 70133 35717 70167 35751
rect 71697 35717 71731 35751
rect 77125 35717 77159 35751
rect 79149 35717 79183 35751
rect 77309 35649 77343 35683
rect 77861 35649 77895 35683
rect 78321 35649 78355 35683
rect 63785 35581 63819 35615
rect 64061 35581 64095 35615
rect 65441 35581 65475 35615
rect 66269 35581 66303 35615
rect 68937 35581 68971 35615
rect 69029 35581 69063 35615
rect 69489 35581 69523 35615
rect 70317 35581 70351 35615
rect 70593 35581 70627 35615
rect 72801 35581 72835 35615
rect 78137 35581 78171 35615
rect 69581 35513 69615 35547
rect 82369 35717 82403 35751
rect 83105 35717 83139 35751
rect 79940 35649 79974 35683
rect 80161 35649 80195 35683
rect 82829 35649 82863 35683
rect 83289 35649 83323 35683
rect 79609 35581 79643 35615
rect 79793 35581 79827 35615
rect 82185 35581 82219 35615
rect 83933 35581 83967 35615
rect 84025 35581 84059 35615
rect 84301 35581 84335 35615
rect 84393 35581 84427 35615
rect 85589 35581 85623 35615
rect 87153 35581 87187 35615
rect 87429 35581 87463 35615
rect 82921 35513 82955 35547
rect 85405 35513 85439 35547
rect 63693 35445 63727 35479
rect 66361 35445 66395 35479
rect 72985 35445 73019 35479
rect 79149 35445 79183 35479
rect 79241 35445 79275 35479
rect 80713 35445 80747 35479
rect 82645 35445 82679 35479
rect 85681 35445 85715 35479
rect 88533 35445 88567 35479
rect 4721 35241 4755 35275
rect 11529 35241 11563 35275
rect 15669 35241 15703 35275
rect 21097 35241 21131 35275
rect 22753 35241 22787 35275
rect 70685 35241 70719 35275
rect 83013 35241 83047 35275
rect 83197 35241 83231 35275
rect 86509 35241 86543 35275
rect 26249 35173 26283 35207
rect 32873 35173 32907 35207
rect 34805 35173 34839 35207
rect 39957 35173 39991 35207
rect 41981 35173 42015 35207
rect 49617 35173 49651 35207
rect 50997 35173 51031 35207
rect 53205 35173 53239 35207
rect 58449 35173 58483 35207
rect 72433 35173 72467 35207
rect 80253 35173 80287 35207
rect 83381 35173 83415 35207
rect 84945 35173 84979 35207
rect 88349 35173 88383 35207
rect 4721 35105 4755 35139
rect 4997 35105 5031 35139
rect 6285 35105 6319 35139
rect 6561 35105 6595 35139
rect 9689 35105 9723 35139
rect 10241 35105 10275 35139
rect 10517 35105 10551 35139
rect 11621 35105 11655 35139
rect 13829 35105 13863 35139
rect 14197 35105 14231 35139
rect 15301 35105 15335 35139
rect 16405 35105 16439 35139
rect 16773 35105 16807 35139
rect 20913 35105 20947 35139
rect 22385 35105 22419 35139
rect 22569 35105 22603 35139
rect 23673 35105 23707 35139
rect 26709 35105 26743 35139
rect 27169 35105 27203 35139
rect 27261 35105 27295 35139
rect 28817 35105 28851 35139
rect 28917 35105 28951 35139
rect 30389 35105 30423 35139
rect 30481 35105 30515 35139
rect 6745 35037 6779 35071
rect 23765 35037 23799 35071
rect 26525 35037 26559 35071
rect 27813 35037 27847 35071
rect 9781 34969 9815 35003
rect 11805 34969 11839 35003
rect 15485 34969 15519 35003
rect 33057 35105 33091 35139
rect 33149 35105 33183 35139
rect 33425 35105 33459 35139
rect 38669 35105 38703 35139
rect 39221 35105 39255 35139
rect 39405 35105 39439 35139
rect 40693 35105 40727 35139
rect 40877 35105 40911 35139
rect 41337 35105 41371 35139
rect 41429 35105 41463 35139
rect 42257 35105 42291 35139
rect 42441 35105 42475 35139
rect 49893 35105 49927 35139
rect 50353 35105 50387 35139
rect 50445 35105 50479 35139
rect 51457 35105 51491 35139
rect 52101 35105 52135 35139
rect 52561 35105 52595 35139
rect 52653 35105 52687 35139
rect 53573 35105 53607 35139
rect 55781 35105 55815 35139
rect 58725 35105 58759 35139
rect 62037 35105 62071 35139
rect 64521 35105 64555 35139
rect 65533 35105 65567 35139
rect 65809 35105 65843 35139
rect 68937 35105 68971 35139
rect 69305 35105 69339 35139
rect 69949 35105 69983 35139
rect 70133 35105 70167 35139
rect 70777 35105 70811 35139
rect 71881 35105 71915 35139
rect 71973 35105 72007 35139
rect 75929 35105 75963 35139
rect 77033 35105 77067 35139
rect 77401 35105 77435 35139
rect 78597 35105 78631 35139
rect 79057 35105 79091 35139
rect 80161 35105 80195 35139
rect 80345 35105 80379 35139
rect 83565 35105 83599 35139
rect 84761 35105 84795 35139
rect 85037 35105 85071 35139
rect 86325 35105 86359 35139
rect 86969 35105 87003 35139
rect 88257 35105 88291 35139
rect 38485 35037 38519 35071
rect 39773 35037 39807 35071
rect 40509 35037 40543 35071
rect 49709 35037 49743 35071
rect 51917 35037 51951 35071
rect 56057 35037 56091 35071
rect 56333 35037 56367 35071
rect 62313 35037 62347 35071
rect 70501 35037 70535 35071
rect 76205 35037 76239 35071
rect 78873 35037 78907 35071
rect 85497 35037 85531 35071
rect 87153 35037 87187 35071
rect 40141 34969 40175 35003
rect 53481 34969 53515 35003
rect 58541 34969 58575 35003
rect 63601 34969 63635 35003
rect 65533 34969 65567 35003
rect 69029 34969 69063 35003
rect 78321 34969 78355 35003
rect 13921 34901 13955 34935
rect 16589 34901 16623 34935
rect 25973 34901 26007 34935
rect 28089 34901 28123 34935
rect 32873 34901 32907 34935
rect 38117 34901 38151 34935
rect 38301 34901 38335 34935
rect 40325 34901 40359 34935
rect 49341 34901 49375 34935
rect 51273 34901 51307 34935
rect 51549 34901 51583 34935
rect 51733 34901 51767 34935
rect 55597 34901 55631 34935
rect 57437 34901 57471 34935
rect 58817 34901 58851 34935
rect 59001 34901 59035 34935
rect 59185 34901 59219 34935
rect 59461 34901 59495 34935
rect 64613 34901 64647 34935
rect 65901 34901 65935 34935
rect 71697 34901 71731 34935
rect 76021 34901 76055 34935
rect 77217 34901 77251 34935
rect 80529 34901 80563 34935
rect 83657 34901 83691 34935
rect 85957 34901 85991 34935
rect 86141 34901 86175 34935
rect 86693 34901 86727 34935
rect 87337 34901 87371 34935
rect 9413 34697 9447 34731
rect 11897 34697 11931 34731
rect 25513 34697 25547 34731
rect 30665 34697 30699 34731
rect 37841 34697 37875 34731
rect 39405 34697 39439 34731
rect 43637 34697 43671 34731
rect 46857 34697 46891 34731
rect 48421 34697 48455 34731
rect 50261 34697 50295 34731
rect 56149 34697 56183 34731
rect 58817 34697 58851 34731
rect 71421 34697 71455 34731
rect 72341 34697 72375 34731
rect 72617 34697 72651 34731
rect 76297 34697 76331 34731
rect 77769 34697 77803 34731
rect 80069 34697 80103 34731
rect 81265 34697 81299 34731
rect 85681 34697 85715 34731
rect 87153 34697 87187 34731
rect 88349 34697 88383 34731
rect 15577 34629 15611 34663
rect 22385 34629 22419 34663
rect 25237 34629 25271 34663
rect 38025 34629 38059 34663
rect 39957 34629 39991 34663
rect 50445 34629 50479 34663
rect 61945 34629 61979 34663
rect 64337 34629 64371 34663
rect 69949 34629 69983 34663
rect 79609 34629 79643 34663
rect 80437 34629 80471 34663
rect 87705 34629 87739 34663
rect 2881 34561 2915 34595
rect 5641 34561 5675 34595
rect 9689 34561 9723 34595
rect 11069 34561 11103 34595
rect 11713 34561 11747 34595
rect 38209 34561 38243 34595
rect 46673 34561 46707 34595
rect 53849 34561 53883 34595
rect 56793 34561 56827 34595
rect 56977 34561 57011 34595
rect 58633 34561 58667 34595
rect 60013 34561 60047 34595
rect 76389 34561 76423 34595
rect 76665 34561 76699 34595
rect 82277 34561 82311 34595
rect 86049 34561 86083 34595
rect 88073 34561 88107 34595
rect 2605 34493 2639 34527
rect 4445 34493 4479 34527
rect 5365 34493 5399 34527
rect 5549 34493 5583 34527
rect 9229 34493 9263 34527
rect 10333 34493 10367 34527
rect 10977 34493 11011 34527
rect 11345 34493 11379 34527
rect 11529 34493 11563 34527
rect 13829 34493 13863 34527
rect 14013 34493 14047 34527
rect 14289 34493 14323 34527
rect 19901 34493 19935 34527
rect 19993 34493 20027 34527
rect 20177 34493 20211 34527
rect 20637 34493 20671 34527
rect 20729 34493 20763 34527
rect 22201 34493 22235 34527
rect 25743 34493 25777 34527
rect 25881 34493 25915 34527
rect 26249 34493 26283 34527
rect 26341 34493 26375 34527
rect 29292 34493 29326 34527
rect 29561 34493 29595 34527
rect 38393 34493 38427 34527
rect 38853 34493 38887 34527
rect 38945 34493 38979 34527
rect 39773 34493 39807 34527
rect 42073 34493 42107 34527
rect 42257 34493 42291 34527
rect 42441 34493 42475 34527
rect 42625 34493 42659 34527
rect 43085 34493 43119 34527
rect 43177 34493 43211 34527
rect 44005 34493 44039 34527
rect 44189 34493 44223 34527
rect 47041 34493 47075 34527
rect 48697 34493 48731 34527
rect 48881 34493 48915 34527
rect 49433 34493 49467 34527
rect 49617 34493 49651 34527
rect 53573 34493 53607 34527
rect 56057 34493 56091 34527
rect 56609 34493 56643 34527
rect 57345 34493 57379 34527
rect 57529 34493 57563 34527
rect 58081 34493 58115 34527
rect 58265 34493 58299 34527
rect 59001 34493 59035 34527
rect 59185 34493 59219 34527
rect 59369 34493 59403 34527
rect 59737 34493 59771 34527
rect 61853 34493 61887 34527
rect 62957 34493 62991 34527
rect 63233 34493 63267 34527
rect 70041 34493 70075 34527
rect 70317 34493 70351 34527
rect 72525 34493 72559 34527
rect 79609 34493 79643 34527
rect 79793 34493 79827 34527
rect 79977 34493 80011 34527
rect 81173 34493 81207 34527
rect 82185 34493 82219 34527
rect 83197 34493 83231 34527
rect 83381 34493 83415 34527
rect 85773 34493 85807 34527
rect 87521 34493 87555 34527
rect 87889 34493 87923 34527
rect 88257 34493 88291 34527
rect 21281 34425 21315 34459
rect 27077 34425 27111 34459
rect 49985 34425 50019 34459
rect 55413 34425 55447 34459
rect 62681 34425 62715 34459
rect 3985 34357 4019 34391
rect 25053 34357 25087 34391
rect 26801 34357 26835 34391
rect 31033 34357 31067 34391
rect 48513 34357 48547 34391
rect 55137 34357 55171 34391
rect 59553 34357 59587 34391
rect 59829 34357 59863 34391
rect 83473 34357 83507 34391
rect 15393 34153 15427 34187
rect 15669 34153 15703 34187
rect 56609 34153 56643 34187
rect 14289 34085 14323 34119
rect 28181 34085 28215 34119
rect 5089 34017 5123 34051
rect 5273 34017 5307 34051
rect 10517 34017 10551 34051
rect 10701 34017 10735 34051
rect 13185 34017 13219 34051
rect 13645 34017 13679 34051
rect 13737 34017 13771 34051
rect 15301 34017 15335 34051
rect 19441 34017 19475 34051
rect 19809 34017 19843 34051
rect 19993 34017 20027 34051
rect 21097 34017 21131 34051
rect 21649 34017 21683 34051
rect 21833 34017 21867 34051
rect 22477 34017 22511 34051
rect 26801 34017 26835 34051
rect 30573 34017 30607 34051
rect 5365 33949 5399 33983
rect 9689 33949 9723 33983
rect 10241 33949 10275 33983
rect 13001 33949 13035 33983
rect 18797 33949 18831 33983
rect 19533 33949 19567 33983
rect 20913 33949 20947 33983
rect 26525 33949 26559 33983
rect 29377 33949 29411 33983
rect 20269 33881 20303 33915
rect 9505 33813 9539 33847
rect 12817 33813 12851 33847
rect 20177 33813 20211 33847
rect 20637 33813 20671 33847
rect 22109 33813 22143 33847
rect 28273 33813 28307 33847
rect 5273 33609 5307 33643
rect 13645 33609 13679 33643
rect 14565 33609 14599 33643
rect 19073 33609 19107 33643
rect 19349 33609 19383 33643
rect 21557 33609 21591 33643
rect 29377 33609 29411 33643
rect 21189 33541 21223 33575
rect 2881 33473 2915 33507
rect 9045 33473 9079 33507
rect 10885 33473 10919 33507
rect 25973 33473 26007 33507
rect 56609 33881 56643 33915
rect 2605 33405 2639 33439
rect 5089 33405 5123 33439
rect 8217 33405 8251 33439
rect 8769 33405 8803 33439
rect 10609 33405 10643 33439
rect 12587 33405 12621 33439
rect 12725 33405 12759 33439
rect 13185 33405 13219 33439
rect 13369 33405 13403 33439
rect 14657 33405 14691 33439
rect 18889 33405 18923 33439
rect 19993 33405 20027 33439
rect 20177 33405 20211 33439
rect 20729 33405 20763 33439
rect 20913 33405 20947 33439
rect 24869 33405 24903 33439
rect 24961 33405 24995 33439
rect 25329 33405 25363 33439
rect 25421 33405 25455 33439
rect 30573 33405 30607 33439
rect 10425 33337 10459 33371
rect 26433 33337 26467 33371
rect 4169 33269 4203 33303
rect 4445 33269 4479 33303
rect 8125 33269 8159 33303
rect 12173 33269 12207 33303
rect 14841 33269 14875 33303
rect 19809 33269 19843 33303
rect 24501 33269 24535 33303
rect 26249 33269 26283 33303
rect 21005 33065 21039 33099
rect 25789 33065 25823 33099
rect 13001 32997 13035 33031
rect 4353 32929 4387 32963
rect 4629 32929 4663 32963
rect 8217 32929 8251 32963
rect 12541 32929 12575 32963
rect 13461 32929 13495 32963
rect 13737 32929 13771 32963
rect 18521 32929 18555 32963
rect 19073 32929 19107 32963
rect 19257 32929 19291 32963
rect 21373 32929 21407 32963
rect 21557 32929 21591 32963
rect 21879 32929 21913 32963
rect 22017 32929 22051 32963
rect 24409 32929 24443 32963
rect 24869 32929 24903 32963
rect 24961 32929 24995 32963
rect 26065 32929 26099 32963
rect 4813 32861 4847 32895
rect 5733 32861 5767 32895
rect 6009 32861 6043 32895
rect 18337 32861 18371 32895
rect 19625 32861 19659 32895
rect 24225 32861 24259 32895
rect 25513 32861 25547 32895
rect 13461 32793 13495 32827
rect 13553 32793 13587 32827
rect 7297 32725 7331 32759
rect 7573 32725 7607 32759
rect 8309 32725 8343 32759
rect 12725 32725 12759 32759
rect 13921 32725 13955 32759
rect 18153 32725 18187 32759
rect 19901 32725 19935 32759
rect 25881 32725 25915 32759
rect 57989 32589 58023 32623
rect 4445 32521 4479 32555
rect 8217 32521 8251 32555
rect 26157 32521 26191 32555
rect 14841 32453 14875 32487
rect 57943 32453 57977 32487
rect 72433 32453 72467 32487
rect 2605 32385 2639 32419
rect 2881 32385 2915 32419
rect 6837 32385 6871 32419
rect 12265 32385 12299 32419
rect 7113 32317 7147 32351
rect 12909 32317 12943 32351
rect 13093 32317 13127 32351
rect 13461 32317 13495 32351
rect 13645 32317 13679 32351
rect 14657 32317 14691 32351
rect 19349 32317 19383 32351
rect 19441 32317 19475 32351
rect 19717 32317 19751 32351
rect 24777 32317 24811 32351
rect 24961 32317 24995 32351
rect 26065 32317 26099 32351
rect 8585 32249 8619 32283
rect 11989 32249 12023 32283
rect 3985 32181 4019 32215
rect 12541 32181 12575 32215
rect 21005 32181 21039 32215
rect 25145 32181 25179 32215
rect 72433 32113 72467 32147
rect 4261 31977 4295 32011
rect 7021 31977 7055 32011
rect 7389 31977 7423 32011
rect 8125 31977 8159 32011
rect 18061 31977 18095 32011
rect 19809 31977 19843 32011
rect 21097 31977 21131 32011
rect 24961 31977 24995 32011
rect 27629 31977 27663 32011
rect 22109 31909 22143 31943
rect 27813 31909 27847 31943
rect 4077 31841 4111 31875
rect 5825 31841 5859 31875
rect 6009 31841 6043 31875
rect 6561 31841 6595 31875
rect 6745 31841 6779 31875
rect 8033 31841 8067 31875
rect 12817 31841 12851 31875
rect 13185 31841 13219 31875
rect 18429 31841 18463 31875
rect 18981 31841 19015 31875
rect 19165 31841 19199 31875
rect 21005 31841 21039 31875
rect 22017 31841 22051 31875
rect 25053 31841 25087 31875
rect 27537 31841 27571 31875
rect 12173 31773 12207 31807
rect 12725 31773 12759 31807
rect 13093 31773 13127 31807
rect 13737 31773 13771 31807
rect 18245 31773 18279 31807
rect 86877 31773 86911 31807
rect 19441 31705 19475 31739
rect 13553 31637 13587 31671
rect 25237 31637 25271 31671
rect 59277 31569 59311 31603
rect 86877 31569 86911 31603
rect 4445 31433 4479 31467
rect 8033 31433 8067 31467
rect 8401 31433 8435 31467
rect 9597 31433 9631 31467
rect 2881 31297 2915 31331
rect 6929 31297 6963 31331
rect 2605 31229 2639 31263
rect 7021 31229 7055 31263
rect 7573 31229 7607 31263
rect 7757 31229 7791 31263
rect 37289 31433 37323 31467
rect 13093 31365 13127 31399
rect 14197 31365 14231 31399
rect 23765 31365 23799 31399
rect 27537 31365 27571 31399
rect 20177 31297 20211 31331
rect 21557 31297 21591 31331
rect 25881 31297 25915 31331
rect 25973 31297 26007 31331
rect 9873 31229 9907 31263
rect 10057 31229 10091 31263
rect 10609 31229 10643 31263
rect 10793 31229 10827 31263
rect 12909 31229 12943 31263
rect 14013 31229 14047 31263
rect 18337 31229 18371 31263
rect 19809 31229 19843 31263
rect 19901 31229 19935 31263
rect 23857 31229 23891 31263
rect 26157 31229 26191 31263
rect 26709 31229 26743 31263
rect 26893 31229 26927 31263
rect 9597 31161 9631 31195
rect 11161 31161 11195 31195
rect 11437 31161 11471 31195
rect 14473 31161 14507 31195
rect 46857 31433 46891 31467
rect 4169 31093 4203 31127
rect 9689 31093 9723 31127
rect 18521 31093 18555 31127
rect 23949 31093 23983 31127
rect 27169 31093 27203 31127
rect 37289 31093 37323 31127
rect 46855 31093 46889 31127
rect 48329 31229 48363 31263
rect 48421 31161 48455 31195
rect 48145 31093 48179 31127
rect 48237 31093 48271 31127
rect 2881 30889 2915 30923
rect 4997 30889 5031 30923
rect 27905 30889 27939 30923
rect 6561 30821 6595 30855
rect 16129 30821 16163 30855
rect 17233 30821 17267 30855
rect 18061 30821 18095 30855
rect 25605 30821 25639 30855
rect 2973 30753 3007 30787
rect 4169 30753 4203 30787
rect 4629 30753 4663 30787
rect 5641 30753 5675 30787
rect 6193 30753 6227 30787
rect 10517 30753 10551 30787
rect 10793 30753 10827 30787
rect 12265 30753 12299 30787
rect 13461 30753 13495 30787
rect 13737 30753 13771 30787
rect 16497 30753 16531 30787
rect 16644 30753 16678 30787
rect 18705 30753 18739 30787
rect 19073 30753 19107 30787
rect 19257 30753 19291 30787
rect 19349 30753 19383 30787
rect 23949 30753 23983 30787
rect 25697 30753 25731 30787
rect 26801 30753 26835 30787
rect 4721 30685 4755 30719
rect 6101 30685 6135 30719
rect 12173 30685 12207 30719
rect 16865 30685 16899 30719
rect 18797 30685 18831 30719
rect 19533 30685 19567 30719
rect 24225 30685 24259 30719
rect 26525 30685 26559 30719
rect 3065 30549 3099 30583
rect 13277 30549 13311 30583
rect 13921 30549 13955 30583
rect 16405 30549 16439 30583
rect 16773 30549 16807 30583
rect 28273 30549 28307 30583
rect 5733 30345 5767 30379
rect 13553 30345 13587 30379
rect 16221 30345 16255 30379
rect 11069 30277 11103 30311
rect 11437 30277 11471 30311
rect 17693 30277 17727 30311
rect 18337 30277 18371 30311
rect 19809 30277 19843 30311
rect 23673 30277 23707 30311
rect 25421 30277 25455 30311
rect 4445 30209 4479 30243
rect 16865 30209 16899 30243
rect 2697 30141 2731 30175
rect 2973 30141 3007 30175
rect 4169 30141 4203 30175
rect 4537 30141 4571 30175
rect 5549 30141 5583 30175
rect 9873 30141 9907 30175
rect 10057 30141 10091 30175
rect 10609 30141 10643 30175
rect 10793 30141 10827 30175
rect 12449 30141 12483 30175
rect 13461 30141 13495 30175
rect 15209 30141 15243 30175
rect 16405 30141 16439 30175
rect 16589 30141 16623 30175
rect 16957 30141 16991 30175
rect 18208 30209 18242 30243
rect 18429 30209 18463 30243
rect 21281 30209 21315 30243
rect 21465 30209 21499 30243
rect 22661 30209 22695 30243
rect 23857 30209 23891 30243
rect 19625 30141 19659 30175
rect 21557 30141 21591 30175
rect 22109 30141 22143 30175
rect 22293 30141 22327 30175
rect 24041 30141 24075 30175
rect 24501 30141 24535 30175
rect 24593 30141 24627 30175
rect 3157 30073 3191 30107
rect 17233 30073 17267 30107
rect 17693 30073 17727 30107
rect 17785 30073 17819 30107
rect 18061 30073 18095 30107
rect 3341 30005 3375 30039
rect 4905 30005 4939 30039
rect 9781 30005 9815 30039
rect 12541 30005 12575 30039
rect 15025 30005 15059 30039
rect 15393 30005 15427 30039
rect 17509 30005 17543 30039
rect 18705 30005 18739 30039
rect 22845 30005 22879 30039
rect 25053 30005 25087 30039
rect 3341 29801 3375 29835
rect 4997 29801 5031 29835
rect 12081 29801 12115 29835
rect 14105 29801 14139 29835
rect 20177 29801 20211 29835
rect 18797 29733 18831 29767
rect 2697 29665 2731 29699
rect 2881 29665 2915 29699
rect 4169 29665 4203 29699
rect 4629 29665 4663 29699
rect 6101 29665 6135 29699
rect 10793 29665 10827 29699
rect 13921 29665 13955 29699
rect 16773 29665 16807 29699
rect 17325 29665 17359 29699
rect 17509 29665 17543 29699
rect 19257 29665 19291 29699
rect 19441 29665 19475 29699
rect 19809 29665 19843 29699
rect 20361 29665 20395 29699
rect 23581 29665 23615 29699
rect 2973 29597 3007 29631
rect 4537 29597 4571 29631
rect 5825 29597 5859 29631
rect 7573 29597 7607 29631
rect 10333 29597 10367 29631
rect 10517 29597 10551 29631
rect 16589 29597 16623 29631
rect 19717 29597 19751 29631
rect 23305 29597 23339 29631
rect 17693 29529 17727 29563
rect 7205 29461 7239 29495
rect 16497 29461 16531 29495
rect 18061 29461 18095 29495
rect 18245 29461 18279 29495
rect 18613 29461 18647 29495
rect 23121 29461 23155 29495
rect 24685 29461 24719 29495
rect 18153 29257 18187 29291
rect 19625 29257 19659 29291
rect 24225 29257 24259 29291
rect 26709 29257 26743 29291
rect 5549 29189 5583 29223
rect 12449 29121 12483 29155
rect 14105 29121 14139 29155
rect 25145 29121 25179 29155
rect 4077 29053 4111 29087
rect 4353 29053 4387 29087
rect 5365 29053 5399 29087
rect 12725 29053 12759 29087
rect 14933 29053 14967 29087
rect 16865 29053 16899 29087
rect 18061 29053 18095 29087
rect 19441 29053 19475 29087
rect 24133 29053 24167 29087
rect 25421 29053 25455 29087
rect 14197 28985 14231 29019
rect 24501 28985 24535 29019
rect 3893 28917 3927 28951
rect 15025 28917 15059 28951
rect 16681 28917 16715 28951
rect 18429 28917 18463 28951
rect 26985 28917 27019 28951
rect 19625 28713 19659 28747
rect 13093 28645 13127 28679
rect 4353 28577 4387 28611
rect 4537 28577 4571 28611
rect 4997 28577 5031 28611
rect 8401 28577 8435 28611
rect 11713 28577 11747 28611
rect 12265 28577 12299 28611
rect 12449 28577 12483 28611
rect 13737 28577 13771 28611
rect 17509 28577 17543 28611
rect 19717 28577 19751 28611
rect 25421 28577 25455 28611
rect 27353 28577 27387 28611
rect 4629 28509 4663 28543
rect 11437 28509 11471 28543
rect 11621 28509 11655 28543
rect 17233 28509 17267 28543
rect 12633 28441 12667 28475
rect 13921 28441 13955 28475
rect 8309 28373 8343 28407
rect 8493 28373 8527 28407
rect 17141 28373 17175 28407
rect 18613 28373 18647 28407
rect 19901 28373 19935 28407
rect 25513 28373 25547 28407
rect 27445 28373 27479 28407
rect 28089 28169 28123 28203
rect 9873 28101 9907 28135
rect 11345 28101 11379 28135
rect 25421 28101 25455 28135
rect 2881 28033 2915 28067
rect 9321 28033 9355 28067
rect 13645 28033 13679 28067
rect 19717 28033 19751 28067
rect 26525 28033 26559 28067
rect 28273 28033 28307 28067
rect 2605 27965 2639 27999
rect 5273 27965 5307 27999
rect 5641 27965 5675 27999
rect 7573 27965 7607 27999
rect 9459 27965 9493 27999
rect 9597 27965 9631 27999
rect 10977 27965 11011 27999
rect 12265 27965 12299 27999
rect 12449 27965 12483 27999
rect 12633 27965 12667 27999
rect 13093 27965 13127 27999
rect 13185 27965 13219 27999
rect 19901 27965 19935 27999
rect 20453 27965 20487 27999
rect 20637 27965 20671 27999
rect 24317 27965 24351 27999
rect 24501 27965 24535 27999
rect 25053 27965 25087 27999
rect 25237 27965 25271 27999
rect 26801 27965 26835 27999
rect 8769 27897 8803 27931
rect 21005 27897 21039 27931
rect 4169 27829 4203 27863
rect 4445 27829 4479 27863
rect 5181 27829 5215 27863
rect 7665 27829 7699 27863
rect 11161 27829 11195 27863
rect 19533 27829 19567 27863
rect 24133 27829 24167 27863
rect 59553 31297 59587 31331
rect 87337 31161 87371 31195
rect 96537 31161 96571 31195
rect 96537 30957 96571 30991
rect 99297 30957 99331 30991
rect 99389 30957 99423 30991
rect 87337 30821 87371 30855
rect 59553 27897 59587 27931
rect 8493 27625 8527 27659
rect 59277 27625 59311 27659
rect 8953 27557 8987 27591
rect 17325 27557 17359 27591
rect 27813 27557 27847 27591
rect 4353 27489 4387 27523
rect 4537 27489 4571 27523
rect 4997 27489 5031 27523
rect 8033 27489 8067 27523
rect 8309 27489 8343 27523
rect 9137 27489 9171 27523
rect 10609 27489 10643 27523
rect 11805 27489 11839 27523
rect 15853 27489 15887 27523
rect 15945 27489 15979 27523
rect 16405 27489 16439 27523
rect 16589 27489 16623 27523
rect 21189 27489 21223 27523
rect 23213 27489 23247 27523
rect 23513 27489 23547 27523
rect 26709 27489 26743 27523
rect 27261 27489 27295 27523
rect 27445 27489 27479 27523
rect 4629 27421 4663 27455
rect 8125 27421 8159 27455
rect 11529 27421 11563 27455
rect 15577 27421 15611 27455
rect 20729 27421 20763 27455
rect 20913 27421 20947 27455
rect 22569 27421 22603 27455
rect 26525 27421 26559 27455
rect 10425 27285 10459 27319
rect 11345 27285 11379 27319
rect 13093 27285 13127 27319
rect 16865 27285 16899 27319
rect 17141 27285 17175 27319
rect 23213 27285 23247 27319
rect 23305 27285 23339 27319
rect 23581 27285 23615 27319
rect 26249 27285 26283 27319
rect 11253 27081 11287 27115
rect 13185 27081 13219 27115
rect 26617 27081 26651 27115
rect 2605 26945 2639 26979
rect 2881 26945 2915 26979
rect 7757 26945 7791 26979
rect 9689 26945 9723 26979
rect 14197 26945 14231 26979
rect 14289 26945 14323 26979
rect 14565 26945 14599 26979
rect 20637 26945 20671 26979
rect 4353 26877 4387 26911
rect 7665 26877 7699 26911
rect 8585 26877 8619 26911
rect 9229 26877 9263 26911
rect 9505 26877 9539 26911
rect 10517 26877 10551 26911
rect 10701 26877 10735 26911
rect 13093 26877 13127 26911
rect 16773 26877 16807 26911
rect 20913 26877 20947 26911
rect 21005 26877 21039 26911
rect 21465 26877 21499 26911
rect 21649 26877 21683 26911
rect 25053 26877 25087 26911
rect 25329 26877 25363 26911
rect 8677 26809 8711 26843
rect 9873 26809 9907 26843
rect 4169 26741 4203 26775
rect 7573 26741 7607 26775
rect 10793 26741 10827 26775
rect 15669 26741 15703 26775
rect 16865 26741 16899 26775
rect 21925 26741 21959 26775
rect 22293 26741 22327 26775
rect 24961 26741 24995 26775
rect 7941 26537 7975 26571
rect 23857 26537 23891 26571
rect 17877 26469 17911 26503
rect 4353 26401 4387 26435
rect 6837 26401 6871 26435
rect 16221 26401 16255 26435
rect 21557 26401 21591 26435
rect 22937 26401 22971 26435
rect 23765 26401 23799 26435
rect 25421 26401 25455 26435
rect 26709 26401 26743 26435
rect 4077 26333 4111 26367
rect 5825 26333 5859 26367
rect 6561 26333 6595 26367
rect 8309 26333 8343 26367
rect 16497 26333 16531 26367
rect 21281 26333 21315 26367
rect 17969 26265 18003 26299
rect 21097 26265 21131 26299
rect 5457 26197 5491 26231
rect 25513 26197 25547 26231
rect 26801 26197 26835 26231
rect 7481 25993 7515 26027
rect 9321 25993 9355 26027
rect 17141 25993 17175 26027
rect 25145 25993 25179 26027
rect 27813 25993 27847 26027
rect 8493 25925 8527 25959
rect 9413 25925 9447 25959
rect 16681 25925 16715 25959
rect 2881 25857 2915 25891
rect 15393 25857 15427 25891
rect 15577 25857 15611 25891
rect 2605 25789 2639 25823
rect 7389 25789 7423 25823
rect 8401 25789 8435 25823
rect 8677 25789 8711 25823
rect 10977 25789 11011 25823
rect 15761 25789 15795 25823
rect 16313 25789 16347 25823
rect 16497 25789 16531 25823
rect 18061 25789 18095 25823
rect 23949 25789 23983 25823
rect 24133 25789 24167 25823
rect 24685 25789 24719 25823
rect 24869 25789 24903 25823
rect 26249 25789 26283 25823
rect 26525 25789 26559 25823
rect 23765 25721 23799 25755
rect 4169 25653 4203 25687
rect 4445 25653 4479 25687
rect 8861 25653 8895 25687
rect 10793 25653 10827 25687
rect 11161 25653 11195 25687
rect 18153 25653 18187 25687
rect 26065 25653 26099 25687
rect 11989 25449 12023 25483
rect 25421 25449 25455 25483
rect 6929 25313 6963 25347
rect 7757 25313 7791 25347
rect 11805 25313 11839 25347
rect 16773 25313 16807 25347
rect 17325 25313 17359 25347
rect 17509 25313 17543 25347
rect 24409 25313 24443 25347
rect 24961 25313 24995 25347
rect 25145 25313 25179 25347
rect 5273 25245 5307 25279
rect 5549 25245 5583 25279
rect 7849 25245 7883 25279
rect 16497 25245 16531 25279
rect 16589 25245 16623 25279
rect 24225 25245 24259 25279
rect 7113 25109 7147 25143
rect 17785 25109 17819 25143
rect 24041 25109 24075 25143
rect 13185 24905 13219 24939
rect 13369 24837 13403 24871
rect 2881 24769 2915 24803
rect 8309 24769 8343 24803
rect 10057 24769 10091 24803
rect 13645 24769 13679 24803
rect 18337 24769 18371 24803
rect 19717 24769 19751 24803
rect 25513 24769 25547 24803
rect 2605 24701 2639 24735
rect 7481 24701 7515 24735
rect 7573 24701 7607 24735
rect 7849 24701 7883 24735
rect 8033 24701 8067 24735
rect 8125 24701 8159 24735
rect 9413 24701 9447 24735
rect 10241 24701 10275 24735
rect 10793 24701 10827 24735
rect 10977 24701 11011 24735
rect 12449 24701 12483 24735
rect 13722 24701 13756 24735
rect 14197 24701 14231 24735
rect 14289 24701 14323 24735
rect 15899 24701 15933 24735
rect 16037 24701 16071 24735
rect 16497 24701 16531 24735
rect 16681 24701 16715 24735
rect 17877 24701 17911 24735
rect 18061 24701 18095 24735
rect 23857 24701 23891 24735
rect 24133 24701 24167 24735
rect 26341 24701 26375 24735
rect 4261 24633 4295 24667
rect 6837 24633 6871 24667
rect 9873 24633 9907 24667
rect 17325 24633 17359 24667
rect 4445 24565 4479 24599
rect 9229 24565 9263 24599
rect 11253 24565 11287 24599
rect 11621 24565 11655 24599
rect 12541 24565 12575 24599
rect 14749 24565 14783 24599
rect 15669 24565 15703 24599
rect 16957 24565 16991 24599
rect 23765 24565 23799 24599
rect 26433 24565 26467 24599
rect 23121 24361 23155 24395
rect 24501 24361 24535 24395
rect 28641 24361 28675 24395
rect 19901 24293 19935 24327
rect 28365 24293 28399 24327
rect 5365 24225 5399 24259
rect 9965 24225 9999 24259
rect 15485 24225 15519 24259
rect 16865 24225 16899 24259
rect 19717 24225 19751 24259
rect 22201 24225 22235 24259
rect 23305 24225 23339 24259
rect 23489 24225 23523 24259
rect 24041 24225 24075 24259
rect 24225 24225 24259 24259
rect 26525 24225 26559 24259
rect 27353 24225 27387 24259
rect 5641 24157 5675 24191
rect 7205 24157 7239 24191
rect 9505 24157 9539 24191
rect 9689 24157 9723 24191
rect 15577 24157 15611 24191
rect 16589 24157 16623 24191
rect 18337 24157 18371 24191
rect 28917 24225 28951 24259
rect 19533 24089 19567 24123
rect 22109 24089 22143 24123
rect 27445 24089 27479 24123
rect 28365 24089 28399 24123
rect 28733 24089 28767 24123
rect 6929 24021 6963 24055
rect 11253 24021 11287 24055
rect 15853 24021 15887 24055
rect 17969 24021 18003 24055
rect 22385 24021 22419 24055
rect 26709 24021 26743 24055
rect 4445 23817 4479 23851
rect 5825 23817 5859 23851
rect 11253 23817 11287 23851
rect 14105 23817 14139 23851
rect 18429 23817 18463 23851
rect 23949 23817 23983 23851
rect 26249 23817 26283 23851
rect 28641 23817 28675 23851
rect 10425 23749 10459 23783
rect 2881 23681 2915 23715
rect 7481 23681 7515 23715
rect 8585 23681 8619 23715
rect 2605 23613 2639 23647
rect 5733 23613 5767 23647
rect 7113 23613 7147 23647
rect 7389 23613 7423 23647
rect 8861 23613 8895 23647
rect 11069 23613 11103 23647
rect 14197 23613 14231 23647
rect 14473 23613 14507 23647
rect 18061 23613 18095 23647
rect 21833 23613 21867 23647
rect 23765 23613 23799 23647
rect 24685 23613 24719 23647
rect 24961 23613 24995 23647
rect 10241 23545 10275 23579
rect 10977 23545 11011 23579
rect 15853 23545 15887 23579
rect 27077 23545 27111 23579
rect 27169 23545 27203 23579
rect 3985 23477 4019 23511
rect 7757 23477 7791 23511
rect 18153 23477 18187 23511
rect 21925 23477 21959 23511
rect 22201 23477 22235 23511
rect 24225 23477 24259 23511
rect 24593 23477 24627 23511
rect 11989 23205 12023 23239
rect 15117 23205 15151 23239
rect 20729 23205 20763 23239
rect 22569 23205 22603 23239
rect 25421 23205 25455 23239
rect 11529 23137 11563 23171
rect 11713 23137 11747 23171
rect 14197 23137 14231 23171
rect 15945 23137 15979 23171
rect 16313 23137 16347 23171
rect 16497 23137 16531 23171
rect 20913 23137 20947 23171
rect 24317 23137 24351 23171
rect 24869 23137 24903 23171
rect 25053 23137 25087 23171
rect 26709 23137 26743 23171
rect 27261 23137 27295 23171
rect 27445 23137 27479 23171
rect 14013 23069 14047 23103
rect 15761 23069 15795 23103
rect 21189 23069 21223 23103
rect 23949 23069 23983 23103
rect 24133 23069 24167 23103
rect 26525 23069 26559 23103
rect 12173 22933 12207 22967
rect 14289 22933 14323 22967
rect 14841 22933 14875 22967
rect 15577 22933 15611 22967
rect 26249 22933 26283 22967
rect 27721 22933 27755 22967
rect 28089 22729 28123 22763
rect 4629 22661 4663 22695
rect 10057 22661 10091 22695
rect 14841 22661 14875 22695
rect 21189 22661 21223 22695
rect 2881 22593 2915 22627
rect 4445 22593 4479 22627
rect 8309 22593 8343 22627
rect 13645 22593 13679 22627
rect 26433 22593 26467 22627
rect 26525 22593 26559 22627
rect 26801 22593 26835 22627
rect 2605 22525 2639 22559
rect 8585 22525 8619 22559
rect 13921 22525 13955 22559
rect 14013 22525 14047 22559
rect 14473 22525 14507 22559
rect 14657 22525 14691 22559
rect 18061 22525 18095 22559
rect 20269 22525 20303 22559
rect 20361 22525 20395 22559
rect 20821 22525 20855 22559
rect 21005 22525 21039 22559
rect 9965 22457 9999 22491
rect 19993 22457 20027 22491
rect 3985 22389 4019 22423
rect 18153 22389 18187 22423
rect 18429 22389 18463 22423
rect 8585 22185 8619 22219
rect 18613 22117 18647 22151
rect 22293 22117 22327 22151
rect 7573 22049 7607 22083
rect 8125 22049 8159 22083
rect 8309 22049 8343 22083
rect 9689 22049 9723 22083
rect 10057 22049 10091 22083
rect 12173 22049 12207 22083
rect 16773 22049 16807 22083
rect 16957 22049 16991 22083
rect 20453 22049 20487 22083
rect 21557 22049 21591 22083
rect 21925 22049 21959 22083
rect 22109 22049 22143 22083
rect 27629 22049 27663 22083
rect 27721 22049 27755 22083
rect 7389 21981 7423 22015
rect 15117 21981 15151 22015
rect 17233 21981 17267 22015
rect 20913 21981 20947 22015
rect 21649 21981 21683 22015
rect 7205 21845 7239 21879
rect 9781 21845 9815 21879
rect 11989 21845 12023 21879
rect 12357 21845 12391 21879
rect 15117 21845 15151 21879
rect 20729 21845 20763 21879
rect 3985 21641 4019 21675
rect 4629 21641 4663 21675
rect 10333 21641 10367 21675
rect 12725 21641 12759 21675
rect 16957 21641 16991 21675
rect 19349 21641 19383 21675
rect 9045 21573 9079 21607
rect 12817 21505 12851 21539
rect 21281 21505 21315 21539
rect 2605 21437 2639 21471
rect 2881 21437 2915 21471
rect 4353 21437 4387 21471
rect 7941 21437 7975 21471
rect 8125 21437 8159 21471
rect 8677 21437 8711 21471
rect 8861 21437 8895 21471
rect 10149 21437 10183 21471
rect 11241 21437 11275 21471
rect 13093 21437 13127 21471
rect 15577 21437 15611 21471
rect 15761 21437 15795 21471
rect 15945 21437 15979 21471
rect 16497 21437 16531 21471
rect 16681 21437 16715 21471
rect 19257 21437 19291 21471
rect 21465 21437 21499 21471
rect 22017 21437 22051 21471
rect 22201 21437 22235 21471
rect 23673 21437 23707 21471
rect 14473 21369 14507 21403
rect 22569 21369 22603 21403
rect 23765 21369 23799 21403
rect 7757 21301 7791 21335
rect 11437 21301 11471 21335
rect 21189 21301 21223 21335
rect 23949 21301 23983 21335
rect 9781 21097 9815 21131
rect 9965 21097 9999 21131
rect 11621 21097 11655 21131
rect 14289 21097 14323 21131
rect 27905 21097 27939 21131
rect 13001 21029 13035 21063
rect 9689 20961 9723 20995
rect 10701 20961 10735 20995
rect 11713 20961 11747 20995
rect 11897 20961 11931 20995
rect 12449 20961 12483 20995
rect 12633 20961 12667 20995
rect 13921 20961 13955 20995
rect 15761 20961 15795 20995
rect 15945 20961 15979 20995
rect 16313 20961 16347 20995
rect 16497 20961 16531 20995
rect 19257 20961 19291 20995
rect 22661 20961 22695 20995
rect 14013 20893 14047 20927
rect 15301 20893 15335 20927
rect 22385 20893 22419 20927
rect 26525 20893 26559 20927
rect 26801 20893 26835 20927
rect 15025 20825 15059 20859
rect 24133 20825 24167 20859
rect 26249 20825 26283 20859
rect 10793 20757 10827 20791
rect 14841 20757 14875 20791
rect 19441 20757 19475 20791
rect 23949 20757 23983 20791
rect 4445 20553 4479 20587
rect 12633 20553 12667 20587
rect 20821 20553 20855 20587
rect 21189 20553 21223 20587
rect 22845 20553 22879 20587
rect 25789 20553 25823 20587
rect 27445 20553 27479 20587
rect 21373 20485 21407 20519
rect 2605 20417 2639 20451
rect 20545 20417 20579 20451
rect 22109 20417 22143 20451
rect 26157 20417 26191 20451
rect 2881 20349 2915 20383
rect 10701 20349 10735 20383
rect 10885 20349 10919 20383
rect 12449 20349 12483 20383
rect 14749 20349 14783 20383
rect 19717 20349 19751 20383
rect 19901 20349 19935 20383
rect 20177 20349 20211 20383
rect 20729 20349 20763 20383
rect 22201 20349 22235 20383
rect 22569 20349 22603 20383
rect 22753 20349 22787 20383
rect 25881 20349 25915 20383
rect 11253 20281 11287 20315
rect 19257 20281 19291 20315
rect 21557 20281 21591 20315
rect 3985 20213 4019 20247
rect 14841 20213 14875 20247
rect 18889 20213 18923 20247
rect 19165 20213 19199 20247
rect 2789 20009 2823 20043
rect 4813 20009 4847 20043
rect 6009 20009 6043 20043
rect 11437 20009 11471 20043
rect 12909 20009 12943 20043
rect 17233 20009 17267 20043
rect 25421 20009 25455 20043
rect 27537 20009 27571 20043
rect 25697 19941 25731 19975
rect 25881 19941 25915 19975
rect 2881 19873 2915 19907
rect 4629 19873 4663 19907
rect 5825 19873 5859 19907
rect 9505 19873 9539 19907
rect 9781 19873 9815 19907
rect 10057 19873 10091 19907
rect 10517 19873 10551 19907
rect 11621 19873 11655 19907
rect 12725 19873 12759 19907
rect 15301 19873 15335 19907
rect 16037 19873 16071 19907
rect 16221 19873 16255 19907
rect 16497 19873 16531 19907
rect 24409 19873 24443 19907
rect 24961 19873 24995 19907
rect 25145 19873 25179 19907
rect 26617 19873 26651 19907
rect 27629 19873 27663 19907
rect 15025 19805 15059 19839
rect 10517 19737 10551 19771
rect 15577 19805 15611 19839
rect 16773 19805 16807 19839
rect 16957 19805 16991 19839
rect 24317 19805 24351 19839
rect 26985 19805 27019 19839
rect 24133 19737 24167 19771
rect 27721 19737 27755 19771
rect 3065 19669 3099 19703
rect 10977 19669 11011 19703
rect 11805 19669 11839 19703
rect 15301 19669 15335 19703
rect 15393 19669 15427 19703
rect 26709 19669 26743 19703
rect 10333 19465 10367 19499
rect 11161 19465 11195 19499
rect 16773 19465 16807 19499
rect 20729 19465 20763 19499
rect 7941 19329 7975 19363
rect 9137 19329 9171 19363
rect 10149 19329 10183 19363
rect 15485 19329 15519 19363
rect 2605 19261 2639 19295
rect 2881 19261 2915 19295
rect 5273 19261 5307 19295
rect 5825 19261 5859 19295
rect 7113 19261 7147 19295
rect 9597 19261 9631 19295
rect 9873 19261 9907 19295
rect 10977 19261 11011 19295
rect 15209 19261 15243 19295
rect 19349 19261 19383 19295
rect 19625 19261 19659 19295
rect 25237 19261 25271 19295
rect 25329 19261 25363 19295
rect 25697 19261 25731 19295
rect 25789 19261 25823 19295
rect 26525 19261 26559 19295
rect 26709 19261 26743 19295
rect 4353 19193 4387 19227
rect 5089 19193 5123 19227
rect 5641 19193 5675 19227
rect 7205 19193 7239 19227
rect 7573 19193 7607 19227
rect 8953 19193 8987 19227
rect 26341 19193 26375 19227
rect 3985 19125 4019 19159
rect 7389 19125 7423 19159
rect 7481 19125 7515 19159
rect 15117 19125 15151 19159
rect 19165 19125 19199 19159
rect 24961 19125 24995 19159
rect 4169 18921 4203 18955
rect 10609 18921 10643 18955
rect 11529 18921 11563 18955
rect 16221 18921 16255 18955
rect 23857 18921 23891 18955
rect 4537 18853 4571 18887
rect 9873 18853 9907 18887
rect 10057 18853 10091 18887
rect 10425 18853 10459 18887
rect 11621 18853 11655 18887
rect 18153 18853 18187 18887
rect 4353 18785 4387 18819
rect 4629 18785 4663 18819
rect 9965 18785 9999 18819
rect 11437 18785 11471 18819
rect 11989 18785 12023 18819
rect 15485 18785 15519 18819
rect 15577 18785 15611 18819
rect 16865 18785 16899 18819
rect 18429 18785 18463 18819
rect 18981 18785 19015 18819
rect 19165 18785 19199 18819
rect 19441 18785 19475 18819
rect 19809 18785 19843 18819
rect 20085 18785 20119 18819
rect 24869 18785 24903 18819
rect 25237 18785 25271 18819
rect 9689 18717 9723 18751
rect 11253 18717 11287 18751
rect 18521 18717 18555 18751
rect 19901 18717 19935 18751
rect 24225 18717 24259 18751
rect 24961 18717 24995 18751
rect 25145 18717 25179 18751
rect 4813 18581 4847 18615
rect 15761 18581 15795 18615
rect 17049 18581 17083 18615
rect 24041 18581 24075 18615
rect 15117 18377 15151 18411
rect 27721 18377 27755 18411
rect 7021 18309 7055 18343
rect 13737 18309 13771 18343
rect 15301 18309 15335 18343
rect 21189 18309 21223 18343
rect 27445 18309 27479 18343
rect 2697 18241 2731 18275
rect 3709 18241 3743 18275
rect 5825 18241 5859 18275
rect 9505 18241 9539 18275
rect 20085 18241 20119 18275
rect 2513 18173 2547 18207
rect 2605 18173 2639 18207
rect 3617 18173 3651 18207
rect 3893 18173 3927 18207
rect 5181 18173 5215 18207
rect 5273 18173 5307 18207
rect 5457 18173 5491 18207
rect 6837 18173 6871 18207
rect 7941 18173 7975 18207
rect 9781 18173 9815 18207
rect 12909 18173 12943 18207
rect 13461 18173 13495 18207
rect 13737 18173 13771 18207
rect 14988 18173 15022 18207
rect 15180 18173 15214 18207
rect 16405 18173 16439 18207
rect 19533 18173 19567 18207
rect 19809 18173 19843 18207
rect 24961 18173 24995 18207
rect 25145 18173 25179 18207
rect 25329 18173 25363 18207
rect 25789 18173 25823 18207
rect 25881 18173 25915 18207
rect 27353 18173 27387 18207
rect 4353 18105 4387 18139
rect 9873 18105 9907 18139
rect 10241 18105 10275 18139
rect 14841 18105 14875 18139
rect 26433 18105 26467 18139
rect 3249 18037 3283 18071
rect 3433 18037 3467 18071
rect 8125 18037 8159 18071
rect 9689 18037 9723 18071
rect 12817 18037 12851 18071
rect 16589 18037 16623 18071
rect 19533 18037 19567 18071
rect 19625 18037 19659 18071
rect 4537 17833 4571 17867
rect 8585 17833 8619 17867
rect 10425 17833 10459 17867
rect 23029 17833 23063 17867
rect 24133 17833 24167 17867
rect 26249 17833 26283 17867
rect 27905 17833 27939 17867
rect 6745 17765 6779 17799
rect 10517 17765 10551 17799
rect 10609 17765 10643 17799
rect 10977 17765 11011 17799
rect 11989 17765 12023 17799
rect 12173 17765 12207 17799
rect 21557 17765 21591 17799
rect 23949 17765 23983 17799
rect 2973 17697 3007 17731
rect 4077 17697 4111 17731
rect 4353 17697 4387 17731
rect 6009 17697 6043 17731
rect 6285 17697 6319 17731
rect 8401 17697 8435 17731
rect 11161 17697 11195 17731
rect 12081 17697 12115 17731
rect 16589 17697 16623 17731
rect 16681 17697 16715 17731
rect 16865 17697 16899 17731
rect 17325 17697 17359 17731
rect 19809 17697 19843 17731
rect 20913 17697 20947 17731
rect 21005 17697 21039 17731
rect 22385 17697 22419 17731
rect 24961 17697 24995 17731
rect 25329 17697 25363 17731
rect 25513 17697 25547 17731
rect 26801 17697 26835 17731
rect 3065 17629 3099 17663
rect 10241 17629 10275 17663
rect 11805 17629 11839 17663
rect 12541 17629 12575 17663
rect 16037 17629 16071 17663
rect 17417 17629 17451 17663
rect 21465 17629 21499 17663
rect 22293 17629 22327 17663
rect 24317 17629 24351 17663
rect 25053 17629 25087 17663
rect 26525 17629 26559 17663
rect 4169 17561 4203 17595
rect 6101 17561 6135 17595
rect 2881 17493 2915 17527
rect 3801 17493 3835 17527
rect 19901 17493 19935 17527
rect 22569 17493 22603 17527
rect 5549 17289 5583 17323
rect 5825 17289 5859 17323
rect 12725 17289 12759 17323
rect 16865 17289 16899 17323
rect 21373 17289 21407 17323
rect 21833 17289 21867 17323
rect 3249 17221 3283 17255
rect 17233 17221 17267 17255
rect 9689 17153 9723 17187
rect 9965 17153 9999 17187
rect 11437 17153 11471 17187
rect 14013 17153 14047 17187
rect 14657 17153 14691 17187
rect 16589 17153 16623 17187
rect 21557 17153 21591 17187
rect 25421 17153 25455 17187
rect 3065 17085 3099 17119
rect 4169 17085 4203 17119
rect 4261 17085 4295 17119
rect 4445 17085 4479 17119
rect 4905 17085 4939 17119
rect 5733 17085 5767 17119
rect 9045 17085 9079 17119
rect 9229 17085 9263 17119
rect 9413 17085 9447 17119
rect 10885 17085 10919 17119
rect 10977 17085 11011 17119
rect 12449 17085 12483 17119
rect 13829 17085 13863 17119
rect 14105 17085 14139 17119
rect 14197 17085 14231 17119
rect 15485 17085 15519 17119
rect 16681 17085 16715 17119
rect 20177 17085 20211 17119
rect 20269 17085 20303 17119
rect 21649 17085 21683 17119
rect 25605 17085 25639 17119
rect 26157 17085 26191 17119
rect 26341 17085 26375 17119
rect 8585 17017 8619 17051
rect 20729 17017 20763 17051
rect 26709 17017 26743 17051
rect 2973 16949 3007 16983
rect 12541 16949 12575 16983
rect 15577 16949 15611 16983
rect 20913 16949 20947 16983
rect 25237 16949 25271 16983
rect 3065 16745 3099 16779
rect 4261 16745 4295 16779
rect 5365 16745 5399 16779
rect 13185 16745 13219 16779
rect 17509 16745 17543 16779
rect 20637 16745 20671 16779
rect 22569 16745 22603 16779
rect 9505 16677 9539 16711
rect 2881 16609 2915 16643
rect 4077 16609 4111 16643
rect 4445 16609 4479 16643
rect 5181 16609 5215 16643
rect 9689 16609 9723 16643
rect 10057 16609 10091 16643
rect 10241 16609 10275 16643
rect 10517 16609 10551 16643
rect 10609 16609 10643 16643
rect 11345 16609 11379 16643
rect 13277 16609 13311 16643
rect 13369 16609 13403 16643
rect 15853 16609 15887 16643
rect 16405 16609 16439 16643
rect 16589 16609 16623 16643
rect 16681 16609 16715 16643
rect 17141 16609 17175 16643
rect 19809 16609 19843 16643
rect 19901 16609 19935 16643
rect 20913 16609 20947 16643
rect 21097 16609 21131 16643
rect 21465 16609 21499 16643
rect 21741 16609 21775 16643
rect 21925 16609 21959 16643
rect 23213 16609 23247 16643
rect 10977 16541 11011 16575
rect 13829 16541 13863 16575
rect 17233 16541 17267 16575
rect 2789 16405 2823 16439
rect 12909 16405 12943 16439
rect 22293 16405 22327 16439
rect 23305 16405 23339 16439
rect 5273 16201 5307 16235
rect 13185 16201 13219 16235
rect 27261 16201 27295 16235
rect 2605 16065 2639 16099
rect 2881 16065 2915 16099
rect 9229 16065 9263 16099
rect 13645 16065 13679 16099
rect 14197 16065 14231 16099
rect 15669 16065 15703 16099
rect 21189 16065 21223 16099
rect 5089 15997 5123 16031
rect 7021 15997 7055 16031
rect 9413 15997 9447 16031
rect 9781 15997 9815 16031
rect 9965 15997 9999 16031
rect 10149 15997 10183 16031
rect 10701 15997 10735 16031
rect 13737 15997 13771 16031
rect 14105 15997 14139 16031
rect 15117 15997 15151 16031
rect 15209 15997 15243 16031
rect 20729 15997 20763 16031
rect 21005 15997 21039 16031
rect 21557 15997 21591 16031
rect 21741 15997 21775 16031
rect 21925 15997 21959 16031
rect 22201 15997 22235 16031
rect 23673 15997 23707 16031
rect 27169 15997 27203 16031
rect 6837 15929 6871 15963
rect 10885 15929 10919 15963
rect 20545 15929 20579 15963
rect 3985 15861 4019 15895
rect 4353 15861 4387 15895
rect 7113 15861 7147 15895
rect 9137 15861 9171 15895
rect 20821 15861 20855 15895
rect 22569 15861 22603 15895
rect 23765 15861 23799 15895
rect 27537 15861 27571 15895
rect 5457 15657 5491 15691
rect 6377 15657 6411 15691
rect 8769 15657 8803 15691
rect 10149 15657 10183 15691
rect 12725 15657 12759 15691
rect 15393 15657 15427 15691
rect 21005 15657 21039 15691
rect 21465 15657 21499 15691
rect 24685 15657 24719 15691
rect 26249 15657 26283 15691
rect 6745 15589 6779 15623
rect 13645 15589 13679 15623
rect 28181 15589 28215 15623
rect 4353 15521 4387 15555
rect 5825 15521 5859 15555
rect 6561 15521 6595 15555
rect 6837 15521 6871 15555
rect 8401 15521 8435 15555
rect 9689 15521 9723 15555
rect 12633 15521 12667 15555
rect 13792 15521 13826 15555
rect 15485 15521 15519 15555
rect 15853 15521 15887 15555
rect 16037 15521 16071 15555
rect 16221 15521 16255 15555
rect 16497 15521 16531 15555
rect 21833 15521 21867 15555
rect 22201 15521 22235 15555
rect 22385 15521 22419 15555
rect 22569 15521 22603 15555
rect 24869 15521 24903 15555
rect 26525 15521 26559 15555
rect 26801 15521 26835 15555
rect 4077 15453 4111 15487
rect 6009 15453 6043 15487
rect 14013 15453 14047 15487
rect 17049 15453 17083 15487
rect 21649 15453 21683 15487
rect 9873 15385 9907 15419
rect 14105 15385 14139 15419
rect 23029 15385 23063 15419
rect 23213 15385 23247 15419
rect 7021 15317 7055 15351
rect 8493 15317 8527 15351
rect 13921 15317 13955 15351
rect 16865 15317 16899 15351
rect 25053 15317 25087 15351
rect 4353 15045 4387 15079
rect 4629 15045 4663 15079
rect 8953 15045 8987 15079
rect 2605 14977 2639 15011
rect 2881 14977 2915 15011
rect 7573 14977 7607 15011
rect 9321 14977 9355 15011
rect 19717 14977 19751 15011
rect 21097 14977 21131 15011
rect 25421 14977 25455 15011
rect 25513 14977 25547 15011
rect 27813 14977 27847 15011
rect 7849 14909 7883 14943
rect 12173 14909 12207 14943
rect 13093 14909 13127 14943
rect 14197 14909 14231 14943
rect 14381 14909 14415 14943
rect 14933 14909 14967 14943
rect 15117 14909 15151 14943
rect 19441 14909 19475 14943
rect 25697 14909 25731 14943
rect 26249 14909 26283 14943
rect 26433 14909 26467 14943
rect 27721 14909 27755 14943
rect 26801 14841 26835 14875
rect 3985 14773 4019 14807
rect 11989 14773 12023 14807
rect 13277 14773 13311 14807
rect 14105 14773 14139 14807
rect 15393 14773 15427 14807
rect 19349 14773 19383 14807
rect 9965 14569 9999 14603
rect 12909 14569 12943 14603
rect 15669 14569 15703 14603
rect 15945 14569 15979 14603
rect 20177 14569 20211 14603
rect 21097 14569 21131 14603
rect 26249 14569 26283 14603
rect 9781 14501 9815 14535
rect 28181 14501 28215 14535
rect 7205 14433 7239 14467
rect 7757 14433 7791 14467
rect 7941 14433 7975 14467
rect 9689 14433 9723 14467
rect 11529 14433 11563 14467
rect 12725 14433 12759 14467
rect 13921 14433 13955 14467
rect 14381 14433 14415 14467
rect 15577 14433 15611 14467
rect 19809 14433 19843 14467
rect 21925 14433 21959 14467
rect 22293 14433 22327 14467
rect 26525 14433 26559 14467
rect 26801 14433 26835 14467
rect 7021 14365 7055 14399
rect 13829 14365 13863 14399
rect 21833 14365 21867 14399
rect 22385 14365 22419 14399
rect 8125 14297 8159 14331
rect 21373 14297 21407 14331
rect 6929 14229 6963 14263
rect 11713 14229 11747 14263
rect 19901 14229 19935 14263
rect 22661 14229 22695 14263
rect 4445 14025 4479 14059
rect 19349 14025 19383 14059
rect 4629 13957 4663 13991
rect 14565 13957 14599 13991
rect 2605 13889 2639 13923
rect 2881 13889 2915 13923
rect 7849 13889 7883 13923
rect 8125 13889 8159 13923
rect 9505 13889 9539 13923
rect 14749 13889 14783 13923
rect 15025 13889 15059 13923
rect 16221 13889 16255 13923
rect 23765 13889 23799 13923
rect 24041 13889 24075 13923
rect 9597 13821 9631 13855
rect 17785 13821 17819 13855
rect 18153 13821 18187 13855
rect 18337 13821 18371 13855
rect 18889 13821 18923 13855
rect 19073 13821 19107 13855
rect 21189 13821 21223 13855
rect 21373 13821 21407 13855
rect 21557 13821 21591 13855
rect 22109 13821 22143 13855
rect 22293 13821 22327 13855
rect 23673 13821 23707 13855
rect 27629 13821 27663 13855
rect 22661 13753 22695 13787
rect 3985 13685 4019 13719
rect 27721 13685 27755 13719
rect 8033 13481 8067 13515
rect 13553 13481 13587 13515
rect 13921 13481 13955 13515
rect 26157 13481 26191 13515
rect 26249 13481 26283 13515
rect 16681 13413 16715 13447
rect 18521 13413 18555 13447
rect 24041 13413 24075 13447
rect 5733 13345 5767 13379
rect 7021 13345 7055 13379
rect 7573 13345 7607 13379
rect 7757 13345 7791 13379
rect 10977 13345 11011 13379
rect 13737 13345 13771 13379
rect 16865 13345 16899 13379
rect 22661 13345 22695 13379
rect 26709 13345 26743 13379
rect 27261 13345 27295 13379
rect 27445 13345 27479 13379
rect 6837 13277 6871 13311
rect 11253 13277 11287 13311
rect 12633 13277 12667 13311
rect 17141 13277 17175 13311
rect 22385 13277 22419 13311
rect 26157 13277 26191 13311
rect 26525 13277 26559 13311
rect 5917 13209 5951 13243
rect 24225 13209 24259 13243
rect 6653 13141 6687 13175
rect 12725 13141 12759 13175
rect 27721 13141 27755 13175
rect 4445 12937 4479 12971
rect 18429 12937 18463 12971
rect 21281 12937 21315 12971
rect 25053 12937 25087 12971
rect 25513 12937 25547 12971
rect 26341 12937 26375 12971
rect 28089 12937 28123 12971
rect 9965 12869 9999 12903
rect 11253 12869 11287 12903
rect 2881 12801 2915 12835
rect 6653 12801 6687 12835
rect 6837 12801 6871 12835
rect 10149 12801 10183 12835
rect 21373 12801 21407 12835
rect 22661 12801 22695 12835
rect 23949 12801 23983 12835
rect 26525 12801 26559 12835
rect 26801 12801 26835 12835
rect 2605 12733 2639 12767
rect 7021 12733 7055 12767
rect 7573 12733 7607 12767
rect 7757 12733 7791 12767
rect 9045 12733 9079 12767
rect 10333 12733 10367 12767
rect 10885 12733 10919 12767
rect 11069 12733 11103 12767
rect 12437 12733 12471 12767
rect 18061 12733 18095 12767
rect 21557 12733 21591 12767
rect 22109 12733 22143 12767
rect 22293 12733 22327 12767
rect 23673 12733 23707 12767
rect 9137 12665 9171 12699
rect 4169 12597 4203 12631
rect 4629 12597 4663 12631
rect 8033 12597 8067 12631
rect 8861 12597 8895 12631
rect 12633 12597 12667 12631
rect 18153 12597 18187 12631
rect 7941 12393 7975 12427
rect 11989 12393 12023 12427
rect 17509 12393 17543 12427
rect 22937 12393 22971 12427
rect 23213 12393 23247 12427
rect 12265 12325 12299 12359
rect 11897 12257 11931 12291
rect 13093 12257 13127 12291
rect 13553 12257 13587 12291
rect 16497 12257 16531 12291
rect 17049 12257 17083 12291
rect 17233 12257 17267 12291
rect 22845 12257 22879 12291
rect 6377 12189 6411 12223
rect 6653 12189 6687 12223
rect 16037 12189 16071 12223
rect 16313 12189 16347 12223
rect 8125 12053 8159 12087
rect 12909 12053 12943 12087
rect 13645 12053 13679 12087
rect 16037 12053 16071 12087
rect 16221 12053 16255 12087
rect 7573 11849 7607 11883
rect 12725 11849 12759 11883
rect 24501 11781 24535 11815
rect 2881 11713 2915 11747
rect 7389 11713 7423 11747
rect 12909 11713 12943 11747
rect 18613 11713 18647 11747
rect 20545 11713 20579 11747
rect 24869 11713 24903 11747
rect 25145 11713 25179 11747
rect 2605 11645 2639 11679
rect 6837 11645 6871 11679
rect 6929 11645 6963 11679
rect 8217 11645 8251 11679
rect 8309 11645 8343 11679
rect 13185 11645 13219 11679
rect 18889 11645 18923 11679
rect 20361 11645 20395 11679
rect 24317 11645 24351 11679
rect 24685 11645 24719 11679
rect 8769 11577 8803 11611
rect 14565 11577 14599 11611
rect 4169 11509 4203 11543
rect 4445 11509 4479 11543
rect 19993 11509 20027 11543
rect 26249 11509 26283 11543
rect 5273 11305 5307 11339
rect 12633 11305 12667 11339
rect 14105 11305 14139 11339
rect 15393 11305 15427 11339
rect 18245 11305 18279 11339
rect 20085 11305 20119 11339
rect 8033 11237 8067 11271
rect 5365 11169 5399 11203
rect 6561 11169 6595 11203
rect 7941 11169 7975 11203
rect 8125 11169 8159 11203
rect 8769 11169 8803 11203
rect 12725 11169 12759 11203
rect 15945 11169 15979 11203
rect 16313 11169 16347 11203
rect 18613 11169 18647 11203
rect 23765 11169 23799 11203
rect 6469 11101 6503 11135
rect 8585 11101 8619 11135
rect 13001 11101 13035 11135
rect 15853 11101 15887 11135
rect 16221 11101 16255 11135
rect 18245 11101 18279 11135
rect 18337 11101 18371 11135
rect 19717 11101 19751 11135
rect 22017 11101 22051 11135
rect 22293 11101 22327 11135
rect 5549 11033 5583 11067
rect 16589 11033 16623 11067
rect 6745 10965 6779 10999
rect 23581 10965 23615 10999
rect 7389 10761 7423 10795
rect 8309 10761 8343 10795
rect 22477 10761 22511 10795
rect 2881 10625 2915 10659
rect 8125 10625 8159 10659
rect 13829 10625 13863 10659
rect 14565 10625 14599 10659
rect 25881 10625 25915 10659
rect 2605 10557 2639 10591
rect 7665 10557 7699 10591
rect 14473 10557 14507 10591
rect 14841 10557 14875 10591
rect 15025 10557 15059 10591
rect 15853 10557 15887 10591
rect 21097 10557 21131 10591
rect 21373 10557 21407 10591
rect 25513 10557 25547 10591
rect 25605 10557 25639 10591
rect 7573 10489 7607 10523
rect 4169 10421 4203 10455
rect 4445 10421 4479 10455
rect 15209 10421 15243 10455
rect 16037 10421 16071 10455
rect 22845 10421 22879 10455
rect 26985 10421 27019 10455
rect 8493 10217 8527 10251
rect 11345 10217 11379 10251
rect 12449 10217 12483 10251
rect 15025 10217 15059 10251
rect 16681 10217 16715 10251
rect 21557 10217 21591 10251
rect 21741 10217 21775 10251
rect 5733 10081 5767 10115
rect 7481 10081 7515 10115
rect 8217 10081 8251 10115
rect 8401 10081 8435 10115
rect 11529 10081 11563 10115
rect 11713 10081 11747 10115
rect 11805 10081 11839 10115
rect 15301 10081 15335 10115
rect 20913 10081 20947 10115
rect 26341 10081 26375 10115
rect 26525 10081 26559 10115
rect 26801 10081 26835 10115
rect 6009 10013 6043 10047
rect 15577 10013 15611 10047
rect 7297 9877 7331 9911
rect 11989 9877 12023 9911
rect 27905 9877 27939 9911
rect 9137 9673 9171 9707
rect 12173 9673 12207 9707
rect 26249 9673 26283 9707
rect 12449 9605 12483 9639
rect 24225 9605 24259 9639
rect 24409 9605 24443 9639
rect 2881 9537 2915 9571
rect 6929 9537 6963 9571
rect 7757 9537 7791 9571
rect 8217 9537 8251 9571
rect 10701 9537 10735 9571
rect 15669 9537 15703 9571
rect 16129 9537 16163 9571
rect 16589 9537 16623 9571
rect 21649 9537 21683 9571
rect 26341 9537 26375 9571
rect 26617 9537 26651 9571
rect 2605 9469 2639 9503
rect 4445 9469 4479 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 7849 9469 7883 9503
rect 9045 9469 9079 9503
rect 10241 9469 10275 9503
rect 12725 9469 12759 9503
rect 16313 9469 16347 9503
rect 16681 9469 16715 9503
rect 24593 9469 24627 9503
rect 8861 9401 8895 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 4169 9333 4203 9367
rect 10425 9333 10459 9367
rect 22293 9333 22327 9367
rect 27721 9333 27755 9367
rect 13737 9129 13771 9163
rect 15485 9129 15519 9163
rect 13461 9061 13495 9095
rect 18245 9061 18279 9095
rect 11897 8993 11931 9027
rect 12081 8993 12115 9027
rect 12449 8993 12483 9027
rect 12541 8993 12575 9027
rect 13645 8993 13679 9027
rect 15393 8993 15427 9027
rect 22293 8993 22327 9027
rect 11437 8925 11471 8959
rect 15761 8925 15795 8959
rect 16589 8925 16623 8959
rect 16865 8925 16899 8959
rect 22845 8925 22879 8959
rect 23121 8925 23155 8959
rect 24225 8925 24259 8959
rect 18337 8789 18371 8823
rect 22109 8789 22143 8823
rect 22753 8789 22787 8823
rect 12725 8585 12759 8619
rect 22661 8585 22695 8619
rect 3985 8449 4019 8483
rect 9229 8449 9263 8483
rect 16405 8449 16439 8483
rect 18061 8449 18095 8483
rect 18521 8449 18555 8483
rect 18981 8449 19015 8483
rect 21097 8449 21131 8483
rect 21373 8449 21407 8483
rect 2605 8381 2639 8415
rect 2881 8381 2915 8415
rect 7573 8381 7607 8415
rect 7849 8381 7883 8415
rect 10057 8381 10091 8415
rect 10517 8381 10551 8415
rect 10701 8381 10735 8415
rect 11069 8381 11103 8415
rect 11253 8381 11287 8415
rect 12449 8381 12483 8415
rect 12633 8381 12667 8415
rect 16589 8381 16623 8415
rect 16928 8381 16962 8415
rect 17141 8381 17175 8415
rect 18705 8381 18739 8415
rect 19073 8381 19107 8415
rect 22937 8313 22971 8347
rect 4445 8245 4479 8279
rect 9413 8245 9447 8279
rect 16221 8245 16255 8279
rect 17509 8041 17543 8075
rect 25053 8041 25087 8075
rect 5825 7973 5859 8007
rect 12541 7973 12575 8007
rect 11161 7905 11195 7939
rect 16405 7905 16439 7939
rect 22109 7905 22143 7939
rect 4169 7837 4203 7871
rect 4445 7837 4479 7871
rect 10885 7837 10919 7871
rect 16129 7837 16163 7871
rect 17969 7837 18003 7871
rect 23673 7837 23707 7871
rect 23949 7837 23983 7871
rect 6009 7701 6043 7735
rect 12725 7701 12759 7735
rect 22753 7701 22787 7735
rect 23581 7701 23615 7735
rect 4629 7497 4663 7531
rect 4905 7497 4939 7531
rect 9229 7497 9263 7531
rect 15301 7497 15335 7531
rect 9413 7429 9447 7463
rect 3065 7361 3099 7395
rect 7665 7361 7699 7395
rect 15485 7361 15519 7395
rect 21741 7361 21775 7395
rect 3341 7293 3375 7327
rect 7941 7293 7975 7327
rect 15761 7293 15795 7327
rect 22385 7293 22419 7327
rect 17049 7157 17083 7191
rect 12725 6953 12759 6987
rect 13185 6953 13219 6987
rect 18429 6953 18463 6987
rect 23949 6953 23983 6987
rect 4721 6817 4755 6851
rect 11345 6817 11379 6851
rect 16681 6817 16715 6851
rect 16957 6817 16991 6851
rect 22845 6817 22879 6851
rect 4077 6749 4111 6783
rect 6653 6749 6687 6783
rect 11621 6749 11655 6783
rect 18061 6749 18095 6783
rect 22477 6749 22511 6783
rect 22569 6749 22603 6783
rect 7297 6681 7331 6715
rect 4445 6409 4479 6443
rect 8401 6409 8435 6443
rect 11437 6409 11471 6443
rect 11713 6409 11747 6443
rect 14381 6341 14415 6375
rect 2881 6273 2915 6307
rect 7113 6273 7147 6307
rect 13737 6273 13771 6307
rect 2605 6205 2639 6239
rect 6837 6205 6871 6239
rect 8677 6205 8711 6239
rect 9873 6205 9907 6239
rect 10149 6205 10183 6239
rect 3985 6069 4019 6103
rect 26801 5729 26835 5763
rect 26249 5661 26283 5695
rect 26525 5661 26559 5695
rect 26157 5593 26191 5627
rect 28089 5525 28123 5559
rect 4445 5321 4479 5355
rect 2881 5185 2915 5219
rect 2605 5117 2639 5151
rect 3985 4981 4019 5015
rect 7665 4777 7699 4811
rect 5917 4641 5951 4675
rect 6193 4573 6227 4607
rect 7297 4437 7331 4471
rect 4813 4233 4847 4267
rect 3157 4097 3191 4131
rect 4721 4097 4755 4131
rect 2881 4029 2915 4063
rect 4261 3893 4295 3927
rect 5089 3145 5123 3179
rect 3617 3009 3651 3043
rect 3341 2941 3375 2975
rect 5273 2941 5307 2975
rect 4721 2805 4755 2839
<< metal1 >>
rect 4062 44140 4068 44192
rect 4120 44180 4126 44192
rect 67266 44180 67272 44192
rect 4120 44152 67272 44180
rect 4120 44140 4126 44152
rect 67266 44140 67272 44152
rect 67324 44140 67330 44192
rect 1104 44090 111136 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 50326 44090
rect 50378 44038 50390 44090
rect 50442 44038 50454 44090
rect 50506 44038 50518 44090
rect 50570 44038 81046 44090
rect 81098 44038 81110 44090
rect 81162 44038 81174 44090
rect 81226 44038 81238 44090
rect 81290 44038 111136 44090
rect 1104 44016 111136 44038
rect 6089 43911 6147 43917
rect 6089 43908 6101 43911
rect 4632 43880 6101 43908
rect 4632 43849 4660 43880
rect 5184 43849 5212 43880
rect 6089 43877 6101 43880
rect 6135 43908 6147 43911
rect 6270 43908 6276 43920
rect 6135 43880 6276 43908
rect 6135 43877 6147 43880
rect 6089 43871 6147 43877
rect 6270 43868 6276 43880
rect 6328 43868 6334 43920
rect 40494 43908 40500 43920
rect 38488 43880 40500 43908
rect 4617 43843 4675 43849
rect 4617 43809 4629 43843
rect 4663 43809 4675 43843
rect 4617 43803 4675 43809
rect 5169 43843 5227 43849
rect 5169 43809 5181 43843
rect 5215 43809 5227 43843
rect 5169 43803 5227 43809
rect 5353 43843 5411 43849
rect 5353 43809 5365 43843
rect 5399 43840 5411 43843
rect 18877 43843 18935 43849
rect 5399 43812 6040 43840
rect 5399 43809 5411 43812
rect 5353 43803 5411 43809
rect 4525 43775 4583 43781
rect 4525 43741 4537 43775
rect 4571 43741 4583 43775
rect 4525 43735 4583 43741
rect 4540 43704 4568 43735
rect 4614 43704 4620 43716
rect 4540 43676 4620 43704
rect 4614 43664 4620 43676
rect 4672 43664 4678 43716
rect 5534 43704 5540 43716
rect 5495 43676 5540 43704
rect 5534 43664 5540 43676
rect 5592 43664 5598 43716
rect 6012 43645 6040 43812
rect 18877 43809 18889 43843
rect 18923 43840 18935 43843
rect 19426 43840 19432 43852
rect 18923 43812 19432 43840
rect 18923 43809 18935 43812
rect 18877 43803 18935 43809
rect 19426 43800 19432 43812
rect 19484 43800 19490 43852
rect 24210 43840 24216 43852
rect 24171 43812 24216 43840
rect 24210 43800 24216 43812
rect 24268 43840 24274 43852
rect 24765 43843 24823 43849
rect 24765 43840 24777 43843
rect 24268 43812 24777 43840
rect 24268 43800 24274 43812
rect 24765 43809 24777 43812
rect 24811 43809 24823 43843
rect 24765 43803 24823 43809
rect 24949 43843 25007 43849
rect 24949 43809 24961 43843
rect 24995 43840 25007 43843
rect 25590 43840 25596 43852
rect 24995 43812 25596 43840
rect 24995 43809 25007 43812
rect 24949 43803 25007 43809
rect 25590 43800 25596 43812
rect 25648 43800 25654 43852
rect 38488 43849 38516 43880
rect 40494 43868 40500 43880
rect 40552 43868 40558 43920
rect 38473 43843 38531 43849
rect 38473 43809 38485 43843
rect 38519 43809 38531 43843
rect 39022 43840 39028 43852
rect 38983 43812 39028 43840
rect 38473 43803 38531 43809
rect 39022 43800 39028 43812
rect 39080 43800 39086 43852
rect 39209 43843 39267 43849
rect 39209 43809 39221 43843
rect 39255 43840 39267 43843
rect 47305 43843 47363 43849
rect 39255 43812 39528 43840
rect 39255 43809 39267 43812
rect 39209 43803 39267 43809
rect 23842 43732 23848 43784
rect 23900 43772 23906 43784
rect 24029 43775 24087 43781
rect 24029 43772 24041 43775
rect 23900 43744 24041 43772
rect 23900 43732 23906 43744
rect 24029 43741 24041 43744
rect 24075 43741 24087 43775
rect 24029 43735 24087 43741
rect 25317 43775 25375 43781
rect 25317 43741 25329 43775
rect 25363 43772 25375 43775
rect 28994 43772 29000 43784
rect 25363 43744 29000 43772
rect 25363 43741 25375 43744
rect 25317 43735 25375 43741
rect 28994 43732 29000 43744
rect 29052 43732 29058 43784
rect 38289 43775 38347 43781
rect 38289 43772 38301 43775
rect 38028 43744 38301 43772
rect 17034 43664 17040 43716
rect 17092 43704 17098 43716
rect 18969 43707 19027 43713
rect 18969 43704 18981 43707
rect 17092 43676 18981 43704
rect 17092 43664 17098 43676
rect 18969 43673 18981 43676
rect 19015 43704 19027 43707
rect 36814 43704 36820 43716
rect 19015 43676 36820 43704
rect 19015 43673 19027 43676
rect 18969 43667 19027 43673
rect 36814 43664 36820 43676
rect 36872 43664 36878 43716
rect 5997 43639 6055 43645
rect 5997 43605 6009 43639
rect 6043 43636 6055 43639
rect 6914 43636 6920 43648
rect 6043 43608 6920 43636
rect 6043 43605 6055 43608
rect 5997 43599 6055 43605
rect 6914 43596 6920 43608
rect 6972 43596 6978 43648
rect 23842 43636 23848 43648
rect 23803 43608 23848 43636
rect 23842 43596 23848 43608
rect 23900 43596 23906 43648
rect 25590 43636 25596 43648
rect 25551 43608 25596 43636
rect 25590 43596 25596 43608
rect 25648 43596 25654 43648
rect 37642 43596 37648 43648
rect 37700 43636 37706 43648
rect 38028 43645 38056 43744
rect 38289 43741 38301 43744
rect 38335 43741 38347 43775
rect 38289 43735 38347 43741
rect 39390 43704 39396 43716
rect 39351 43676 39396 43704
rect 39390 43664 39396 43676
rect 39448 43664 39454 43716
rect 37829 43639 37887 43645
rect 37829 43636 37841 43639
rect 37700 43608 37841 43636
rect 37700 43596 37706 43608
rect 37829 43605 37841 43608
rect 37875 43636 37887 43639
rect 38013 43639 38071 43645
rect 38013 43636 38025 43639
rect 37875 43608 38025 43636
rect 37875 43605 37887 43608
rect 37829 43599 37887 43605
rect 38013 43605 38025 43608
rect 38059 43636 38071 43639
rect 39500 43636 39528 43812
rect 47305 43809 47317 43843
rect 47351 43840 47363 43843
rect 48038 43840 48044 43852
rect 47351 43812 48044 43840
rect 47351 43809 47363 43812
rect 47305 43803 47363 43809
rect 48038 43800 48044 43812
rect 48096 43800 48102 43852
rect 48501 43843 48559 43849
rect 48501 43809 48513 43843
rect 48547 43809 48559 43843
rect 48501 43803 48559 43809
rect 49697 43843 49755 43849
rect 49697 43809 49709 43843
rect 49743 43840 49755 43843
rect 49786 43840 49792 43852
rect 49743 43812 49792 43840
rect 49743 43809 49755 43812
rect 49697 43803 49755 43809
rect 47670 43732 47676 43784
rect 47728 43772 47734 43784
rect 48516 43772 48544 43803
rect 49786 43800 49792 43812
rect 49844 43800 49850 43852
rect 49881 43843 49939 43849
rect 49881 43809 49893 43843
rect 49927 43809 49939 43843
rect 61930 43840 61936 43852
rect 61891 43812 61936 43840
rect 49881 43803 49939 43809
rect 47728 43744 48544 43772
rect 48593 43775 48651 43781
rect 47728 43732 47734 43744
rect 48593 43741 48605 43775
rect 48639 43772 48651 43775
rect 49142 43772 49148 43784
rect 48639 43744 49148 43772
rect 48639 43741 48651 43744
rect 48593 43735 48651 43741
rect 49142 43732 49148 43744
rect 49200 43772 49206 43784
rect 49896 43772 49924 43803
rect 61930 43800 61936 43812
rect 61988 43800 61994 43852
rect 62025 43843 62083 43849
rect 62025 43809 62037 43843
rect 62071 43840 62083 43843
rect 63034 43840 63040 43852
rect 62071 43812 63040 43840
rect 62071 43809 62083 43812
rect 62025 43803 62083 43809
rect 63034 43800 63040 43812
rect 63092 43800 63098 43852
rect 69106 43800 69112 43852
rect 69164 43840 69170 43852
rect 69661 43843 69719 43849
rect 69661 43840 69673 43843
rect 69164 43812 69673 43840
rect 69164 43800 69170 43812
rect 69661 43809 69673 43812
rect 69707 43840 69719 43843
rect 69937 43843 69995 43849
rect 69937 43840 69949 43843
rect 69707 43812 69949 43840
rect 69707 43809 69719 43812
rect 69661 43803 69719 43809
rect 69937 43809 69949 43812
rect 69983 43840 69995 43843
rect 70302 43840 70308 43852
rect 69983 43812 70308 43840
rect 69983 43809 69995 43812
rect 69937 43803 69995 43809
rect 70302 43800 70308 43812
rect 70360 43800 70366 43852
rect 49200 43744 49924 43772
rect 49200 43732 49206 43744
rect 61749 43707 61807 43713
rect 61749 43673 61761 43707
rect 61795 43704 61807 43707
rect 62577 43707 62635 43713
rect 62577 43704 62589 43707
rect 61795 43676 62589 43704
rect 61795 43673 61807 43676
rect 61749 43667 61807 43673
rect 62577 43673 62589 43676
rect 62623 43704 62635 43707
rect 63494 43704 63500 43716
rect 62623 43676 63500 43704
rect 62623 43673 62635 43676
rect 62577 43667 62635 43673
rect 63494 43664 63500 43676
rect 63552 43664 63558 43716
rect 38059 43608 39528 43636
rect 38059 43605 38071 43608
rect 38013 43599 38071 43605
rect 46750 43596 46756 43648
rect 46808 43636 46814 43648
rect 47397 43639 47455 43645
rect 47397 43636 47409 43639
rect 46808 43608 47409 43636
rect 46808 43596 46814 43608
rect 47397 43605 47409 43608
rect 47443 43605 47455 43639
rect 47397 43599 47455 43605
rect 49234 43596 49240 43648
rect 49292 43636 49298 43648
rect 49973 43639 50031 43645
rect 49973 43636 49985 43639
rect 49292 43608 49985 43636
rect 49292 43596 49298 43608
rect 49973 43605 49985 43608
rect 50019 43605 50031 43639
rect 62206 43636 62212 43648
rect 62167 43608 62212 43636
rect 49973 43599 50031 43605
rect 62206 43596 62212 43608
rect 62264 43596 62270 43648
rect 69750 43636 69756 43648
rect 69711 43608 69756 43636
rect 69750 43596 69756 43608
rect 69808 43596 69814 43648
rect 1104 43546 111136 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 65686 43546
rect 65738 43494 65750 43546
rect 65802 43494 65814 43546
rect 65866 43494 65878 43546
rect 65930 43494 96406 43546
rect 96458 43494 96470 43546
rect 96522 43494 96534 43546
rect 96586 43494 96598 43546
rect 96650 43494 111136 43546
rect 1104 43472 111136 43494
rect 19426 43432 19432 43444
rect 19387 43404 19432 43432
rect 19426 43392 19432 43404
rect 19484 43392 19490 43444
rect 36814 43432 36820 43444
rect 36775 43404 36820 43432
rect 36814 43392 36820 43404
rect 36872 43432 36878 43444
rect 37001 43435 37059 43441
rect 37001 43432 37013 43435
rect 36872 43404 37013 43432
rect 36872 43392 36878 43404
rect 37001 43401 37013 43404
rect 37047 43401 37059 43435
rect 37001 43395 37059 43401
rect 3697 43299 3755 43305
rect 3697 43265 3709 43299
rect 3743 43296 3755 43299
rect 4798 43296 4804 43308
rect 3743 43268 4804 43296
rect 3743 43265 3755 43268
rect 3697 43259 3755 43265
rect 4798 43256 4804 43268
rect 4856 43256 4862 43308
rect 18230 43256 18236 43308
rect 18288 43296 18294 43308
rect 24949 43299 25007 43305
rect 18288 43268 23888 43296
rect 18288 43256 18294 43268
rect 3973 43231 4031 43237
rect 3973 43197 3985 43231
rect 4019 43228 4031 43231
rect 5074 43228 5080 43240
rect 4019 43200 5080 43228
rect 4019 43197 4031 43200
rect 3973 43191 4031 43197
rect 5074 43188 5080 43200
rect 5132 43188 5138 43240
rect 6454 43188 6460 43240
rect 6512 43228 6518 43240
rect 6825 43231 6883 43237
rect 6825 43228 6837 43231
rect 6512 43200 6837 43228
rect 6512 43188 6518 43200
rect 6825 43197 6837 43200
rect 6871 43197 6883 43231
rect 6825 43191 6883 43197
rect 9868 43231 9926 43237
rect 9868 43197 9880 43231
rect 9914 43228 9926 43231
rect 10137 43231 10195 43237
rect 9914 43200 9996 43228
rect 9914 43197 9926 43200
rect 9868 43191 9926 43197
rect 4798 43120 4804 43172
rect 4856 43160 4862 43172
rect 5537 43163 5595 43169
rect 5537 43160 5549 43163
rect 4856 43132 5549 43160
rect 4856 43120 4862 43132
rect 5537 43129 5549 43132
rect 5583 43160 5595 43163
rect 6638 43160 6644 43172
rect 5583 43132 6644 43160
rect 5583 43129 5595 43132
rect 5537 43123 5595 43129
rect 6638 43120 6644 43132
rect 6696 43160 6702 43172
rect 9674 43160 9680 43172
rect 6696 43132 9680 43160
rect 6696 43120 6702 43132
rect 9674 43120 9680 43132
rect 9732 43160 9738 43172
rect 9968 43160 9996 43200
rect 10137 43197 10149 43231
rect 10183 43228 10195 43231
rect 10778 43228 10784 43240
rect 10183 43200 10784 43228
rect 10183 43197 10195 43200
rect 10137 43191 10195 43197
rect 10778 43188 10784 43200
rect 10836 43188 10842 43240
rect 18049 43231 18107 43237
rect 18049 43197 18061 43231
rect 18095 43197 18107 43231
rect 18322 43228 18328 43240
rect 18283 43200 18328 43228
rect 18049 43191 18107 43197
rect 9732 43132 9996 43160
rect 11517 43163 11575 43169
rect 9732 43120 9738 43132
rect 11517 43129 11529 43163
rect 11563 43160 11575 43163
rect 12618 43160 12624 43172
rect 11563 43132 12624 43160
rect 11563 43129 11575 43132
rect 11517 43123 11575 43129
rect 12618 43120 12624 43132
rect 12676 43120 12682 43172
rect 5258 43092 5264 43104
rect 5219 43064 5264 43092
rect 5258 43052 5264 43064
rect 5316 43052 5322 43104
rect 6914 43092 6920 43104
rect 6827 43064 6920 43092
rect 6914 43052 6920 43064
rect 6972 43092 6978 43104
rect 8018 43092 8024 43104
rect 6972 43064 8024 43092
rect 6972 43052 6978 43064
rect 8018 43052 8024 43064
rect 8076 43052 8082 43104
rect 11698 43092 11704 43104
rect 11659 43064 11704 43092
rect 11698 43052 11704 43064
rect 11756 43052 11762 43104
rect 17678 43052 17684 43104
rect 17736 43092 17742 43104
rect 18064 43092 18092 43191
rect 18322 43188 18328 43200
rect 18380 43188 18386 43240
rect 23860 43237 23888 43268
rect 24949 43265 24961 43299
rect 24995 43296 25007 43299
rect 29086 43296 29092 43308
rect 24995 43268 29092 43296
rect 24995 43265 25007 43268
rect 24949 43259 25007 43265
rect 29086 43256 29092 43268
rect 29144 43256 29150 43308
rect 30466 43256 30472 43308
rect 30524 43296 30530 43308
rect 32585 43299 32643 43305
rect 32585 43296 32597 43299
rect 30524 43268 32597 43296
rect 30524 43256 30530 43268
rect 32585 43265 32597 43268
rect 32631 43265 32643 43299
rect 37016 43296 37044 43395
rect 45462 43392 45468 43444
rect 45520 43432 45526 43444
rect 49421 43435 49479 43441
rect 49421 43432 49433 43435
rect 45520 43404 49433 43432
rect 45520 43392 45526 43404
rect 49421 43401 49433 43404
rect 49467 43401 49479 43435
rect 49421 43395 49479 43401
rect 70302 43392 70308 43444
rect 70360 43432 70366 43444
rect 70489 43435 70547 43441
rect 70489 43432 70501 43435
rect 70360 43404 70501 43432
rect 70360 43392 70366 43404
rect 70489 43401 70501 43404
rect 70535 43401 70547 43435
rect 70489 43395 70547 43401
rect 48682 43324 48688 43376
rect 48740 43364 48746 43376
rect 50617 43367 50675 43373
rect 50617 43364 50629 43367
rect 48740 43336 50629 43364
rect 48740 43324 48746 43336
rect 50617 43333 50629 43336
rect 50663 43333 50675 43367
rect 66254 43364 66260 43376
rect 66215 43336 66260 43364
rect 50617 43327 50675 43333
rect 66254 43324 66260 43336
rect 66312 43324 66318 43376
rect 37185 43299 37243 43305
rect 37185 43296 37197 43299
rect 37016 43268 37197 43296
rect 32585 43259 32643 43265
rect 37185 43265 37197 43268
rect 37231 43296 37243 43299
rect 46750 43296 46756 43308
rect 37231 43268 37504 43296
rect 46711 43268 46756 43296
rect 37231 43265 37243 43268
rect 37185 43259 37243 43265
rect 23661 43231 23719 43237
rect 23661 43228 23673 43231
rect 23492 43200 23673 43228
rect 23492 43104 23520 43200
rect 23661 43197 23673 43200
rect 23707 43197 23719 43231
rect 23661 43191 23719 43197
rect 23845 43231 23903 43237
rect 23845 43197 23857 43231
rect 23891 43197 23903 43231
rect 23845 43191 23903 43197
rect 24397 43231 24455 43237
rect 24397 43197 24409 43231
rect 24443 43197 24455 43231
rect 24397 43191 24455 43197
rect 24581 43231 24639 43237
rect 24581 43197 24593 43231
rect 24627 43228 24639 43231
rect 26697 43231 26755 43237
rect 26697 43228 26709 43231
rect 24627 43200 25268 43228
rect 24627 43197 24639 43200
rect 24581 43191 24639 43197
rect 23860 43160 23888 43191
rect 24210 43160 24216 43172
rect 23860 43132 24216 43160
rect 24210 43120 24216 43132
rect 24268 43160 24274 43172
rect 24412 43160 24440 43191
rect 24268 43132 24440 43160
rect 24268 43120 24274 43132
rect 25240 43104 25268 43200
rect 26528 43200 26709 43228
rect 26528 43104 26556 43200
rect 26697 43197 26709 43200
rect 26743 43197 26755 43231
rect 26970 43228 26976 43240
rect 26931 43200 26976 43228
rect 26697 43191 26755 43197
rect 26970 43188 26976 43200
rect 27028 43188 27034 43240
rect 32309 43231 32367 43237
rect 32309 43197 32321 43231
rect 32355 43197 32367 43231
rect 32309 43191 32367 43197
rect 37369 43231 37427 43237
rect 37369 43197 37381 43231
rect 37415 43197 37427 43231
rect 37476 43228 37504 43268
rect 46750 43256 46756 43268
rect 46808 43256 46814 43308
rect 59265 43299 59323 43305
rect 59265 43265 59277 43299
rect 59311 43296 59323 43299
rect 61102 43296 61108 43308
rect 59311 43268 61108 43296
rect 59311 43265 59323 43268
rect 59265 43259 59323 43265
rect 61102 43256 61108 43268
rect 61160 43256 61166 43308
rect 37829 43231 37887 43237
rect 37829 43228 37841 43231
rect 37476 43200 37841 43228
rect 37369 43191 37427 43197
rect 37829 43197 37841 43200
rect 37875 43197 37887 43231
rect 37829 43191 37887 43197
rect 37921 43231 37979 43237
rect 37921 43197 37933 43231
rect 37967 43228 37979 43231
rect 39022 43228 39028 43240
rect 37967 43200 39028 43228
rect 37967 43197 37979 43200
rect 37921 43191 37979 43197
rect 28353 43163 28411 43169
rect 28353 43129 28365 43163
rect 28399 43160 28411 43163
rect 29730 43160 29736 43172
rect 28399 43132 29736 43160
rect 28399 43129 28411 43132
rect 28353 43123 28411 43129
rect 29730 43120 29736 43132
rect 29788 43120 29794 43172
rect 19242 43092 19248 43104
rect 17736 43064 19248 43092
rect 17736 43052 17742 43064
rect 19242 43052 19248 43064
rect 19300 43092 19306 43104
rect 19797 43095 19855 43101
rect 19797 43092 19809 43095
rect 19300 43064 19809 43092
rect 19300 43052 19306 43064
rect 19797 43061 19809 43064
rect 19843 43061 19855 43095
rect 23474 43092 23480 43104
rect 23435 43064 23480 43092
rect 19797 43055 19855 43061
rect 23474 43052 23480 43064
rect 23532 43052 23538 43104
rect 25222 43092 25228 43104
rect 25183 43064 25228 43092
rect 25222 43052 25228 43064
rect 25280 43052 25286 43104
rect 26510 43092 26516 43104
rect 26471 43064 26516 43092
rect 26510 43052 26516 43064
rect 26568 43052 26574 43104
rect 32324 43092 32352 43191
rect 33965 43163 34023 43169
rect 33965 43129 33977 43163
rect 34011 43160 34023 43163
rect 34790 43160 34796 43172
rect 34011 43132 34796 43160
rect 34011 43129 34023 43132
rect 33965 43123 34023 43129
rect 34790 43120 34796 43132
rect 34848 43120 34854 43172
rect 37384 43160 37412 43191
rect 37936 43160 37964 43191
rect 39022 43188 39028 43200
rect 39080 43188 39086 43240
rect 40494 43228 40500 43240
rect 40455 43200 40500 43228
rect 40494 43188 40500 43200
rect 40552 43188 40558 43240
rect 42337 43231 42395 43237
rect 42337 43197 42349 43231
rect 42383 43197 42395 43231
rect 42337 43191 42395 43197
rect 42613 43231 42671 43237
rect 42613 43197 42625 43231
rect 42659 43228 42671 43231
rect 43438 43228 43444 43240
rect 42659 43200 43444 43228
rect 42659 43197 42671 43200
rect 42613 43191 42671 43197
rect 38470 43160 38476 43172
rect 37384 43132 37964 43160
rect 38431 43132 38476 43160
rect 38470 43120 38476 43132
rect 38528 43120 38534 43172
rect 38562 43120 38568 43172
rect 38620 43160 38626 43172
rect 42153 43163 42211 43169
rect 42153 43160 42165 43163
rect 38620 43132 42165 43160
rect 38620 43120 38626 43132
rect 42153 43129 42165 43132
rect 42199 43160 42211 43163
rect 42352 43160 42380 43191
rect 43438 43188 43444 43200
rect 43496 43188 43502 43240
rect 46477 43231 46535 43237
rect 46477 43197 46489 43231
rect 46523 43228 46535 43231
rect 48317 43231 48375 43237
rect 48317 43228 48329 43231
rect 46523 43200 48329 43228
rect 46523 43197 46535 43200
rect 46477 43191 46535 43197
rect 48317 43197 48329 43200
rect 48363 43228 48375 43231
rect 48958 43228 48964 43240
rect 48363 43200 48964 43228
rect 48363 43197 48375 43200
rect 48317 43191 48375 43197
rect 48958 43188 48964 43200
rect 49016 43188 49022 43240
rect 49053 43231 49111 43237
rect 49053 43197 49065 43231
rect 49099 43197 49111 43231
rect 49234 43228 49240 43240
rect 49195 43200 49240 43228
rect 49053 43191 49111 43197
rect 42199 43132 42380 43160
rect 43640 43132 46612 43160
rect 42199 43129 42211 43132
rect 42153 43123 42211 43129
rect 34146 43092 34152 43104
rect 32324 43064 34152 43092
rect 34146 43052 34152 43064
rect 34204 43052 34210 43104
rect 39022 43052 39028 43104
rect 39080 43092 39086 43104
rect 40681 43095 40739 43101
rect 40681 43092 40693 43095
rect 39080 43064 40693 43092
rect 39080 43052 39086 43064
rect 40681 43061 40693 43064
rect 40727 43092 40739 43095
rect 43640 43092 43668 43132
rect 40727 43064 43668 43092
rect 40727 43061 40739 43064
rect 40681 43055 40739 43061
rect 43714 43052 43720 43104
rect 43772 43092 43778 43104
rect 46584 43092 46612 43132
rect 47670 43092 47676 43104
rect 43772 43064 43817 43092
rect 46584 43064 47676 43092
rect 43772 43052 43778 43064
rect 47670 43052 47676 43064
rect 47728 43052 47734 43104
rect 47854 43092 47860 43104
rect 47815 43064 47860 43092
rect 47854 43052 47860 43064
rect 47912 43052 47918 43104
rect 49068 43092 49096 43191
rect 49234 43188 49240 43200
rect 49292 43188 49298 43240
rect 49786 43188 49792 43240
rect 49844 43228 49850 43240
rect 50525 43231 50583 43237
rect 50525 43228 50537 43231
rect 49844 43200 50537 43228
rect 49844 43188 49850 43200
rect 50525 43197 50537 43200
rect 50571 43228 50583 43231
rect 50798 43228 50804 43240
rect 50571 43200 50804 43228
rect 50571 43197 50583 43200
rect 50525 43191 50583 43197
rect 50798 43188 50804 43200
rect 50856 43188 50862 43240
rect 55766 43228 55772 43240
rect 55727 43200 55772 43228
rect 55766 43188 55772 43200
rect 55824 43188 55830 43240
rect 56045 43231 56103 43237
rect 56045 43197 56057 43231
rect 56091 43197 56103 43231
rect 56226 43228 56232 43240
rect 56187 43200 56232 43228
rect 56045 43191 56103 43197
rect 49145 43163 49203 43169
rect 49145 43129 49157 43163
rect 49191 43160 49203 43163
rect 49326 43160 49332 43172
rect 49191 43132 49332 43160
rect 49191 43129 49203 43132
rect 49145 43123 49203 43129
rect 49326 43120 49332 43132
rect 49384 43120 49390 43172
rect 55214 43160 55220 43172
rect 55175 43132 55220 43160
rect 55214 43120 55220 43132
rect 55272 43120 55278 43172
rect 56060 43160 56088 43191
rect 56226 43188 56232 43200
rect 56284 43188 56290 43240
rect 59538 43228 59544 43240
rect 59499 43200 59544 43228
rect 59538 43188 59544 43200
rect 59596 43188 59602 43240
rect 66165 43231 66223 43237
rect 66165 43197 66177 43231
rect 66211 43197 66223 43231
rect 66530 43228 66536 43240
rect 66491 43200 66536 43228
rect 66165 43191 66223 43197
rect 56594 43160 56600 43172
rect 56060 43132 56600 43160
rect 56594 43120 56600 43132
rect 56652 43160 56658 43172
rect 57882 43160 57888 43172
rect 56652 43132 57888 43160
rect 56652 43120 56658 43132
rect 57882 43120 57888 43132
rect 57940 43120 57946 43172
rect 66180 43104 66208 43191
rect 66530 43188 66536 43200
rect 66588 43188 66594 43240
rect 66898 43228 66904 43240
rect 66859 43200 66904 43228
rect 66898 43188 66904 43200
rect 66956 43188 66962 43240
rect 69109 43231 69167 43237
rect 69109 43197 69121 43231
rect 69155 43197 69167 43231
rect 69382 43228 69388 43240
rect 69343 43200 69388 43228
rect 69109 43191 69167 43197
rect 66548 43160 66576 43188
rect 67177 43163 67235 43169
rect 67177 43160 67189 43163
rect 66548 43132 67189 43160
rect 67177 43129 67189 43132
rect 67223 43129 67235 43163
rect 67177 43123 67235 43129
rect 49881 43095 49939 43101
rect 49881 43092 49893 43095
rect 49068 43064 49893 43092
rect 49881 43061 49893 43064
rect 49927 43092 49939 43095
rect 49970 43092 49976 43104
rect 49927 43064 49976 43092
rect 49927 43061 49939 43064
rect 49881 43055 49939 43061
rect 49970 43052 49976 43064
rect 50028 43052 50034 43104
rect 60826 43092 60832 43104
rect 60787 43064 60832 43092
rect 60826 43052 60832 43064
rect 60884 43052 60890 43104
rect 61102 43092 61108 43104
rect 61063 43064 61108 43092
rect 61102 43052 61108 43064
rect 61160 43052 61166 43104
rect 66162 43052 66168 43104
rect 66220 43092 66226 43104
rect 67361 43095 67419 43101
rect 67361 43092 67373 43095
rect 66220 43064 67373 43092
rect 66220 43052 66226 43064
rect 67361 43061 67373 43064
rect 67407 43061 67419 43095
rect 67361 43055 67419 43061
rect 69017 43095 69075 43101
rect 69017 43061 69029 43095
rect 69063 43092 69075 43095
rect 69124 43092 69152 43191
rect 69382 43188 69388 43200
rect 69440 43188 69446 43240
rect 69658 43092 69664 43104
rect 69063 43064 69664 43092
rect 69063 43061 69075 43064
rect 69017 43055 69075 43061
rect 69658 43052 69664 43064
rect 69716 43052 69722 43104
rect 1104 43002 111136 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 50326 43002
rect 50378 42950 50390 43002
rect 50442 42950 50454 43002
rect 50506 42950 50518 43002
rect 50570 42950 81046 43002
rect 81098 42950 81110 43002
rect 81162 42950 81174 43002
rect 81226 42950 81238 43002
rect 81290 42950 111136 43002
rect 1104 42928 111136 42950
rect 6638 42888 6644 42900
rect 6599 42860 6644 42888
rect 6638 42848 6644 42860
rect 6696 42848 6702 42900
rect 18414 42888 18420 42900
rect 16316 42860 18420 42888
rect 6454 42820 6460 42832
rect 6415 42792 6460 42820
rect 6454 42780 6460 42792
rect 6512 42780 6518 42832
rect 15488 42792 15792 42820
rect 4798 42752 4804 42764
rect 4759 42724 4804 42752
rect 4798 42712 4804 42724
rect 4856 42712 4862 42764
rect 5077 42755 5135 42761
rect 5077 42721 5089 42755
rect 5123 42752 5135 42755
rect 5534 42752 5540 42764
rect 5123 42724 5540 42752
rect 5123 42721 5135 42724
rect 5077 42715 5135 42721
rect 5534 42712 5540 42724
rect 5592 42712 5598 42764
rect 9674 42712 9680 42764
rect 9732 42752 9738 42764
rect 10413 42755 10471 42761
rect 10413 42752 10425 42755
rect 9732 42724 10425 42752
rect 9732 42712 9738 42724
rect 10413 42721 10425 42724
rect 10459 42752 10471 42755
rect 12069 42755 12127 42761
rect 10459 42724 11744 42752
rect 10459 42721 10471 42724
rect 10413 42715 10471 42721
rect 11716 42696 11744 42724
rect 12069 42721 12081 42755
rect 12115 42752 12127 42755
rect 12897 42755 12955 42761
rect 12897 42752 12909 42755
rect 12115 42724 12909 42752
rect 12115 42721 12127 42724
rect 12069 42715 12127 42721
rect 12897 42721 12909 42724
rect 12943 42721 12955 42755
rect 12897 42715 12955 42721
rect 14090 42712 14096 42764
rect 14148 42752 14154 42764
rect 15381 42755 15439 42761
rect 15381 42752 15393 42755
rect 14148 42724 15393 42752
rect 14148 42712 14154 42724
rect 15381 42721 15393 42724
rect 15427 42752 15439 42755
rect 15488 42752 15516 42792
rect 15654 42752 15660 42764
rect 15427 42724 15516 42752
rect 15615 42724 15660 42752
rect 15427 42721 15439 42724
rect 15381 42715 15439 42721
rect 15654 42712 15660 42724
rect 15712 42712 15718 42764
rect 15764 42752 15792 42792
rect 16209 42755 16267 42761
rect 16209 42752 16221 42755
rect 15764 42724 16221 42752
rect 16209 42721 16221 42724
rect 16255 42752 16267 42755
rect 16316 42752 16344 42860
rect 18414 42848 18420 42860
rect 18472 42848 18478 42900
rect 19978 42848 19984 42900
rect 20036 42888 20042 42900
rect 25222 42888 25228 42900
rect 20036 42860 25228 42888
rect 20036 42848 20042 42860
rect 25222 42848 25228 42860
rect 25280 42848 25286 42900
rect 28445 42891 28503 42897
rect 28445 42857 28457 42891
rect 28491 42888 28503 42891
rect 38562 42888 38568 42900
rect 28491 42860 38568 42888
rect 28491 42857 28503 42860
rect 28445 42851 28503 42857
rect 38562 42848 38568 42860
rect 38620 42848 38626 42900
rect 40405 42891 40463 42897
rect 40405 42857 40417 42891
rect 40451 42888 40463 42891
rect 40494 42888 40500 42900
rect 40451 42860 40500 42888
rect 40451 42857 40463 42860
rect 40405 42851 40463 42857
rect 40494 42848 40500 42860
rect 40552 42848 40558 42900
rect 44910 42848 44916 42900
rect 44968 42888 44974 42900
rect 49421 42891 49479 42897
rect 49421 42888 49433 42891
rect 44968 42860 49433 42888
rect 44968 42848 44974 42860
rect 49421 42857 49433 42860
rect 49467 42857 49479 42891
rect 50798 42888 50804 42900
rect 50759 42860 50804 42888
rect 49421 42851 49479 42857
rect 50798 42848 50804 42860
rect 50856 42848 50862 42900
rect 55766 42848 55772 42900
rect 55824 42888 55830 42900
rect 57333 42891 57391 42897
rect 57333 42888 57345 42891
rect 55824 42860 57345 42888
rect 55824 42848 55830 42860
rect 57333 42857 57345 42860
rect 57379 42857 57391 42891
rect 57333 42851 57391 42857
rect 17034 42820 17040 42832
rect 16592 42792 17040 42820
rect 16255 42724 16344 42752
rect 16393 42755 16451 42761
rect 16255 42721 16267 42724
rect 16209 42715 16267 42721
rect 16393 42721 16405 42755
rect 16439 42752 16451 42755
rect 16592 42752 16620 42792
rect 17034 42780 17040 42792
rect 17092 42780 17098 42832
rect 25590 42820 25596 42832
rect 23492 42792 25596 42820
rect 18322 42752 18328 42764
rect 16439 42724 16620 42752
rect 16776 42724 18328 42752
rect 16439 42721 16451 42724
rect 16393 42715 16451 42721
rect 10686 42684 10692 42696
rect 10647 42656 10692 42684
rect 10686 42644 10692 42656
rect 10744 42644 10750 42696
rect 11698 42644 11704 42696
rect 11756 42684 11762 42696
rect 12253 42687 12311 42693
rect 12253 42684 12265 42687
rect 11756 42656 12265 42684
rect 11756 42644 11762 42656
rect 12253 42653 12265 42656
rect 12299 42653 12311 42687
rect 12253 42647 12311 42653
rect 12268 42616 12296 42647
rect 15010 42644 15016 42696
rect 15068 42684 15074 42696
rect 16776 42693 16804 42724
rect 18322 42712 18328 42724
rect 18380 42712 18386 42764
rect 23106 42712 23112 42764
rect 23164 42752 23170 42764
rect 23492 42752 23520 42792
rect 25590 42780 25596 42792
rect 25648 42780 25654 42832
rect 49326 42820 49332 42832
rect 45112 42792 45508 42820
rect 23937 42755 23995 42761
rect 23937 42752 23949 42755
rect 23164 42724 23520 42752
rect 23584 42724 23949 42752
rect 23164 42712 23170 42724
rect 15105 42687 15163 42693
rect 15105 42684 15117 42687
rect 15068 42656 15117 42684
rect 15068 42644 15074 42656
rect 15105 42653 15117 42656
rect 15151 42684 15163 42687
rect 15473 42687 15531 42693
rect 15473 42684 15485 42687
rect 15151 42656 15485 42684
rect 15151 42653 15163 42656
rect 15105 42647 15163 42653
rect 15473 42653 15485 42656
rect 15519 42653 15531 42687
rect 15473 42647 15531 42653
rect 16761 42687 16819 42693
rect 16761 42653 16773 42687
rect 16807 42653 16819 42687
rect 17034 42684 17040 42696
rect 16995 42656 17040 42684
rect 16761 42647 16819 42653
rect 17034 42644 17040 42656
rect 17092 42644 17098 42696
rect 17678 42684 17684 42696
rect 17639 42656 17684 42684
rect 17678 42644 17684 42656
rect 17736 42644 17742 42696
rect 17954 42684 17960 42696
rect 17915 42656 17960 42684
rect 17954 42644 17960 42656
rect 18012 42644 18018 42696
rect 19334 42684 19340 42696
rect 19295 42656 19340 42684
rect 19334 42644 19340 42656
rect 19392 42644 19398 42696
rect 23382 42684 23388 42696
rect 23308 42656 23388 42684
rect 17696 42616 17724 42644
rect 23308 42616 23336 42656
rect 23382 42644 23388 42656
rect 23440 42644 23446 42696
rect 23584 42616 23612 42724
rect 23937 42721 23949 42724
rect 23983 42752 23995 42755
rect 24489 42755 24547 42761
rect 24489 42752 24501 42755
rect 23983 42724 24501 42752
rect 23983 42721 23995 42724
rect 23937 42715 23995 42721
rect 24489 42721 24501 42724
rect 24535 42721 24547 42755
rect 24489 42715 24547 42721
rect 24673 42755 24731 42761
rect 24673 42721 24685 42755
rect 24719 42752 24731 42755
rect 24719 42724 24992 42752
rect 24719 42721 24731 42724
rect 24673 42715 24731 42721
rect 23661 42687 23719 42693
rect 23661 42653 23673 42687
rect 23707 42684 23719 42687
rect 23842 42684 23848 42696
rect 23707 42656 23848 42684
rect 23707 42653 23719 42656
rect 23661 42647 23719 42653
rect 23842 42644 23848 42656
rect 23900 42644 23906 42696
rect 12268 42588 17724 42616
rect 19444 42588 23336 42616
rect 23400 42588 23612 42616
rect 24964 42616 24992 42724
rect 25222 42712 25228 42764
rect 25280 42752 25286 42764
rect 28994 42752 29000 42764
rect 25280 42724 28856 42752
rect 28955 42724 29000 42752
rect 25280 42712 25286 42724
rect 25041 42687 25099 42693
rect 25041 42653 25053 42687
rect 25087 42684 25099 42687
rect 26970 42684 26976 42696
rect 25087 42656 26976 42684
rect 25087 42653 25099 42656
rect 25041 42647 25099 42653
rect 26970 42644 26976 42656
rect 27028 42644 27034 42696
rect 28445 42687 28503 42693
rect 28445 42653 28457 42687
rect 28491 42684 28503 42687
rect 28721 42687 28779 42693
rect 28721 42684 28733 42687
rect 28491 42656 28733 42684
rect 28491 42653 28503 42656
rect 28445 42647 28503 42653
rect 28721 42653 28733 42656
rect 28767 42653 28779 42687
rect 28828 42684 28856 42724
rect 28994 42712 29000 42724
rect 29052 42712 29058 42764
rect 29086 42712 29092 42764
rect 29144 42752 29150 42764
rect 32953 42755 33011 42761
rect 32953 42752 32965 42755
rect 29144 42724 32965 42752
rect 29144 42712 29150 42724
rect 32953 42721 32965 42724
rect 32999 42721 33011 42755
rect 32953 42715 33011 42721
rect 34333 42755 34391 42761
rect 34333 42721 34345 42755
rect 34379 42752 34391 42755
rect 35161 42755 35219 42761
rect 35161 42752 35173 42755
rect 34379 42724 35173 42752
rect 34379 42721 34391 42724
rect 34333 42715 34391 42721
rect 35161 42721 35173 42724
rect 35207 42752 35219 42755
rect 35434 42752 35440 42764
rect 35207 42724 35440 42752
rect 35207 42721 35219 42724
rect 35161 42715 35219 42721
rect 35434 42712 35440 42724
rect 35492 42712 35498 42764
rect 37461 42755 37519 42761
rect 37461 42721 37473 42755
rect 37507 42752 37519 42755
rect 37553 42755 37611 42761
rect 37553 42752 37565 42755
rect 37507 42724 37565 42752
rect 37507 42721 37519 42724
rect 37461 42715 37519 42721
rect 37553 42721 37565 42724
rect 37599 42721 37611 42755
rect 37553 42715 37611 42721
rect 43349 42755 43407 42761
rect 43349 42721 43361 42755
rect 43395 42752 43407 42755
rect 44082 42752 44088 42764
rect 43395 42724 44088 42752
rect 43395 42721 43407 42724
rect 43349 42715 43407 42721
rect 44082 42712 44088 42724
rect 44140 42712 44146 42764
rect 44358 42712 44364 42764
rect 44416 42752 44422 42764
rect 45112 42752 45140 42792
rect 45278 42752 45284 42764
rect 44416 42724 45140 42752
rect 45239 42724 45284 42752
rect 44416 42712 44422 42724
rect 45278 42712 45284 42724
rect 45336 42712 45342 42764
rect 45373 42755 45431 42761
rect 45373 42721 45385 42755
rect 45419 42721 45431 42755
rect 45480 42752 45508 42792
rect 48424 42792 49332 42820
rect 46750 42752 46756 42764
rect 45480 42724 46756 42752
rect 45373 42715 45431 42721
rect 30374 42684 30380 42696
rect 28828 42656 29684 42684
rect 30335 42656 30380 42684
rect 28721 42647 28779 42653
rect 25317 42619 25375 42625
rect 25317 42616 25329 42619
rect 24964 42588 25329 42616
rect 6914 42508 6920 42560
rect 6972 42548 6978 42560
rect 12158 42548 12164 42560
rect 6972 42520 12164 42548
rect 6972 42508 6978 42520
rect 12158 42508 12164 42520
rect 12216 42508 12222 42560
rect 12250 42508 12256 42560
rect 12308 42548 12314 42560
rect 12989 42551 13047 42557
rect 12989 42548 13001 42551
rect 12308 42520 13001 42548
rect 12308 42508 12314 42520
rect 12989 42517 13001 42520
rect 13035 42548 13047 42551
rect 17586 42548 17592 42560
rect 13035 42520 17592 42548
rect 13035 42517 13047 42520
rect 12989 42511 13047 42517
rect 17586 42508 17592 42520
rect 17644 42508 17650 42560
rect 19242 42508 19248 42560
rect 19300 42548 19306 42560
rect 19444 42557 19472 42588
rect 19429 42551 19487 42557
rect 19429 42548 19441 42551
rect 19300 42520 19441 42548
rect 19300 42508 19306 42520
rect 19429 42517 19441 42520
rect 19475 42517 19487 42551
rect 23290 42548 23296 42560
rect 23251 42520 23296 42548
rect 19429 42511 19487 42517
rect 23290 42508 23296 42520
rect 23348 42548 23354 42560
rect 23400 42557 23428 42588
rect 23385 42551 23443 42557
rect 23385 42548 23397 42551
rect 23348 42520 23397 42548
rect 23348 42508 23354 42520
rect 23385 42517 23397 42520
rect 23431 42517 23443 42551
rect 23385 42511 23443 42517
rect 23566 42508 23572 42560
rect 23624 42548 23630 42560
rect 24964 42548 24992 42588
rect 25317 42585 25329 42588
rect 25363 42616 25375 42619
rect 29656 42616 29684 42656
rect 30374 42644 30380 42656
rect 30432 42644 30438 42696
rect 32677 42687 32735 42693
rect 32677 42653 32689 42687
rect 32723 42684 32735 42687
rect 34146 42684 34152 42696
rect 32723 42656 34152 42684
rect 32723 42653 32735 42656
rect 32677 42647 32735 42653
rect 34146 42644 34152 42656
rect 34204 42684 34210 42696
rect 34422 42684 34428 42696
rect 34204 42656 34428 42684
rect 34204 42644 34210 42656
rect 34422 42644 34428 42656
rect 34480 42684 34486 42696
rect 34517 42687 34575 42693
rect 34517 42684 34529 42687
rect 34480 42656 34529 42684
rect 34480 42644 34486 42656
rect 34517 42653 34529 42656
rect 34563 42684 34575 42687
rect 39025 42687 39083 42693
rect 39025 42684 39037 42687
rect 34563 42656 39037 42684
rect 34563 42653 34575 42656
rect 34517 42647 34575 42653
rect 39025 42653 39037 42656
rect 39071 42653 39083 42687
rect 39025 42647 39083 42653
rect 39301 42687 39359 42693
rect 39301 42653 39313 42687
rect 39347 42684 39359 42687
rect 43438 42684 43444 42696
rect 39347 42656 43300 42684
rect 43399 42656 43444 42684
rect 39347 42653 39359 42656
rect 39301 42647 39359 42653
rect 35526 42616 35532 42628
rect 25363 42588 28672 42616
rect 29656 42588 32720 42616
rect 25363 42585 25375 42588
rect 25317 42579 25375 42585
rect 23624 42520 24992 42548
rect 23624 42508 23630 42520
rect 26510 42508 26516 42560
rect 26568 42548 26574 42560
rect 28445 42551 28503 42557
rect 28445 42548 28457 42551
rect 26568 42520 28457 42548
rect 26568 42508 26574 42520
rect 28445 42517 28457 42520
rect 28491 42548 28503 42551
rect 28537 42551 28595 42557
rect 28537 42548 28549 42551
rect 28491 42520 28549 42548
rect 28491 42517 28503 42520
rect 28445 42511 28503 42517
rect 28537 42517 28549 42520
rect 28583 42517 28595 42551
rect 28644 42548 28672 42588
rect 31570 42548 31576 42560
rect 28644 42520 31576 42548
rect 28537 42511 28595 42517
rect 31570 42508 31576 42520
rect 31628 42508 31634 42560
rect 32692 42548 32720 42588
rect 35268 42588 35532 42616
rect 35268 42557 35296 42588
rect 35526 42576 35532 42588
rect 35584 42576 35590 42628
rect 35253 42551 35311 42557
rect 35253 42548 35265 42551
rect 32692 42520 35265 42548
rect 35253 42517 35265 42520
rect 35299 42517 35311 42551
rect 35253 42511 35311 42517
rect 35342 42508 35348 42560
rect 35400 42548 35406 42560
rect 37277 42551 37335 42557
rect 37277 42548 37289 42551
rect 35400 42520 37289 42548
rect 35400 42508 35406 42520
rect 37277 42517 37289 42520
rect 37323 42517 37335 42551
rect 37277 42511 37335 42517
rect 37553 42551 37611 42557
rect 37553 42517 37565 42551
rect 37599 42548 37611 42551
rect 37826 42548 37832 42560
rect 37599 42520 37832 42548
rect 37599 42517 37611 42520
rect 37553 42511 37611 42517
rect 37826 42508 37832 42520
rect 37884 42508 37890 42560
rect 38933 42551 38991 42557
rect 38933 42517 38945 42551
rect 38979 42548 38991 42551
rect 39040 42548 39068 42647
rect 43272 42616 43300 42656
rect 43438 42644 43444 42656
rect 43496 42644 43502 42696
rect 43898 42644 43904 42696
rect 43956 42684 43962 42696
rect 45388 42684 45416 42715
rect 46750 42712 46756 42724
rect 46808 42712 46814 42764
rect 47489 42755 47547 42761
rect 47489 42721 47501 42755
rect 47535 42721 47547 42755
rect 47670 42752 47676 42764
rect 47631 42724 47676 42752
rect 47489 42715 47547 42721
rect 45830 42684 45836 42696
rect 43956 42656 45416 42684
rect 45791 42656 45836 42684
rect 43956 42644 43962 42656
rect 45830 42644 45836 42656
rect 45888 42644 45894 42696
rect 47504 42684 47532 42715
rect 47670 42712 47676 42724
rect 47728 42712 47734 42764
rect 48041 42755 48099 42761
rect 48041 42721 48053 42755
rect 48087 42752 48099 42755
rect 48424 42752 48452 42792
rect 49326 42780 49332 42792
rect 49384 42780 49390 42832
rect 57348 42792 57560 42820
rect 48087 42724 48452 42752
rect 48961 42755 49019 42761
rect 48087 42721 48099 42724
rect 48041 42715 48099 42721
rect 48961 42721 48973 42755
rect 49007 42721 49019 42755
rect 48961 42715 49019 42721
rect 48682 42684 48688 42696
rect 47504 42656 48688 42684
rect 48682 42644 48688 42656
rect 48740 42644 48746 42696
rect 48976 42684 49004 42715
rect 49050 42712 49056 42764
rect 49108 42752 49114 42764
rect 49237 42755 49295 42761
rect 49237 42752 49249 42755
rect 49108 42724 49249 42752
rect 49108 42712 49114 42724
rect 49237 42721 49249 42724
rect 49283 42752 49295 42755
rect 50525 42755 50583 42761
rect 49283 42724 49556 42752
rect 49283 42721 49295 42724
rect 49237 42715 49295 42721
rect 49326 42684 49332 42696
rect 48976 42656 49332 42684
rect 49326 42644 49332 42656
rect 49384 42644 49390 42696
rect 49528 42684 49556 42724
rect 50525 42721 50537 42755
rect 50571 42752 50583 42755
rect 50614 42752 50620 42764
rect 50571 42724 50620 42752
rect 50571 42721 50583 42724
rect 50525 42715 50583 42721
rect 50614 42712 50620 42724
rect 50672 42712 50678 42764
rect 50709 42755 50767 42761
rect 50709 42721 50721 42755
rect 50755 42721 50767 42755
rect 50709 42715 50767 42721
rect 54772 42724 55352 42752
rect 50724 42684 50752 42715
rect 49528 42656 50752 42684
rect 53742 42644 53748 42696
rect 53800 42684 53806 42696
rect 54772 42693 54800 42724
rect 54757 42687 54815 42693
rect 54757 42684 54769 42687
rect 53800 42656 54769 42684
rect 53800 42644 53806 42656
rect 54757 42653 54769 42656
rect 54803 42653 54815 42687
rect 54757 42647 54815 42653
rect 55033 42687 55091 42693
rect 55033 42653 55045 42687
rect 55079 42684 55091 42687
rect 55214 42684 55220 42696
rect 55079 42656 55220 42684
rect 55079 42653 55091 42656
rect 55033 42647 55091 42653
rect 55214 42644 55220 42656
rect 55272 42644 55278 42696
rect 55324 42684 55352 42724
rect 56226 42712 56232 42764
rect 56284 42752 56290 42764
rect 57348 42752 57376 42792
rect 56284 42724 57376 42752
rect 57425 42755 57483 42761
rect 56284 42712 56290 42724
rect 57425 42721 57437 42755
rect 57471 42721 57483 42755
rect 57532 42752 57560 42792
rect 57793 42755 57851 42761
rect 57793 42752 57805 42755
rect 57532 42724 57805 42752
rect 57425 42715 57483 42721
rect 57793 42721 57805 42724
rect 57839 42721 57851 42755
rect 57793 42715 57851 42721
rect 56505 42687 56563 42693
rect 56505 42684 56517 42687
rect 55324 42656 56517 42684
rect 56505 42653 56517 42656
rect 56551 42653 56563 42687
rect 57440 42684 57468 42715
rect 57882 42712 57888 42764
rect 57940 42752 57946 42764
rect 58069 42755 58127 42761
rect 58069 42752 58081 42755
rect 57940 42724 58081 42752
rect 57940 42712 57946 42724
rect 58069 42721 58081 42724
rect 58115 42721 58127 42755
rect 58069 42715 58127 42721
rect 60277 42755 60335 42761
rect 60277 42721 60289 42755
rect 60323 42752 60335 42755
rect 60826 42752 60832 42764
rect 60323 42724 60832 42752
rect 60323 42721 60335 42724
rect 60277 42715 60335 42721
rect 60826 42712 60832 42724
rect 60884 42712 60890 42764
rect 61565 42755 61623 42761
rect 61565 42721 61577 42755
rect 61611 42752 61623 42755
rect 62206 42752 62212 42764
rect 61611 42724 62212 42752
rect 61611 42721 61623 42724
rect 61565 42715 61623 42721
rect 62206 42712 62212 42724
rect 62264 42712 62270 42764
rect 63494 42712 63500 42764
rect 63552 42752 63558 42764
rect 64598 42752 64604 42764
rect 63552 42724 64604 42752
rect 63552 42712 63558 42724
rect 64598 42712 64604 42724
rect 64656 42752 64662 42764
rect 69017 42755 69075 42761
rect 69017 42752 69029 42755
rect 64656 42724 69029 42752
rect 64656 42712 64662 42724
rect 69017 42721 69029 42724
rect 69063 42721 69075 42755
rect 69198 42752 69204 42764
rect 69159 42724 69204 42752
rect 69017 42715 69075 42721
rect 58526 42684 58532 42696
rect 57440 42656 58532 42684
rect 56505 42647 56563 42653
rect 58526 42644 58532 42656
rect 58584 42644 58590 42696
rect 61102 42644 61108 42696
rect 61160 42684 61166 42696
rect 61289 42687 61347 42693
rect 61289 42684 61301 42687
rect 61160 42656 61301 42684
rect 61160 42644 61166 42656
rect 61289 42653 61301 42656
rect 61335 42684 61347 42687
rect 63129 42687 63187 42693
rect 63129 42684 63141 42687
rect 61335 42656 63141 42684
rect 61335 42653 61347 42656
rect 61289 42647 61347 42653
rect 63129 42653 63141 42656
rect 63175 42684 63187 42687
rect 65797 42687 65855 42693
rect 65797 42684 65809 42687
rect 63175 42656 65809 42684
rect 63175 42653 63187 42656
rect 63129 42647 63187 42653
rect 65797 42653 65809 42656
rect 65843 42653 65855 42687
rect 66070 42684 66076 42696
rect 66031 42656 66076 42684
rect 65797 42647 65855 42653
rect 45462 42616 45468 42628
rect 43272 42588 45468 42616
rect 45462 42576 45468 42588
rect 45520 42576 45526 42628
rect 49053 42619 49111 42625
rect 49053 42585 49065 42619
rect 49099 42616 49111 42619
rect 49142 42616 49148 42628
rect 49099 42588 49148 42616
rect 49099 42585 49111 42588
rect 49053 42579 49111 42585
rect 49142 42576 49148 42588
rect 49200 42576 49206 42628
rect 59446 42616 59452 42628
rect 55692 42588 59452 42616
rect 44542 42548 44548 42560
rect 38979 42520 44548 42548
rect 38979 42517 38991 42520
rect 38933 42511 38991 42517
rect 44542 42508 44548 42520
rect 44600 42508 44606 42560
rect 45097 42551 45155 42557
rect 45097 42517 45109 42551
rect 45143 42548 45155 42551
rect 46017 42551 46075 42557
rect 46017 42548 46029 42551
rect 45143 42520 46029 42548
rect 45143 42517 45155 42520
rect 45097 42511 45155 42517
rect 46017 42517 46029 42520
rect 46063 42548 46075 42551
rect 49970 42548 49976 42560
rect 46063 42520 49976 42548
rect 46063 42517 46075 42520
rect 46017 42511 46075 42517
rect 49970 42508 49976 42520
rect 50028 42508 50034 42560
rect 51074 42508 51080 42560
rect 51132 42548 51138 42560
rect 55692 42548 55720 42588
rect 59446 42576 59452 42588
rect 59504 42576 59510 42628
rect 51132 42520 55720 42548
rect 51132 42508 51138 42520
rect 55950 42508 55956 42560
rect 56008 42548 56014 42560
rect 56137 42551 56195 42557
rect 56137 42548 56149 42551
rect 56008 42520 56149 42548
rect 56008 42508 56014 42520
rect 56137 42517 56149 42520
rect 56183 42517 56195 42551
rect 58526 42548 58532 42560
rect 58487 42520 58532 42548
rect 56137 42511 56195 42517
rect 58526 42508 58532 42520
rect 58584 42508 58590 42560
rect 60366 42548 60372 42560
rect 60327 42520 60372 42548
rect 60366 42508 60372 42520
rect 60424 42508 60430 42560
rect 60826 42508 60832 42560
rect 60884 42548 60890 42560
rect 62669 42551 62727 42557
rect 62669 42548 62681 42551
rect 60884 42520 62681 42548
rect 60884 42508 60890 42520
rect 62669 42517 62681 42520
rect 62715 42517 62727 42551
rect 65812 42548 65840 42647
rect 66070 42644 66076 42656
rect 66128 42644 66134 42696
rect 69032 42684 69060 42715
rect 69198 42712 69204 42724
rect 69256 42712 69262 42764
rect 69290 42712 69296 42764
rect 69348 42752 69354 42764
rect 71406 42752 71412 42764
rect 69348 42724 69393 42752
rect 71367 42724 71412 42752
rect 69348 42712 69354 42724
rect 71406 42712 71412 42724
rect 71464 42712 71470 42764
rect 69845 42687 69903 42693
rect 69845 42684 69857 42687
rect 69032 42656 69857 42684
rect 69845 42653 69857 42656
rect 69891 42684 69903 42687
rect 70394 42684 70400 42696
rect 69891 42656 70400 42684
rect 69891 42653 69903 42656
rect 69845 42647 69903 42653
rect 70394 42644 70400 42656
rect 70452 42644 70458 42696
rect 66806 42576 66812 42628
rect 66864 42616 66870 42628
rect 67637 42619 67695 42625
rect 67637 42616 67649 42619
rect 66864 42588 67649 42616
rect 66864 42576 66870 42588
rect 67637 42585 67649 42588
rect 67683 42616 67695 42619
rect 69658 42616 69664 42628
rect 67683 42588 69664 42616
rect 67683 42585 67695 42588
rect 67637 42579 67695 42585
rect 69658 42576 69664 42588
rect 69716 42576 69722 42628
rect 66824 42548 66852 42576
rect 65812 42520 66852 42548
rect 62669 42511 62727 42517
rect 66990 42508 66996 42560
rect 67048 42548 67054 42560
rect 67177 42551 67235 42557
rect 67177 42548 67189 42551
rect 67048 42520 67189 42548
rect 67048 42508 67054 42520
rect 67177 42517 67189 42520
rect 67223 42517 67235 42551
rect 67177 42511 67235 42517
rect 69382 42508 69388 42560
rect 69440 42548 69446 42560
rect 69477 42551 69535 42557
rect 69477 42548 69489 42551
rect 69440 42520 69489 42548
rect 69440 42508 69446 42520
rect 69477 42517 69489 42520
rect 69523 42517 69535 42551
rect 69477 42511 69535 42517
rect 70026 42508 70032 42560
rect 70084 42548 70090 42560
rect 71501 42551 71559 42557
rect 71501 42548 71513 42551
rect 70084 42520 71513 42548
rect 70084 42508 70090 42520
rect 71501 42517 71513 42520
rect 71547 42517 71559 42551
rect 71501 42511 71559 42517
rect 1104 42458 111136 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 65686 42458
rect 65738 42406 65750 42458
rect 65802 42406 65814 42458
rect 65866 42406 65878 42458
rect 65930 42406 96406 42458
rect 96458 42406 96470 42458
rect 96522 42406 96534 42458
rect 96586 42406 96598 42458
rect 96650 42406 111136 42458
rect 1104 42384 111136 42406
rect 2406 42344 2412 42356
rect 2367 42316 2412 42344
rect 2406 42304 2412 42316
rect 2464 42304 2470 42356
rect 4433 42347 4491 42353
rect 4433 42313 4445 42347
rect 4479 42344 4491 42347
rect 4798 42344 4804 42356
rect 4479 42316 4804 42344
rect 4479 42313 4491 42316
rect 4433 42307 4491 42313
rect 2593 42211 2651 42217
rect 2593 42177 2605 42211
rect 2639 42208 2651 42211
rect 4448 42208 4476 42307
rect 4798 42304 4804 42316
rect 4856 42304 4862 42356
rect 10060 42316 10916 42344
rect 6270 42236 6276 42288
rect 6328 42276 6334 42288
rect 9950 42276 9956 42288
rect 6328 42248 9956 42276
rect 6328 42236 6334 42248
rect 9950 42236 9956 42248
rect 10008 42236 10014 42288
rect 2639 42180 4476 42208
rect 2639 42177 2651 42180
rect 2593 42171 2651 42177
rect 6086 42168 6092 42220
rect 6144 42208 6150 42220
rect 10060 42208 10088 42316
rect 10778 42276 10784 42288
rect 10739 42248 10784 42276
rect 10778 42236 10784 42248
rect 10836 42236 10842 42288
rect 6144 42180 10088 42208
rect 10888 42208 10916 42316
rect 12526 42304 12532 42356
rect 12584 42344 12590 42356
rect 12584 42316 16988 42344
rect 12584 42304 12590 42316
rect 16960 42276 16988 42316
rect 18414 42304 18420 42356
rect 18472 42344 18478 42356
rect 23109 42347 23167 42353
rect 23109 42344 23121 42347
rect 18472 42316 23121 42344
rect 18472 42304 18478 42316
rect 23109 42313 23121 42316
rect 23155 42344 23167 42347
rect 23290 42344 23296 42356
rect 23155 42316 23296 42344
rect 23155 42313 23167 42316
rect 23109 42307 23167 42313
rect 23290 42304 23296 42316
rect 23348 42304 23354 42356
rect 23658 42304 23664 42356
rect 23716 42344 23722 42356
rect 24578 42344 24584 42356
rect 23716 42316 24584 42344
rect 23716 42304 23722 42316
rect 24578 42304 24584 42316
rect 24636 42304 24642 42356
rect 25406 42304 25412 42356
rect 25464 42344 25470 42356
rect 51074 42344 51080 42356
rect 25464 42316 51080 42344
rect 25464 42304 25470 42316
rect 51074 42304 51080 42316
rect 51132 42304 51138 42356
rect 63034 42344 63040 42356
rect 51184 42316 52776 42344
rect 62995 42316 63040 42344
rect 22925 42279 22983 42285
rect 22925 42276 22937 42279
rect 16960 42248 22937 42276
rect 22925 42245 22937 42248
rect 22971 42276 22983 42279
rect 23474 42276 23480 42288
rect 22971 42248 23480 42276
rect 22971 42245 22983 42248
rect 22925 42239 22983 42245
rect 23474 42236 23480 42248
rect 23532 42276 23538 42288
rect 23532 42248 23704 42276
rect 23532 42236 23538 42248
rect 10888 42180 13584 42208
rect 6144 42168 6150 42180
rect 2406 42100 2412 42152
rect 2464 42140 2470 42152
rect 2866 42140 2872 42152
rect 2464 42112 2872 42140
rect 2464 42100 2470 42112
rect 2866 42100 2872 42112
rect 2924 42100 2930 42152
rect 5258 42140 5264 42152
rect 5219 42112 5264 42140
rect 5258 42100 5264 42112
rect 5316 42100 5322 42152
rect 9677 42143 9735 42149
rect 9677 42109 9689 42143
rect 9723 42109 9735 42143
rect 9677 42103 9735 42109
rect 9846 42143 9904 42149
rect 9846 42109 9858 42143
rect 9892 42140 9904 42143
rect 10410 42140 10416 42152
rect 9892 42112 10416 42140
rect 9892 42109 9904 42112
rect 9846 42103 9904 42109
rect 8018 42032 8024 42084
rect 8076 42072 8082 42084
rect 9582 42072 9588 42084
rect 8076 42044 9588 42072
rect 8076 42032 8082 42044
rect 9582 42032 9588 42044
rect 9640 42032 9646 42084
rect 3970 42004 3976 42016
rect 3931 41976 3976 42004
rect 3970 41964 3976 41976
rect 4028 41964 4034 42016
rect 5166 41964 5172 42016
rect 5224 42004 5230 42016
rect 5353 42007 5411 42013
rect 5353 42004 5365 42007
rect 5224 41976 5365 42004
rect 5224 41964 5230 41976
rect 5353 41973 5365 41976
rect 5399 41973 5411 42007
rect 9490 42004 9496 42016
rect 9451 41976 9496 42004
rect 5353 41967 5411 41973
rect 9490 41964 9496 41976
rect 9548 42004 9554 42016
rect 9692 42004 9720 42103
rect 10410 42100 10416 42112
rect 10468 42100 10474 42152
rect 10588 42143 10646 42149
rect 10588 42140 10600 42143
rect 10520 42112 10600 42140
rect 9548 41976 9720 42004
rect 9548 41964 9554 41976
rect 10226 41964 10232 42016
rect 10284 42004 10290 42016
rect 10520 42004 10548 42112
rect 10588 42109 10600 42112
rect 10634 42109 10646 42143
rect 10588 42103 10646 42109
rect 12429 42143 12487 42149
rect 12429 42109 12441 42143
rect 12475 42140 12487 42143
rect 12618 42140 12624 42152
rect 12475 42112 12624 42140
rect 12475 42109 12487 42112
rect 12429 42103 12487 42109
rect 12618 42100 12624 42112
rect 12676 42100 12682 42152
rect 13556 42140 13584 42180
rect 13630 42168 13636 42220
rect 13688 42208 13694 42220
rect 15749 42211 15807 42217
rect 15749 42208 15761 42211
rect 13688 42180 15761 42208
rect 13688 42168 13694 42180
rect 15749 42177 15761 42180
rect 15795 42208 15807 42211
rect 16850 42208 16856 42220
rect 15795 42180 16856 42208
rect 15795 42177 15807 42180
rect 15749 42171 15807 42177
rect 16850 42168 16856 42180
rect 16908 42208 16914 42220
rect 17218 42208 17224 42220
rect 16908 42180 16988 42208
rect 16908 42168 16914 42180
rect 16390 42140 16396 42152
rect 13556 42112 16068 42140
rect 16351 42112 16396 42140
rect 15286 42032 15292 42084
rect 15344 42072 15350 42084
rect 15933 42075 15991 42081
rect 15933 42072 15945 42075
rect 15344 42044 15945 42072
rect 15344 42032 15350 42044
rect 15933 42041 15945 42044
rect 15979 42041 15991 42075
rect 16040 42072 16068 42112
rect 16390 42100 16396 42112
rect 16448 42100 16454 42152
rect 16574 42140 16580 42152
rect 16535 42112 16580 42140
rect 16574 42100 16580 42112
rect 16632 42100 16638 42152
rect 16960 42149 16988 42180
rect 17052 42180 17224 42208
rect 17052 42149 17080 42180
rect 17218 42168 17224 42180
rect 17276 42168 17282 42220
rect 17494 42208 17500 42220
rect 17407 42180 17500 42208
rect 17494 42168 17500 42180
rect 17552 42208 17558 42220
rect 18322 42208 18328 42220
rect 17552 42180 18328 42208
rect 17552 42168 17558 42180
rect 18322 42168 18328 42180
rect 18380 42168 18386 42220
rect 18785 42211 18843 42217
rect 18785 42177 18797 42211
rect 18831 42208 18843 42211
rect 19429 42211 19487 42217
rect 19429 42208 19441 42211
rect 18831 42180 19196 42208
rect 18831 42177 18843 42180
rect 18785 42171 18843 42177
rect 16945 42143 17003 42149
rect 16945 42109 16957 42143
rect 16991 42109 17003 42143
rect 16945 42103 17003 42109
rect 17037 42143 17095 42149
rect 17037 42109 17049 42143
rect 17083 42109 17095 42143
rect 17037 42103 17095 42109
rect 17678 42100 17684 42152
rect 17736 42140 17742 42152
rect 18693 42143 18751 42149
rect 18693 42140 18705 42143
rect 17736 42112 18705 42140
rect 17736 42100 17742 42112
rect 18693 42109 18705 42112
rect 18739 42109 18751 42143
rect 18693 42103 18751 42109
rect 19061 42143 19119 42149
rect 19061 42109 19073 42143
rect 19107 42109 19119 42143
rect 19061 42103 19119 42109
rect 18049 42075 18107 42081
rect 18049 42072 18061 42075
rect 16040 42044 18061 42072
rect 15933 42035 15991 42041
rect 18049 42041 18061 42044
rect 18095 42041 18107 42075
rect 18049 42035 18107 42041
rect 11241 42007 11299 42013
rect 11241 42004 11253 42007
rect 10284 41976 11253 42004
rect 10284 41964 10290 41976
rect 11241 41973 11253 41976
rect 11287 42004 11299 42007
rect 12526 42004 12532 42016
rect 11287 41976 12532 42004
rect 11287 41973 11299 41976
rect 11241 41967 11299 41973
rect 12526 41964 12532 41976
rect 12584 41964 12590 42016
rect 15194 41964 15200 42016
rect 15252 42004 15258 42016
rect 15565 42007 15623 42013
rect 15565 42004 15577 42007
rect 15252 41976 15577 42004
rect 15252 41964 15258 41976
rect 15565 41973 15577 41976
rect 15611 42004 15623 42007
rect 16574 42004 16580 42016
rect 15611 41976 16580 42004
rect 15611 41973 15623 41976
rect 15565 41967 15623 41973
rect 16574 41964 16580 41976
rect 16632 42004 16638 42016
rect 17586 42004 17592 42016
rect 16632 41976 17592 42004
rect 16632 41964 16638 41976
rect 17586 41964 17592 41976
rect 17644 41964 17650 42016
rect 17770 42004 17776 42016
rect 17731 41976 17776 42004
rect 17770 41964 17776 41976
rect 17828 42004 17834 42016
rect 19076 42004 19104 42103
rect 17828 41976 19104 42004
rect 19168 42004 19196 42180
rect 19260 42180 19441 42208
rect 19260 42149 19288 42180
rect 19429 42177 19441 42180
rect 19475 42208 19487 42211
rect 23566 42208 23572 42220
rect 19475 42180 23572 42208
rect 19475 42177 19487 42180
rect 19429 42171 19487 42177
rect 23566 42168 23572 42180
rect 23624 42168 23630 42220
rect 23676 42217 23704 42248
rect 23934 42236 23940 42288
rect 23992 42276 23998 42288
rect 29457 42279 29515 42285
rect 29457 42276 29469 42279
rect 23992 42248 29469 42276
rect 23992 42236 23998 42248
rect 29457 42245 29469 42248
rect 29503 42276 29515 42279
rect 29641 42279 29699 42285
rect 29641 42276 29653 42279
rect 29503 42248 29653 42276
rect 29503 42245 29515 42248
rect 29457 42239 29515 42245
rect 29641 42245 29653 42248
rect 29687 42276 29699 42279
rect 44082 42276 44088 42288
rect 29687 42248 29868 42276
rect 29687 42245 29699 42248
rect 29641 42239 29699 42245
rect 23661 42211 23719 42217
rect 23661 42177 23673 42211
rect 23707 42177 23719 42211
rect 23661 42171 23719 42177
rect 24949 42211 25007 42217
rect 24949 42177 24961 42211
rect 24995 42208 25007 42211
rect 25866 42208 25872 42220
rect 24995 42180 25872 42208
rect 24995 42177 25007 42180
rect 24949 42171 25007 42177
rect 25866 42168 25872 42180
rect 25924 42168 25930 42220
rect 29840 42217 29868 42248
rect 31496 42248 37596 42276
rect 44043 42248 44088 42276
rect 29825 42211 29883 42217
rect 25976 42180 26280 42208
rect 19245 42143 19303 42149
rect 19245 42109 19257 42143
rect 19291 42109 19303 42143
rect 19245 42103 19303 42109
rect 19334 42100 19340 42152
rect 19392 42140 19398 42152
rect 20073 42143 20131 42149
rect 20073 42140 20085 42143
rect 19392 42112 20085 42140
rect 19392 42100 19398 42112
rect 20073 42109 20085 42112
rect 20119 42109 20131 42143
rect 20073 42103 20131 42109
rect 23290 42100 23296 42152
rect 23348 42140 23354 42152
rect 23845 42143 23903 42149
rect 23845 42140 23857 42143
rect 23348 42112 23857 42140
rect 23348 42100 23354 42112
rect 23845 42109 23857 42112
rect 23891 42140 23903 42143
rect 24397 42143 24455 42149
rect 24397 42140 24409 42143
rect 23891 42112 24409 42140
rect 23891 42109 23903 42112
rect 23845 42103 23903 42109
rect 24397 42109 24409 42112
rect 24443 42109 24455 42143
rect 24578 42140 24584 42152
rect 24491 42112 24584 42140
rect 24397 42103 24455 42109
rect 24578 42100 24584 42112
rect 24636 42140 24642 42152
rect 25682 42140 25688 42152
rect 24636 42112 25688 42140
rect 24636 42100 24642 42112
rect 25682 42100 25688 42112
rect 25740 42100 25746 42152
rect 25976 42149 26004 42180
rect 25961 42143 26019 42149
rect 25961 42109 25973 42143
rect 26007 42109 26019 42143
rect 25961 42103 26019 42109
rect 26145 42143 26203 42149
rect 26145 42109 26157 42143
rect 26191 42109 26203 42143
rect 26252 42140 26280 42180
rect 29825 42177 29837 42211
rect 29871 42208 29883 42211
rect 29871 42180 30144 42208
rect 29871 42177 29883 42180
rect 29825 42171 29883 42177
rect 26605 42143 26663 42149
rect 26605 42140 26617 42143
rect 26252 42112 26617 42140
rect 26145 42103 26203 42109
rect 26605 42109 26617 42112
rect 26651 42109 26663 42143
rect 26605 42103 26663 42109
rect 26697 42143 26755 42149
rect 26697 42109 26709 42143
rect 26743 42140 26755 42143
rect 27433 42143 27491 42149
rect 27433 42140 27445 42143
rect 26743 42112 27445 42140
rect 26743 42109 26755 42112
rect 26697 42103 26755 42109
rect 27433 42109 27445 42112
rect 27479 42140 27491 42143
rect 27617 42143 27675 42149
rect 27617 42140 27629 42143
rect 27479 42112 27629 42140
rect 27479 42109 27491 42112
rect 27433 42103 27491 42109
rect 27617 42109 27629 42112
rect 27663 42140 27675 42143
rect 30009 42143 30067 42149
rect 30009 42140 30021 42143
rect 27663 42112 30021 42140
rect 27663 42109 27675 42112
rect 27617 42103 27675 42109
rect 30009 42109 30021 42112
rect 30055 42109 30067 42143
rect 30116 42140 30144 42180
rect 31496 42149 31524 42248
rect 31570 42168 31576 42220
rect 31628 42208 31634 42220
rect 36265 42211 36323 42217
rect 36265 42208 36277 42211
rect 31628 42180 36277 42208
rect 31628 42168 31634 42180
rect 36265 42177 36277 42180
rect 36311 42208 36323 42211
rect 37568 42208 37596 42248
rect 44082 42236 44088 42248
rect 44140 42236 44146 42288
rect 45094 42276 45100 42288
rect 44652 42248 45100 42276
rect 44652 42208 44680 42248
rect 45094 42236 45100 42248
rect 45152 42236 45158 42288
rect 45296 42248 48820 42276
rect 45296 42217 45324 42248
rect 36311 42180 36860 42208
rect 37568 42180 44680 42208
rect 44729 42211 44787 42217
rect 36311 42177 36323 42180
rect 36265 42171 36323 42177
rect 30469 42143 30527 42149
rect 30469 42140 30481 42143
rect 30116 42112 30481 42140
rect 30009 42103 30067 42109
rect 30469 42109 30481 42112
rect 30515 42109 30527 42143
rect 30469 42103 30527 42109
rect 30561 42143 30619 42149
rect 30561 42109 30573 42143
rect 30607 42140 30619 42143
rect 31297 42143 31355 42149
rect 31297 42140 31309 42143
rect 30607 42112 31309 42140
rect 30607 42109 30619 42112
rect 30561 42103 30619 42109
rect 31297 42109 31309 42112
rect 31343 42140 31355 42143
rect 31481 42143 31539 42149
rect 31481 42140 31493 42143
rect 31343 42112 31493 42140
rect 31343 42109 31355 42112
rect 31297 42103 31355 42109
rect 31481 42109 31493 42112
rect 31527 42109 31539 42143
rect 31481 42103 31539 42109
rect 20165 42075 20223 42081
rect 20165 42041 20177 42075
rect 20211 42072 20223 42075
rect 20254 42072 20260 42084
rect 20211 42044 20260 42072
rect 20211 42041 20223 42044
rect 20165 42035 20223 42041
rect 20254 42032 20260 42044
rect 20312 42072 20318 42084
rect 23750 42072 23756 42084
rect 20312 42044 23756 42072
rect 20312 42032 20318 42044
rect 23750 42032 23756 42044
rect 23808 42032 23814 42084
rect 25593 42075 25651 42081
rect 25593 42072 25605 42075
rect 25148 42044 25605 42072
rect 19613 42007 19671 42013
rect 19613 42004 19625 42007
rect 19168 41976 19625 42004
rect 17828 41964 17834 41976
rect 19613 41973 19625 41976
rect 19659 42004 19671 42007
rect 23106 42004 23112 42016
rect 19659 41976 23112 42004
rect 19659 41973 19671 41976
rect 19613 41967 19671 41973
rect 23106 41964 23112 41976
rect 23164 41964 23170 42016
rect 23566 41964 23572 42016
rect 23624 42004 23630 42016
rect 25148 42004 25176 42044
rect 25593 42041 25605 42044
rect 25639 42072 25651 42075
rect 25777 42075 25835 42081
rect 25777 42072 25789 42075
rect 25639 42044 25789 42072
rect 25639 42041 25651 42044
rect 25593 42035 25651 42041
rect 25777 42041 25789 42044
rect 25823 42072 25835 42075
rect 25976 42072 26004 42103
rect 25823 42044 26004 42072
rect 26160 42072 26188 42103
rect 26712 42072 26740 42103
rect 27246 42072 27252 42084
rect 26160 42044 26740 42072
rect 27207 42044 27252 42072
rect 25823 42041 25835 42044
rect 25777 42035 25835 42041
rect 27246 42032 27252 42044
rect 27304 42032 27310 42084
rect 30024 42072 30052 42103
rect 30576 42072 30604 42103
rect 34790 42100 34796 42152
rect 34848 42140 34854 42152
rect 34885 42143 34943 42149
rect 34885 42140 34897 42143
rect 34848 42112 34897 42140
rect 34848 42100 34854 42112
rect 34885 42109 34897 42112
rect 34931 42109 34943 42143
rect 34885 42103 34943 42109
rect 36449 42143 36507 42149
rect 36449 42109 36461 42143
rect 36495 42109 36507 42143
rect 36449 42103 36507 42109
rect 36633 42143 36691 42149
rect 36633 42109 36645 42143
rect 36679 42140 36691 42143
rect 36722 42140 36728 42152
rect 36679 42112 36728 42140
rect 36679 42109 36691 42112
rect 36633 42103 36691 42109
rect 30024 42044 30604 42072
rect 31113 42075 31171 42081
rect 31113 42041 31125 42075
rect 31159 42072 31171 42075
rect 32582 42072 32588 42084
rect 31159 42044 32588 42072
rect 31159 42041 31171 42044
rect 31113 42035 31171 42041
rect 32582 42032 32588 42044
rect 32640 42032 32646 42084
rect 35894 42032 35900 42084
rect 35952 42072 35958 42084
rect 36081 42075 36139 42081
rect 36081 42072 36093 42075
rect 35952 42044 36093 42072
rect 35952 42032 35958 42044
rect 36081 42041 36093 42044
rect 36127 42072 36139 42075
rect 36464 42072 36492 42103
rect 36722 42100 36728 42112
rect 36780 42100 36786 42152
rect 36832 42140 36860 42180
rect 44729 42177 44741 42211
rect 44775 42208 44787 42211
rect 45281 42211 45339 42217
rect 45281 42208 45293 42211
rect 44775 42180 45293 42208
rect 44775 42177 44787 42180
rect 44729 42171 44787 42177
rect 45281 42177 45293 42180
rect 45327 42177 45339 42211
rect 48038 42208 48044 42220
rect 47999 42180 48044 42208
rect 45281 42171 45339 42177
rect 48038 42168 48044 42180
rect 48096 42168 48102 42220
rect 37093 42143 37151 42149
rect 37093 42140 37105 42143
rect 36832 42112 37105 42140
rect 37093 42109 37105 42112
rect 37139 42109 37151 42143
rect 37093 42103 37151 42109
rect 37185 42143 37243 42149
rect 37185 42109 37197 42143
rect 37231 42140 37243 42143
rect 37274 42140 37280 42152
rect 37231 42112 37280 42140
rect 37231 42109 37243 42112
rect 37185 42103 37243 42109
rect 37274 42100 37280 42112
rect 37332 42100 37338 42152
rect 39758 42140 39764 42152
rect 37384 42112 39764 42140
rect 37384 42072 37412 42112
rect 39758 42100 39764 42112
rect 39816 42100 39822 42152
rect 44358 42140 44364 42152
rect 43548 42112 44364 42140
rect 37734 42072 37740 42084
rect 36127 42044 36492 42072
rect 36832 42044 37412 42072
rect 37695 42044 37740 42072
rect 36127 42041 36139 42044
rect 36081 42035 36139 42041
rect 23624 41976 25176 42004
rect 25225 42007 25283 42013
rect 23624 41964 23630 41976
rect 25225 41973 25237 42007
rect 25271 42004 25283 42007
rect 25682 42004 25688 42016
rect 25271 41976 25688 42004
rect 25271 41973 25283 41976
rect 25225 41967 25283 41973
rect 25682 41964 25688 41976
rect 25740 41964 25746 42016
rect 25866 41964 25872 42016
rect 25924 42004 25930 42016
rect 30466 42004 30472 42016
rect 25924 41976 30472 42004
rect 25924 41964 25930 41976
rect 30466 41964 30472 41976
rect 30524 41964 30530 42016
rect 30558 41964 30564 42016
rect 30616 42004 30622 42016
rect 34977 42007 35035 42013
rect 34977 42004 34989 42007
rect 30616 41976 34989 42004
rect 30616 41964 30622 41976
rect 34977 41973 34989 41976
rect 35023 42004 35035 42007
rect 36832 42004 36860 42044
rect 37734 42032 37740 42044
rect 37792 42032 37798 42084
rect 37826 42032 37832 42084
rect 37884 42072 37890 42084
rect 43548 42072 43576 42112
rect 44358 42100 44364 42112
rect 44416 42100 44422 42152
rect 44450 42100 44456 42152
rect 44508 42140 44514 42152
rect 44637 42143 44695 42149
rect 44637 42140 44649 42143
rect 44508 42112 44649 42140
rect 44508 42100 44514 42112
rect 44637 42109 44649 42112
rect 44683 42109 44695 42143
rect 44637 42103 44695 42109
rect 44818 42100 44824 42152
rect 44876 42140 44882 42152
rect 45005 42143 45063 42149
rect 45005 42140 45017 42143
rect 44876 42112 45017 42140
rect 44876 42100 44882 42112
rect 45005 42109 45017 42112
rect 45051 42109 45063 42143
rect 45005 42103 45063 42109
rect 45097 42143 45155 42149
rect 45097 42109 45109 42143
rect 45143 42109 45155 42143
rect 45097 42103 45155 42109
rect 37884 42044 43576 42072
rect 43640 42044 43944 42072
rect 37884 42032 37890 42044
rect 35023 41976 36860 42004
rect 35023 41973 35035 41976
rect 34977 41967 35035 41973
rect 36906 41964 36912 42016
rect 36964 42004 36970 42016
rect 38013 42007 38071 42013
rect 38013 42004 38025 42007
rect 36964 41976 38025 42004
rect 36964 41964 36970 41976
rect 38013 41973 38025 41976
rect 38059 42004 38071 42007
rect 38930 42004 38936 42016
rect 38059 41976 38936 42004
rect 38059 41973 38071 41976
rect 38013 41967 38071 41973
rect 38930 41964 38936 41976
rect 38988 42004 38994 42016
rect 43640 42004 43668 42044
rect 43806 42004 43812 42016
rect 38988 41976 43668 42004
rect 43767 41976 43812 42004
rect 38988 41964 38994 41976
rect 43806 41964 43812 41976
rect 43864 41964 43870 42016
rect 43916 42004 43944 42044
rect 44910 42032 44916 42084
rect 44968 42072 44974 42084
rect 45112 42072 45140 42103
rect 45462 42100 45468 42152
rect 45520 42140 45526 42152
rect 46109 42143 46167 42149
rect 46109 42140 46121 42143
rect 45520 42112 46121 42140
rect 45520 42100 45526 42112
rect 46109 42109 46121 42112
rect 46155 42109 46167 42143
rect 48682 42140 48688 42152
rect 48643 42112 48688 42140
rect 46109 42103 46167 42109
rect 48682 42100 48688 42112
rect 48740 42100 48746 42152
rect 48792 42149 48820 42248
rect 49142 42236 49148 42288
rect 49200 42276 49206 42288
rect 51184 42276 51212 42316
rect 49200 42248 51212 42276
rect 52748 42276 52776 42316
rect 63034 42304 63040 42316
rect 63092 42304 63098 42356
rect 69290 42344 69296 42356
rect 69251 42316 69296 42344
rect 69290 42304 69296 42316
rect 69348 42304 69354 42356
rect 59170 42276 59176 42288
rect 52748 42248 59176 42276
rect 49200 42236 49206 42248
rect 59170 42236 59176 42248
rect 59228 42276 59234 42288
rect 59357 42279 59415 42285
rect 59357 42276 59369 42279
rect 59228 42248 59369 42276
rect 59228 42236 59234 42248
rect 59357 42245 59369 42248
rect 59403 42245 59415 42279
rect 59357 42239 59415 42245
rect 48958 42168 48964 42220
rect 49016 42208 49022 42220
rect 51721 42211 51779 42217
rect 51721 42208 51733 42211
rect 49016 42180 51733 42208
rect 49016 42168 49022 42180
rect 51721 42177 51733 42180
rect 51767 42208 51779 42211
rect 53469 42211 53527 42217
rect 53469 42208 53481 42211
rect 51767 42180 53481 42208
rect 51767 42177 51779 42180
rect 51721 42171 51779 42177
rect 53469 42177 53481 42180
rect 53515 42208 53527 42211
rect 53742 42208 53748 42220
rect 53515 42180 53748 42208
rect 53515 42177 53527 42180
rect 53469 42171 53527 42177
rect 53742 42168 53748 42180
rect 53800 42168 53806 42220
rect 56134 42208 56140 42220
rect 54956 42180 56140 42208
rect 48777 42143 48835 42149
rect 48777 42109 48789 42143
rect 48823 42109 48835 42143
rect 49050 42140 49056 42152
rect 49011 42112 49056 42140
rect 48777 42103 48835 42109
rect 44968 42044 45140 42072
rect 44968 42032 44974 42044
rect 45186 42032 45192 42084
rect 45244 42072 45250 42084
rect 46201 42075 46259 42081
rect 46201 42072 46213 42075
rect 45244 42044 46213 42072
rect 45244 42032 45250 42044
rect 46201 42041 46213 42044
rect 46247 42041 46259 42075
rect 48792 42072 48820 42103
rect 49050 42100 49056 42112
rect 49108 42100 49114 42152
rect 49237 42143 49295 42149
rect 49237 42109 49249 42143
rect 49283 42140 49295 42143
rect 49326 42140 49332 42152
rect 49283 42112 49332 42140
rect 49283 42109 49295 42112
rect 49237 42103 49295 42109
rect 49326 42100 49332 42112
rect 49384 42140 49390 42152
rect 50614 42140 50620 42152
rect 49384 42112 50620 42140
rect 49384 42100 49390 42112
rect 50614 42100 50620 42112
rect 50672 42100 50678 42152
rect 51994 42140 52000 42152
rect 51955 42112 52000 42140
rect 51994 42100 52000 42112
rect 52052 42100 52058 42152
rect 54956 42149 54984 42180
rect 56134 42168 56140 42180
rect 56192 42168 56198 42220
rect 59372 42208 59400 42239
rect 59446 42236 59452 42288
rect 59504 42276 59510 42288
rect 65702 42276 65708 42288
rect 59504 42248 65708 42276
rect 59504 42236 59510 42248
rect 65702 42236 65708 42248
rect 65760 42236 65766 42288
rect 60553 42211 60611 42217
rect 59372 42180 60136 42208
rect 54941 42143 54999 42149
rect 54941 42109 54953 42143
rect 54987 42109 54999 42143
rect 55950 42140 55956 42152
rect 55911 42112 55956 42140
rect 54941 42103 54999 42109
rect 55950 42100 55956 42112
rect 56008 42140 56014 42152
rect 56229 42143 56287 42149
rect 56229 42140 56241 42143
rect 56008 42112 56241 42140
rect 56008 42100 56014 42112
rect 56229 42109 56241 42112
rect 56275 42109 56287 42143
rect 56229 42103 56287 42109
rect 58526 42100 58532 42152
rect 58584 42140 58590 42152
rect 60108 42149 60136 42180
rect 60553 42177 60565 42211
rect 60599 42208 60611 42211
rect 61010 42208 61016 42220
rect 60599 42180 61016 42208
rect 60599 42177 60611 42180
rect 60553 42171 60611 42177
rect 61010 42168 61016 42180
rect 61068 42208 61074 42220
rect 61930 42208 61936 42220
rect 61068 42180 61936 42208
rect 61068 42168 61074 42180
rect 61930 42168 61936 42180
rect 61988 42168 61994 42220
rect 63862 42208 63868 42220
rect 62960 42180 63868 42208
rect 59725 42143 59783 42149
rect 59725 42140 59737 42143
rect 58584 42112 59737 42140
rect 58584 42100 58590 42112
rect 59725 42109 59737 42112
rect 59771 42109 59783 42143
rect 59725 42103 59783 42109
rect 60093 42143 60151 42149
rect 60093 42109 60105 42143
rect 60139 42109 60151 42143
rect 60093 42103 60151 42109
rect 61473 42143 61531 42149
rect 61473 42109 61485 42143
rect 61519 42140 61531 42143
rect 61562 42140 61568 42152
rect 61519 42112 61568 42140
rect 61519 42109 61531 42112
rect 61473 42103 61531 42109
rect 49418 42072 49424 42084
rect 48792 42044 49424 42072
rect 46201 42035 46259 42041
rect 49418 42032 49424 42044
rect 49476 42032 49482 42084
rect 55030 42072 55036 42084
rect 54991 42044 55036 42072
rect 55030 42032 55036 42044
rect 55088 42032 55094 42084
rect 59740 42072 59768 42103
rect 61562 42100 61568 42112
rect 61620 42100 61626 42152
rect 61658 42143 61716 42149
rect 61658 42109 61670 42143
rect 61704 42109 61716 42143
rect 61658 42103 61716 42109
rect 61672 42072 61700 42103
rect 61746 42100 61752 42152
rect 61804 42140 61810 42152
rect 62960 42149 62988 42180
rect 63862 42168 63868 42180
rect 63920 42168 63926 42220
rect 65797 42211 65855 42217
rect 65797 42177 65809 42211
rect 65843 42208 65855 42211
rect 66070 42208 66076 42220
rect 65843 42180 66076 42208
rect 65843 42177 65855 42180
rect 65797 42171 65855 42177
rect 66070 42168 66076 42180
rect 66128 42168 66134 42220
rect 66254 42168 66260 42220
rect 66312 42208 66318 42220
rect 66349 42211 66407 42217
rect 66349 42208 66361 42211
rect 66312 42180 66361 42208
rect 66312 42168 66318 42180
rect 66349 42177 66361 42180
rect 66395 42177 66407 42211
rect 66898 42208 66904 42220
rect 66349 42171 66407 42177
rect 66640 42180 66904 42208
rect 66640 42149 66668 42180
rect 66898 42168 66904 42180
rect 66956 42208 66962 42220
rect 69198 42208 69204 42220
rect 66956 42180 69204 42208
rect 66956 42168 66962 42180
rect 69198 42168 69204 42180
rect 69256 42168 69262 42220
rect 69658 42168 69664 42220
rect 69716 42208 69722 42220
rect 70765 42211 70823 42217
rect 70765 42208 70777 42211
rect 69716 42180 70777 42208
rect 69716 42168 69722 42180
rect 70765 42177 70777 42180
rect 70811 42208 70823 42211
rect 70857 42211 70915 42217
rect 70857 42208 70869 42211
rect 70811 42180 70869 42208
rect 70811 42177 70823 42180
rect 70765 42171 70823 42177
rect 70857 42177 70869 42180
rect 70903 42208 70915 42211
rect 72510 42208 72516 42220
rect 70903 42180 72516 42208
rect 70903 42177 70915 42180
rect 70857 42171 70915 42177
rect 72510 42168 72516 42180
rect 72568 42168 72574 42220
rect 62945 42143 63003 42149
rect 62945 42140 62957 42143
rect 61804 42112 62957 42140
rect 61804 42100 61810 42112
rect 62945 42109 62957 42112
rect 62991 42109 63003 42143
rect 62945 42103 63003 42109
rect 63497 42143 63555 42149
rect 63497 42109 63509 42143
rect 63543 42109 63555 42143
rect 63497 42103 63555 42109
rect 66625 42143 66683 42149
rect 66625 42109 66637 42143
rect 66671 42109 66683 42143
rect 66625 42103 66683 42109
rect 66809 42143 66867 42149
rect 66809 42109 66821 42143
rect 66855 42109 66867 42143
rect 66809 42103 66867 42109
rect 69477 42143 69535 42149
rect 69477 42109 69489 42143
rect 69523 42109 69535 42143
rect 69750 42140 69756 42152
rect 69711 42112 69756 42140
rect 69477 42103 69535 42109
rect 62022 42072 62028 42084
rect 59740 42044 60872 42072
rect 61672 42044 62028 42072
rect 49142 42004 49148 42016
rect 43916 41976 49148 42004
rect 49142 41964 49148 41976
rect 49200 41964 49206 42016
rect 52270 41964 52276 42016
rect 52328 42004 52334 42016
rect 53101 42007 53159 42013
rect 53101 42004 53113 42007
rect 52328 41976 53113 42004
rect 52328 41964 52334 41976
rect 53101 41973 53113 41976
rect 53147 41973 53159 42007
rect 53101 41967 53159 41973
rect 55398 41964 55404 42016
rect 55456 42004 55462 42016
rect 56045 42007 56103 42013
rect 56045 42004 56057 42007
rect 55456 41976 56057 42004
rect 55456 41964 55462 41976
rect 56045 41973 56057 41976
rect 56091 42004 56103 42007
rect 56226 42004 56232 42016
rect 56091 41976 56232 42004
rect 56091 41973 56103 41976
rect 56045 41967 56103 41973
rect 56226 41964 56232 41976
rect 56284 41964 56290 42016
rect 59630 42004 59636 42016
rect 59591 41976 59636 42004
rect 59630 41964 59636 41976
rect 59688 41964 59694 42016
rect 60844 42013 60872 42044
rect 62022 42032 62028 42044
rect 62080 42072 62086 42084
rect 63512 42072 63540 42103
rect 62080 42044 63540 42072
rect 62080 42032 62086 42044
rect 65978 42032 65984 42084
rect 66036 42072 66042 42084
rect 66530 42072 66536 42084
rect 66036 42044 66536 42072
rect 66036 42032 66042 42044
rect 66530 42032 66536 42044
rect 66588 42072 66594 42084
rect 66824 42072 66852 42103
rect 66901 42075 66959 42081
rect 66901 42072 66913 42075
rect 66588 42044 66913 42072
rect 66588 42032 66594 42044
rect 66901 42041 66913 42044
rect 66947 42041 66959 42075
rect 69492 42072 69520 42103
rect 69750 42100 69756 42112
rect 69808 42100 69814 42152
rect 71130 42140 71136 42152
rect 71091 42112 71136 42140
rect 71130 42100 71136 42112
rect 71188 42100 71194 42152
rect 70302 42072 70308 42084
rect 69492 42044 70308 42072
rect 66901 42035 66959 42041
rect 70302 42032 70308 42044
rect 70360 42032 70366 42084
rect 60829 42007 60887 42013
rect 60829 41973 60841 42007
rect 60875 42004 60887 42007
rect 66162 42004 66168 42016
rect 60875 41976 66168 42004
rect 60875 41973 60887 41976
rect 60829 41967 60887 41973
rect 66162 41964 66168 41976
rect 66220 41964 66226 42016
rect 71406 41964 71412 42016
rect 71464 42004 71470 42016
rect 72237 42007 72295 42013
rect 72237 42004 72249 42007
rect 71464 41976 72249 42004
rect 71464 41964 71470 41976
rect 72237 41973 72249 41976
rect 72283 41973 72295 42007
rect 72237 41967 72295 41973
rect 1104 41914 111136 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 50326 41914
rect 50378 41862 50390 41914
rect 50442 41862 50454 41914
rect 50506 41862 50518 41914
rect 50570 41862 81046 41914
rect 81098 41862 81110 41914
rect 81162 41862 81174 41914
rect 81226 41862 81238 41914
rect 81290 41862 111136 41914
rect 1104 41840 111136 41862
rect 5074 41760 5080 41812
rect 5132 41800 5138 41812
rect 5261 41803 5319 41809
rect 5261 41800 5273 41803
rect 5132 41772 5273 41800
rect 5132 41760 5138 41772
rect 5261 41769 5273 41772
rect 5307 41769 5319 41803
rect 10410 41800 10416 41812
rect 5261 41763 5319 41769
rect 5368 41772 10416 41800
rect 5368 41732 5396 41772
rect 10410 41760 10416 41772
rect 10468 41760 10474 41812
rect 10686 41760 10692 41812
rect 10744 41800 10750 41812
rect 10873 41803 10931 41809
rect 10873 41800 10885 41803
rect 10744 41772 10885 41800
rect 10744 41760 10750 41772
rect 10873 41769 10885 41772
rect 10919 41769 10931 41803
rect 10873 41763 10931 41769
rect 10962 41760 10968 41812
rect 11020 41800 11026 41812
rect 11241 41803 11299 41809
rect 11241 41800 11253 41803
rect 11020 41772 11253 41800
rect 11020 41760 11026 41772
rect 11241 41769 11253 41772
rect 11287 41800 11299 41803
rect 12250 41800 12256 41812
rect 11287 41772 12256 41800
rect 11287 41769 11299 41772
rect 11241 41763 11299 41769
rect 12250 41760 12256 41772
rect 12308 41760 12314 41812
rect 14752 41772 14964 41800
rect 4264 41704 5396 41732
rect 4264 41673 4292 41704
rect 4249 41667 4307 41673
rect 4249 41633 4261 41667
rect 4295 41633 4307 41667
rect 4249 41627 4307 41633
rect 4341 41667 4399 41673
rect 4341 41633 4353 41667
rect 4387 41664 4399 41667
rect 4614 41664 4620 41676
rect 4387 41636 4620 41664
rect 4387 41633 4399 41636
rect 4341 41627 4399 41633
rect 4614 41624 4620 41636
rect 4672 41624 4678 41676
rect 4816 41673 4844 41704
rect 8110 41692 8116 41744
rect 8168 41732 8174 41744
rect 9401 41735 9459 41741
rect 9401 41732 9413 41735
rect 8168 41704 9413 41732
rect 8168 41692 8174 41704
rect 9401 41701 9413 41704
rect 9447 41732 9459 41735
rect 9490 41732 9496 41744
rect 9447 41704 9496 41732
rect 9447 41701 9459 41704
rect 9401 41695 9459 41701
rect 9490 41692 9496 41704
rect 9548 41732 9554 41744
rect 9548 41704 9720 41732
rect 9548 41692 9554 41704
rect 4801 41667 4859 41673
rect 4801 41633 4813 41667
rect 4847 41633 4859 41667
rect 4801 41627 4859 41633
rect 4985 41667 5043 41673
rect 4985 41633 4997 41667
rect 5031 41664 5043 41667
rect 5166 41664 5172 41676
rect 5031 41636 5172 41664
rect 5031 41633 5043 41636
rect 4985 41627 5043 41633
rect 5166 41624 5172 41636
rect 5224 41624 5230 41676
rect 7285 41667 7343 41673
rect 7285 41633 7297 41667
rect 7331 41664 7343 41667
rect 8018 41664 8024 41676
rect 7331 41636 8024 41664
rect 7331 41633 7343 41636
rect 7285 41627 7343 41633
rect 8018 41624 8024 41636
rect 8076 41624 8082 41676
rect 8205 41667 8263 41673
rect 8205 41633 8217 41667
rect 8251 41664 8263 41667
rect 8294 41664 8300 41676
rect 8251 41636 8300 41664
rect 8251 41633 8263 41636
rect 8205 41627 8263 41633
rect 8294 41624 8300 41636
rect 8352 41624 8358 41676
rect 8573 41667 8631 41673
rect 8573 41633 8585 41667
rect 8619 41664 8631 41667
rect 8662 41664 8668 41676
rect 8619 41636 8668 41664
rect 8619 41633 8631 41636
rect 8573 41627 8631 41633
rect 8662 41624 8668 41636
rect 8720 41624 8726 41676
rect 9692 41673 9720 41704
rect 9766 41692 9772 41744
rect 9824 41732 9830 41744
rect 9824 41704 11100 41732
rect 9824 41692 9830 41704
rect 8757 41667 8815 41673
rect 8757 41633 8769 41667
rect 8803 41633 8815 41667
rect 8757 41627 8815 41633
rect 9677 41667 9735 41673
rect 9677 41633 9689 41667
rect 9723 41633 9735 41667
rect 9677 41627 9735 41633
rect 9861 41667 9919 41673
rect 9861 41633 9873 41667
rect 9907 41664 9919 41667
rect 9950 41664 9956 41676
rect 9907 41636 9956 41664
rect 9907 41633 9919 41636
rect 9861 41627 9919 41633
rect 5184 41528 5212 41624
rect 5350 41556 5356 41608
rect 5408 41596 5414 41608
rect 7561 41599 7619 41605
rect 7561 41596 7573 41599
rect 5408 41568 7573 41596
rect 5408 41556 5414 41568
rect 7561 41565 7573 41568
rect 7607 41565 7619 41599
rect 8772 41596 8800 41627
rect 9950 41624 9956 41636
rect 10008 41664 10014 41676
rect 10410 41664 10416 41676
rect 10008 41636 10416 41664
rect 10008 41624 10014 41636
rect 10410 41624 10416 41636
rect 10468 41624 10474 41676
rect 10597 41667 10655 41673
rect 10597 41633 10609 41667
rect 10643 41664 10655 41667
rect 10962 41664 10968 41676
rect 10643 41636 10968 41664
rect 10643 41633 10655 41636
rect 10597 41627 10655 41633
rect 10962 41624 10968 41636
rect 11020 41624 11026 41676
rect 11072 41596 11100 41704
rect 11514 41692 11520 41744
rect 11572 41732 11578 41744
rect 14642 41732 14648 41744
rect 11572 41704 14648 41732
rect 11572 41692 11578 41704
rect 14642 41692 14648 41704
rect 14700 41692 14706 41744
rect 13814 41624 13820 41676
rect 13872 41664 13878 41676
rect 14001 41667 14059 41673
rect 14001 41664 14013 41667
rect 13872 41636 14013 41664
rect 13872 41624 13878 41636
rect 14001 41633 14013 41636
rect 14047 41633 14059 41667
rect 14001 41627 14059 41633
rect 14752 41596 14780 41772
rect 14936 41732 14964 41772
rect 15010 41760 15016 41812
rect 15068 41800 15074 41812
rect 16485 41803 16543 41809
rect 16485 41800 16497 41803
rect 15068 41772 16497 41800
rect 15068 41760 15074 41772
rect 16485 41769 16497 41772
rect 16531 41800 16543 41803
rect 16577 41803 16635 41809
rect 16577 41800 16589 41803
rect 16531 41772 16589 41800
rect 16531 41769 16543 41772
rect 16485 41763 16543 41769
rect 16577 41769 16589 41772
rect 16623 41769 16635 41803
rect 16577 41763 16635 41769
rect 16850 41760 16856 41812
rect 16908 41800 16914 41812
rect 17770 41800 17776 41812
rect 16908 41772 17776 41800
rect 16908 41760 16914 41772
rect 17770 41760 17776 41772
rect 17828 41760 17834 41812
rect 17954 41800 17960 41812
rect 17915 41772 17960 41800
rect 17954 41760 17960 41772
rect 18012 41760 18018 41812
rect 18322 41800 18328 41812
rect 18235 41772 18328 41800
rect 18322 41760 18328 41772
rect 18380 41800 18386 41812
rect 20254 41800 20260 41812
rect 18380 41772 20260 41800
rect 18380 41760 18386 41772
rect 20254 41760 20260 41772
rect 20312 41760 20318 41812
rect 23750 41760 23756 41812
rect 23808 41800 23814 41812
rect 23808 41772 37228 41800
rect 23808 41760 23814 41772
rect 23934 41732 23940 41744
rect 14936 41704 23940 41732
rect 23934 41692 23940 41704
rect 23992 41692 23998 41744
rect 24670 41732 24676 41744
rect 24044 41704 24676 41732
rect 16485 41667 16543 41673
rect 16485 41633 16497 41667
rect 16531 41664 16543 41667
rect 16761 41667 16819 41673
rect 16761 41664 16773 41667
rect 16531 41636 16773 41664
rect 16531 41633 16543 41636
rect 16485 41627 16543 41633
rect 16761 41633 16773 41636
rect 16807 41633 16819 41667
rect 16761 41627 16819 41633
rect 16945 41667 17003 41673
rect 16945 41633 16957 41667
rect 16991 41664 17003 41667
rect 17310 41664 17316 41676
rect 16991 41636 17316 41664
rect 16991 41633 17003 41636
rect 16945 41627 17003 41633
rect 7561 41559 7619 41565
rect 7668 41568 10088 41596
rect 11072 41568 14780 41596
rect 5629 41531 5687 41537
rect 5629 41528 5641 41531
rect 5184 41500 5641 41528
rect 5629 41497 5641 41500
rect 5675 41528 5687 41531
rect 7469 41531 7527 41537
rect 7469 41528 7481 41531
rect 5675 41500 7481 41528
rect 5675 41497 5687 41500
rect 5629 41491 5687 41497
rect 7469 41497 7481 41500
rect 7515 41528 7527 41531
rect 7668 41528 7696 41568
rect 7515 41500 7696 41528
rect 7515 41497 7527 41500
rect 7469 41491 7527 41497
rect 8846 41488 8852 41540
rect 8904 41528 8910 41540
rect 8941 41531 8999 41537
rect 8941 41528 8953 41531
rect 8904 41500 8953 41528
rect 8904 41488 8910 41500
rect 8941 41497 8953 41500
rect 8987 41528 8999 41531
rect 9950 41528 9956 41540
rect 8987 41500 9956 41528
rect 8987 41497 8999 41500
rect 8941 41491 8999 41497
rect 9950 41488 9956 41500
rect 10008 41488 10014 41540
rect 10060 41528 10088 41568
rect 14918 41556 14924 41608
rect 14976 41596 14982 41608
rect 16960 41596 16988 41627
rect 17310 41624 17316 41636
rect 17368 41624 17374 41676
rect 17494 41664 17500 41676
rect 17455 41636 17500 41664
rect 17494 41624 17500 41636
rect 17552 41624 17558 41676
rect 17586 41624 17592 41676
rect 17644 41664 17650 41676
rect 17681 41667 17739 41673
rect 17681 41664 17693 41667
rect 17644 41636 17693 41664
rect 17644 41624 17650 41636
rect 17681 41633 17693 41636
rect 17727 41633 17739 41667
rect 17681 41627 17739 41633
rect 17862 41624 17868 41676
rect 17920 41664 17926 41676
rect 23382 41664 23388 41676
rect 17920 41636 23388 41664
rect 17920 41624 17926 41636
rect 23382 41624 23388 41636
rect 23440 41624 23446 41676
rect 23474 41624 23480 41676
rect 23532 41664 23538 41676
rect 24044 41673 24072 41704
rect 24670 41692 24676 41704
rect 24728 41692 24734 41744
rect 25682 41692 25688 41744
rect 25740 41732 25746 41744
rect 30558 41732 30564 41744
rect 25740 41704 30564 41732
rect 25740 41692 25746 41704
rect 30558 41692 30564 41704
rect 30616 41692 30622 41744
rect 31662 41692 31668 41744
rect 31720 41732 31726 41744
rect 35342 41732 35348 41744
rect 31720 41704 35348 41732
rect 31720 41692 31726 41704
rect 35342 41692 35348 41704
rect 35400 41692 35406 41744
rect 36909 41735 36967 41741
rect 36909 41732 36921 41735
rect 36188 41704 36921 41732
rect 24029 41667 24087 41673
rect 23532 41636 23980 41664
rect 23532 41624 23538 41636
rect 23566 41596 23572 41608
rect 14976 41568 16988 41596
rect 17880 41568 23572 41596
rect 14976 41556 14982 41568
rect 17880 41528 17908 41568
rect 23566 41556 23572 41568
rect 23624 41556 23630 41608
rect 23845 41599 23903 41605
rect 23845 41565 23857 41599
rect 23891 41565 23903 41599
rect 23952 41596 23980 41636
rect 24029 41633 24041 41667
rect 24075 41633 24087 41667
rect 24486 41664 24492 41676
rect 24447 41636 24492 41664
rect 24029 41627 24087 41633
rect 24486 41624 24492 41636
rect 24544 41624 24550 41676
rect 24581 41667 24639 41673
rect 24581 41633 24593 41667
rect 24627 41664 24639 41667
rect 25406 41664 25412 41676
rect 24627 41636 25412 41664
rect 24627 41633 24639 41636
rect 24581 41627 24639 41633
rect 25406 41624 25412 41636
rect 25464 41624 25470 41676
rect 26234 41664 26240 41676
rect 26195 41636 26240 41664
rect 26234 41624 26240 41636
rect 26292 41624 26298 41676
rect 29730 41624 29736 41676
rect 29788 41664 29794 41676
rect 29825 41667 29883 41673
rect 29825 41664 29837 41667
rect 29788 41636 29837 41664
rect 29788 41624 29794 41636
rect 29825 41633 29837 41636
rect 29871 41633 29883 41667
rect 29825 41627 29883 41633
rect 30374 41624 30380 41676
rect 30432 41664 30438 41676
rect 30837 41667 30895 41673
rect 30837 41664 30849 41667
rect 30432 41636 30849 41664
rect 30432 41624 30438 41636
rect 30837 41633 30849 41636
rect 30883 41664 30895 41667
rect 30926 41664 30932 41676
rect 30883 41636 30932 41664
rect 30883 41633 30895 41636
rect 30837 41627 30895 41633
rect 30926 41624 30932 41636
rect 30984 41624 30990 41676
rect 35434 41664 35440 41676
rect 35395 41636 35440 41664
rect 35434 41624 35440 41636
rect 35492 41624 35498 41676
rect 35621 41667 35679 41673
rect 35621 41633 35633 41667
rect 35667 41664 35679 41667
rect 35986 41664 35992 41676
rect 35667 41636 35992 41664
rect 35667 41633 35679 41636
rect 35621 41627 35679 41633
rect 35986 41624 35992 41636
rect 36044 41624 36050 41676
rect 36188 41673 36216 41704
rect 36909 41701 36921 41704
rect 36955 41732 36967 41735
rect 37090 41732 37096 41744
rect 36955 41704 37096 41732
rect 36955 41701 36967 41704
rect 36909 41695 36967 41701
rect 37090 41692 37096 41704
rect 37148 41692 37154 41744
rect 37200 41732 37228 41772
rect 37274 41760 37280 41812
rect 37332 41800 37338 41812
rect 43714 41800 43720 41812
rect 37332 41772 38792 41800
rect 37332 41760 37338 41772
rect 37642 41732 37648 41744
rect 37200 41704 37648 41732
rect 37642 41692 37648 41704
rect 37700 41692 37706 41744
rect 38102 41732 38108 41744
rect 37936 41704 38108 41732
rect 36173 41667 36231 41673
rect 36173 41633 36185 41667
rect 36219 41633 36231 41667
rect 36173 41627 36231 41633
rect 36262 41624 36268 41676
rect 36320 41664 36326 41676
rect 37936 41673 37964 41704
rect 38102 41692 38108 41704
rect 38160 41692 38166 41744
rect 38654 41732 38660 41744
rect 38396 41704 38660 41732
rect 38396 41673 38424 41704
rect 38654 41692 38660 41704
rect 38712 41692 38718 41744
rect 36357 41667 36415 41673
rect 36357 41664 36369 41667
rect 36320 41636 36369 41664
rect 36320 41624 36326 41636
rect 36357 41633 36369 41636
rect 36403 41633 36415 41667
rect 36357 41627 36415 41633
rect 37921 41667 37979 41673
rect 37921 41633 37933 41667
rect 37967 41633 37979 41667
rect 37921 41627 37979 41633
rect 38381 41667 38439 41673
rect 38381 41633 38393 41667
rect 38427 41633 38439 41667
rect 38381 41627 38439 41633
rect 38473 41667 38531 41673
rect 38473 41633 38485 41667
rect 38519 41664 38531 41667
rect 38764 41664 38792 41772
rect 40696 41772 43720 41800
rect 40696 41664 40724 41772
rect 43714 41760 43720 41772
rect 43772 41760 43778 41812
rect 44542 41800 44548 41812
rect 44503 41772 44548 41800
rect 44542 41760 44548 41772
rect 44600 41760 44606 41812
rect 45094 41760 45100 41812
rect 45152 41800 45158 41812
rect 49050 41800 49056 41812
rect 45152 41772 45692 41800
rect 49011 41772 49056 41800
rect 45152 41760 45158 41772
rect 43349 41735 43407 41741
rect 43349 41701 43361 41735
rect 43395 41732 43407 41735
rect 44726 41732 44732 41744
rect 43395 41704 44732 41732
rect 43395 41701 43407 41704
rect 43349 41695 43407 41701
rect 44726 41692 44732 41704
rect 44784 41692 44790 41744
rect 45664 41732 45692 41772
rect 49050 41760 49056 41772
rect 49108 41760 49114 41812
rect 51626 41760 51632 41812
rect 51684 41760 51690 41812
rect 51721 41803 51779 41809
rect 51721 41769 51733 41803
rect 51767 41800 51779 41803
rect 51994 41800 52000 41812
rect 51767 41772 52000 41800
rect 51767 41769 51779 41772
rect 51721 41763 51779 41769
rect 51994 41760 52000 41772
rect 52052 41760 52058 41812
rect 54205 41803 54263 41809
rect 54205 41769 54217 41803
rect 54251 41800 54263 41803
rect 58802 41800 58808 41812
rect 54251 41772 58808 41800
rect 54251 41769 54263 41772
rect 54205 41763 54263 41769
rect 58802 41760 58808 41772
rect 58860 41760 58866 41812
rect 59170 41800 59176 41812
rect 59131 41772 59176 41800
rect 59170 41760 59176 41772
rect 59228 41800 59234 41812
rect 59909 41803 59967 41809
rect 59909 41800 59921 41803
rect 59228 41772 59921 41800
rect 59228 41760 59234 41772
rect 59909 41769 59921 41772
rect 59955 41800 59967 41803
rect 63862 41800 63868 41812
rect 59955 41772 61240 41800
rect 63823 41772 63868 41800
rect 59955 41769 59967 41772
rect 59909 41763 59967 41769
rect 51442 41732 51448 41744
rect 45664 41704 51448 41732
rect 51442 41692 51448 41704
rect 51500 41692 51506 41744
rect 43530 41664 43536 41676
rect 38519 41636 40724 41664
rect 43491 41636 43536 41664
rect 38519 41633 38531 41636
rect 38473 41627 38531 41633
rect 43530 41624 43536 41636
rect 43588 41624 43594 41676
rect 43898 41664 43904 41676
rect 43859 41636 43904 41664
rect 43898 41624 43904 41636
rect 43956 41624 43962 41676
rect 45005 41667 45063 41673
rect 44008 41636 44864 41664
rect 25133 41599 25191 41605
rect 23952 41568 24256 41596
rect 23845 41559 23903 41565
rect 10060 41500 16896 41528
rect 9122 41460 9128 41472
rect 9083 41432 9128 41460
rect 9122 41420 9128 41432
rect 9180 41420 9186 41472
rect 10410 41420 10416 41472
rect 10468 41460 10474 41472
rect 11333 41463 11391 41469
rect 11333 41460 11345 41463
rect 10468 41432 11345 41460
rect 10468 41420 10474 41432
rect 11333 41429 11345 41432
rect 11379 41460 11391 41463
rect 11514 41460 11520 41472
rect 11379 41432 11520 41460
rect 11379 41429 11391 41432
rect 11333 41423 11391 41429
rect 11514 41420 11520 41432
rect 11572 41420 11578 41472
rect 13354 41420 13360 41472
rect 13412 41460 13418 41472
rect 13722 41460 13728 41472
rect 13412 41432 13728 41460
rect 13412 41420 13418 41432
rect 13722 41420 13728 41432
rect 13780 41460 13786 41472
rect 13817 41463 13875 41469
rect 13817 41460 13829 41463
rect 13780 41432 13829 41460
rect 13780 41420 13786 41432
rect 13817 41429 13829 41432
rect 13863 41429 13875 41463
rect 14182 41460 14188 41472
rect 14095 41432 14188 41460
rect 13817 41423 13875 41429
rect 14182 41420 14188 41432
rect 14240 41460 14246 41472
rect 15654 41460 15660 41472
rect 14240 41432 15660 41460
rect 14240 41420 14246 41432
rect 15654 41420 15660 41432
rect 15712 41420 15718 41472
rect 16868 41460 16896 41500
rect 17236 41500 17908 41528
rect 17236 41460 17264 41500
rect 18046 41488 18052 41540
rect 18104 41528 18110 41540
rect 23661 41531 23719 41537
rect 23661 41528 23673 41531
rect 18104 41500 23673 41528
rect 18104 41488 18110 41500
rect 23661 41497 23673 41500
rect 23707 41528 23719 41531
rect 23860 41528 23888 41559
rect 23934 41528 23940 41540
rect 23707 41500 23940 41528
rect 23707 41497 23719 41500
rect 23661 41491 23719 41497
rect 23934 41488 23940 41500
rect 23992 41488 23998 41540
rect 24228 41528 24256 41568
rect 25133 41565 25145 41599
rect 25179 41596 25191 41599
rect 26786 41596 26792 41608
rect 25179 41568 26792 41596
rect 25179 41565 25191 41568
rect 25133 41559 25191 41565
rect 26786 41556 26792 41568
rect 26844 41556 26850 41608
rect 29917 41599 29975 41605
rect 29917 41565 29929 41599
rect 29963 41596 29975 41599
rect 31570 41596 31576 41608
rect 29963 41568 31576 41596
rect 29963 41565 29975 41568
rect 29917 41559 29975 41565
rect 31570 41556 31576 41568
rect 31628 41556 31634 41608
rect 37274 41596 37280 41608
rect 36556 41568 37280 41596
rect 26053 41531 26111 41537
rect 26053 41528 26065 41531
rect 24228 41500 26065 41528
rect 26053 41497 26065 41500
rect 26099 41528 26111 41531
rect 26510 41528 26516 41540
rect 26099 41500 26516 41528
rect 26099 41497 26111 41500
rect 26053 41491 26111 41497
rect 26510 41488 26516 41500
rect 26568 41488 26574 41540
rect 30929 41531 30987 41537
rect 30929 41497 30941 41531
rect 30975 41528 30987 41531
rect 36556 41528 36584 41568
rect 37274 41556 37280 41568
rect 37332 41596 37338 41608
rect 37737 41599 37795 41605
rect 37332 41568 37377 41596
rect 37332 41556 37338 41568
rect 37737 41565 37749 41599
rect 37783 41565 37795 41599
rect 37737 41559 37795 41565
rect 39301 41599 39359 41605
rect 39301 41565 39313 41599
rect 39347 41596 39359 41599
rect 44008 41596 44036 41636
rect 39347 41568 44036 41596
rect 44729 41599 44787 41605
rect 39347 41565 39359 41568
rect 39301 41559 39359 41565
rect 44729 41565 44741 41599
rect 44775 41565 44787 41599
rect 44836 41596 44864 41636
rect 45005 41633 45017 41667
rect 45051 41664 45063 41667
rect 45830 41664 45836 41676
rect 45051 41636 45836 41664
rect 45051 41633 45063 41636
rect 45005 41627 45063 41633
rect 45830 41624 45836 41636
rect 45888 41624 45894 41676
rect 45922 41624 45928 41676
rect 45980 41664 45986 41676
rect 47854 41664 47860 41676
rect 45980 41636 47860 41664
rect 45980 41624 45986 41636
rect 47854 41624 47860 41636
rect 47912 41664 47918 41676
rect 51644 41673 51672 41760
rect 59357 41735 59415 41741
rect 59357 41732 59369 41735
rect 52196 41704 59369 41732
rect 48961 41667 49019 41673
rect 48961 41664 48973 41667
rect 47912 41636 48973 41664
rect 47912 41624 47918 41636
rect 48961 41633 48973 41636
rect 49007 41664 49019 41667
rect 49237 41667 49295 41673
rect 49237 41664 49249 41667
rect 49007 41636 49249 41664
rect 49007 41633 49019 41636
rect 48961 41627 49019 41633
rect 49237 41633 49249 41636
rect 49283 41633 49295 41667
rect 49237 41627 49295 41633
rect 51629 41667 51687 41673
rect 51629 41633 51641 41667
rect 51675 41633 51687 41667
rect 51629 41627 51687 41633
rect 51718 41624 51724 41676
rect 51776 41664 51782 41676
rect 52196 41664 52224 41704
rect 51776 41636 52224 41664
rect 53101 41667 53159 41673
rect 51776 41624 51782 41636
rect 53101 41633 53113 41667
rect 53147 41664 53159 41667
rect 53282 41664 53288 41676
rect 53147 41636 53288 41664
rect 53147 41633 53159 41636
rect 53101 41627 53159 41633
rect 53282 41624 53288 41636
rect 53340 41624 53346 41676
rect 54389 41667 54447 41673
rect 54389 41664 54401 41667
rect 54036 41636 54401 41664
rect 51534 41596 51540 41608
rect 44836 41568 51540 41596
rect 44729 41559 44787 41565
rect 30975 41500 36584 41528
rect 36633 41531 36691 41537
rect 30975 41497 30987 41500
rect 30929 41491 30987 41497
rect 36633 41497 36645 41531
rect 36679 41528 36691 41531
rect 37642 41528 37648 41540
rect 36679 41500 37648 41528
rect 36679 41497 36691 41500
rect 36633 41491 36691 41497
rect 16868 41432 17264 41460
rect 17310 41420 17316 41472
rect 17368 41460 17374 41472
rect 17954 41460 17960 41472
rect 17368 41432 17960 41460
rect 17368 41420 17374 41432
rect 17954 41420 17960 41432
rect 18012 41420 18018 41472
rect 18506 41460 18512 41472
rect 18467 41432 18512 41460
rect 18506 41420 18512 41432
rect 18564 41420 18570 41472
rect 23474 41420 23480 41472
rect 23532 41460 23538 41472
rect 23569 41463 23627 41469
rect 23569 41460 23581 41463
rect 23532 41432 23581 41460
rect 23532 41420 23538 41432
rect 23569 41429 23581 41432
rect 23615 41460 23627 41463
rect 24486 41460 24492 41472
rect 23615 41432 24492 41460
rect 23615 41429 23627 41432
rect 23569 41423 23627 41429
rect 24486 41420 24492 41432
rect 24544 41420 24550 41472
rect 25498 41460 25504 41472
rect 25459 41432 25504 41460
rect 25498 41420 25504 41432
rect 25556 41420 25562 41472
rect 25590 41420 25596 41472
rect 25648 41460 25654 41472
rect 30944 41460 30972 41491
rect 37642 41488 37648 41500
rect 37700 41488 37706 41540
rect 37458 41460 37464 41472
rect 25648 41432 30972 41460
rect 37419 41432 37464 41460
rect 25648 41420 25654 41432
rect 37458 41420 37464 41432
rect 37516 41460 37522 41472
rect 37752 41460 37780 41559
rect 38286 41488 38292 41540
rect 38344 41528 38350 41540
rect 38841 41531 38899 41537
rect 38841 41528 38853 41531
rect 38344 41500 38853 41528
rect 38344 41488 38350 41500
rect 38841 41497 38853 41500
rect 38887 41497 38899 41531
rect 38841 41491 38899 41497
rect 37516 41432 37780 41460
rect 37516 41420 37522 41432
rect 38102 41420 38108 41472
rect 38160 41460 38166 41472
rect 39316 41460 39344 41559
rect 44542 41488 44548 41540
rect 44600 41528 44606 41540
rect 44744 41528 44772 41559
rect 51534 41556 51540 41568
rect 51592 41556 51598 41608
rect 52178 41556 52184 41608
rect 52236 41596 52242 41608
rect 54036 41605 54064 41636
rect 54389 41633 54401 41636
rect 54435 41633 54447 41667
rect 54570 41664 54576 41676
rect 54483 41636 54576 41664
rect 54389 41627 54447 41633
rect 54570 41624 54576 41636
rect 54628 41664 54634 41676
rect 57146 41664 57152 41676
rect 54628 41636 57152 41664
rect 54628 41624 54634 41636
rect 57146 41624 57152 41636
rect 57204 41624 57210 41676
rect 59004 41673 59032 41704
rect 59357 41701 59369 41704
rect 59403 41701 59415 41735
rect 59357 41695 59415 41701
rect 58989 41667 59047 41673
rect 58989 41633 59001 41667
rect 59035 41633 59047 41667
rect 58989 41627 59047 41633
rect 54021 41599 54079 41605
rect 54021 41596 54033 41599
rect 52236 41568 54033 41596
rect 52236 41556 52242 41568
rect 54021 41565 54033 41568
rect 54067 41565 54079 41599
rect 54021 41559 54079 41565
rect 54941 41599 54999 41605
rect 54941 41565 54953 41599
rect 54987 41596 54999 41599
rect 59372 41596 59400 41695
rect 59538 41692 59544 41744
rect 59596 41732 59602 41744
rect 60185 41735 60243 41741
rect 60185 41732 60197 41735
rect 59596 41704 60197 41732
rect 59596 41692 59602 41704
rect 60185 41701 60197 41704
rect 60231 41701 60243 41735
rect 60185 41695 60243 41701
rect 59630 41624 59636 41676
rect 59688 41664 59694 41676
rect 60737 41667 60795 41673
rect 60737 41664 60749 41667
rect 59688 41636 60749 41664
rect 59688 41624 59694 41636
rect 60737 41633 60749 41636
rect 60783 41633 60795 41667
rect 61010 41664 61016 41676
rect 60971 41636 61016 41664
rect 60737 41627 60795 41633
rect 61010 41624 61016 41636
rect 61068 41624 61074 41676
rect 61212 41673 61240 41772
rect 63862 41760 63868 41772
rect 63920 41760 63926 41812
rect 69750 41732 69756 41744
rect 68664 41704 69756 41732
rect 68664 41676 68692 41704
rect 69750 41692 69756 41704
rect 69808 41692 69814 41744
rect 61197 41667 61255 41673
rect 61197 41633 61209 41667
rect 61243 41633 61255 41667
rect 62025 41667 62083 41673
rect 62025 41664 62037 41667
rect 61197 41627 61255 41633
rect 61856 41636 62037 41664
rect 60366 41596 60372 41608
rect 54987 41568 55536 41596
rect 59372 41568 60372 41596
rect 54987 41565 54999 41568
rect 54941 41559 54999 41565
rect 44600 41500 44772 41528
rect 44600 41488 44606 41500
rect 50614 41488 50620 41540
rect 50672 41528 50678 41540
rect 55033 41531 55091 41537
rect 55033 41528 55045 41531
rect 50672 41500 55045 41528
rect 50672 41488 50678 41500
rect 55033 41497 55045 41500
rect 55079 41497 55091 41531
rect 55033 41491 55091 41497
rect 55508 41472 55536 41568
rect 60366 41556 60372 41568
rect 60424 41596 60430 41608
rect 61856 41605 61884 41636
rect 62025 41633 62037 41636
rect 62071 41633 62083 41667
rect 63586 41664 63592 41676
rect 63547 41636 63592 41664
rect 62025 41627 62083 41633
rect 63586 41624 63592 41636
rect 63644 41624 63650 41676
rect 63773 41667 63831 41673
rect 63773 41633 63785 41667
rect 63819 41633 63831 41667
rect 63773 41627 63831 41633
rect 61841 41599 61899 41605
rect 61841 41596 61853 41599
rect 60424 41568 61853 41596
rect 60424 41556 60430 41568
rect 61841 41565 61853 41568
rect 61887 41565 61899 41599
rect 61841 41559 61899 41565
rect 62393 41599 62451 41605
rect 62393 41565 62405 41599
rect 62439 41596 62451 41599
rect 62574 41596 62580 41608
rect 62439 41568 62580 41596
rect 62439 41565 62451 41568
rect 62393 41559 62451 41565
rect 62574 41556 62580 41568
rect 62632 41556 62638 41608
rect 62022 41488 62028 41540
rect 62080 41528 62086 41540
rect 62163 41531 62221 41537
rect 62163 41528 62175 41531
rect 62080 41500 62175 41528
rect 62080 41488 62086 41500
rect 62163 41497 62175 41500
rect 62209 41497 62221 41531
rect 62163 41491 62221 41497
rect 62301 41531 62359 41537
rect 62301 41497 62313 41531
rect 62347 41528 62359 41531
rect 63788 41528 63816 41627
rect 65702 41624 65708 41676
rect 65760 41664 65766 41676
rect 65797 41667 65855 41673
rect 65797 41664 65809 41667
rect 65760 41636 65809 41664
rect 65760 41624 65766 41636
rect 65797 41633 65809 41636
rect 65843 41664 65855 41667
rect 66165 41667 66223 41673
rect 66165 41664 66177 41667
rect 65843 41636 66177 41664
rect 65843 41633 65855 41636
rect 65797 41627 65855 41633
rect 66165 41633 66177 41636
rect 66211 41633 66223 41667
rect 66990 41664 66996 41676
rect 66951 41636 66996 41664
rect 66165 41627 66223 41633
rect 66180 41596 66208 41627
rect 66990 41624 66996 41636
rect 67048 41624 67054 41676
rect 68465 41667 68523 41673
rect 68465 41633 68477 41667
rect 68511 41633 68523 41667
rect 68646 41664 68652 41676
rect 68559 41636 68652 41664
rect 68465 41627 68523 41633
rect 67085 41599 67143 41605
rect 67085 41596 67097 41599
rect 66180 41568 67097 41596
rect 67085 41565 67097 41568
rect 67131 41596 67143 41599
rect 68094 41596 68100 41608
rect 67131 41568 68100 41596
rect 67131 41565 67143 41568
rect 67085 41559 67143 41565
rect 68094 41556 68100 41568
rect 68152 41556 68158 41608
rect 68480 41596 68508 41627
rect 68646 41624 68652 41636
rect 68704 41624 68710 41676
rect 69017 41667 69075 41673
rect 69017 41633 69029 41667
rect 69063 41664 69075 41667
rect 69198 41664 69204 41676
rect 69063 41636 69204 41664
rect 69063 41633 69075 41636
rect 69017 41627 69075 41633
rect 69198 41624 69204 41636
rect 69256 41624 69262 41676
rect 69842 41664 69848 41676
rect 69803 41636 69848 41664
rect 69842 41624 69848 41636
rect 69900 41624 69906 41676
rect 70026 41664 70032 41676
rect 69987 41636 70032 41664
rect 70026 41624 70032 41636
rect 70084 41624 70090 41676
rect 71406 41664 71412 41676
rect 71367 41636 71412 41664
rect 71406 41624 71412 41636
rect 71464 41624 71470 41676
rect 70302 41596 70308 41608
rect 68480 41568 70308 41596
rect 70302 41556 70308 41568
rect 70360 41556 70366 41608
rect 77941 41599 77999 41605
rect 77941 41565 77953 41599
rect 77987 41565 77999 41599
rect 78214 41596 78220 41608
rect 78175 41568 78220 41596
rect 77941 41559 77999 41565
rect 64506 41528 64512 41540
rect 62347 41500 64512 41528
rect 62347 41497 62359 41500
rect 62301 41491 62359 41497
rect 64506 41488 64512 41500
rect 64564 41488 64570 41540
rect 77956 41472 77984 41559
rect 78214 41556 78220 41568
rect 78272 41556 78278 41608
rect 38160 41432 39344 41460
rect 38160 41420 38166 41432
rect 45002 41420 45008 41472
rect 45060 41460 45066 41472
rect 46109 41463 46167 41469
rect 46109 41460 46121 41463
rect 45060 41432 46121 41460
rect 45060 41420 45066 41432
rect 46109 41429 46121 41432
rect 46155 41429 46167 41463
rect 46109 41423 46167 41429
rect 46750 41420 46756 41472
rect 46808 41460 46814 41472
rect 52178 41460 52184 41472
rect 46808 41432 52184 41460
rect 46808 41420 46814 41432
rect 52178 41420 52184 41432
rect 52236 41420 52242 41472
rect 52546 41420 52552 41472
rect 52604 41460 52610 41472
rect 53193 41463 53251 41469
rect 53193 41460 53205 41463
rect 52604 41432 53205 41460
rect 52604 41420 52610 41432
rect 53193 41429 53205 41432
rect 53239 41429 53251 41463
rect 53193 41423 53251 41429
rect 54662 41420 54668 41472
rect 54720 41469 54726 41472
rect 54720 41463 54769 41469
rect 54720 41429 54723 41463
rect 54757 41429 54769 41463
rect 54720 41423 54769 41429
rect 54849 41463 54907 41469
rect 54849 41429 54861 41463
rect 54895 41460 54907 41463
rect 55398 41460 55404 41472
rect 54895 41432 55404 41460
rect 54895 41429 54907 41432
rect 54849 41423 54907 41429
rect 54720 41420 54726 41423
rect 55398 41420 55404 41432
rect 55456 41420 55462 41472
rect 55490 41420 55496 41472
rect 55548 41460 55554 41472
rect 62669 41463 62727 41469
rect 55548 41432 55593 41460
rect 55548 41420 55554 41432
rect 62669 41429 62681 41463
rect 62715 41460 62727 41463
rect 63034 41460 63040 41472
rect 62715 41432 63040 41460
rect 62715 41429 62727 41432
rect 62669 41423 62727 41429
rect 63034 41420 63040 41432
rect 63092 41420 63098 41472
rect 65978 41460 65984 41472
rect 65939 41432 65984 41460
rect 65978 41420 65984 41432
rect 66036 41420 66042 41472
rect 69014 41420 69020 41472
rect 69072 41460 69078 41472
rect 70026 41460 70032 41472
rect 69072 41432 70032 41460
rect 69072 41420 69078 41432
rect 70026 41420 70032 41432
rect 70084 41420 70090 41472
rect 71590 41460 71596 41472
rect 71551 41432 71596 41460
rect 71590 41420 71596 41432
rect 71648 41420 71654 41472
rect 72510 41420 72516 41472
rect 72568 41460 72574 41472
rect 77849 41463 77907 41469
rect 77849 41460 77861 41463
rect 72568 41432 77861 41460
rect 72568 41420 72574 41432
rect 77849 41429 77861 41432
rect 77895 41460 77907 41463
rect 77938 41460 77944 41472
rect 77895 41432 77944 41460
rect 77895 41429 77907 41432
rect 77849 41423 77907 41429
rect 77938 41420 77944 41432
rect 77996 41420 78002 41472
rect 79505 41463 79563 41469
rect 79505 41429 79517 41463
rect 79551 41460 79563 41463
rect 79778 41460 79784 41472
rect 79551 41432 79784 41460
rect 79551 41429 79563 41432
rect 79505 41423 79563 41429
rect 79778 41420 79784 41432
rect 79836 41420 79842 41472
rect 1104 41370 111136 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 65686 41370
rect 65738 41318 65750 41370
rect 65802 41318 65814 41370
rect 65866 41318 65878 41370
rect 65930 41318 96406 41370
rect 96458 41318 96470 41370
rect 96522 41318 96534 41370
rect 96586 41318 96598 41370
rect 96650 41318 111136 41370
rect 1104 41296 111136 41318
rect 10226 41256 10232 41268
rect 10187 41228 10232 41256
rect 10226 41216 10232 41228
rect 10284 41216 10290 41268
rect 10781 41259 10839 41265
rect 10781 41225 10793 41259
rect 10827 41256 10839 41259
rect 13078 41256 13084 41268
rect 10827 41228 13084 41256
rect 10827 41225 10839 41228
rect 10781 41219 10839 41225
rect 3145 41123 3203 41129
rect 3145 41089 3157 41123
rect 3191 41120 3203 41123
rect 9585 41123 9643 41129
rect 3191 41092 3556 41120
rect 3191 41089 3203 41092
rect 3145 41083 3203 41089
rect 3528 41061 3556 41092
rect 9585 41089 9597 41123
rect 9631 41089 9643 41123
rect 9585 41083 9643 41089
rect 3421 41055 3479 41061
rect 3421 41021 3433 41055
rect 3467 41021 3479 41055
rect 3421 41015 3479 41021
rect 3513 41055 3571 41061
rect 3513 41021 3525 41055
rect 3559 41052 3571 41055
rect 3602 41052 3608 41064
rect 3559 41024 3608 41052
rect 3559 41021 3571 41024
rect 3513 41015 3571 41021
rect 3436 40984 3464 41015
rect 3602 41012 3608 41024
rect 3660 41012 3666 41064
rect 3878 41052 3884 41064
rect 3839 41024 3884 41052
rect 3878 41012 3884 41024
rect 3936 41012 3942 41064
rect 3973 41055 4031 41061
rect 3973 41021 3985 41055
rect 4019 41052 4031 41055
rect 5442 41052 5448 41064
rect 4019 41024 5028 41052
rect 5403 41024 5448 41052
rect 4019 41021 4031 41024
rect 3973 41015 4031 41021
rect 3988 40984 4016 41015
rect 3436 40956 4016 40984
rect 4525 40987 4583 40993
rect 4525 40953 4537 40987
rect 4571 40984 4583 40987
rect 4614 40984 4620 40996
rect 4571 40956 4620 40984
rect 4571 40953 4583 40956
rect 4525 40947 4583 40953
rect 4614 40944 4620 40956
rect 4672 40944 4678 40996
rect 5000 40993 5028 41024
rect 5442 41012 5448 41024
rect 5500 41012 5506 41064
rect 8294 41012 8300 41064
rect 8352 41052 8358 41064
rect 9122 41052 9128 41064
rect 8352 41024 9128 41052
rect 8352 41012 8358 41024
rect 9122 41012 9128 41024
rect 9180 41052 9186 41064
rect 9493 41055 9551 41061
rect 9493 41052 9505 41055
rect 9180 41024 9505 41052
rect 9180 41012 9186 41024
rect 9493 41021 9505 41024
rect 9539 41021 9551 41055
rect 9493 41015 9551 41021
rect 4985 40987 5043 40993
rect 4985 40953 4997 40987
rect 5031 40984 5043 40987
rect 5169 40987 5227 40993
rect 5169 40984 5181 40987
rect 5031 40956 5181 40984
rect 5031 40953 5043 40956
rect 4985 40947 5043 40953
rect 5169 40953 5181 40956
rect 5215 40984 5227 40987
rect 7282 40984 7288 40996
rect 5215 40956 7288 40984
rect 5215 40953 5227 40956
rect 5169 40947 5227 40953
rect 7282 40944 7288 40956
rect 7340 40944 7346 40996
rect 8846 40984 8852 40996
rect 8807 40956 8852 40984
rect 8846 40944 8852 40956
rect 8904 40944 8910 40996
rect 3878 40876 3884 40928
rect 3936 40916 3942 40928
rect 4801 40919 4859 40925
rect 4801 40916 4813 40919
rect 3936 40888 4813 40916
rect 3936 40876 3942 40888
rect 4801 40885 4813 40888
rect 4847 40916 4859 40919
rect 5537 40919 5595 40925
rect 5537 40916 5549 40919
rect 4847 40888 5549 40916
rect 4847 40885 4859 40888
rect 4801 40879 4859 40885
rect 5537 40885 5549 40888
rect 5583 40916 5595 40919
rect 8018 40916 8024 40928
rect 5583 40888 8024 40916
rect 5583 40885 5595 40888
rect 5537 40879 5595 40885
rect 8018 40876 8024 40888
rect 8076 40876 8082 40928
rect 9508 40916 9536 41015
rect 9600 40984 9628 41083
rect 9861 41055 9919 41061
rect 9861 41021 9873 41055
rect 9907 41052 9919 41055
rect 9950 41052 9956 41064
rect 9907 41024 9956 41052
rect 9907 41021 9919 41024
rect 9861 41015 9919 41021
rect 9950 41012 9956 41024
rect 10008 41012 10014 41064
rect 10045 41055 10103 41061
rect 10045 41021 10057 41055
rect 10091 41052 10103 41055
rect 10244 41052 10272 41216
rect 10413 41191 10471 41197
rect 10413 41157 10425 41191
rect 10459 41188 10471 41191
rect 10962 41188 10968 41200
rect 10459 41160 10968 41188
rect 10459 41157 10471 41160
rect 10413 41151 10471 41157
rect 10428 41052 10456 41151
rect 10962 41148 10968 41160
rect 11020 41148 11026 41200
rect 10091 41024 10272 41052
rect 10336 41024 10456 41052
rect 10091 41021 10103 41024
rect 10045 41015 10103 41021
rect 10336 40984 10364 41024
rect 11072 40984 11100 41228
rect 13078 41216 13084 41228
rect 13136 41256 13142 41268
rect 15194 41256 15200 41268
rect 13136 41228 15200 41256
rect 13136 41216 13142 41228
rect 15194 41216 15200 41228
rect 15252 41216 15258 41268
rect 17494 41216 17500 41268
rect 17552 41256 17558 41268
rect 18230 41256 18236 41268
rect 17552 41228 18236 41256
rect 17552 41216 17558 41228
rect 18230 41216 18236 41228
rect 18288 41216 18294 41268
rect 18506 41216 18512 41268
rect 18564 41256 18570 41268
rect 19337 41259 19395 41265
rect 19337 41256 19349 41259
rect 18564 41228 19349 41256
rect 18564 41216 18570 41228
rect 19337 41225 19349 41228
rect 19383 41225 19395 41259
rect 19337 41219 19395 41225
rect 23382 41216 23388 41268
rect 23440 41256 23446 41268
rect 23753 41259 23811 41265
rect 23753 41256 23765 41259
rect 23440 41228 23765 41256
rect 23440 41216 23446 41228
rect 23753 41225 23765 41228
rect 23799 41225 23811 41259
rect 23753 41219 23811 41225
rect 17954 41148 17960 41200
rect 18012 41188 18018 41200
rect 18524 41188 18552 41216
rect 18012 41160 18552 41188
rect 23768 41188 23796 41219
rect 23934 41216 23940 41268
rect 23992 41256 23998 41268
rect 29822 41256 29828 41268
rect 23992 41228 29828 41256
rect 23992 41216 23998 41228
rect 29822 41216 29828 41228
rect 29880 41216 29886 41268
rect 31570 41256 31576 41268
rect 29932 41228 31576 41256
rect 23768 41160 24072 41188
rect 18012 41148 18018 41160
rect 12437 41123 12495 41129
rect 12437 41089 12449 41123
rect 12483 41120 12495 41123
rect 12802 41120 12808 41132
rect 12483 41092 12808 41120
rect 12483 41089 12495 41092
rect 12437 41083 12495 41089
rect 12802 41080 12808 41092
rect 12860 41120 12866 41132
rect 24044 41120 24072 41160
rect 26234 41148 26240 41200
rect 26292 41188 26298 41200
rect 27249 41191 27307 41197
rect 27249 41188 27261 41191
rect 26292 41160 27261 41188
rect 26292 41148 26298 41160
rect 27249 41157 27261 41160
rect 27295 41157 27307 41191
rect 27525 41191 27583 41197
rect 27525 41188 27537 41191
rect 27249 41151 27307 41157
rect 27448 41160 27537 41188
rect 12860 41092 14320 41120
rect 24044 41092 24256 41120
rect 12860 41080 12866 41092
rect 12710 41052 12716 41064
rect 12671 41024 12716 41052
rect 12710 41012 12716 41024
rect 12768 41012 12774 41064
rect 9600 40956 10364 40984
rect 10428 40956 11100 40984
rect 10428 40916 10456 40956
rect 9508 40888 10456 40916
rect 10502 40876 10508 40928
rect 10560 40916 10566 40928
rect 13630 40916 13636 40928
rect 10560 40888 13636 40916
rect 10560 40876 10566 40888
rect 13630 40876 13636 40888
rect 13688 40876 13694 40928
rect 13998 40916 14004 40928
rect 13959 40888 14004 40916
rect 13998 40876 14004 40888
rect 14056 40876 14062 40928
rect 14292 40925 14320 41092
rect 16942 41012 16948 41064
rect 17000 41052 17006 41064
rect 18049 41055 18107 41061
rect 18049 41052 18061 41055
rect 17000 41024 18061 41052
rect 17000 41012 17006 41024
rect 18049 41021 18061 41024
rect 18095 41052 18107 41055
rect 18417 41055 18475 41061
rect 18417 41052 18429 41055
rect 18095 41024 18429 41052
rect 18095 41021 18107 41024
rect 18049 41015 18107 41021
rect 18417 41021 18429 41024
rect 18463 41021 18475 41055
rect 18417 41015 18475 41021
rect 19153 41055 19211 41061
rect 19153 41021 19165 41055
rect 19199 41052 19211 41055
rect 19521 41055 19579 41061
rect 19521 41052 19533 41055
rect 19199 41024 19533 41052
rect 19199 41021 19211 41024
rect 19153 41015 19211 41021
rect 19521 41021 19533 41024
rect 19567 41052 19579 41055
rect 20898 41052 20904 41064
rect 19567 41024 20904 41052
rect 19567 41021 19579 41024
rect 19521 41015 19579 41021
rect 20898 41012 20904 41024
rect 20956 41012 20962 41064
rect 23658 41012 23664 41064
rect 23716 41052 23722 41064
rect 23937 41055 23995 41061
rect 23937 41052 23949 41055
rect 23716 41024 23949 41052
rect 23716 41012 23722 41024
rect 23937 41021 23949 41024
rect 23983 41021 23995 41055
rect 24118 41052 24124 41064
rect 24079 41024 24124 41052
rect 23937 41015 23995 41021
rect 24118 41012 24124 41024
rect 24176 41012 24182 41064
rect 24228 41052 24256 41092
rect 25498 41080 25504 41132
rect 25556 41120 25562 41132
rect 25685 41123 25743 41129
rect 25685 41120 25697 41123
rect 25556 41092 25697 41120
rect 25556 41080 25562 41092
rect 25685 41089 25697 41092
rect 25731 41120 25743 41123
rect 27338 41120 27344 41132
rect 25731 41092 27344 41120
rect 25731 41089 25743 41092
rect 25685 41083 25743 41089
rect 27338 41080 27344 41092
rect 27396 41080 27402 41132
rect 24581 41055 24639 41061
rect 24581 41052 24593 41055
rect 24228 41024 24593 41052
rect 24581 41021 24593 41024
rect 24627 41021 24639 41055
rect 24581 41015 24639 41021
rect 24670 41012 24676 41064
rect 24728 41052 24734 41064
rect 25516 41052 25544 41080
rect 24728 41024 25544 41052
rect 24728 41012 24734 41024
rect 26234 41012 26240 41064
rect 26292 41052 26298 41064
rect 27448 41061 27476 41160
rect 27525 41157 27537 41160
rect 27571 41188 27583 41191
rect 29932 41188 29960 41228
rect 31570 41216 31576 41228
rect 31628 41216 31634 41268
rect 31665 41259 31723 41265
rect 31665 41225 31677 41259
rect 31711 41256 31723 41259
rect 44634 41256 44640 41268
rect 31711 41228 44640 41256
rect 31711 41225 31723 41228
rect 31665 41219 31723 41225
rect 31680 41188 31708 41219
rect 44634 41216 44640 41228
rect 44692 41216 44698 41268
rect 44726 41216 44732 41268
rect 44784 41256 44790 41268
rect 44913 41259 44971 41265
rect 44913 41256 44925 41259
rect 44784 41228 44925 41256
rect 44784 41216 44790 41228
rect 44913 41225 44925 41228
rect 44959 41256 44971 41259
rect 45462 41256 45468 41268
rect 44959 41228 45468 41256
rect 44959 41225 44971 41228
rect 44913 41219 44971 41225
rect 45462 41216 45468 41228
rect 45520 41216 45526 41268
rect 51810 41216 51816 41268
rect 51868 41256 51874 41268
rect 51997 41259 52055 41265
rect 51997 41256 52009 41259
rect 51868 41228 52009 41256
rect 51868 41216 51874 41228
rect 51997 41225 52009 41228
rect 52043 41225 52055 41259
rect 51997 41219 52055 41225
rect 53098 41216 53104 41268
rect 53156 41256 53162 41268
rect 54570 41256 54576 41268
rect 53156 41228 54576 41256
rect 53156 41216 53162 41228
rect 54570 41216 54576 41228
rect 54628 41216 54634 41268
rect 63494 41216 63500 41268
rect 63552 41256 63558 41268
rect 63865 41259 63923 41265
rect 63865 41256 63877 41259
rect 63552 41228 63877 41256
rect 63552 41216 63558 41228
rect 63865 41225 63877 41228
rect 63911 41256 63923 41259
rect 64690 41256 64696 41268
rect 63911 41228 64696 41256
rect 63911 41225 63923 41228
rect 63865 41219 63923 41225
rect 64690 41216 64696 41228
rect 64748 41216 64754 41268
rect 68094 41256 68100 41268
rect 68055 41228 68100 41256
rect 68094 41216 68100 41228
rect 68152 41216 68158 41268
rect 68646 41216 68652 41268
rect 68704 41265 68710 41268
rect 68704 41259 68753 41265
rect 68704 41225 68707 41259
rect 68741 41225 68753 41259
rect 68704 41219 68753 41225
rect 68833 41259 68891 41265
rect 68833 41225 68845 41259
rect 68879 41256 68891 41259
rect 69014 41256 69020 41268
rect 68879 41228 69020 41256
rect 68879 41225 68891 41228
rect 68833 41219 68891 41225
rect 68704 41216 68710 41219
rect 69014 41216 69020 41228
rect 69072 41216 69078 41268
rect 69216 41228 77708 41256
rect 27571 41160 29960 41188
rect 30024 41160 31708 41188
rect 27571 41157 27583 41160
rect 27525 41151 27583 41157
rect 27614 41080 27620 41132
rect 27672 41120 27678 41132
rect 30024 41120 30052 41160
rect 27672 41092 30052 41120
rect 30101 41123 30159 41129
rect 27672 41080 27678 41092
rect 30101 41089 30113 41123
rect 30147 41089 30159 41123
rect 30101 41083 30159 41089
rect 26329 41055 26387 41061
rect 26329 41052 26341 41055
rect 26292 41024 26341 41052
rect 26292 41012 26298 41024
rect 26329 41021 26341 41024
rect 26375 41021 26387 41055
rect 26329 41015 26387 41021
rect 27433 41055 27491 41061
rect 27433 41021 27445 41055
rect 27479 41021 27491 41055
rect 27433 41015 27491 41021
rect 30006 40984 30012 40996
rect 22112 40956 30012 40984
rect 14277 40919 14335 40925
rect 14277 40885 14289 40919
rect 14323 40916 14335 40919
rect 16390 40916 16396 40928
rect 14323 40888 16396 40916
rect 14323 40885 14335 40888
rect 14277 40879 14335 40885
rect 16390 40876 16396 40888
rect 16448 40876 16454 40928
rect 21726 40876 21732 40928
rect 21784 40916 21790 40928
rect 22112 40916 22140 40956
rect 30006 40944 30012 40956
rect 30064 40984 30070 40996
rect 30116 40984 30144 41083
rect 30193 41055 30251 41061
rect 30193 41021 30205 41055
rect 30239 41021 30251 41055
rect 30650 41052 30656 41064
rect 30611 41024 30656 41052
rect 30193 41015 30251 41021
rect 30064 40956 30144 40984
rect 30064 40944 30070 40956
rect 21784 40888 22140 40916
rect 21784 40876 21790 40888
rect 24118 40876 24124 40928
rect 24176 40916 24182 40928
rect 24578 40916 24584 40928
rect 24176 40888 24584 40916
rect 24176 40876 24182 40888
rect 24578 40876 24584 40888
rect 24636 40876 24642 40928
rect 25133 40919 25191 40925
rect 25133 40885 25145 40919
rect 25179 40916 25191 40919
rect 25222 40916 25228 40928
rect 25179 40888 25228 40916
rect 25179 40885 25191 40888
rect 25133 40879 25191 40885
rect 25222 40876 25228 40888
rect 25280 40876 25286 40928
rect 25501 40919 25559 40925
rect 25501 40885 25513 40919
rect 25547 40916 25559 40919
rect 25682 40916 25688 40928
rect 25547 40888 25688 40916
rect 25547 40885 25559 40888
rect 25501 40879 25559 40885
rect 25682 40876 25688 40888
rect 25740 40876 25746 40928
rect 25866 40876 25872 40928
rect 25924 40916 25930 40928
rect 26145 40919 26203 40925
rect 26145 40916 26157 40919
rect 25924 40888 26157 40916
rect 25924 40876 25930 40888
rect 26145 40885 26157 40888
rect 26191 40885 26203 40919
rect 30208 40916 30236 41015
rect 30650 41012 30656 41024
rect 30708 41012 30714 41064
rect 30745 41055 30803 41061
rect 30745 41021 30757 41055
rect 30791 41052 30803 41055
rect 31128 41052 31156 41160
rect 36170 41148 36176 41200
rect 36228 41188 36234 41200
rect 38381 41191 38439 41197
rect 38381 41188 38393 41191
rect 36228 41160 38393 41188
rect 36228 41148 36234 41160
rect 38381 41157 38393 41160
rect 38427 41157 38439 41191
rect 38381 41151 38439 41157
rect 38562 41148 38568 41200
rect 38620 41188 38626 41200
rect 60642 41188 60648 41200
rect 38620 41160 60648 41188
rect 38620 41148 38626 41160
rect 60642 41148 60648 41160
rect 60700 41148 60706 41200
rect 60829 41191 60887 41197
rect 60829 41157 60841 41191
rect 60875 41188 60887 41191
rect 62022 41188 62028 41200
rect 60875 41160 62028 41188
rect 60875 41157 60887 41160
rect 60829 41151 60887 41157
rect 62022 41148 62028 41160
rect 62080 41148 62086 41200
rect 63034 41188 63040 41200
rect 62995 41160 63040 41188
rect 63034 41148 63040 41160
rect 63092 41148 63098 41200
rect 63126 41148 63132 41200
rect 63184 41188 63190 41200
rect 69216 41188 69244 41228
rect 71225 41191 71283 41197
rect 71225 41188 71237 41191
rect 63184 41160 69244 41188
rect 70964 41160 71237 41188
rect 63184 41148 63190 41160
rect 34790 41080 34796 41132
rect 34848 41120 34854 41132
rect 35897 41123 35955 41129
rect 35897 41120 35909 41123
rect 34848 41092 35909 41120
rect 34848 41080 34854 41092
rect 35897 41089 35909 41092
rect 35943 41089 35955 41123
rect 35897 41083 35955 41089
rect 35986 41080 35992 41132
rect 36044 41120 36050 41132
rect 37185 41123 37243 41129
rect 36044 41092 36124 41120
rect 36044 41080 36050 41092
rect 36096 41061 36124 41092
rect 37185 41089 37197 41123
rect 37231 41120 37243 41123
rect 38252 41123 38310 41129
rect 38252 41120 38264 41123
rect 37231 41092 38264 41120
rect 37231 41089 37243 41092
rect 37185 41083 37243 41089
rect 38252 41089 38264 41092
rect 38298 41089 38310 41123
rect 38470 41120 38476 41132
rect 38431 41092 38476 41120
rect 38252 41083 38310 41089
rect 38470 41080 38476 41092
rect 38528 41080 38534 41132
rect 38654 41120 38660 41132
rect 38580 41092 38660 41120
rect 36081 41055 36139 41061
rect 30791 41024 31156 41052
rect 31220 41024 36032 41052
rect 30791 41021 30803 41024
rect 30745 41015 30803 41021
rect 31220 40916 31248 41024
rect 31297 40987 31355 40993
rect 31297 40953 31309 40987
rect 31343 40984 31355 40987
rect 32674 40984 32680 40996
rect 31343 40956 32680 40984
rect 31343 40953 31355 40956
rect 31297 40947 31355 40953
rect 32674 40944 32680 40956
rect 32732 40944 32738 40996
rect 36004 40984 36032 41024
rect 36081 41021 36093 41055
rect 36127 41052 36139 41055
rect 36262 41052 36268 41064
rect 36127 41024 36268 41052
rect 36127 41021 36139 41024
rect 36081 41015 36139 41021
rect 36262 41012 36268 41024
rect 36320 41012 36326 41064
rect 36446 41012 36452 41064
rect 36504 41052 36510 41064
rect 36541 41055 36599 41061
rect 36541 41052 36553 41055
rect 36504 41024 36553 41052
rect 36504 41012 36510 41024
rect 36541 41021 36553 41024
rect 36587 41021 36599 41055
rect 36541 41015 36599 41021
rect 36630 41012 36636 41064
rect 36688 41052 36694 41064
rect 36688 41024 36733 41052
rect 36688 41012 36694 41024
rect 37734 41012 37740 41064
rect 37792 41052 37798 41064
rect 38105 41055 38163 41061
rect 38105 41052 38117 41055
rect 37792 41024 38117 41052
rect 37792 41012 37798 41024
rect 38105 41021 38117 41024
rect 38151 41021 38163 41055
rect 38105 41015 38163 41021
rect 38580 40984 38608 41092
rect 38654 41080 38660 41092
rect 38712 41080 38718 41132
rect 39022 41080 39028 41132
rect 39080 41120 39086 41132
rect 68925 41123 68983 41129
rect 39080 41092 68784 41120
rect 39080 41080 39086 41092
rect 43165 41055 43223 41061
rect 43165 41021 43177 41055
rect 43211 41052 43223 41055
rect 43714 41052 43720 41064
rect 43211 41024 43720 41052
rect 43211 41021 43223 41024
rect 43165 41015 43223 41021
rect 43714 41012 43720 41024
rect 43772 41012 43778 41064
rect 43806 41012 43812 41064
rect 43864 41052 43870 41064
rect 44818 41052 44824 41064
rect 43864 41024 44824 41052
rect 43864 41012 43870 41024
rect 44818 41012 44824 41024
rect 44876 41012 44882 41064
rect 52454 41012 52460 41064
rect 52512 41052 52518 41064
rect 52549 41055 52607 41061
rect 52549 41052 52561 41055
rect 52512 41024 52561 41052
rect 52512 41012 52518 41024
rect 52549 41021 52561 41024
rect 52595 41021 52607 41055
rect 52549 41015 52607 41021
rect 52641 41055 52699 41061
rect 52641 41021 52653 41055
rect 52687 41021 52699 41055
rect 52914 41052 52920 41064
rect 52875 41024 52920 41052
rect 52641 41015 52699 41021
rect 36004 40956 38608 40984
rect 38841 40987 38899 40993
rect 38841 40953 38853 40987
rect 38887 40984 38899 40987
rect 39942 40984 39948 40996
rect 38887 40956 39948 40984
rect 38887 40953 38899 40956
rect 38841 40947 38899 40953
rect 39942 40944 39948 40956
rect 40000 40944 40006 40996
rect 40034 40944 40040 40996
rect 40092 40984 40098 40996
rect 42886 40984 42892 40996
rect 40092 40956 42892 40984
rect 40092 40944 40098 40956
rect 42886 40944 42892 40956
rect 42944 40944 42950 40996
rect 44637 40987 44695 40993
rect 44637 40953 44649 40987
rect 44683 40984 44695 40987
rect 45094 40984 45100 40996
rect 44683 40956 45100 40984
rect 44683 40953 44695 40956
rect 44637 40947 44695 40953
rect 45094 40944 45100 40956
rect 45152 40944 45158 40996
rect 49418 40944 49424 40996
rect 49476 40984 49482 40996
rect 52656 40984 52684 41015
rect 52914 41012 52920 41024
rect 52972 41012 52978 41064
rect 53098 41052 53104 41064
rect 53059 41024 53104 41052
rect 53098 41012 53104 41024
rect 53156 41012 53162 41064
rect 54113 41055 54171 41061
rect 54113 41052 54125 41055
rect 53208 41024 54125 41052
rect 49476 40956 52684 40984
rect 52932 40984 52960 41012
rect 53208 40984 53236 41024
rect 54113 41021 54125 41024
rect 54159 41021 54171 41055
rect 54478 41052 54484 41064
rect 54439 41024 54484 41052
rect 54113 41015 54171 41021
rect 54478 41012 54484 41024
rect 54536 41012 54542 41064
rect 55490 41052 55496 41064
rect 55403 41024 55496 41052
rect 55490 41012 55496 41024
rect 55548 41012 55554 41064
rect 60737 41055 60795 41061
rect 60737 41021 60749 41055
rect 60783 41052 60795 41055
rect 60826 41052 60832 41064
rect 60783 41024 60832 41052
rect 60783 41021 60795 41024
rect 60737 41015 60795 41021
rect 60826 41012 60832 41024
rect 60884 41052 60890 41064
rect 61013 41055 61071 41061
rect 61013 41052 61025 41055
rect 60884 41024 61025 41052
rect 60884 41012 60890 41024
rect 61013 41021 61025 41024
rect 61059 41021 61071 41055
rect 61013 41015 61071 41021
rect 61562 41012 61568 41064
rect 61620 41052 61626 41064
rect 61749 41055 61807 41061
rect 61749 41052 61761 41055
rect 61620 41024 61761 41052
rect 61620 41012 61626 41024
rect 61749 41021 61761 41024
rect 61795 41021 61807 41055
rect 61749 41015 61807 41021
rect 62761 41055 62819 41061
rect 62761 41021 62773 41055
rect 62807 41052 62819 41055
rect 62945 41055 63003 41061
rect 62945 41052 62957 41055
rect 62807 41024 62957 41052
rect 62807 41021 62819 41024
rect 62761 41015 62819 41021
rect 62945 41021 62957 41024
rect 62991 41021 63003 41055
rect 62945 41015 63003 41021
rect 63034 41012 63040 41064
rect 63092 41052 63098 41064
rect 63221 41055 63279 41061
rect 63221 41052 63233 41055
rect 63092 41024 63233 41052
rect 63092 41012 63098 41024
rect 63221 41021 63233 41024
rect 63267 41052 63279 41055
rect 64230 41052 64236 41064
rect 63267 41024 64236 41052
rect 63267 41021 63279 41024
rect 63221 41015 63279 41021
rect 64230 41012 64236 41024
rect 64288 41012 64294 41064
rect 64693 41055 64751 41061
rect 64693 41052 64705 41055
rect 64340 41024 64705 41052
rect 52932 40956 53236 40984
rect 49476 40944 49482 40956
rect 31481 40919 31539 40925
rect 31481 40916 31493 40919
rect 30208 40888 31493 40916
rect 26145 40879 26203 40885
rect 31481 40885 31493 40888
rect 31527 40885 31539 40919
rect 31481 40879 31539 40885
rect 31570 40876 31576 40928
rect 31628 40916 31634 40928
rect 36538 40916 36544 40928
rect 31628 40888 36544 40916
rect 31628 40876 31634 40888
rect 36538 40876 36544 40888
rect 36596 40876 36602 40928
rect 36630 40876 36636 40928
rect 36688 40916 36694 40928
rect 37090 40916 37096 40928
rect 36688 40888 37096 40916
rect 36688 40876 36694 40888
rect 37090 40876 37096 40888
rect 37148 40916 37154 40928
rect 37461 40919 37519 40925
rect 37461 40916 37473 40919
rect 37148 40888 37473 40916
rect 37148 40876 37154 40888
rect 37461 40885 37473 40888
rect 37507 40916 37519 40919
rect 39022 40916 39028 40928
rect 37507 40888 39028 40916
rect 37507 40885 37519 40888
rect 37461 40879 37519 40885
rect 39022 40876 39028 40888
rect 39080 40876 39086 40928
rect 39114 40876 39120 40928
rect 39172 40916 39178 40928
rect 42794 40916 42800 40928
rect 39172 40888 42800 40916
rect 39172 40876 39178 40888
rect 42794 40876 42800 40888
rect 42852 40876 42858 40928
rect 42978 40876 42984 40928
rect 43036 40916 43042 40928
rect 43257 40919 43315 40925
rect 43257 40916 43269 40919
rect 43036 40888 43269 40916
rect 43036 40876 43042 40888
rect 43257 40885 43269 40888
rect 43303 40916 43315 40919
rect 43806 40916 43812 40928
rect 43303 40888 43812 40916
rect 43303 40885 43315 40888
rect 43257 40879 43315 40885
rect 43806 40876 43812 40888
rect 43864 40916 43870 40928
rect 44453 40919 44511 40925
rect 44453 40916 44465 40919
rect 43864 40888 44465 40916
rect 43864 40876 43870 40888
rect 44453 40885 44465 40888
rect 44499 40885 44511 40919
rect 52656 40916 52684 40956
rect 53466 40944 53472 40996
rect 53524 40984 53530 40996
rect 53929 40987 53987 40993
rect 53929 40984 53941 40987
rect 53524 40956 53941 40984
rect 53524 40944 53530 40956
rect 53929 40953 53941 40956
rect 53975 40953 53987 40987
rect 53929 40947 53987 40953
rect 55122 40944 55128 40996
rect 55180 40984 55186 40996
rect 55309 40987 55367 40993
rect 55309 40984 55321 40987
rect 55180 40956 55321 40984
rect 55180 40944 55186 40956
rect 55309 40953 55321 40956
rect 55355 40953 55367 40987
rect 55309 40947 55367 40953
rect 53285 40919 53343 40925
rect 53285 40916 53297 40919
rect 52656 40888 53297 40916
rect 44453 40879 44511 40885
rect 53285 40885 53297 40888
rect 53331 40916 53343 40919
rect 53374 40916 53380 40928
rect 53331 40888 53380 40916
rect 53331 40885 53343 40888
rect 53285 40879 53343 40885
rect 53374 40876 53380 40888
rect 53432 40876 53438 40928
rect 55508 40916 55536 41012
rect 55861 40987 55919 40993
rect 55861 40953 55873 40987
rect 55907 40984 55919 40987
rect 56594 40984 56600 40996
rect 55907 40956 56600 40984
rect 55907 40953 55919 40956
rect 55861 40947 55919 40953
rect 56594 40944 56600 40956
rect 56652 40984 56658 40996
rect 57054 40984 57060 40996
rect 56652 40956 57060 40984
rect 56652 40944 56658 40956
rect 57054 40944 57060 40956
rect 57112 40944 57118 40996
rect 57146 40944 57152 40996
rect 57204 40984 57210 40996
rect 57204 40956 63448 40984
rect 57204 40944 57210 40956
rect 55950 40916 55956 40928
rect 55508 40888 55956 40916
rect 55950 40876 55956 40888
rect 56008 40876 56014 40928
rect 61562 40916 61568 40928
rect 61523 40888 61568 40916
rect 61562 40876 61568 40888
rect 61620 40876 61626 40928
rect 61838 40916 61844 40928
rect 61799 40888 61844 40916
rect 61838 40876 61844 40888
rect 61896 40916 61902 40928
rect 62574 40916 62580 40928
rect 61896 40888 62580 40916
rect 61896 40876 61902 40888
rect 62574 40876 62580 40888
rect 62632 40876 62638 40928
rect 62761 40919 62819 40925
rect 62761 40885 62773 40919
rect 62807 40916 62819 40919
rect 63310 40916 63316 40928
rect 62807 40888 63316 40916
rect 62807 40885 62819 40888
rect 62761 40879 62819 40885
rect 63310 40876 63316 40888
rect 63368 40876 63374 40928
rect 63420 40925 63448 40956
rect 64340 40928 64368 41024
rect 64693 41021 64705 41024
rect 64739 41021 64751 41055
rect 64693 41015 64751 41021
rect 68094 41012 68100 41064
rect 68152 41052 68158 41064
rect 68557 41055 68615 41061
rect 68557 41052 68569 41055
rect 68152 41024 68569 41052
rect 68152 41012 68158 41024
rect 68557 41021 68569 41024
rect 68603 41021 68615 41055
rect 68756 41052 68784 41092
rect 68925 41089 68937 41123
rect 68971 41120 68983 41123
rect 69382 41120 69388 41132
rect 68971 41092 69388 41120
rect 68971 41089 68983 41092
rect 68925 41083 68983 41089
rect 69382 41080 69388 41092
rect 69440 41080 69446 41132
rect 70394 41080 70400 41132
rect 70452 41120 70458 41132
rect 70964 41120 70992 41160
rect 71225 41157 71237 41160
rect 71271 41188 71283 41191
rect 71682 41188 71688 41200
rect 71271 41160 71688 41188
rect 71271 41157 71283 41160
rect 71225 41151 71283 41157
rect 71682 41148 71688 41160
rect 71740 41148 71746 41200
rect 71130 41120 71136 41132
rect 70452 41092 70992 41120
rect 71091 41092 71136 41120
rect 70452 41080 70458 41092
rect 71130 41080 71136 41092
rect 71188 41080 71194 41132
rect 72421 41123 72479 41129
rect 72421 41120 72433 41123
rect 71424 41092 72433 41120
rect 70486 41052 70492 41064
rect 68756 41024 70492 41052
rect 68557 41015 68615 41021
rect 70486 41012 70492 41024
rect 70544 41012 70550 41064
rect 70673 41055 70731 41061
rect 70673 41021 70685 41055
rect 70719 41052 70731 41055
rect 71424 41052 71452 41092
rect 72421 41089 72433 41092
rect 72467 41089 72479 41123
rect 72421 41083 72479 41089
rect 77680 41120 77708 41228
rect 78122 41120 78128 41132
rect 77680 41092 78128 41120
rect 77680 41061 77708 41092
rect 78122 41080 78128 41092
rect 78180 41120 78186 41132
rect 78309 41123 78367 41129
rect 78309 41120 78321 41123
rect 78180 41092 78321 41120
rect 78180 41080 78186 41092
rect 78309 41089 78321 41092
rect 78355 41089 78367 41123
rect 78309 41083 78367 41089
rect 70719 41024 71452 41052
rect 72145 41055 72203 41061
rect 70719 41021 70731 41024
rect 70673 41015 70731 41021
rect 72145 41021 72157 41055
rect 72191 41021 72203 41055
rect 77113 41055 77171 41061
rect 77113 41052 77125 41055
rect 72145 41015 72203 41021
rect 76944 41024 77125 41052
rect 64414 40944 64420 40996
rect 64472 40984 64478 40996
rect 69293 40987 69351 40993
rect 69293 40984 69305 40987
rect 64472 40956 69305 40984
rect 64472 40944 64478 40956
rect 69293 40953 69305 40956
rect 69339 40953 69351 40987
rect 69293 40947 69351 40953
rect 70302 40944 70308 40996
rect 70360 40984 70366 40996
rect 70581 40987 70639 40993
rect 70581 40984 70593 40987
rect 70360 40956 70593 40984
rect 70360 40944 70366 40956
rect 70581 40953 70593 40956
rect 70627 40953 70639 40987
rect 71958 40984 71964 40996
rect 71919 40956 71964 40984
rect 70581 40947 70639 40953
rect 71958 40944 71964 40956
rect 72016 40944 72022 40996
rect 63405 40919 63463 40925
rect 63405 40885 63417 40919
rect 63451 40885 63463 40919
rect 64322 40916 64328 40928
rect 64283 40888 64328 40916
rect 63405 40879 63463 40885
rect 64322 40876 64328 40888
rect 64380 40876 64386 40928
rect 64509 40919 64567 40925
rect 64509 40885 64521 40919
rect 64555 40916 64567 40919
rect 66714 40916 66720 40928
rect 64555 40888 66720 40916
rect 64555 40885 64567 40888
rect 64509 40879 64567 40885
rect 66714 40876 66720 40888
rect 66772 40876 66778 40928
rect 68370 40916 68376 40928
rect 68331 40888 68376 40916
rect 68370 40876 68376 40888
rect 68428 40876 68434 40928
rect 69014 40876 69020 40928
rect 69072 40916 69078 40928
rect 71590 40916 71596 40928
rect 69072 40888 71596 40916
rect 69072 40876 69078 40888
rect 71590 40876 71596 40888
rect 71648 40916 71654 40928
rect 71777 40919 71835 40925
rect 71777 40916 71789 40919
rect 71648 40888 71789 40916
rect 71648 40876 71654 40888
rect 71777 40885 71789 40888
rect 71823 40916 71835 40919
rect 72160 40916 72188 41015
rect 71823 40888 72188 40916
rect 71823 40885 71835 40888
rect 71777 40879 71835 40885
rect 74258 40876 74264 40928
rect 74316 40916 74322 40928
rect 76834 40916 76840 40928
rect 74316 40888 76840 40916
rect 74316 40876 74322 40888
rect 76834 40876 76840 40888
rect 76892 40916 76898 40928
rect 76944 40925 76972 41024
rect 77113 41021 77125 41024
rect 77159 41021 77171 41055
rect 77113 41015 77171 41021
rect 77665 41055 77723 41061
rect 77665 41021 77677 41055
rect 77711 41021 77723 41055
rect 77665 41015 77723 41021
rect 77846 41012 77852 41064
rect 77904 41052 77910 41064
rect 77941 41055 77999 41061
rect 77941 41052 77953 41055
rect 77904 41024 77953 41052
rect 77904 41012 77910 41024
rect 77941 41021 77953 41024
rect 77987 41021 77999 41055
rect 79778 41052 79784 41064
rect 79739 41024 79784 41052
rect 77941 41015 77999 41021
rect 79778 41012 79784 41024
rect 79836 41012 79842 41064
rect 76929 40919 76987 40925
rect 76929 40916 76941 40919
rect 76892 40888 76941 40916
rect 76892 40876 76898 40888
rect 76929 40885 76941 40888
rect 76975 40885 76987 40919
rect 76929 40879 76987 40885
rect 77205 40919 77263 40925
rect 77205 40885 77217 40919
rect 77251 40916 77263 40919
rect 77570 40916 77576 40928
rect 77251 40888 77576 40916
rect 77251 40885 77263 40888
rect 77205 40879 77263 40885
rect 77570 40876 77576 40888
rect 77628 40876 77634 40928
rect 79870 40916 79876 40928
rect 79831 40888 79876 40916
rect 79870 40876 79876 40888
rect 79928 40876 79934 40928
rect 1104 40826 111136 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 50326 40826
rect 50378 40774 50390 40826
rect 50442 40774 50454 40826
rect 50506 40774 50518 40826
rect 50570 40774 81046 40826
rect 81098 40774 81110 40826
rect 81162 40774 81174 40826
rect 81226 40774 81238 40826
rect 81290 40774 111136 40826
rect 1104 40752 111136 40774
rect 9950 40672 9956 40724
rect 10008 40712 10014 40724
rect 10502 40712 10508 40724
rect 10008 40684 10508 40712
rect 10008 40672 10014 40684
rect 10502 40672 10508 40684
rect 10560 40672 10566 40724
rect 12713 40715 12771 40721
rect 12713 40712 12725 40715
rect 10888 40684 12725 40712
rect 4706 40536 4712 40588
rect 4764 40576 4770 40588
rect 10888 40585 10916 40684
rect 12713 40681 12725 40684
rect 12759 40712 12771 40715
rect 12802 40712 12808 40724
rect 12759 40684 12808 40712
rect 12759 40681 12771 40684
rect 12713 40675 12771 40681
rect 12802 40672 12808 40684
rect 12860 40672 12866 40724
rect 13725 40715 13783 40721
rect 13725 40681 13737 40715
rect 13771 40712 13783 40715
rect 13998 40712 14004 40724
rect 13771 40684 14004 40712
rect 13771 40681 13783 40684
rect 13725 40675 13783 40681
rect 4801 40579 4859 40585
rect 4801 40576 4813 40579
rect 4764 40548 4813 40576
rect 4764 40536 4770 40548
rect 4801 40545 4813 40548
rect 4847 40576 4859 40579
rect 6641 40579 6699 40585
rect 6641 40576 6653 40579
rect 4847 40548 6653 40576
rect 4847 40545 4859 40548
rect 4801 40539 4859 40545
rect 6641 40545 6653 40548
rect 6687 40576 6699 40579
rect 10873 40579 10931 40585
rect 10873 40576 10885 40579
rect 6687 40548 10885 40576
rect 6687 40545 6699 40548
rect 6641 40539 6699 40545
rect 10873 40545 10885 40548
rect 10919 40545 10931 40579
rect 10873 40539 10931 40545
rect 13357 40579 13415 40585
rect 13357 40545 13369 40579
rect 13403 40576 13415 40579
rect 13740 40576 13768 40675
rect 13998 40672 14004 40684
rect 14056 40712 14062 40724
rect 28626 40712 28632 40724
rect 14056 40684 28632 40712
rect 14056 40672 14062 40684
rect 28626 40672 28632 40684
rect 28684 40672 28690 40724
rect 36170 40712 36176 40724
rect 36131 40684 36176 40712
rect 36170 40672 36176 40684
rect 36228 40672 36234 40724
rect 36262 40672 36268 40724
rect 36320 40712 36326 40724
rect 38933 40715 38991 40721
rect 36320 40684 38424 40712
rect 36320 40672 36326 40684
rect 23658 40604 23664 40656
rect 23716 40644 23722 40656
rect 25682 40644 25688 40656
rect 23716 40616 24532 40644
rect 23716 40604 23722 40616
rect 13403 40548 13768 40576
rect 13403 40545 13415 40548
rect 13357 40539 13415 40545
rect 16482 40536 16488 40588
rect 16540 40576 16546 40588
rect 24504 40585 24532 40616
rect 25148 40616 25688 40644
rect 16945 40579 17003 40585
rect 16945 40576 16957 40579
rect 16540 40548 16957 40576
rect 16540 40536 16546 40548
rect 16945 40545 16957 40548
rect 16991 40545 17003 40579
rect 16945 40539 17003 40545
rect 24029 40579 24087 40585
rect 24029 40545 24041 40579
rect 24075 40576 24087 40579
rect 24489 40579 24547 40585
rect 24075 40548 24256 40576
rect 24075 40545 24087 40548
rect 24029 40539 24087 40545
rect 5077 40511 5135 40517
rect 5077 40477 5089 40511
rect 5123 40508 5135 40511
rect 5534 40508 5540 40520
rect 5123 40480 5540 40508
rect 5123 40477 5135 40480
rect 5077 40471 5135 40477
rect 5534 40468 5540 40480
rect 5592 40468 5598 40520
rect 11146 40508 11152 40520
rect 11107 40480 11152 40508
rect 11146 40468 11152 40480
rect 11204 40468 11210 40520
rect 12529 40511 12587 40517
rect 12529 40477 12541 40511
rect 12575 40508 12587 40511
rect 12894 40508 12900 40520
rect 12575 40480 12900 40508
rect 12575 40477 12587 40480
rect 12529 40471 12587 40477
rect 12894 40468 12900 40480
rect 12952 40468 12958 40520
rect 16390 40468 16396 40520
rect 16448 40508 16454 40520
rect 16669 40511 16727 40517
rect 16669 40508 16681 40511
rect 16448 40480 16681 40508
rect 16448 40468 16454 40480
rect 16669 40477 16681 40480
rect 16715 40508 16727 40511
rect 23845 40511 23903 40517
rect 16715 40480 18460 40508
rect 16715 40477 16727 40480
rect 16669 40471 16727 40477
rect 18432 40384 18460 40480
rect 23845 40477 23857 40511
rect 23891 40477 23903 40511
rect 23845 40471 23903 40477
rect 5718 40332 5724 40384
rect 5776 40372 5782 40384
rect 6181 40375 6239 40381
rect 6181 40372 6193 40375
rect 5776 40344 6193 40372
rect 5776 40332 5782 40344
rect 6181 40341 6193 40344
rect 6227 40341 6239 40375
rect 6181 40335 6239 40341
rect 12618 40332 12624 40384
rect 12676 40372 12682 40384
rect 13449 40375 13507 40381
rect 13449 40372 13461 40375
rect 12676 40344 13461 40372
rect 12676 40332 12682 40344
rect 13449 40341 13461 40344
rect 13495 40341 13507 40375
rect 18230 40372 18236 40384
rect 18191 40344 18236 40372
rect 13449 40335 13507 40341
rect 18230 40332 18236 40344
rect 18288 40332 18294 40384
rect 18414 40372 18420 40384
rect 18375 40344 18420 40372
rect 18414 40332 18420 40344
rect 18472 40332 18478 40384
rect 23753 40375 23811 40381
rect 23753 40341 23765 40375
rect 23799 40372 23811 40375
rect 23860 40372 23888 40471
rect 24228 40440 24256 40548
rect 24489 40545 24501 40579
rect 24535 40545 24547 40579
rect 24489 40539 24547 40545
rect 24578 40536 24584 40588
rect 24636 40576 24642 40588
rect 25148 40576 25176 40616
rect 25682 40604 25688 40616
rect 25740 40604 25746 40656
rect 27246 40604 27252 40656
rect 27304 40644 27310 40656
rect 27340 40647 27398 40653
rect 27340 40644 27352 40647
rect 27304 40616 27352 40644
rect 27304 40604 27310 40616
rect 27340 40613 27352 40616
rect 27386 40613 27398 40647
rect 27340 40607 27398 40613
rect 29089 40647 29147 40653
rect 29089 40613 29101 40647
rect 29135 40644 29147 40647
rect 34606 40644 34612 40656
rect 29135 40616 30144 40644
rect 34567 40616 34612 40644
rect 29135 40613 29147 40616
rect 29089 40607 29147 40613
rect 24636 40548 25176 40576
rect 24636 40536 24642 40548
rect 25222 40536 25228 40588
rect 25280 40576 25286 40588
rect 27488 40579 27546 40585
rect 27488 40576 27500 40579
rect 25280 40548 27500 40576
rect 25280 40536 25286 40548
rect 27488 40545 27500 40548
rect 27534 40545 27546 40579
rect 27488 40539 27546 40545
rect 27614 40536 27620 40588
rect 27672 40576 27678 40588
rect 29181 40579 29239 40585
rect 29181 40576 29193 40579
rect 27672 40548 29193 40576
rect 27672 40536 27678 40548
rect 29181 40545 29193 40548
rect 29227 40576 29239 40579
rect 29365 40579 29423 40585
rect 29365 40576 29377 40579
rect 29227 40548 29377 40576
rect 29227 40545 29239 40548
rect 29181 40539 29239 40545
rect 29365 40545 29377 40548
rect 29411 40545 29423 40579
rect 29365 40539 29423 40545
rect 29549 40579 29607 40585
rect 29549 40545 29561 40579
rect 29595 40576 29607 40579
rect 30006 40576 30012 40588
rect 29595 40548 29776 40576
rect 29967 40548 30012 40576
rect 29595 40545 29607 40548
rect 29549 40539 29607 40545
rect 25133 40511 25191 40517
rect 25133 40477 25145 40511
rect 25179 40508 25191 40511
rect 27709 40511 27767 40517
rect 27709 40508 27721 40511
rect 25179 40480 27721 40508
rect 25179 40477 25191 40480
rect 25133 40471 25191 40477
rect 27709 40477 27721 40480
rect 27755 40477 27767 40511
rect 27709 40471 27767 40477
rect 28077 40511 28135 40517
rect 28077 40477 28089 40511
rect 28123 40508 28135 40511
rect 28718 40508 28724 40520
rect 28123 40480 28724 40508
rect 28123 40477 28135 40480
rect 28077 40471 28135 40477
rect 28718 40468 28724 40480
rect 28776 40468 28782 40520
rect 28810 40468 28816 40520
rect 28868 40508 28874 40520
rect 28994 40508 29000 40520
rect 28868 40480 29000 40508
rect 28868 40468 28874 40480
rect 28994 40468 29000 40480
rect 29052 40468 29058 40520
rect 25409 40443 25467 40449
rect 24228 40412 25084 40440
rect 25056 40384 25084 40412
rect 25409 40409 25421 40443
rect 25455 40440 25467 40443
rect 25682 40440 25688 40452
rect 25455 40412 25688 40440
rect 25455 40409 25467 40412
rect 25409 40403 25467 40409
rect 25682 40400 25688 40412
rect 25740 40440 25746 40452
rect 29089 40443 29147 40449
rect 29089 40440 29101 40443
rect 25740 40412 29101 40440
rect 25740 40400 25746 40412
rect 29089 40409 29101 40412
rect 29135 40409 29147 40443
rect 29089 40403 29147 40409
rect 23934 40372 23940 40384
rect 23799 40344 23940 40372
rect 23799 40341 23811 40344
rect 23753 40335 23811 40341
rect 23934 40332 23940 40344
rect 23992 40332 23998 40384
rect 25038 40332 25044 40384
rect 25096 40372 25102 40384
rect 25593 40375 25651 40381
rect 25593 40372 25605 40375
rect 25096 40344 25605 40372
rect 25096 40332 25102 40344
rect 25593 40341 25605 40344
rect 25639 40372 25651 40375
rect 26602 40372 26608 40384
rect 25639 40344 26608 40372
rect 25639 40341 25651 40344
rect 25593 40335 25651 40341
rect 26602 40332 26608 40344
rect 26660 40332 26666 40384
rect 27617 40375 27675 40381
rect 27617 40341 27629 40375
rect 27663 40372 27675 40375
rect 28258 40372 28264 40384
rect 27663 40344 28264 40372
rect 27663 40341 27675 40344
rect 27617 40335 27675 40341
rect 28258 40332 28264 40344
rect 28316 40332 28322 40384
rect 28350 40332 28356 40384
rect 28408 40372 28414 40384
rect 29748 40372 29776 40548
rect 30006 40536 30012 40548
rect 30064 40536 30070 40588
rect 30116 40585 30144 40616
rect 34606 40604 34612 40616
rect 34664 40644 34670 40656
rect 34664 40616 35020 40644
rect 34664 40604 34670 40616
rect 34992 40585 35020 40616
rect 35084 40616 36124 40644
rect 30101 40579 30159 40585
rect 30101 40545 30113 40579
rect 30147 40576 30159 40579
rect 34977 40579 35035 40585
rect 30147 40548 30604 40576
rect 30147 40545 30159 40548
rect 30101 40539 30159 40545
rect 30576 40440 30604 40548
rect 34977 40545 34989 40579
rect 35023 40545 35035 40579
rect 34977 40539 35035 40545
rect 30653 40511 30711 40517
rect 30653 40477 30665 40511
rect 30699 40508 30711 40511
rect 32950 40508 32956 40520
rect 30699 40480 32956 40508
rect 30699 40477 30711 40480
rect 30653 40471 30711 40477
rect 32950 40468 32956 40480
rect 33008 40468 33014 40520
rect 35084 40508 35112 40616
rect 35161 40579 35219 40585
rect 35161 40545 35173 40579
rect 35207 40576 35219 40579
rect 35342 40576 35348 40588
rect 35207 40548 35348 40576
rect 35207 40545 35219 40548
rect 35161 40539 35219 40545
rect 35342 40536 35348 40548
rect 35400 40536 35406 40588
rect 35618 40576 35624 40588
rect 35579 40548 35624 40576
rect 35618 40536 35624 40548
rect 35676 40536 35682 40588
rect 35710 40536 35716 40588
rect 35768 40576 35774 40588
rect 35768 40548 35813 40576
rect 35768 40536 35774 40548
rect 33060 40480 35112 40508
rect 36096 40508 36124 40616
rect 36538 40604 36544 40656
rect 36596 40644 36602 40656
rect 37458 40644 37464 40656
rect 36596 40616 37464 40644
rect 36596 40604 36602 40616
rect 37458 40604 37464 40616
rect 37516 40644 37522 40656
rect 37918 40644 37924 40656
rect 37516 40616 37924 40644
rect 37516 40604 37522 40616
rect 37918 40604 37924 40616
rect 37976 40604 37982 40656
rect 38286 40644 38292 40656
rect 38247 40616 38292 40644
rect 38286 40604 38292 40616
rect 38344 40604 38350 40656
rect 38396 40644 38424 40684
rect 38933 40681 38945 40715
rect 38979 40712 38991 40715
rect 39114 40712 39120 40724
rect 38979 40684 39120 40712
rect 38979 40681 38991 40684
rect 38933 40675 38991 40681
rect 39114 40672 39120 40684
rect 39172 40672 39178 40724
rect 40144 40684 46244 40712
rect 40034 40644 40040 40656
rect 38396 40616 40040 40644
rect 40034 40604 40040 40616
rect 40092 40604 40098 40656
rect 36449 40579 36507 40585
rect 36449 40545 36461 40579
rect 36495 40576 36507 40579
rect 36630 40576 36636 40588
rect 36495 40548 36636 40576
rect 36495 40545 36507 40548
rect 36449 40539 36507 40545
rect 36630 40536 36636 40548
rect 36688 40576 36694 40588
rect 40144 40576 40172 40684
rect 41049 40647 41107 40653
rect 41049 40613 41061 40647
rect 41095 40644 41107 40647
rect 42610 40644 42616 40656
rect 41095 40616 42616 40644
rect 41095 40613 41107 40616
rect 41049 40607 41107 40613
rect 42610 40604 42616 40616
rect 42668 40604 42674 40656
rect 42886 40604 42892 40656
rect 42944 40644 42950 40656
rect 43530 40644 43536 40656
rect 42944 40616 43536 40644
rect 42944 40604 42950 40616
rect 43530 40604 43536 40616
rect 43588 40644 43594 40656
rect 43717 40647 43775 40653
rect 43717 40644 43729 40647
rect 43588 40616 43729 40644
rect 43588 40604 43594 40616
rect 43717 40613 43729 40616
rect 43763 40613 43775 40647
rect 43717 40607 43775 40613
rect 44450 40604 44456 40656
rect 44508 40644 44514 40656
rect 44821 40647 44879 40653
rect 44821 40644 44833 40647
rect 44508 40616 44833 40644
rect 44508 40604 44514 40616
rect 44821 40613 44833 40616
rect 44867 40644 44879 40647
rect 45186 40644 45192 40656
rect 44867 40616 45192 40644
rect 44867 40613 44879 40616
rect 44821 40607 44879 40613
rect 45186 40604 45192 40616
rect 45244 40604 45250 40656
rect 45370 40644 45376 40656
rect 45331 40616 45376 40644
rect 45370 40604 45376 40616
rect 45428 40604 45434 40656
rect 46216 40644 46244 40684
rect 46290 40672 46296 40724
rect 46348 40712 46354 40724
rect 72510 40712 72516 40724
rect 46348 40684 72372 40712
rect 72471 40684 72516 40712
rect 46348 40672 46354 40684
rect 55766 40644 55772 40656
rect 46216 40616 55772 40644
rect 55766 40604 55772 40616
rect 55824 40604 55830 40656
rect 57054 40644 57060 40656
rect 57015 40616 57060 40644
rect 57054 40604 57060 40616
rect 57112 40604 57118 40656
rect 60734 40604 60740 40656
rect 60792 40644 60798 40656
rect 62942 40644 62948 40656
rect 60792 40616 60837 40644
rect 62408 40616 62948 40644
rect 60792 40604 60798 40616
rect 36688 40548 40172 40576
rect 36688 40536 36694 40548
rect 41230 40536 41236 40588
rect 41288 40576 41294 40588
rect 41288 40548 41552 40576
rect 41288 40536 41294 40548
rect 38470 40508 38476 40520
rect 36096 40480 38476 40508
rect 30929 40443 30987 40449
rect 30929 40440 30941 40443
rect 30576 40412 30941 40440
rect 30929 40409 30941 40412
rect 30975 40440 30987 40443
rect 33060 40440 33088 40480
rect 38470 40468 38476 40480
rect 38528 40468 38534 40520
rect 38657 40511 38715 40517
rect 38657 40477 38669 40511
rect 38703 40508 38715 40511
rect 39390 40508 39396 40520
rect 38703 40480 39396 40508
rect 38703 40477 38715 40480
rect 38657 40471 38715 40477
rect 39390 40468 39396 40480
rect 39448 40468 39454 40520
rect 40954 40468 40960 40520
rect 41012 40508 41018 40520
rect 41524 40517 41552 40548
rect 43346 40536 43352 40588
rect 43404 40576 43410 40588
rect 43625 40579 43683 40585
rect 43625 40576 43637 40579
rect 43404 40548 43637 40576
rect 43404 40536 43410 40548
rect 43625 40545 43637 40548
rect 43671 40576 43683 40579
rect 45002 40576 45008 40588
rect 43671 40548 45008 40576
rect 43671 40545 43683 40548
rect 43625 40539 43683 40545
rect 45002 40536 45008 40548
rect 45060 40536 45066 40588
rect 51997 40579 52055 40585
rect 51997 40545 52009 40579
rect 52043 40576 52055 40579
rect 52270 40576 52276 40588
rect 52043 40548 52276 40576
rect 52043 40545 52055 40548
rect 51997 40539 52055 40545
rect 52270 40536 52276 40548
rect 52328 40536 52334 40588
rect 53009 40579 53067 40585
rect 53009 40545 53021 40579
rect 53055 40576 53067 40579
rect 53098 40576 53104 40588
rect 53055 40548 53104 40576
rect 53055 40545 53067 40548
rect 53009 40539 53067 40545
rect 53098 40536 53104 40548
rect 53156 40536 53162 40588
rect 53193 40579 53251 40585
rect 53193 40545 53205 40579
rect 53239 40545 53251 40579
rect 53193 40539 53251 40545
rect 41417 40511 41475 40517
rect 41417 40508 41429 40511
rect 41012 40480 41429 40508
rect 41012 40468 41018 40480
rect 41417 40477 41429 40480
rect 41463 40477 41475 40511
rect 41417 40471 41475 40477
rect 41509 40511 41567 40517
rect 41509 40477 41521 40511
rect 41555 40477 41567 40511
rect 41509 40471 41567 40477
rect 52089 40511 52147 40517
rect 52089 40477 52101 40511
rect 52135 40508 52147 40511
rect 52914 40508 52920 40520
rect 52135 40480 52920 40508
rect 52135 40477 52147 40480
rect 52089 40471 52147 40477
rect 52914 40468 52920 40480
rect 52972 40508 52978 40520
rect 53208 40508 53236 40539
rect 54754 40536 54760 40588
rect 54812 40576 54818 40588
rect 55122 40576 55128 40588
rect 54812 40548 55128 40576
rect 54812 40536 54818 40548
rect 55122 40536 55128 40548
rect 55180 40576 55186 40588
rect 55309 40579 55367 40585
rect 55309 40576 55321 40579
rect 55180 40548 55321 40576
rect 55180 40536 55186 40548
rect 55309 40545 55321 40548
rect 55355 40545 55367 40579
rect 55858 40576 55864 40588
rect 55819 40548 55864 40576
rect 55309 40539 55367 40545
rect 55858 40536 55864 40548
rect 55916 40576 55922 40588
rect 56137 40579 56195 40585
rect 56137 40576 56149 40579
rect 55916 40548 56149 40576
rect 55916 40536 55922 40548
rect 56137 40545 56149 40548
rect 56183 40545 56195 40579
rect 56137 40539 56195 40545
rect 57149 40579 57207 40585
rect 57149 40545 57161 40579
rect 57195 40545 57207 40579
rect 57149 40539 57207 40545
rect 60645 40579 60703 40585
rect 60645 40545 60657 40579
rect 60691 40576 60703 40579
rect 61657 40579 61715 40585
rect 61657 40576 61669 40579
rect 60691 40548 61669 40576
rect 60691 40545 60703 40548
rect 60645 40539 60703 40545
rect 61657 40545 61669 40548
rect 61703 40545 61715 40579
rect 62298 40576 62304 40588
rect 62259 40548 62304 40576
rect 61657 40539 61715 40545
rect 52972 40480 53236 40508
rect 55677 40511 55735 40517
rect 52972 40468 52978 40480
rect 55677 40477 55689 40511
rect 55723 40508 55735 40511
rect 57164 40508 57192 40539
rect 62298 40536 62304 40548
rect 62356 40536 62362 40588
rect 62408 40585 62436 40616
rect 62942 40604 62948 40616
rect 63000 40604 63006 40656
rect 63862 40644 63868 40656
rect 63823 40616 63868 40644
rect 63862 40604 63868 40616
rect 63920 40604 63926 40656
rect 64598 40644 64604 40656
rect 64559 40616 64604 40644
rect 64598 40604 64604 40616
rect 64656 40604 64662 40656
rect 64690 40604 64696 40656
rect 64748 40644 64754 40656
rect 69569 40647 69627 40653
rect 69569 40644 69581 40647
rect 64748 40616 69581 40644
rect 64748 40604 64754 40616
rect 69569 40613 69581 40616
rect 69615 40644 69627 40647
rect 70118 40644 70124 40656
rect 69615 40616 70124 40644
rect 69615 40613 69627 40616
rect 69569 40607 69627 40613
rect 70118 40604 70124 40616
rect 70176 40644 70182 40656
rect 70213 40647 70271 40653
rect 70213 40644 70225 40647
rect 70176 40616 70225 40644
rect 70176 40604 70182 40616
rect 70213 40613 70225 40616
rect 70259 40613 70271 40647
rect 70213 40607 70271 40613
rect 62393 40579 62451 40585
rect 62393 40545 62405 40579
rect 62439 40545 62451 40579
rect 62393 40539 62451 40545
rect 55723 40480 57192 40508
rect 55723 40477 55735 40480
rect 55677 40471 55735 40477
rect 57238 40468 57244 40520
rect 57296 40508 57302 40520
rect 62408 40508 62436 40539
rect 62574 40536 62580 40588
rect 62632 40585 62638 40588
rect 62632 40579 62693 40585
rect 62632 40545 62647 40579
rect 62681 40545 62693 40579
rect 62632 40539 62693 40545
rect 62853 40579 62911 40585
rect 62853 40545 62865 40579
rect 62899 40545 62911 40579
rect 62853 40539 62911 40545
rect 62632 40536 62638 40539
rect 57296 40480 62436 40508
rect 57296 40468 57302 40480
rect 62758 40468 62764 40520
rect 62816 40508 62822 40520
rect 62868 40508 62896 40539
rect 63770 40536 63776 40588
rect 63828 40576 63834 40588
rect 63957 40579 64015 40585
rect 63957 40576 63969 40579
rect 63828 40548 63969 40576
rect 63828 40536 63834 40548
rect 63957 40545 63969 40548
rect 64003 40545 64015 40579
rect 64414 40576 64420 40588
rect 64375 40548 64420 40576
rect 63957 40539 64015 40545
rect 64414 40536 64420 40548
rect 64472 40536 64478 40588
rect 62816 40480 62896 40508
rect 63681 40511 63739 40517
rect 62816 40468 62822 40480
rect 63681 40477 63693 40511
rect 63727 40508 63739 40511
rect 64616 40508 64644 40604
rect 66714 40576 66720 40588
rect 66675 40548 66720 40576
rect 66714 40536 66720 40548
rect 66772 40536 66778 40588
rect 68462 40576 68468 40588
rect 68423 40548 68468 40576
rect 68462 40536 68468 40548
rect 68520 40536 68526 40588
rect 69382 40536 69388 40588
rect 69440 40576 69446 40588
rect 69753 40579 69811 40585
rect 69753 40576 69765 40579
rect 69440 40548 69765 40576
rect 69440 40536 69446 40548
rect 69753 40545 69765 40548
rect 69799 40545 69811 40579
rect 69753 40539 69811 40545
rect 63727 40480 64644 40508
rect 69768 40508 69796 40539
rect 69842 40536 69848 40588
rect 69900 40576 69906 40588
rect 71409 40579 71467 40585
rect 71409 40576 71421 40579
rect 69900 40548 71421 40576
rect 69900 40536 69906 40548
rect 71409 40545 71421 40548
rect 71455 40545 71467 40579
rect 71409 40539 71467 40545
rect 70394 40508 70400 40520
rect 69768 40480 70400 40508
rect 63727 40477 63739 40480
rect 63681 40471 63739 40477
rect 70394 40468 70400 40480
rect 70452 40468 70458 40520
rect 72344 40508 72372 40684
rect 72510 40672 72516 40684
rect 72568 40672 72574 40724
rect 77938 40672 77944 40724
rect 77996 40712 78002 40724
rect 78677 40715 78735 40721
rect 78677 40712 78689 40715
rect 77996 40684 78689 40712
rect 77996 40672 78002 40684
rect 78677 40681 78689 40684
rect 78723 40681 78735 40715
rect 78677 40675 78735 40681
rect 72528 40576 72556 40672
rect 77021 40647 77079 40653
rect 77021 40613 77033 40647
rect 77067 40644 77079 40647
rect 78214 40644 78220 40656
rect 77067 40616 78220 40644
rect 77067 40613 77079 40616
rect 77021 40607 77079 40613
rect 78214 40604 78220 40616
rect 78272 40604 78278 40656
rect 72605 40579 72663 40585
rect 72605 40576 72617 40579
rect 72528 40548 72617 40576
rect 72605 40545 72617 40548
rect 72651 40545 72663 40579
rect 75822 40576 75828 40588
rect 72605 40539 72663 40545
rect 72804 40548 75828 40576
rect 72804 40508 72832 40548
rect 75822 40536 75828 40548
rect 75880 40536 75886 40588
rect 77570 40576 77576 40588
rect 77531 40548 77576 40576
rect 77570 40536 77576 40548
rect 77628 40536 77634 40588
rect 77662 40536 77668 40588
rect 77720 40576 77726 40588
rect 77846 40576 77852 40588
rect 77720 40548 77852 40576
rect 77720 40536 77726 40548
rect 77846 40536 77852 40548
rect 77904 40536 77910 40588
rect 78033 40579 78091 40585
rect 78033 40545 78045 40579
rect 78079 40576 78091 40579
rect 78122 40576 78128 40588
rect 78079 40548 78128 40576
rect 78079 40545 78091 40548
rect 78033 40539 78091 40545
rect 78122 40536 78128 40548
rect 78180 40536 78186 40588
rect 78692 40576 78720 40675
rect 78861 40579 78919 40585
rect 78861 40576 78873 40579
rect 78692 40548 78873 40576
rect 78861 40545 78873 40548
rect 78907 40576 78919 40579
rect 83185 40579 83243 40585
rect 83185 40576 83197 40579
rect 78907 40548 83197 40576
rect 78907 40545 78919 40548
rect 78861 40539 78919 40545
rect 83185 40545 83197 40548
rect 83231 40576 83243 40579
rect 83369 40579 83427 40585
rect 83369 40576 83381 40579
rect 83231 40548 83381 40576
rect 83231 40545 83243 40548
rect 83185 40539 83243 40545
rect 83369 40545 83381 40548
rect 83415 40545 83427 40579
rect 83369 40539 83427 40545
rect 72344 40480 72832 40508
rect 72881 40511 72939 40517
rect 72881 40477 72893 40511
rect 72927 40508 72939 40511
rect 74442 40508 74448 40520
rect 72927 40480 74448 40508
rect 72927 40477 72939 40480
rect 72881 40471 72939 40477
rect 74442 40468 74448 40480
rect 74500 40468 74506 40520
rect 79137 40511 79195 40517
rect 79137 40477 79149 40511
rect 79183 40508 79195 40511
rect 80790 40508 80796 40520
rect 79183 40480 80796 40508
rect 79183 40477 79195 40480
rect 79137 40471 79195 40477
rect 80790 40468 80796 40480
rect 80848 40468 80854 40520
rect 83642 40508 83648 40520
rect 83603 40480 83648 40508
rect 83642 40468 83648 40480
rect 83700 40468 83706 40520
rect 62666 40440 62672 40452
rect 30975 40412 33088 40440
rect 33152 40412 62672 40440
rect 30975 40409 30987 40412
rect 30929 40403 30987 40409
rect 31113 40375 31171 40381
rect 31113 40372 31125 40375
rect 28408 40344 31125 40372
rect 28408 40332 28414 40344
rect 31113 40341 31125 40344
rect 31159 40372 31171 40375
rect 33152 40372 33180 40412
rect 62666 40400 62672 40412
rect 62724 40400 62730 40452
rect 66533 40443 66591 40449
rect 66533 40409 66545 40443
rect 66579 40440 66591 40443
rect 66806 40440 66812 40452
rect 66579 40412 66812 40440
rect 66579 40409 66591 40412
rect 66533 40403 66591 40409
rect 66806 40400 66812 40412
rect 66864 40400 66870 40452
rect 31159 40344 33180 40372
rect 31159 40341 31171 40344
rect 31113 40335 31171 40341
rect 34790 40332 34796 40384
rect 34848 40372 34854 40384
rect 34848 40344 34893 40372
rect 34848 40332 34854 40344
rect 35710 40332 35716 40384
rect 35768 40372 35774 40384
rect 36633 40375 36691 40381
rect 36633 40372 36645 40375
rect 35768 40344 36645 40372
rect 35768 40332 35774 40344
rect 36633 40341 36645 40344
rect 36679 40372 36691 40375
rect 36814 40372 36820 40384
rect 36679 40344 36820 40372
rect 36679 40341 36691 40344
rect 36633 40335 36691 40341
rect 36814 40332 36820 40344
rect 36872 40332 36878 40384
rect 37642 40332 37648 40384
rect 37700 40372 37706 40384
rect 38427 40375 38485 40381
rect 38427 40372 38439 40375
rect 37700 40344 38439 40372
rect 37700 40332 37706 40344
rect 38427 40341 38439 40344
rect 38473 40341 38485 40375
rect 38562 40372 38568 40384
rect 38523 40344 38568 40372
rect 38427 40335 38485 40341
rect 38562 40332 38568 40344
rect 38620 40332 38626 40384
rect 38654 40332 38660 40384
rect 38712 40372 38718 40384
rect 41187 40375 41245 40381
rect 41187 40372 41199 40375
rect 38712 40344 41199 40372
rect 38712 40332 38718 40344
rect 41187 40341 41199 40344
rect 41233 40341 41245 40375
rect 41187 40335 41245 40341
rect 41325 40375 41383 40381
rect 41325 40341 41337 40375
rect 41371 40372 41383 40375
rect 42702 40372 42708 40384
rect 41371 40344 42708 40372
rect 41371 40341 41383 40344
rect 41325 40335 41383 40341
rect 42702 40332 42708 40344
rect 42760 40332 42766 40384
rect 42794 40332 42800 40384
rect 42852 40372 42858 40384
rect 43622 40372 43628 40384
rect 42852 40344 43628 40372
rect 42852 40332 42858 40344
rect 43622 40332 43628 40344
rect 43680 40332 43686 40384
rect 53282 40372 53288 40384
rect 53243 40344 53288 40372
rect 53282 40332 53288 40344
rect 53340 40332 53346 40384
rect 56870 40372 56876 40384
rect 56831 40344 56876 40372
rect 56870 40332 56876 40344
rect 56928 40332 56934 40384
rect 57330 40372 57336 40384
rect 57291 40344 57336 40372
rect 57330 40332 57336 40344
rect 57388 40332 57394 40384
rect 57790 40372 57796 40384
rect 57751 40344 57796 40372
rect 57790 40332 57796 40344
rect 57848 40332 57854 40384
rect 62942 40332 62948 40384
rect 63000 40372 63006 40384
rect 63037 40375 63095 40381
rect 63037 40372 63049 40375
rect 63000 40344 63049 40372
rect 63000 40332 63006 40344
rect 63037 40341 63049 40344
rect 63083 40372 63095 40375
rect 68646 40372 68652 40384
rect 63083 40344 68652 40372
rect 63083 40341 63095 40344
rect 63037 40335 63095 40341
rect 68646 40332 68652 40344
rect 68704 40332 68710 40384
rect 69382 40372 69388 40384
rect 69343 40344 69388 40372
rect 69382 40332 69388 40344
rect 69440 40332 69446 40384
rect 69842 40372 69848 40384
rect 69803 40344 69848 40372
rect 69842 40332 69848 40344
rect 69900 40332 69906 40384
rect 70026 40332 70032 40384
rect 70084 40372 70090 40384
rect 71501 40375 71559 40381
rect 71501 40372 71513 40375
rect 70084 40344 71513 40372
rect 70084 40332 70090 40344
rect 71501 40341 71513 40344
rect 71547 40372 71559 40375
rect 71958 40372 71964 40384
rect 71547 40344 71964 40372
rect 71547 40341 71559 40344
rect 71501 40335 71559 40341
rect 71958 40332 71964 40344
rect 72016 40332 72022 40384
rect 73982 40372 73988 40384
rect 73943 40344 73988 40372
rect 73982 40332 73988 40344
rect 74040 40332 74046 40384
rect 75822 40332 75828 40384
rect 75880 40372 75886 40384
rect 78030 40372 78036 40384
rect 75880 40344 78036 40372
rect 75880 40332 75886 40344
rect 78030 40332 78036 40344
rect 78088 40332 78094 40384
rect 80238 40372 80244 40384
rect 80199 40344 80244 40372
rect 80238 40332 80244 40344
rect 80296 40332 80302 40384
rect 84746 40372 84752 40384
rect 84707 40344 84752 40372
rect 84746 40332 84752 40344
rect 84804 40332 84810 40384
rect 1104 40282 111136 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 65686 40282
rect 65738 40230 65750 40282
rect 65802 40230 65814 40282
rect 65866 40230 65878 40282
rect 65930 40230 96406 40282
rect 96458 40230 96470 40282
rect 96522 40230 96534 40282
rect 96586 40230 96598 40282
rect 96650 40230 111136 40282
rect 1104 40208 111136 40230
rect 4433 40171 4491 40177
rect 4433 40137 4445 40171
rect 4479 40168 4491 40171
rect 5442 40168 5448 40180
rect 4479 40140 5448 40168
rect 4479 40137 4491 40140
rect 4433 40131 4491 40137
rect 5442 40128 5448 40140
rect 5500 40128 5506 40180
rect 6914 40168 6920 40180
rect 6875 40140 6920 40168
rect 6914 40128 6920 40140
rect 6972 40128 6978 40180
rect 11146 40168 11152 40180
rect 11107 40140 11152 40168
rect 11146 40128 11152 40140
rect 11204 40128 11210 40180
rect 12894 40128 12900 40180
rect 12952 40168 12958 40180
rect 31570 40168 31576 40180
rect 12952 40140 31576 40168
rect 12952 40128 12958 40140
rect 31570 40128 31576 40140
rect 31628 40128 31634 40180
rect 35713 40171 35771 40177
rect 35713 40168 35725 40171
rect 32784 40140 35725 40168
rect 4706 40100 4712 40112
rect 4667 40072 4712 40100
rect 4706 40060 4712 40072
rect 4764 40060 4770 40112
rect 10686 40100 10692 40112
rect 10336 40072 10692 40100
rect 3145 40035 3203 40041
rect 3145 40001 3157 40035
rect 3191 40032 3203 40035
rect 4614 40032 4620 40044
rect 3191 40004 4620 40032
rect 3191 40001 3203 40004
rect 3145 39995 3203 40001
rect 4614 39992 4620 40004
rect 4672 39992 4678 40044
rect 2869 39967 2927 39973
rect 2869 39933 2881 39967
rect 2915 39964 2927 39967
rect 4724 39964 4752 40060
rect 9766 39992 9772 40044
rect 9824 40032 9830 40044
rect 9953 40035 10011 40041
rect 9953 40032 9965 40035
rect 9824 40004 9965 40032
rect 9824 39992 9830 40004
rect 9953 40001 9965 40004
rect 9999 40001 10011 40035
rect 9953 39995 10011 40001
rect 5718 39964 5724 39976
rect 2915 39936 4752 39964
rect 5679 39936 5724 39964
rect 2915 39933 2927 39936
rect 2869 39927 2927 39933
rect 5718 39924 5724 39936
rect 5776 39924 5782 39976
rect 7098 39973 7104 39976
rect 7093 39927 7104 39973
rect 7156 39964 7162 39976
rect 7156 39936 7193 39964
rect 7098 39924 7104 39927
rect 7156 39924 7162 39936
rect 7282 39924 7288 39976
rect 7340 39964 7346 39976
rect 10137 39967 10195 39973
rect 10137 39964 10149 39967
rect 7340 39936 10149 39964
rect 7340 39924 7346 39936
rect 10137 39933 10149 39936
rect 10183 39964 10195 39967
rect 10336 39964 10364 40072
rect 10686 40060 10692 40072
rect 10744 40100 10750 40112
rect 11517 40103 11575 40109
rect 11517 40100 11529 40103
rect 10744 40072 11529 40100
rect 10744 40060 10750 40072
rect 11517 40069 11529 40072
rect 11563 40100 11575 40103
rect 11701 40103 11759 40109
rect 11701 40100 11713 40103
rect 11563 40072 11713 40100
rect 11563 40069 11575 40072
rect 11517 40063 11575 40069
rect 11701 40069 11713 40072
rect 11747 40100 11759 40103
rect 14182 40100 14188 40112
rect 11747 40072 14188 40100
rect 11747 40069 11759 40072
rect 11701 40063 11759 40069
rect 14182 40060 14188 40072
rect 14240 40060 14246 40112
rect 16850 40060 16856 40112
rect 16908 40100 16914 40112
rect 17773 40103 17831 40109
rect 17773 40100 17785 40103
rect 16908 40072 17785 40100
rect 16908 40060 16914 40072
rect 17773 40069 17785 40072
rect 17819 40100 17831 40103
rect 19613 40103 19671 40109
rect 17819 40072 19104 40100
rect 17819 40069 17831 40072
rect 17773 40063 17831 40069
rect 17678 40032 17684 40044
rect 17639 40004 17684 40032
rect 17678 39992 17684 40004
rect 17736 39992 17742 40044
rect 18785 40035 18843 40041
rect 18785 40001 18797 40035
rect 18831 40001 18843 40035
rect 18785 39995 18843 40001
rect 10183 39936 10364 39964
rect 10183 39933 10195 39936
rect 10137 39927 10195 39933
rect 10686 39924 10692 39976
rect 10744 39964 10750 39976
rect 10744 39936 10789 39964
rect 10744 39924 10750 39936
rect 10870 39924 10876 39976
rect 10928 39964 10934 39976
rect 12986 39964 12992 39976
rect 10928 39936 12992 39964
rect 10928 39924 10934 39936
rect 12986 39924 12992 39936
rect 13044 39924 13050 39976
rect 13081 39967 13139 39973
rect 13081 39933 13093 39967
rect 13127 39964 13139 39967
rect 13354 39964 13360 39976
rect 13127 39936 13360 39964
rect 13127 39933 13139 39936
rect 13081 39927 13139 39933
rect 13354 39924 13360 39936
rect 13412 39924 13418 39976
rect 17696 39964 17724 39992
rect 18693 39967 18751 39973
rect 18693 39964 18705 39967
rect 17696 39936 18705 39964
rect 18693 39933 18705 39936
rect 18739 39933 18751 39967
rect 18693 39927 18751 39933
rect 4062 39856 4068 39908
rect 4120 39896 4126 39908
rect 18800 39896 18828 39995
rect 19076 39973 19104 40072
rect 19613 40069 19625 40103
rect 19659 40100 19671 40103
rect 19978 40100 19984 40112
rect 19659 40072 19984 40100
rect 19659 40069 19671 40072
rect 19613 40063 19671 40069
rect 19978 40060 19984 40072
rect 20036 40060 20042 40112
rect 23201 40103 23259 40109
rect 23201 40069 23213 40103
rect 23247 40100 23259 40103
rect 23382 40100 23388 40112
rect 23247 40072 23388 40100
rect 23247 40069 23259 40072
rect 23201 40063 23259 40069
rect 23382 40060 23388 40072
rect 23440 40100 23446 40112
rect 25409 40103 25467 40109
rect 25409 40100 25421 40103
rect 23440 40072 23704 40100
rect 23440 40060 23446 40072
rect 19429 40035 19487 40041
rect 19429 40032 19441 40035
rect 19260 40004 19441 40032
rect 19260 39973 19288 40004
rect 19429 40001 19441 40004
rect 19475 40032 19487 40035
rect 23566 40032 23572 40044
rect 19475 40004 23572 40032
rect 19475 40001 19487 40004
rect 19429 39995 19487 40001
rect 23566 39992 23572 40004
rect 23624 39992 23630 40044
rect 23676 40041 23704 40072
rect 23952 40072 25421 40100
rect 23661 40035 23719 40041
rect 23661 40001 23673 40035
rect 23707 40001 23719 40035
rect 23952 40032 23980 40072
rect 25409 40069 25421 40072
rect 25455 40100 25467 40103
rect 25498 40100 25504 40112
rect 25455 40072 25504 40100
rect 25455 40069 25467 40072
rect 25409 40063 25467 40069
rect 25498 40060 25504 40072
rect 25556 40060 25562 40112
rect 25682 40060 25688 40112
rect 25740 40100 25746 40112
rect 25777 40103 25835 40109
rect 25777 40100 25789 40103
rect 25740 40072 25789 40100
rect 25740 40060 25746 40072
rect 25777 40069 25789 40072
rect 25823 40100 25835 40103
rect 26510 40100 26516 40112
rect 25823 40072 26516 40100
rect 25823 40069 25835 40072
rect 25777 40063 25835 40069
rect 26510 40060 26516 40072
rect 26568 40100 26574 40112
rect 27522 40100 27528 40112
rect 26568 40072 27528 40100
rect 26568 40060 26574 40072
rect 27522 40060 27528 40072
rect 27580 40060 27586 40112
rect 27617 40103 27675 40109
rect 27617 40069 27629 40103
rect 27663 40100 27675 40103
rect 28350 40100 28356 40112
rect 27663 40072 28356 40100
rect 27663 40069 27675 40072
rect 27617 40063 27675 40069
rect 23661 39995 23719 40001
rect 23860 40004 23980 40032
rect 19061 39967 19119 39973
rect 19061 39933 19073 39967
rect 19107 39933 19119 39967
rect 19061 39927 19119 39933
rect 19245 39967 19303 39973
rect 19245 39933 19257 39967
rect 19291 39933 19303 39967
rect 19245 39927 19303 39933
rect 19334 39924 19340 39976
rect 19392 39964 19398 39976
rect 23474 39964 23480 39976
rect 19392 39936 23480 39964
rect 19392 39924 19398 39936
rect 23474 39924 23480 39936
rect 23532 39924 23538 39976
rect 23860 39973 23888 40004
rect 24854 39992 24860 40044
rect 24912 40032 24918 40044
rect 25225 40035 25283 40041
rect 25225 40032 25237 40035
rect 24912 40004 25237 40032
rect 24912 39992 24918 40004
rect 25225 40001 25237 40004
rect 25271 40032 25283 40035
rect 25271 40004 26096 40032
rect 25271 40001 25283 40004
rect 25225 39995 25283 40001
rect 23845 39967 23903 39973
rect 23845 39933 23857 39967
rect 23891 39933 23903 39967
rect 23845 39927 23903 39933
rect 24305 39967 24363 39973
rect 24305 39933 24317 39967
rect 24351 39933 24363 39967
rect 24305 39927 24363 39933
rect 24397 39967 24455 39973
rect 24397 39933 24409 39967
rect 24443 39933 24455 39967
rect 24397 39927 24455 39933
rect 19978 39896 19984 39908
rect 4120 39868 10732 39896
rect 4120 39856 4126 39868
rect 5810 39828 5816 39840
rect 5771 39800 5816 39828
rect 5810 39788 5816 39800
rect 5868 39788 5874 39840
rect 7193 39831 7251 39837
rect 7193 39797 7205 39831
rect 7239 39828 7251 39831
rect 7834 39828 7840 39840
rect 7239 39800 7840 39828
rect 7239 39797 7251 39800
rect 7193 39791 7251 39797
rect 7834 39788 7840 39800
rect 7892 39788 7898 39840
rect 9766 39828 9772 39840
rect 9727 39800 9772 39828
rect 9766 39788 9772 39800
rect 9824 39788 9830 39840
rect 10704 39828 10732 39868
rect 11072 39868 18276 39896
rect 18800 39868 19984 39896
rect 11072 39828 11100 39868
rect 10704 39800 11100 39828
rect 11698 39788 11704 39840
rect 11756 39828 11762 39840
rect 13262 39828 13268 39840
rect 11756 39800 13268 39828
rect 11756 39788 11762 39800
rect 13262 39788 13268 39800
rect 13320 39788 13326 39840
rect 13354 39788 13360 39840
rect 13412 39828 13418 39840
rect 13449 39831 13507 39837
rect 13449 39828 13461 39831
rect 13412 39800 13461 39828
rect 13412 39788 13418 39800
rect 13449 39797 13461 39800
rect 13495 39797 13507 39831
rect 13449 39791 13507 39797
rect 14642 39788 14648 39840
rect 14700 39828 14706 39840
rect 18141 39831 18199 39837
rect 18141 39828 18153 39831
rect 14700 39800 18153 39828
rect 14700 39788 14706 39800
rect 18141 39797 18153 39800
rect 18187 39797 18199 39831
rect 18248 39828 18276 39868
rect 19978 39856 19984 39868
rect 20036 39856 20042 39908
rect 23385 39899 23443 39905
rect 23385 39865 23397 39899
rect 23431 39896 23443 39899
rect 23566 39896 23572 39908
rect 23431 39868 23572 39896
rect 23431 39865 23443 39868
rect 23385 39859 23443 39865
rect 23566 39856 23572 39868
rect 23624 39896 23630 39908
rect 24320 39896 24348 39927
rect 23624 39868 24348 39896
rect 24412 39896 24440 39927
rect 24578 39924 24584 39976
rect 24636 39964 24642 39976
rect 26068 39973 26096 40004
rect 25501 39967 25559 39973
rect 25501 39964 25513 39967
rect 24636 39936 25513 39964
rect 24636 39924 24642 39936
rect 25501 39933 25513 39936
rect 25547 39964 25559 39967
rect 25869 39967 25927 39973
rect 25869 39964 25881 39967
rect 25547 39936 25881 39964
rect 25547 39933 25559 39936
rect 25501 39927 25559 39933
rect 25869 39933 25881 39936
rect 25915 39933 25927 39967
rect 25869 39927 25927 39933
rect 26053 39967 26111 39973
rect 26053 39933 26065 39967
rect 26099 39964 26111 39967
rect 26510 39964 26516 39976
rect 26099 39936 26188 39964
rect 26471 39936 26516 39964
rect 26099 39933 26111 39936
rect 26053 39927 26111 39933
rect 24854 39896 24860 39908
rect 24412 39868 24860 39896
rect 23624 39856 23630 39868
rect 20438 39828 20444 39840
rect 18248 39800 20444 39828
rect 18141 39791 18199 39797
rect 20438 39788 20444 39800
rect 20496 39788 20502 39840
rect 23290 39788 23296 39840
rect 23348 39828 23354 39840
rect 24412 39828 24440 39868
rect 24854 39856 24860 39868
rect 24912 39856 24918 39908
rect 24949 39899 25007 39905
rect 24949 39865 24961 39899
rect 24995 39896 25007 39899
rect 26160 39896 26188 39936
rect 26510 39924 26516 39936
rect 26568 39924 26574 39976
rect 26602 39924 26608 39976
rect 26660 39964 26666 39976
rect 27632 39964 27660 40063
rect 28350 40060 28356 40072
rect 28408 40060 28414 40112
rect 28626 40060 28632 40112
rect 28684 40100 28690 40112
rect 32784 40100 32812 40140
rect 35713 40137 35725 40140
rect 35759 40168 35771 40171
rect 35894 40168 35900 40180
rect 35759 40140 35900 40168
rect 35759 40137 35771 40140
rect 35713 40131 35771 40137
rect 35894 40128 35900 40140
rect 35952 40168 35958 40180
rect 37185 40171 37243 40177
rect 35952 40140 36400 40168
rect 35952 40128 35958 40140
rect 28684 40072 32812 40100
rect 32861 40103 32919 40109
rect 28684 40060 28690 40072
rect 32861 40069 32873 40103
rect 32907 40100 32919 40103
rect 32907 40072 33548 40100
rect 32907 40069 32919 40072
rect 32861 40063 32919 40069
rect 32125 40035 32183 40041
rect 32125 40001 32137 40035
rect 32171 40032 32183 40035
rect 32214 40032 32220 40044
rect 32171 40004 32220 40032
rect 32171 40001 32183 40004
rect 32125 39995 32183 40001
rect 32214 39992 32220 40004
rect 32272 39992 32278 40044
rect 32674 39992 32680 40044
rect 32732 40041 32738 40044
rect 32732 40035 32790 40041
rect 32732 40001 32744 40035
rect 32778 40001 32790 40035
rect 32950 40032 32956 40044
rect 32911 40004 32956 40032
rect 32732 39995 32790 40001
rect 32732 39992 32738 39995
rect 32950 39992 32956 40004
rect 33008 39992 33014 40044
rect 30558 39964 30564 39976
rect 26660 39936 27660 39964
rect 30519 39936 30564 39964
rect 26660 39924 26666 39936
rect 30558 39924 30564 39936
rect 30616 39924 30622 39976
rect 30653 39967 30711 39973
rect 30653 39933 30665 39967
rect 30699 39964 30711 39967
rect 30742 39964 30748 39976
rect 30699 39936 30748 39964
rect 30699 39933 30711 39936
rect 30653 39927 30711 39933
rect 30742 39924 30748 39936
rect 30800 39924 30806 39976
rect 30926 39924 30932 39976
rect 30984 39964 30990 39976
rect 31021 39967 31079 39973
rect 31021 39964 31033 39967
rect 30984 39936 31033 39964
rect 30984 39924 30990 39936
rect 31021 39933 31033 39936
rect 31067 39933 31079 39967
rect 31021 39927 31079 39933
rect 31110 39924 31116 39976
rect 31168 39964 31174 39976
rect 32582 39964 32588 39976
rect 31168 39936 31213 39964
rect 31312 39936 32444 39964
rect 32543 39936 32588 39964
rect 31168 39924 31174 39936
rect 27433 39899 27491 39905
rect 27433 39896 27445 39899
rect 24995 39868 26096 39896
rect 26160 39868 27445 39896
rect 24995 39865 25007 39868
rect 24949 39859 25007 39865
rect 23348 39800 24440 39828
rect 26068 39828 26096 39868
rect 27433 39865 27445 39868
rect 27479 39896 27491 39899
rect 31312 39896 31340 39936
rect 27479 39868 31340 39896
rect 31665 39899 31723 39905
rect 27479 39865 27491 39868
rect 27433 39859 27491 39865
rect 31665 39865 31677 39899
rect 31711 39896 31723 39899
rect 32122 39896 32128 39908
rect 31711 39868 32128 39896
rect 31711 39865 31723 39868
rect 31665 39859 31723 39865
rect 32122 39856 32128 39868
rect 32180 39856 32186 39908
rect 32416 39896 32444 39936
rect 32582 39924 32588 39936
rect 32640 39924 32646 39976
rect 33321 39967 33379 39973
rect 33321 39933 33333 39967
rect 33367 39964 33379 39967
rect 33410 39964 33416 39976
rect 33367 39936 33416 39964
rect 33367 39933 33379 39936
rect 33321 39927 33379 39933
rect 33410 39924 33416 39936
rect 33468 39924 33474 39976
rect 33520 39905 33548 40072
rect 34790 40060 34796 40112
rect 34848 40100 34854 40112
rect 35618 40100 35624 40112
rect 34848 40072 35624 40100
rect 34848 40060 34854 40072
rect 35618 40060 35624 40072
rect 35676 40100 35682 40112
rect 35805 40103 35863 40109
rect 35805 40100 35817 40103
rect 35676 40072 35817 40100
rect 35676 40060 35682 40072
rect 35805 40069 35817 40072
rect 35851 40069 35863 40103
rect 35805 40063 35863 40069
rect 34054 39992 34060 40044
rect 34112 40032 34118 40044
rect 35342 40032 35348 40044
rect 34112 40004 35348 40032
rect 34112 39992 34118 40004
rect 35342 39992 35348 40004
rect 35400 39992 35406 40044
rect 35820 40032 35848 40063
rect 35989 40035 36047 40041
rect 35989 40032 36001 40035
rect 35820 40004 36001 40032
rect 35989 40001 36001 40004
rect 36035 40001 36047 40035
rect 35989 39995 36047 40001
rect 35710 39924 35716 39976
rect 35768 39964 35774 39976
rect 36127 39967 36185 39973
rect 36127 39964 36139 39967
rect 35768 39936 36139 39964
rect 35768 39924 35774 39936
rect 36127 39933 36139 39936
rect 36173 39933 36185 39967
rect 36372 39964 36400 40140
rect 37185 40137 37197 40171
rect 37231 40168 37243 40171
rect 38654 40168 38660 40180
rect 37231 40140 38660 40168
rect 37231 40137 37243 40140
rect 37185 40131 37243 40137
rect 38654 40128 38660 40140
rect 38712 40128 38718 40180
rect 39393 40171 39451 40177
rect 39393 40137 39405 40171
rect 39439 40168 39451 40171
rect 43855 40171 43913 40177
rect 43855 40168 43867 40171
rect 39439 40140 43867 40168
rect 39439 40137 39451 40140
rect 39393 40131 39451 40137
rect 43855 40137 43867 40140
rect 43901 40137 43913 40171
rect 43855 40131 43913 40137
rect 52641 40171 52699 40177
rect 52641 40137 52653 40171
rect 52687 40168 52699 40171
rect 54846 40168 54852 40180
rect 52687 40140 54852 40168
rect 52687 40137 52699 40140
rect 52641 40131 52699 40137
rect 54846 40128 54852 40140
rect 54904 40128 54910 40180
rect 55766 40128 55772 40180
rect 55824 40168 55830 40180
rect 61562 40168 61568 40180
rect 55824 40140 61568 40168
rect 55824 40128 55830 40140
rect 61562 40128 61568 40140
rect 61620 40128 61626 40180
rect 62666 40128 62672 40180
rect 62724 40168 62730 40180
rect 69106 40168 69112 40180
rect 62724 40140 69112 40168
rect 62724 40128 62730 40140
rect 69106 40128 69112 40140
rect 69164 40128 69170 40180
rect 70118 40128 70124 40180
rect 70176 40168 70182 40180
rect 70302 40168 70308 40180
rect 70176 40140 70308 40168
rect 70176 40128 70182 40140
rect 70302 40128 70308 40140
rect 70360 40128 70366 40180
rect 70486 40128 70492 40180
rect 70544 40168 70550 40180
rect 70544 40140 77800 40168
rect 70544 40128 70550 40140
rect 36814 40060 36820 40112
rect 36872 40100 36878 40112
rect 37918 40100 37924 40112
rect 36872 40072 37228 40100
rect 37831 40072 37924 40100
rect 36872 40060 36878 40072
rect 37200 40032 37228 40072
rect 37918 40060 37924 40072
rect 37976 40100 37982 40112
rect 42242 40100 42248 40112
rect 37976 40072 38516 40100
rect 37976 40060 37982 40072
rect 37737 40035 37795 40041
rect 37737 40032 37749 40035
rect 37200 40004 37749 40032
rect 37737 40001 37749 40004
rect 37783 40032 37795 40035
rect 37783 40004 38424 40032
rect 37783 40001 37795 40004
rect 37737 39995 37795 40001
rect 38396 39976 38424 40004
rect 36633 39967 36691 39973
rect 36633 39964 36645 39967
rect 36372 39936 36645 39964
rect 36127 39927 36185 39933
rect 36633 39933 36645 39936
rect 36679 39933 36691 39967
rect 36633 39927 36691 39933
rect 36725 39967 36783 39973
rect 36725 39933 36737 39967
rect 36771 39964 36783 39967
rect 36906 39964 36912 39976
rect 36771 39936 36912 39964
rect 36771 39933 36783 39936
rect 36725 39927 36783 39933
rect 36906 39924 36912 39936
rect 36964 39964 36970 39976
rect 37461 39967 37519 39973
rect 37461 39964 37473 39967
rect 36964 39936 37473 39964
rect 36964 39924 36970 39936
rect 37461 39933 37473 39936
rect 37507 39933 37519 39967
rect 38194 39964 38200 39976
rect 38155 39936 38200 39964
rect 37461 39927 37519 39933
rect 38194 39924 38200 39936
rect 38252 39924 38258 39976
rect 38378 39964 38384 39976
rect 38339 39936 38384 39964
rect 38378 39924 38384 39936
rect 38436 39924 38442 39976
rect 38488 39964 38516 40072
rect 41800 40072 42248 40100
rect 38841 39967 38899 39973
rect 38841 39964 38853 39967
rect 38488 39936 38853 39964
rect 38841 39933 38853 39936
rect 38887 39933 38899 39967
rect 38841 39927 38899 39933
rect 38930 39924 38936 39976
rect 38988 39964 38994 39976
rect 39669 39967 39727 39973
rect 39669 39964 39681 39967
rect 38988 39936 39681 39964
rect 38988 39924 38994 39936
rect 39669 39933 39681 39936
rect 39715 39933 39727 39967
rect 39669 39927 39727 39933
rect 40034 39924 40040 39976
rect 40092 39964 40098 39976
rect 41141 39967 41199 39973
rect 41141 39964 41153 39967
rect 40092 39936 41153 39964
rect 40092 39924 40098 39936
rect 41141 39933 41153 39936
rect 41187 39964 41199 39967
rect 41325 39967 41383 39973
rect 41325 39964 41337 39967
rect 41187 39936 41337 39964
rect 41187 39933 41199 39936
rect 41141 39927 41199 39933
rect 41325 39933 41337 39936
rect 41371 39964 41383 39967
rect 41506 39964 41512 39976
rect 41371 39936 41512 39964
rect 41371 39933 41383 39936
rect 41325 39927 41383 39933
rect 41506 39924 41512 39936
rect 41564 39924 41570 39976
rect 41693 39967 41751 39973
rect 41693 39933 41705 39967
rect 41739 39964 41751 39967
rect 41800 39964 41828 40072
rect 42242 40060 42248 40072
rect 42300 40060 42306 40112
rect 43993 40103 44051 40109
rect 43993 40069 44005 40103
rect 44039 40100 44051 40103
rect 44634 40100 44640 40112
rect 44039 40072 44640 40100
rect 44039 40069 44051 40072
rect 43993 40063 44051 40069
rect 44634 40060 44640 40072
rect 44692 40060 44698 40112
rect 47780 40072 48544 40100
rect 42702 40032 42708 40044
rect 42663 40004 42708 40032
rect 42702 39992 42708 40004
rect 42760 39992 42766 40044
rect 44085 40035 44143 40041
rect 44085 40001 44097 40035
rect 44131 40001 44143 40035
rect 47780 40032 47808 40072
rect 44085 39995 44143 40001
rect 47596 40004 47808 40032
rect 48516 40032 48544 40072
rect 56870 40060 56876 40112
rect 56928 40100 56934 40112
rect 57790 40100 57796 40112
rect 56928 40072 57796 40100
rect 56928 40060 56934 40072
rect 57790 40060 57796 40072
rect 57848 40060 57854 40112
rect 66162 40060 66168 40112
rect 66220 40100 66226 40112
rect 71593 40103 71651 40109
rect 71593 40100 71605 40103
rect 66220 40072 71605 40100
rect 66220 40060 66226 40072
rect 71593 40069 71605 40072
rect 71639 40100 71651 40103
rect 74258 40100 74264 40112
rect 71639 40072 74264 40100
rect 71639 40069 71651 40072
rect 71593 40063 71651 40069
rect 74258 40060 74264 40072
rect 74316 40060 74322 40112
rect 74460 40072 75040 40100
rect 48866 40032 48872 40044
rect 48516 40004 48872 40032
rect 42153 39967 42211 39973
rect 42153 39964 42165 39967
rect 41739 39936 41828 39964
rect 41892 39936 42165 39964
rect 41739 39933 41751 39936
rect 41693 39927 41751 39933
rect 33505 39899 33563 39905
rect 32416 39868 33364 39896
rect 26142 39828 26148 39840
rect 26068 39800 26148 39828
rect 23348 39788 23354 39800
rect 26142 39788 26148 39800
rect 26200 39788 26206 39840
rect 26510 39788 26516 39840
rect 26568 39828 26574 39840
rect 27065 39831 27123 39837
rect 27065 39828 27077 39831
rect 26568 39800 27077 39828
rect 26568 39788 26574 39800
rect 27065 39797 27077 39800
rect 27111 39797 27123 39831
rect 27065 39791 27123 39797
rect 31110 39788 31116 39840
rect 31168 39828 31174 39840
rect 31754 39828 31760 39840
rect 31168 39800 31760 39828
rect 31168 39788 31174 39800
rect 31754 39788 31760 39800
rect 31812 39828 31818 39840
rect 31849 39831 31907 39837
rect 31849 39828 31861 39831
rect 31812 39800 31861 39828
rect 31812 39788 31818 39800
rect 31849 39797 31861 39800
rect 31895 39797 31907 39831
rect 33336 39828 33364 39868
rect 33505 39865 33517 39899
rect 33551 39896 33563 39899
rect 38102 39896 38108 39908
rect 33551 39868 38108 39896
rect 33551 39865 33563 39868
rect 33505 39859 33563 39865
rect 38102 39856 38108 39868
rect 38160 39856 38166 39908
rect 35526 39828 35532 39840
rect 33336 39800 35532 39828
rect 31849 39791 31907 39797
rect 35526 39788 35532 39800
rect 35584 39788 35590 39840
rect 35802 39788 35808 39840
rect 35860 39828 35866 39840
rect 38013 39831 38071 39837
rect 38013 39828 38025 39831
rect 35860 39800 38025 39828
rect 35860 39788 35866 39800
rect 38013 39797 38025 39800
rect 38059 39828 38071 39831
rect 38194 39828 38200 39840
rect 38059 39800 38200 39828
rect 38059 39797 38071 39800
rect 38013 39791 38071 39797
rect 38194 39788 38200 39800
rect 38252 39788 38258 39840
rect 38378 39788 38384 39840
rect 38436 39828 38442 39840
rect 39945 39831 40003 39837
rect 39945 39828 39957 39831
rect 38436 39800 39957 39828
rect 38436 39788 38442 39800
rect 39945 39797 39957 39800
rect 39991 39828 40003 39831
rect 41046 39828 41052 39840
rect 39991 39800 41052 39828
rect 39991 39797 40003 39800
rect 39945 39791 40003 39797
rect 41046 39788 41052 39800
rect 41104 39788 41110 39840
rect 41506 39788 41512 39840
rect 41564 39828 41570 39840
rect 41892 39828 41920 39936
rect 42153 39933 42165 39936
rect 42199 39933 42211 39967
rect 42153 39927 42211 39933
rect 42242 39924 42248 39976
rect 42300 39964 42306 39976
rect 43257 39967 43315 39973
rect 43257 39964 43269 39967
rect 42300 39936 43269 39964
rect 42300 39924 42306 39936
rect 43257 39933 43269 39936
rect 43303 39964 43315 39967
rect 43441 39967 43499 39973
rect 43441 39964 43453 39967
rect 43303 39936 43453 39964
rect 43303 39933 43315 39936
rect 43257 39927 43315 39933
rect 43441 39933 43453 39936
rect 43487 39964 43499 39967
rect 43530 39964 43536 39976
rect 43487 39936 43536 39964
rect 43487 39933 43499 39936
rect 43441 39927 43499 39933
rect 43530 39924 43536 39936
rect 43588 39924 43594 39976
rect 43990 39924 43996 39976
rect 44048 39964 44054 39976
rect 44100 39964 44128 39995
rect 47596 39973 47624 40004
rect 48866 39992 48872 40004
rect 48924 40032 48930 40044
rect 48961 40035 49019 40041
rect 48961 40032 48973 40035
rect 48924 40004 48973 40032
rect 48924 39992 48930 40004
rect 48961 40001 48973 40004
rect 49007 40032 49019 40035
rect 49007 40004 55628 40032
rect 49007 40001 49019 40004
rect 48961 39995 49019 40001
rect 44048 39936 44128 39964
rect 47581 39967 47639 39973
rect 44048 39924 44054 39936
rect 47581 39933 47593 39967
rect 47627 39933 47639 39967
rect 47581 39927 47639 39933
rect 47670 39924 47676 39976
rect 47728 39964 47734 39976
rect 48041 39967 48099 39973
rect 47728 39936 47773 39964
rect 47728 39924 47734 39936
rect 48041 39933 48053 39967
rect 48087 39933 48099 39967
rect 48041 39927 48099 39933
rect 43714 39896 43720 39908
rect 42904 39868 43576 39896
rect 43675 39868 43720 39896
rect 41564 39800 41920 39828
rect 41564 39788 41570 39800
rect 42242 39788 42248 39840
rect 42300 39828 42306 39840
rect 42904 39828 42932 39868
rect 43070 39828 43076 39840
rect 42300 39800 42932 39828
rect 43031 39800 43076 39828
rect 42300 39788 42306 39800
rect 43070 39788 43076 39800
rect 43128 39788 43134 39840
rect 43548 39828 43576 39868
rect 43714 39856 43720 39868
rect 43772 39856 43778 39908
rect 47213 39899 47271 39905
rect 47213 39896 47225 39899
rect 44008 39868 47225 39896
rect 44008 39828 44036 39868
rect 47213 39865 47225 39868
rect 47259 39896 47271 39899
rect 48056 39896 48084 39927
rect 48130 39924 48136 39976
rect 48188 39964 48194 39976
rect 49142 39964 49148 39976
rect 48188 39936 49148 39964
rect 48188 39924 48194 39936
rect 49142 39924 49148 39936
rect 49200 39924 49206 39976
rect 52365 39967 52423 39973
rect 52365 39933 52377 39967
rect 52411 39964 52423 39967
rect 52454 39964 52460 39976
rect 52411 39936 52460 39964
rect 52411 39933 52423 39936
rect 52365 39927 52423 39933
rect 52454 39924 52460 39936
rect 52512 39924 52518 39976
rect 52546 39924 52552 39976
rect 52604 39964 52610 39976
rect 53742 39964 53748 39976
rect 52604 39936 52649 39964
rect 53703 39936 53748 39964
rect 52604 39924 52610 39936
rect 53742 39924 53748 39936
rect 53800 39924 53806 39976
rect 54018 39964 54024 39976
rect 53979 39936 54024 39964
rect 54018 39924 54024 39936
rect 54076 39924 54082 39976
rect 54110 39924 54116 39976
rect 54168 39964 54174 39976
rect 55490 39964 55496 39976
rect 54168 39936 55496 39964
rect 54168 39924 54174 39936
rect 55490 39924 55496 39936
rect 55548 39924 55554 39976
rect 52178 39896 52184 39908
rect 47259 39868 48084 39896
rect 48148 39868 52184 39896
rect 47259 39865 47271 39868
rect 47213 39859 47271 39865
rect 43548 39800 44036 39828
rect 44266 39788 44272 39840
rect 44324 39828 44330 39840
rect 44361 39831 44419 39837
rect 44361 39828 44373 39831
rect 44324 39800 44373 39828
rect 44324 39788 44330 39800
rect 44361 39797 44373 39800
rect 44407 39797 44419 39831
rect 44361 39791 44419 39797
rect 44542 39788 44548 39840
rect 44600 39828 44606 39840
rect 48148 39828 48176 39868
rect 52178 39856 52184 39868
rect 52236 39856 52242 39908
rect 48590 39828 48596 39840
rect 44600 39800 48176 39828
rect 48551 39800 48596 39828
rect 44600 39788 44606 39800
rect 48590 39788 48596 39800
rect 48648 39788 48654 39840
rect 48682 39788 48688 39840
rect 48740 39828 48746 39840
rect 52270 39828 52276 39840
rect 48740 39800 52276 39828
rect 48740 39788 48746 39800
rect 52270 39788 52276 39800
rect 52328 39788 52334 39840
rect 52546 39788 52552 39840
rect 52604 39828 52610 39840
rect 55125 39831 55183 39837
rect 55125 39828 55137 39831
rect 52604 39800 55137 39828
rect 52604 39788 52610 39800
rect 55125 39797 55137 39800
rect 55171 39797 55183 39831
rect 55600 39828 55628 40004
rect 56042 39992 56048 40044
rect 56100 40032 56106 40044
rect 56888 40032 56916 40060
rect 56100 40004 56916 40032
rect 60185 40035 60243 40041
rect 56100 39992 56106 40004
rect 60185 40001 60197 40035
rect 60231 40032 60243 40035
rect 61930 40032 61936 40044
rect 60231 40004 61936 40032
rect 60231 40001 60243 40004
rect 60185 39995 60243 40001
rect 61930 39992 61936 40004
rect 61988 39992 61994 40044
rect 63957 40035 64015 40041
rect 63957 40001 63969 40035
rect 64003 40032 64015 40035
rect 64414 40032 64420 40044
rect 64003 40004 64420 40032
rect 64003 40001 64015 40004
rect 63957 39995 64015 40001
rect 64414 39992 64420 40004
rect 64472 39992 64478 40044
rect 65521 40035 65579 40041
rect 65521 40001 65533 40035
rect 65567 40032 65579 40035
rect 66806 40032 66812 40044
rect 65567 40004 66812 40032
rect 65567 40001 65579 40004
rect 65521 39995 65579 40001
rect 60461 39967 60519 39973
rect 60461 39933 60473 39967
rect 60507 39964 60519 39967
rect 60734 39964 60740 39976
rect 60507 39936 60740 39964
rect 60507 39933 60519 39936
rect 60461 39927 60519 39933
rect 60734 39924 60740 39936
rect 60792 39924 60798 39976
rect 63681 39967 63739 39973
rect 63681 39933 63693 39967
rect 63727 39964 63739 39967
rect 65536 39964 65564 39995
rect 66806 39992 66812 40004
rect 66864 39992 66870 40044
rect 67266 40032 67272 40044
rect 67227 40004 67272 40032
rect 67266 39992 67272 40004
rect 67324 39992 67330 40044
rect 67726 39992 67732 40044
rect 67784 40032 67790 40044
rect 68370 40032 68376 40044
rect 67784 40004 68376 40032
rect 67784 39992 67790 40004
rect 68370 39992 68376 40004
rect 68428 40032 68434 40044
rect 69201 40035 69259 40041
rect 69201 40032 69213 40035
rect 68428 40004 69213 40032
rect 68428 39992 68434 40004
rect 69201 40001 69213 40004
rect 69247 40032 69259 40035
rect 69382 40032 69388 40044
rect 69247 40004 69388 40032
rect 69247 40001 69259 40004
rect 69201 39995 69259 40001
rect 69382 39992 69388 40004
rect 69440 39992 69446 40044
rect 69934 40032 69940 40044
rect 69895 40004 69940 40032
rect 69934 39992 69940 40004
rect 69992 39992 69998 40044
rect 70302 39992 70308 40044
rect 70360 40032 70366 40044
rect 70489 40035 70547 40041
rect 70489 40032 70501 40035
rect 70360 40004 70501 40032
rect 70360 39992 70366 40004
rect 70489 40001 70501 40004
rect 70535 40032 70547 40035
rect 70765 40035 70823 40041
rect 70765 40032 70777 40035
rect 70535 40004 70777 40032
rect 70535 40001 70547 40004
rect 70489 39995 70547 40001
rect 70765 40001 70777 40004
rect 70811 40032 70823 40035
rect 74460 40032 74488 40072
rect 70811 40004 74304 40032
rect 70811 40001 70823 40004
rect 70765 39995 70823 40001
rect 63727 39936 65564 39964
rect 67284 39964 67312 39992
rect 67453 39967 67511 39973
rect 67453 39964 67465 39967
rect 67284 39936 67465 39964
rect 63727 39933 63739 39936
rect 63681 39927 63739 39933
rect 67453 39933 67465 39936
rect 67499 39933 67511 39967
rect 67453 39927 67511 39933
rect 67545 39967 67603 39973
rect 67545 39933 67557 39967
rect 67591 39964 67603 39967
rect 68462 39964 68468 39976
rect 67591 39936 68468 39964
rect 67591 39933 67603 39936
rect 67545 39927 67603 39933
rect 68462 39924 68468 39936
rect 68520 39924 68526 39976
rect 70026 39924 70032 39976
rect 70084 39964 70090 39976
rect 70084 39936 70129 39964
rect 70084 39924 70090 39936
rect 70394 39924 70400 39976
rect 70452 39964 70458 39976
rect 71406 39964 71412 39976
rect 70452 39936 70497 39964
rect 71367 39936 71412 39964
rect 70452 39924 70458 39936
rect 71406 39924 71412 39936
rect 71464 39924 71470 39976
rect 71866 39924 71872 39976
rect 71924 39964 71930 39976
rect 72881 39967 72939 39973
rect 72881 39964 72893 39967
rect 71924 39936 72893 39964
rect 71924 39924 71930 39936
rect 72881 39933 72893 39936
rect 72927 39933 72939 39967
rect 74169 39967 74227 39973
rect 74169 39964 74181 39967
rect 72881 39927 72939 39933
rect 73908 39936 74181 39964
rect 68554 39896 68560 39908
rect 64708 39868 68560 39896
rect 64708 39828 64736 39868
rect 68554 39856 68560 39868
rect 68612 39856 68618 39908
rect 69382 39896 69388 39908
rect 69343 39868 69388 39896
rect 69382 39856 69388 39868
rect 69440 39856 69446 39908
rect 55600 39800 64736 39828
rect 55125 39791 55183 39797
rect 64782 39788 64788 39840
rect 64840 39828 64846 39840
rect 65061 39831 65119 39837
rect 65061 39828 65073 39831
rect 64840 39800 65073 39828
rect 64840 39788 64846 39800
rect 65061 39797 65073 39800
rect 65107 39797 65119 39831
rect 65061 39791 65119 39797
rect 67174 39788 67180 39840
rect 67232 39828 67238 39840
rect 69658 39828 69664 39840
rect 67232 39800 69664 39828
rect 67232 39788 67238 39800
rect 69658 39788 69664 39800
rect 69716 39788 69722 39840
rect 70946 39828 70952 39840
rect 70907 39800 70952 39828
rect 70946 39788 70952 39800
rect 71004 39788 71010 39840
rect 71682 39788 71688 39840
rect 71740 39828 71746 39840
rect 73908 39837 73936 39936
rect 74169 39933 74181 39936
rect 74215 39933 74227 39967
rect 74169 39927 74227 39933
rect 73065 39831 73123 39837
rect 73065 39828 73077 39831
rect 71740 39800 73077 39828
rect 71740 39788 71746 39800
rect 73065 39797 73077 39800
rect 73111 39828 73123 39831
rect 73893 39831 73951 39837
rect 73893 39828 73905 39831
rect 73111 39800 73905 39828
rect 73111 39797 73123 39800
rect 73065 39791 73123 39797
rect 73893 39797 73905 39800
rect 73939 39797 73951 39831
rect 74276 39828 74304 40004
rect 74368 40004 74488 40032
rect 74368 39973 74396 40004
rect 74534 39992 74540 40044
rect 74592 40032 74598 40044
rect 74905 40035 74963 40041
rect 74905 40032 74917 40035
rect 74592 40004 74917 40032
rect 74592 39992 74598 40004
rect 74905 40001 74917 40004
rect 74951 40001 74963 40035
rect 75012 40032 75040 40072
rect 77662 40032 77668 40044
rect 75012 40004 77668 40032
rect 74905 39995 74963 40001
rect 77662 39992 77668 40004
rect 77720 39992 77726 40044
rect 74353 39967 74411 39973
rect 74353 39933 74365 39967
rect 74399 39933 74411 39967
rect 74353 39927 74411 39933
rect 74445 39967 74503 39973
rect 74445 39933 74457 39967
rect 74491 39964 74503 39967
rect 75178 39964 75184 39976
rect 74491 39936 75184 39964
rect 74491 39933 74503 39936
rect 74445 39927 74503 39933
rect 75178 39924 75184 39936
rect 75236 39924 75242 39976
rect 75822 39964 75828 39976
rect 75783 39936 75828 39964
rect 75822 39924 75828 39936
rect 75880 39964 75886 39976
rect 76101 39967 76159 39973
rect 76101 39964 76113 39967
rect 75880 39936 76113 39964
rect 75880 39924 75886 39936
rect 76101 39933 76113 39936
rect 76147 39933 76159 39967
rect 77021 39967 77079 39973
rect 77021 39964 77033 39967
rect 76101 39927 76159 39933
rect 76668 39936 77033 39964
rect 76190 39896 76196 39908
rect 74460 39868 76196 39896
rect 74460 39828 74488 39868
rect 76190 39856 76196 39868
rect 76248 39856 76254 39908
rect 76668 39840 76696 39936
rect 77021 39933 77033 39936
rect 77067 39933 77079 39967
rect 77772 39964 77800 40140
rect 78122 40128 78128 40180
rect 78180 40168 78186 40180
rect 78401 40171 78459 40177
rect 78401 40168 78413 40171
rect 78180 40140 78413 40168
rect 78180 40128 78186 40140
rect 78401 40137 78413 40140
rect 78447 40137 78459 40171
rect 78401 40131 78459 40137
rect 83642 40128 83648 40180
rect 83700 40168 83706 40180
rect 83921 40171 83979 40177
rect 83921 40168 83933 40171
rect 83700 40140 83933 40168
rect 83700 40128 83706 40140
rect 83921 40137 83933 40140
rect 83967 40137 83979 40171
rect 83921 40131 83979 40137
rect 78030 40060 78036 40112
rect 78088 40100 78094 40112
rect 84746 40100 84752 40112
rect 78088 40072 84752 40100
rect 78088 40060 78094 40072
rect 84746 40060 84752 40072
rect 84804 40060 84810 40112
rect 78217 39967 78275 39973
rect 78217 39964 78229 39967
rect 77772 39936 78229 39964
rect 77021 39927 77079 39933
rect 78217 39933 78229 39936
rect 78263 39964 78275 39967
rect 78585 39967 78643 39973
rect 78585 39964 78597 39967
rect 78263 39936 78597 39964
rect 78263 39933 78275 39936
rect 78217 39927 78275 39933
rect 78585 39933 78597 39936
rect 78631 39964 78643 39967
rect 79870 39964 79876 39976
rect 78631 39936 79876 39964
rect 78631 39933 78643 39936
rect 78585 39927 78643 39933
rect 79870 39924 79876 39936
rect 79928 39924 79934 39976
rect 79965 39967 80023 39973
rect 79965 39933 79977 39967
rect 80011 39964 80023 39967
rect 80238 39964 80244 39976
rect 80011 39936 80244 39964
rect 80011 39933 80023 39936
rect 79965 39927 80023 39933
rect 80238 39924 80244 39936
rect 80296 39924 80302 39976
rect 83734 39924 83740 39976
rect 83792 39964 83798 39976
rect 83829 39967 83887 39973
rect 83829 39964 83841 39967
rect 83792 39936 83841 39964
rect 83792 39924 83798 39936
rect 83829 39933 83841 39936
rect 83875 39933 83887 39967
rect 83829 39927 83887 39933
rect 85206 39924 85212 39976
rect 85264 39964 85270 39976
rect 85577 39967 85635 39973
rect 85577 39964 85589 39967
rect 85264 39936 85589 39964
rect 85264 39924 85270 39936
rect 85577 39933 85589 39936
rect 85623 39964 85635 39967
rect 86037 39967 86095 39973
rect 86037 39964 86049 39967
rect 85623 39936 86049 39964
rect 85623 39933 85635 39936
rect 85577 39927 85635 39933
rect 86037 39933 86049 39936
rect 86083 39933 86095 39967
rect 86037 39927 86095 39933
rect 76837 39899 76895 39905
rect 76837 39865 76849 39899
rect 76883 39865 76895 39899
rect 77386 39896 77392 39908
rect 77347 39868 77392 39896
rect 76837 39859 76895 39865
rect 74276 39800 74488 39828
rect 73893 39791 73951 39797
rect 75822 39788 75828 39840
rect 75880 39828 75886 39840
rect 75917 39831 75975 39837
rect 75917 39828 75929 39831
rect 75880 39800 75929 39828
rect 75880 39788 75886 39800
rect 75917 39797 75929 39800
rect 75963 39797 75975 39831
rect 76650 39828 76656 39840
rect 76611 39800 76656 39828
rect 75917 39791 75975 39797
rect 76650 39788 76656 39800
rect 76708 39788 76714 39840
rect 76852 39828 76880 39859
rect 77386 39856 77392 39868
rect 77444 39856 77450 39908
rect 85390 39896 85396 39908
rect 85351 39868 85396 39896
rect 85390 39856 85396 39868
rect 85448 39856 85454 39908
rect 85942 39896 85948 39908
rect 85903 39868 85948 39896
rect 85942 39856 85948 39868
rect 86000 39856 86006 39908
rect 77018 39828 77024 39840
rect 76852 39800 77024 39828
rect 77018 39788 77024 39800
rect 77076 39788 77082 39840
rect 79594 39788 79600 39840
rect 79652 39828 79658 39840
rect 80057 39831 80115 39837
rect 80057 39828 80069 39831
rect 79652 39800 80069 39828
rect 79652 39788 79658 39800
rect 80057 39797 80069 39800
rect 80103 39797 80115 39831
rect 80057 39791 80115 39797
rect 1104 39738 111136 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 50326 39738
rect 50378 39686 50390 39738
rect 50442 39686 50454 39738
rect 50506 39686 50518 39738
rect 50570 39686 81046 39738
rect 81098 39686 81110 39738
rect 81162 39686 81174 39738
rect 81226 39686 81238 39738
rect 81290 39686 111136 39738
rect 1104 39664 111136 39686
rect 5534 39584 5540 39636
rect 5592 39624 5598 39636
rect 5629 39627 5687 39633
rect 5629 39624 5641 39627
rect 5592 39596 5641 39624
rect 5592 39584 5598 39596
rect 5629 39593 5641 39596
rect 5675 39593 5687 39627
rect 5629 39587 5687 39593
rect 8018 39584 8024 39636
rect 8076 39624 8082 39636
rect 8076 39596 26924 39624
rect 8076 39584 8082 39596
rect 11698 39556 11704 39568
rect 5184 39528 10916 39556
rect 5184 39497 5212 39528
rect 4617 39491 4675 39497
rect 4617 39457 4629 39491
rect 4663 39488 4675 39491
rect 5169 39491 5227 39497
rect 5169 39488 5181 39491
rect 4663 39460 5181 39488
rect 4663 39457 4675 39460
rect 4617 39451 4675 39457
rect 5169 39457 5181 39460
rect 5215 39457 5227 39491
rect 5169 39451 5227 39457
rect 5353 39491 5411 39497
rect 5353 39457 5365 39491
rect 5399 39488 5411 39491
rect 5810 39488 5816 39500
rect 5399 39460 5816 39488
rect 5399 39457 5411 39460
rect 5353 39451 5411 39457
rect 5810 39448 5816 39460
rect 5868 39488 5874 39500
rect 10888 39497 10916 39528
rect 11440 39528 11704 39556
rect 11440 39497 11468 39528
rect 11698 39516 11704 39528
rect 11756 39516 11762 39568
rect 11977 39559 12035 39565
rect 11977 39525 11989 39559
rect 12023 39556 12035 39559
rect 12710 39556 12716 39568
rect 12023 39528 12716 39556
rect 12023 39525 12035 39528
rect 11977 39519 12035 39525
rect 12710 39516 12716 39528
rect 12768 39516 12774 39568
rect 12986 39556 12992 39568
rect 12947 39528 12992 39556
rect 12986 39516 12992 39528
rect 13044 39516 13050 39568
rect 17402 39516 17408 39568
rect 17460 39556 17466 39568
rect 18969 39559 19027 39565
rect 18969 39556 18981 39559
rect 17460 39528 18981 39556
rect 17460 39516 17466 39528
rect 18969 39525 18981 39528
rect 19015 39556 19027 39559
rect 26510 39556 26516 39568
rect 19015 39528 26372 39556
rect 26471 39528 26516 39556
rect 19015 39525 19027 39528
rect 18969 39519 19027 39525
rect 10873 39491 10931 39497
rect 5868 39460 6040 39488
rect 5868 39448 5874 39460
rect 4433 39423 4491 39429
rect 4433 39420 4445 39423
rect 4264 39392 4445 39420
rect 3602 39244 3608 39296
rect 3660 39284 3666 39296
rect 4264 39293 4292 39392
rect 4433 39389 4445 39392
rect 4479 39389 4491 39423
rect 4433 39383 4491 39389
rect 6012 39361 6040 39460
rect 10873 39457 10885 39491
rect 10919 39488 10931 39491
rect 11425 39491 11483 39497
rect 11425 39488 11437 39491
rect 10919 39460 11437 39488
rect 10919 39457 10931 39460
rect 10873 39451 10931 39457
rect 11425 39457 11437 39460
rect 11471 39457 11483 39491
rect 11425 39451 11483 39457
rect 11609 39491 11667 39497
rect 11609 39457 11621 39491
rect 11655 39488 11667 39491
rect 12618 39488 12624 39500
rect 11655 39460 12624 39488
rect 11655 39457 11667 39460
rect 11609 39451 11667 39457
rect 12618 39448 12624 39460
rect 12676 39448 12682 39500
rect 12894 39488 12900 39500
rect 12855 39460 12900 39488
rect 12894 39448 12900 39460
rect 12952 39448 12958 39500
rect 16390 39488 16396 39500
rect 16351 39460 16396 39488
rect 16390 39448 16396 39460
rect 16448 39448 16454 39500
rect 16500 39460 16804 39488
rect 9766 39380 9772 39432
rect 9824 39420 9830 39432
rect 10505 39423 10563 39429
rect 10505 39420 10517 39423
rect 9824 39392 10517 39420
rect 9824 39380 9830 39392
rect 10505 39389 10517 39392
rect 10551 39420 10563 39423
rect 10689 39423 10747 39429
rect 10689 39420 10701 39423
rect 10551 39392 10701 39420
rect 10551 39389 10563 39392
rect 10505 39383 10563 39389
rect 10689 39389 10701 39392
rect 10735 39389 10747 39423
rect 10689 39383 10747 39389
rect 12713 39423 12771 39429
rect 12713 39389 12725 39423
rect 12759 39420 12771 39423
rect 12912 39420 12940 39448
rect 12759 39392 12940 39420
rect 12759 39389 12771 39392
rect 12713 39383 12771 39389
rect 15746 39380 15752 39432
rect 15804 39420 15810 39432
rect 16500 39420 16528 39460
rect 16666 39420 16672 39432
rect 15804 39392 16528 39420
rect 16627 39392 16672 39420
rect 15804 39380 15810 39392
rect 16666 39380 16672 39392
rect 16724 39380 16730 39432
rect 16776 39420 16804 39460
rect 18230 39448 18236 39500
rect 18288 39488 18294 39500
rect 18877 39491 18935 39497
rect 18877 39488 18889 39491
rect 18288 39460 18889 39488
rect 18288 39448 18294 39460
rect 18877 39457 18889 39460
rect 18923 39457 18935 39491
rect 18877 39451 18935 39457
rect 23290 39448 23296 39500
rect 23348 39488 23354 39500
rect 23431 39491 23489 39497
rect 23431 39488 23443 39491
rect 23348 39460 23443 39488
rect 23348 39448 23354 39460
rect 23431 39457 23443 39460
rect 23477 39457 23489 39491
rect 23566 39488 23572 39500
rect 23527 39460 23572 39488
rect 23431 39451 23489 39457
rect 23566 39448 23572 39460
rect 23624 39448 23630 39500
rect 23934 39488 23940 39500
rect 23895 39460 23940 39488
rect 23934 39448 23940 39460
rect 23992 39448 23998 39500
rect 24029 39491 24087 39497
rect 24029 39457 24041 39491
rect 24075 39488 24087 39491
rect 24075 39460 24808 39488
rect 24075 39457 24087 39460
rect 24029 39451 24087 39457
rect 19334 39420 19340 39432
rect 16776 39392 19340 39420
rect 19334 39380 19340 39392
rect 19392 39380 19398 39432
rect 22922 39380 22928 39432
rect 22980 39420 22986 39432
rect 23017 39423 23075 39429
rect 23017 39420 23029 39423
rect 22980 39392 23029 39420
rect 22980 39380 22986 39392
rect 23017 39389 23029 39392
rect 23063 39420 23075 39423
rect 23584 39420 23612 39448
rect 23063 39392 23612 39420
rect 24780 39420 24808 39460
rect 24854 39448 24860 39500
rect 24912 39488 24918 39500
rect 25038 39488 25044 39500
rect 24912 39460 24957 39488
rect 24999 39460 25044 39488
rect 24912 39448 24918 39460
rect 25038 39448 25044 39460
rect 25096 39448 25102 39500
rect 26344 39488 26372 39528
rect 26510 39516 26516 39528
rect 26568 39516 26574 39568
rect 26896 39556 26924 39596
rect 29822 39584 29828 39636
rect 29880 39624 29886 39636
rect 30558 39624 30564 39636
rect 29880 39596 30564 39624
rect 29880 39584 29886 39596
rect 30558 39584 30564 39596
rect 30616 39624 30622 39636
rect 30616 39596 31340 39624
rect 30616 39584 30622 39596
rect 31018 39556 31024 39568
rect 26896 39528 31024 39556
rect 31018 39516 31024 39528
rect 31076 39516 31082 39568
rect 31312 39556 31340 39596
rect 31386 39584 31392 39636
rect 31444 39624 31450 39636
rect 34793 39627 34851 39633
rect 34793 39624 34805 39627
rect 31444 39596 34805 39624
rect 31444 39584 31450 39596
rect 34793 39593 34805 39596
rect 34839 39593 34851 39627
rect 34793 39587 34851 39593
rect 31312 39528 31432 39556
rect 26970 39488 26976 39500
rect 26344 39460 26976 39488
rect 26970 39448 26976 39460
rect 27028 39448 27034 39500
rect 29822 39488 29828 39500
rect 29783 39460 29828 39488
rect 29822 39448 29828 39460
rect 29880 39448 29886 39500
rect 29914 39448 29920 39500
rect 29972 39488 29978 39500
rect 30285 39491 30343 39497
rect 30285 39488 30297 39491
rect 29972 39460 30297 39488
rect 29972 39448 29978 39460
rect 30285 39457 30297 39460
rect 30331 39457 30343 39491
rect 30285 39451 30343 39457
rect 30377 39491 30435 39497
rect 30377 39457 30389 39491
rect 30423 39488 30435 39491
rect 31110 39488 31116 39500
rect 30423 39460 31116 39488
rect 30423 39457 30435 39460
rect 30377 39451 30435 39457
rect 31110 39448 31116 39460
rect 31168 39448 31174 39500
rect 31404 39497 31432 39528
rect 31389 39491 31447 39497
rect 31389 39457 31401 39491
rect 31435 39488 31447 39491
rect 32214 39488 32220 39500
rect 31435 39460 32220 39488
rect 31435 39457 31447 39460
rect 31389 39451 31447 39457
rect 32214 39448 32220 39460
rect 32272 39448 32278 39500
rect 34808 39488 34836 39587
rect 36170 39584 36176 39636
rect 36228 39624 36234 39636
rect 36814 39624 36820 39636
rect 36228 39596 36820 39624
rect 36228 39584 36234 39596
rect 36814 39584 36820 39596
rect 36872 39584 36878 39636
rect 38470 39584 38476 39636
rect 38528 39624 38534 39636
rect 38528 39596 69612 39624
rect 38528 39584 38534 39596
rect 35526 39516 35532 39568
rect 35584 39556 35590 39568
rect 36449 39559 36507 39565
rect 35584 39528 36216 39556
rect 35584 39516 35590 39528
rect 35161 39491 35219 39497
rect 35161 39488 35173 39491
rect 34808 39460 35173 39488
rect 35161 39457 35173 39460
rect 35207 39457 35219 39491
rect 35342 39488 35348 39500
rect 35303 39460 35348 39488
rect 35161 39451 35219 39457
rect 35342 39448 35348 39460
rect 35400 39448 35406 39500
rect 35802 39488 35808 39500
rect 35452 39460 35808 39488
rect 25056 39420 25084 39448
rect 26878 39420 26884 39432
rect 24780 39392 25084 39420
rect 26839 39392 26884 39420
rect 23063 39389 23075 39392
rect 23017 39383 23075 39389
rect 26878 39380 26884 39392
rect 26936 39380 26942 39432
rect 27246 39420 27252 39432
rect 27207 39392 27252 39420
rect 27246 39380 27252 39392
rect 27304 39380 27310 39432
rect 29730 39420 29736 39432
rect 29691 39392 29736 39420
rect 29730 39380 29736 39392
rect 29788 39380 29794 39432
rect 31205 39423 31263 39429
rect 31205 39389 31217 39423
rect 31251 39420 31263 39423
rect 31754 39420 31760 39432
rect 31251 39392 31760 39420
rect 31251 39389 31263 39392
rect 31205 39383 31263 39389
rect 31754 39380 31760 39392
rect 31812 39420 31818 39432
rect 34146 39420 34152 39432
rect 31812 39392 34152 39420
rect 31812 39380 31818 39392
rect 34146 39380 34152 39392
rect 34204 39380 34210 39432
rect 35452 39420 35480 39460
rect 35802 39448 35808 39460
rect 35860 39448 35866 39500
rect 35897 39491 35955 39497
rect 35897 39457 35909 39491
rect 35943 39488 35955 39491
rect 36078 39488 36084 39500
rect 35943 39460 36084 39488
rect 35943 39457 35955 39460
rect 35897 39451 35955 39457
rect 36078 39448 36084 39460
rect 36136 39448 36142 39500
rect 36188 39488 36216 39528
rect 36449 39525 36461 39559
rect 36495 39556 36507 39559
rect 38562 39556 38568 39568
rect 36495 39528 38568 39556
rect 36495 39525 36507 39528
rect 36449 39519 36507 39525
rect 38562 39516 38568 39528
rect 38620 39516 38626 39568
rect 42337 39559 42395 39565
rect 42337 39525 42349 39559
rect 42383 39556 42395 39559
rect 43714 39556 43720 39568
rect 42383 39528 43720 39556
rect 42383 39525 42395 39528
rect 42337 39519 42395 39525
rect 43714 39516 43720 39528
rect 43772 39516 43778 39568
rect 43806 39516 43812 39568
rect 43864 39556 43870 39568
rect 44634 39556 44640 39568
rect 43864 39528 44404 39556
rect 44595 39528 44640 39556
rect 43864 39516 43870 39528
rect 40862 39488 40868 39500
rect 36188 39460 40868 39488
rect 40862 39448 40868 39460
rect 40920 39448 40926 39500
rect 41233 39491 41291 39497
rect 41233 39457 41245 39491
rect 41279 39488 41291 39491
rect 41690 39488 41696 39500
rect 41279 39460 41460 39488
rect 41651 39460 41696 39488
rect 41279 39457 41291 39460
rect 41233 39451 41291 39457
rect 36630 39420 36636 39432
rect 34992 39392 35480 39420
rect 36591 39392 36636 39420
rect 5997 39355 6055 39361
rect 5997 39321 6009 39355
rect 6043 39352 6055 39355
rect 8754 39352 8760 39364
rect 6043 39324 8760 39352
rect 6043 39321 6055 39324
rect 5997 39315 6055 39321
rect 8754 39312 8760 39324
rect 8812 39352 8818 39364
rect 8812 39324 10548 39352
rect 8812 39312 8818 39324
rect 4249 39287 4307 39293
rect 4249 39284 4261 39287
rect 3660 39256 4261 39284
rect 3660 39244 3666 39256
rect 4249 39253 4261 39256
rect 4295 39253 4307 39287
rect 10520 39284 10548 39324
rect 10594 39312 10600 39364
rect 10652 39352 10658 39364
rect 10870 39352 10876 39364
rect 10652 39324 10876 39352
rect 10652 39312 10658 39324
rect 10870 39312 10876 39324
rect 10928 39312 10934 39364
rect 34606 39352 34612 39364
rect 17328 39324 34612 39352
rect 17328 39284 17356 39324
rect 34606 39312 34612 39324
rect 34664 39312 34670 39364
rect 10520 39256 17356 39284
rect 17957 39287 18015 39293
rect 4249 39247 4307 39253
rect 17957 39253 17969 39287
rect 18003 39284 18015 39287
rect 18046 39284 18052 39296
rect 18003 39256 18052 39284
rect 18003 39253 18015 39256
rect 17957 39247 18015 39253
rect 18046 39244 18052 39256
rect 18104 39244 18110 39296
rect 18233 39287 18291 39293
rect 18233 39253 18245 39287
rect 18279 39284 18291 39287
rect 18414 39284 18420 39296
rect 18279 39256 18420 39284
rect 18279 39253 18291 39256
rect 18233 39247 18291 39253
rect 18414 39244 18420 39256
rect 18472 39284 18478 39296
rect 18966 39284 18972 39296
rect 18472 39256 18972 39284
rect 18472 39244 18478 39256
rect 18966 39244 18972 39256
rect 19024 39244 19030 39296
rect 23201 39287 23259 39293
rect 23201 39253 23213 39287
rect 23247 39284 23259 39287
rect 23750 39284 23756 39296
rect 23247 39256 23756 39284
rect 23247 39253 23259 39256
rect 23201 39247 23259 39253
rect 23750 39244 23756 39256
rect 23808 39284 23814 39296
rect 23934 39284 23940 39296
rect 23808 39256 23940 39284
rect 23808 39244 23814 39256
rect 23934 39244 23940 39256
rect 23992 39244 23998 39296
rect 24489 39287 24547 39293
rect 24489 39253 24501 39287
rect 24535 39284 24547 39287
rect 25774 39284 25780 39296
rect 24535 39256 25780 39284
rect 24535 39253 24547 39256
rect 24489 39247 24547 39253
rect 25774 39244 25780 39256
rect 25832 39244 25838 39296
rect 26326 39244 26332 39296
rect 26384 39284 26390 39296
rect 26651 39287 26709 39293
rect 26651 39284 26663 39287
rect 26384 39256 26663 39284
rect 26384 39244 26390 39256
rect 26651 39253 26663 39256
rect 26697 39253 26709 39287
rect 26786 39284 26792 39296
rect 26747 39256 26792 39284
rect 26651 39247 26709 39253
rect 26786 39244 26792 39256
rect 26844 39244 26850 39296
rect 30834 39284 30840 39296
rect 30795 39256 30840 39284
rect 30834 39244 30840 39256
rect 30892 39244 30898 39296
rect 34698 39244 34704 39296
rect 34756 39284 34762 39296
rect 34992 39293 35020 39392
rect 36630 39380 36636 39392
rect 36688 39380 36694 39432
rect 37734 39380 37740 39432
rect 37792 39420 37798 39432
rect 40954 39420 40960 39432
rect 37792 39392 40960 39420
rect 37792 39380 37798 39392
rect 40954 39380 40960 39392
rect 41012 39380 41018 39432
rect 41141 39423 41199 39429
rect 41141 39389 41153 39423
rect 41187 39389 41199 39423
rect 41141 39383 41199 39389
rect 35066 39312 35072 39364
rect 35124 39352 35130 39364
rect 40865 39355 40923 39361
rect 40865 39352 40877 39355
rect 35124 39324 40877 39352
rect 35124 39312 35130 39324
rect 40865 39321 40877 39324
rect 40911 39352 40923 39355
rect 41156 39352 41184 39383
rect 40911 39324 41184 39352
rect 41432 39352 41460 39460
rect 41690 39448 41696 39460
rect 41748 39448 41754 39500
rect 41785 39491 41843 39497
rect 41785 39457 41797 39491
rect 41831 39488 41843 39491
rect 41831 39460 42288 39488
rect 41831 39457 41843 39460
rect 41785 39451 41843 39457
rect 42260 39432 42288 39460
rect 42426 39448 42432 39500
rect 42484 39488 42490 39500
rect 42484 39460 43484 39488
rect 42484 39448 42490 39460
rect 42242 39380 42248 39432
rect 42300 39380 42306 39432
rect 42797 39423 42855 39429
rect 42797 39389 42809 39423
rect 42843 39420 42855 39423
rect 42843 39392 43208 39420
rect 42843 39389 42855 39392
rect 42797 39383 42855 39389
rect 43180 39364 43208 39392
rect 43254 39380 43260 39432
rect 43312 39420 43318 39432
rect 43349 39423 43407 39429
rect 43349 39420 43361 39423
rect 43312 39392 43361 39420
rect 43312 39380 43318 39392
rect 43349 39389 43361 39392
rect 43395 39389 43407 39423
rect 43456 39420 43484 39460
rect 43530 39448 43536 39500
rect 43588 39488 43594 39500
rect 44082 39488 44088 39500
rect 43588 39460 44088 39488
rect 43588 39448 43594 39460
rect 44082 39448 44088 39460
rect 44140 39448 44146 39500
rect 44174 39448 44180 39500
rect 44232 39488 44238 39500
rect 44269 39491 44327 39497
rect 44269 39488 44281 39491
rect 44232 39460 44281 39488
rect 44232 39448 44238 39460
rect 44269 39457 44281 39460
rect 44315 39457 44327 39491
rect 44376 39488 44404 39528
rect 44634 39516 44640 39528
rect 44692 39516 44698 39568
rect 48682 39556 48688 39568
rect 44744 39528 48688 39556
rect 44744 39488 44772 39528
rect 48682 39516 48688 39528
rect 48740 39516 48746 39568
rect 49970 39516 49976 39568
rect 50028 39556 50034 39568
rect 51994 39556 52000 39568
rect 50028 39528 52000 39556
rect 50028 39516 50034 39528
rect 51994 39516 52000 39528
rect 52052 39516 52058 39568
rect 52181 39559 52239 39565
rect 52181 39525 52193 39559
rect 52227 39556 52239 39559
rect 53101 39559 53159 39565
rect 52227 39528 53052 39556
rect 52227 39525 52239 39528
rect 52181 39519 52239 39525
rect 44376 39460 44772 39488
rect 44269 39451 44327 39457
rect 44818 39448 44824 39500
rect 44876 39488 44882 39500
rect 44913 39491 44971 39497
rect 44913 39488 44925 39491
rect 44876 39460 44925 39488
rect 44876 39448 44882 39460
rect 44913 39457 44925 39460
rect 44959 39488 44971 39491
rect 45097 39491 45155 39497
rect 45097 39488 45109 39491
rect 44959 39460 45109 39488
rect 44959 39457 44971 39460
rect 44913 39451 44971 39457
rect 45097 39457 45109 39460
rect 45143 39488 45155 39491
rect 48774 39488 48780 39500
rect 45143 39460 48780 39488
rect 45143 39457 45155 39460
rect 45097 39451 45155 39457
rect 48774 39448 48780 39460
rect 48832 39448 48838 39500
rect 48958 39488 48964 39500
rect 48919 39460 48964 39488
rect 48958 39448 48964 39460
rect 49016 39488 49022 39500
rect 50709 39491 50767 39497
rect 50709 39488 50721 39491
rect 49016 39460 50721 39488
rect 49016 39448 49022 39460
rect 50709 39457 50721 39460
rect 50755 39488 50767 39491
rect 50982 39488 50988 39500
rect 50755 39460 50988 39488
rect 50755 39457 50767 39460
rect 50709 39451 50767 39457
rect 50982 39448 50988 39460
rect 51040 39448 51046 39500
rect 51718 39448 51724 39500
rect 51776 39488 51782 39500
rect 52089 39491 52147 39497
rect 52089 39488 52101 39491
rect 51776 39460 52101 39488
rect 51776 39448 51782 39460
rect 52089 39457 52101 39460
rect 52135 39488 52147 39491
rect 52546 39488 52552 39500
rect 52135 39460 52552 39488
rect 52135 39457 52147 39460
rect 52089 39451 52147 39457
rect 52546 39448 52552 39460
rect 52604 39488 52610 39500
rect 52822 39488 52828 39500
rect 52604 39460 52828 39488
rect 52604 39448 52610 39460
rect 52822 39448 52828 39460
rect 52880 39448 52886 39500
rect 53024 39488 53052 39528
rect 53101 39525 53113 39559
rect 53147 39556 53159 39559
rect 53190 39556 53196 39568
rect 53147 39528 53196 39556
rect 53147 39525 53159 39528
rect 53101 39519 53159 39525
rect 53190 39516 53196 39528
rect 53248 39516 53254 39568
rect 54018 39516 54024 39568
rect 54076 39556 54082 39568
rect 55309 39559 55367 39565
rect 55309 39556 55321 39559
rect 54076 39528 55321 39556
rect 54076 39516 54082 39528
rect 55309 39525 55321 39528
rect 55355 39525 55367 39559
rect 55309 39519 55367 39525
rect 55398 39516 55404 39568
rect 55456 39556 55462 39568
rect 55493 39559 55551 39565
rect 55493 39556 55505 39559
rect 55456 39528 55505 39556
rect 55456 39516 55462 39528
rect 55493 39525 55505 39528
rect 55539 39556 55551 39559
rect 56042 39556 56048 39568
rect 55539 39528 56048 39556
rect 55539 39525 55551 39528
rect 55493 39519 55551 39525
rect 56042 39516 56048 39528
rect 56100 39516 56106 39568
rect 61654 39556 61660 39568
rect 61615 39528 61660 39556
rect 61654 39516 61660 39528
rect 61712 39516 61718 39568
rect 66530 39516 66536 39568
rect 66588 39556 66594 39568
rect 68465 39559 68523 39565
rect 68465 39556 68477 39559
rect 66588 39528 68477 39556
rect 66588 39516 66594 39528
rect 68465 39525 68477 39528
rect 68511 39556 68523 39559
rect 69584 39556 69612 39596
rect 69658 39584 69664 39636
rect 69716 39624 69722 39636
rect 69716 39596 76144 39624
rect 69716 39584 69722 39596
rect 68511 39528 68692 39556
rect 69584 39528 75500 39556
rect 68511 39525 68523 39528
rect 68465 39519 68523 39525
rect 53285 39491 53343 39497
rect 53285 39488 53297 39491
rect 53024 39460 53297 39488
rect 53285 39457 53297 39460
rect 53331 39488 53343 39491
rect 53466 39488 53472 39500
rect 53331 39460 53472 39488
rect 53331 39457 53343 39460
rect 53285 39451 53343 39457
rect 53466 39448 53472 39460
rect 53524 39448 53530 39500
rect 53653 39491 53711 39497
rect 53653 39457 53665 39491
rect 53699 39488 53711 39491
rect 54754 39488 54760 39500
rect 53699 39460 54760 39488
rect 53699 39457 53711 39460
rect 53653 39451 53711 39457
rect 54754 39448 54760 39460
rect 54812 39448 54818 39500
rect 54846 39448 54852 39500
rect 54904 39488 54910 39500
rect 56413 39491 56471 39497
rect 54904 39460 54949 39488
rect 55876 39460 56272 39488
rect 54904 39448 54910 39460
rect 43714 39420 43720 39432
rect 43456 39392 43720 39420
rect 43349 39383 43407 39389
rect 43714 39380 43720 39392
rect 43772 39380 43778 39432
rect 44634 39380 44640 39432
rect 44692 39420 44698 39432
rect 48682 39420 48688 39432
rect 44692 39392 48688 39420
rect 44692 39380 44698 39392
rect 48682 39380 48688 39392
rect 48740 39380 48746 39432
rect 49234 39420 49240 39432
rect 49195 39392 49240 39420
rect 49234 39380 49240 39392
rect 49292 39380 49298 39432
rect 49326 39380 49332 39432
rect 49384 39420 49390 39432
rect 55876 39420 55904 39460
rect 56137 39423 56195 39429
rect 56137 39420 56149 39423
rect 49384 39392 55904 39420
rect 55968 39392 56149 39420
rect 49384 39380 49390 39392
rect 41598 39352 41604 39364
rect 41432 39324 41604 39352
rect 40911 39321 40923 39324
rect 40865 39315 40923 39321
rect 34977 39287 35035 39293
rect 34977 39284 34989 39287
rect 34756 39256 34989 39284
rect 34756 39244 34762 39256
rect 34977 39253 34989 39256
rect 35023 39253 35035 39287
rect 34977 39247 35035 39253
rect 35342 39244 35348 39296
rect 35400 39284 35406 39296
rect 36630 39284 36636 39296
rect 35400 39256 36636 39284
rect 35400 39244 35406 39256
rect 36630 39244 36636 39256
rect 36688 39244 36694 39296
rect 36906 39244 36912 39296
rect 36964 39284 36970 39296
rect 40954 39284 40960 39296
rect 36964 39256 40960 39284
rect 36964 39244 36970 39256
rect 40954 39244 40960 39256
rect 41012 39244 41018 39296
rect 41156 39284 41184 39324
rect 41598 39312 41604 39324
rect 41656 39352 41662 39364
rect 43162 39352 43168 39364
rect 41656 39324 42932 39352
rect 43075 39324 43168 39352
rect 41656 39312 41662 39324
rect 42904 39296 42932 39324
rect 43162 39312 43168 39324
rect 43220 39352 43226 39364
rect 43990 39352 43996 39364
rect 43220 39324 43996 39352
rect 43220 39312 43226 39324
rect 43990 39312 43996 39324
rect 44048 39312 44054 39364
rect 44082 39312 44088 39364
rect 44140 39352 44146 39364
rect 44818 39352 44824 39364
rect 44140 39324 44824 39352
rect 44140 39312 44146 39324
rect 44818 39312 44824 39324
rect 44876 39312 44882 39364
rect 55858 39352 55864 39364
rect 49896 39324 55864 39352
rect 41874 39284 41880 39296
rect 41156 39256 41880 39284
rect 41874 39244 41880 39256
rect 41932 39244 41938 39296
rect 42518 39244 42524 39296
rect 42576 39284 42582 39296
rect 42886 39284 42892 39296
rect 42576 39256 42621 39284
rect 42847 39256 42892 39284
rect 42576 39244 42582 39256
rect 42886 39244 42892 39256
rect 42944 39244 42950 39296
rect 43070 39284 43076 39296
rect 43031 39256 43076 39284
rect 43070 39244 43076 39256
rect 43128 39244 43134 39296
rect 44450 39244 44456 39296
rect 44508 39284 44514 39296
rect 49896 39284 49924 39324
rect 55858 39312 55864 39324
rect 55916 39312 55922 39364
rect 44508 39256 49924 39284
rect 44508 39244 44514 39256
rect 50154 39244 50160 39296
rect 50212 39284 50218 39296
rect 50341 39287 50399 39293
rect 50341 39284 50353 39287
rect 50212 39256 50353 39284
rect 50212 39244 50218 39256
rect 50341 39253 50353 39256
rect 50387 39253 50399 39287
rect 50341 39247 50399 39253
rect 54570 39244 54576 39296
rect 54628 39284 54634 39296
rect 55398 39284 55404 39296
rect 54628 39256 55404 39284
rect 54628 39244 54634 39256
rect 55398 39244 55404 39256
rect 55456 39244 55462 39296
rect 55490 39244 55496 39296
rect 55548 39284 55554 39296
rect 55968 39293 55996 39392
rect 56137 39389 56149 39392
rect 56183 39389 56195 39423
rect 56244 39420 56272 39460
rect 56413 39457 56425 39491
rect 56459 39488 56471 39491
rect 57330 39488 57336 39500
rect 56459 39460 57336 39488
rect 56459 39457 56471 39460
rect 56413 39451 56471 39457
rect 57330 39448 57336 39460
rect 57388 39448 57394 39500
rect 61838 39488 61844 39500
rect 61799 39460 61844 39488
rect 61838 39448 61844 39460
rect 61896 39448 61902 39500
rect 62206 39488 62212 39500
rect 62167 39460 62212 39488
rect 62206 39448 62212 39460
rect 62264 39448 62270 39500
rect 63034 39448 63040 39500
rect 63092 39488 63098 39500
rect 63221 39491 63279 39497
rect 63092 39460 63137 39488
rect 63092 39448 63098 39460
rect 63221 39457 63233 39491
rect 63267 39488 63279 39491
rect 63494 39488 63500 39500
rect 63267 39460 63500 39488
rect 63267 39457 63279 39460
rect 63221 39451 63279 39457
rect 63494 39448 63500 39460
rect 63552 39448 63558 39500
rect 64441 39491 64499 39497
rect 64441 39457 64453 39491
rect 64487 39488 64499 39491
rect 64598 39488 64604 39500
rect 64487 39460 64604 39488
rect 64487 39457 64499 39460
rect 64441 39451 64499 39457
rect 64598 39448 64604 39460
rect 64656 39448 64662 39500
rect 66714 39488 66720 39500
rect 66675 39460 66720 39488
rect 66714 39448 66720 39460
rect 66772 39448 66778 39500
rect 67634 39488 67640 39500
rect 67595 39460 67640 39488
rect 67634 39448 67640 39460
rect 67692 39488 67698 39500
rect 68664 39497 68692 39528
rect 67913 39491 67971 39497
rect 67913 39488 67925 39491
rect 67692 39460 67925 39488
rect 67692 39448 67698 39460
rect 67913 39457 67925 39460
rect 67959 39457 67971 39491
rect 67913 39451 67971 39457
rect 68649 39491 68707 39497
rect 68649 39457 68661 39491
rect 68695 39488 68707 39491
rect 69014 39488 69020 39500
rect 68695 39460 69020 39488
rect 68695 39457 68707 39460
rect 68649 39451 68707 39457
rect 65518 39420 65524 39432
rect 56244 39392 65524 39420
rect 56137 39383 56195 39389
rect 65518 39380 65524 39392
rect 65576 39380 65582 39432
rect 63218 39312 63224 39364
rect 63276 39352 63282 39364
rect 64509 39355 64567 39361
rect 64509 39352 64521 39355
rect 63276 39324 64521 39352
rect 63276 39312 63282 39324
rect 64509 39321 64521 39324
rect 64555 39321 64567 39355
rect 66530 39352 66536 39364
rect 66491 39324 66536 39352
rect 64509 39315 64567 39321
rect 66530 39312 66536 39324
rect 66588 39312 66594 39364
rect 67928 39352 67956 39451
rect 69014 39448 69020 39460
rect 69072 39448 69078 39500
rect 69382 39448 69388 39500
rect 69440 39488 69446 39500
rect 71409 39491 71467 39497
rect 71409 39488 71421 39491
rect 69440 39460 71421 39488
rect 69440 39448 69446 39460
rect 71409 39457 71421 39460
rect 71455 39457 71467 39491
rect 71409 39451 71467 39457
rect 68925 39423 68983 39429
rect 68925 39389 68937 39423
rect 68971 39420 68983 39423
rect 71501 39423 71559 39429
rect 71501 39420 71513 39423
rect 68971 39392 71513 39420
rect 68971 39389 68983 39392
rect 68925 39383 68983 39389
rect 71501 39389 71513 39392
rect 71547 39389 71559 39423
rect 71501 39383 71559 39389
rect 67928 39324 68600 39352
rect 55953 39287 56011 39293
rect 55953 39284 55965 39287
rect 55548 39256 55965 39284
rect 55548 39244 55554 39256
rect 55953 39253 55965 39256
rect 55999 39253 56011 39287
rect 55953 39247 56011 39253
rect 56042 39244 56048 39296
rect 56100 39284 56106 39296
rect 57517 39287 57575 39293
rect 57517 39284 57529 39287
rect 56100 39256 57529 39284
rect 56100 39244 56106 39256
rect 57517 39253 57529 39256
rect 57563 39253 57575 39287
rect 57517 39247 57575 39253
rect 61654 39244 61660 39296
rect 61712 39284 61718 39296
rect 62758 39284 62764 39296
rect 61712 39256 62764 39284
rect 61712 39244 61718 39256
rect 62758 39244 62764 39256
rect 62816 39284 62822 39296
rect 63313 39287 63371 39293
rect 63313 39284 63325 39287
rect 62816 39256 63325 39284
rect 62816 39244 62822 39256
rect 63313 39253 63325 39256
rect 63359 39253 63371 39287
rect 63313 39247 63371 39253
rect 63494 39244 63500 39296
rect 63552 39284 63558 39296
rect 63773 39287 63831 39293
rect 63773 39284 63785 39287
rect 63552 39256 63785 39284
rect 63552 39244 63558 39256
rect 63773 39253 63785 39256
rect 63819 39284 63831 39287
rect 64690 39284 64696 39296
rect 63819 39256 64696 39284
rect 63819 39253 63831 39256
rect 63773 39247 63831 39253
rect 64690 39244 64696 39256
rect 64748 39244 64754 39296
rect 67726 39284 67732 39296
rect 67687 39256 67732 39284
rect 67726 39244 67732 39256
rect 67784 39244 67790 39296
rect 68572 39284 68600 39324
rect 69934 39312 69940 39364
rect 69992 39352 69998 39364
rect 70946 39352 70952 39364
rect 69992 39324 70952 39352
rect 69992 39312 69998 39324
rect 70946 39312 70952 39324
rect 71004 39312 71010 39364
rect 75472 39352 75500 39528
rect 75822 39488 75828 39500
rect 75735 39460 75828 39488
rect 75822 39448 75828 39460
rect 75880 39448 75886 39500
rect 76116 39488 76144 39596
rect 76190 39584 76196 39636
rect 76248 39624 76254 39636
rect 79597 39627 79655 39633
rect 79597 39624 79609 39627
rect 76248 39596 79609 39624
rect 76248 39584 76254 39596
rect 79597 39593 79609 39596
rect 79643 39593 79655 39627
rect 80790 39624 80796 39636
rect 80751 39596 80796 39624
rect 79597 39587 79655 39593
rect 80790 39584 80796 39596
rect 80848 39584 80854 39636
rect 83568 39596 84792 39624
rect 76466 39516 76472 39568
rect 76524 39556 76530 39568
rect 83458 39556 83464 39568
rect 76524 39528 83464 39556
rect 76524 39516 76530 39528
rect 83458 39516 83464 39528
rect 83516 39556 83522 39568
rect 83568 39565 83596 39596
rect 83553 39559 83611 39565
rect 83553 39556 83565 39559
rect 83516 39528 83565 39556
rect 83516 39516 83522 39528
rect 83553 39525 83565 39528
rect 83599 39525 83611 39559
rect 83734 39556 83740 39568
rect 83695 39528 83740 39556
rect 83553 39519 83611 39525
rect 83734 39516 83740 39528
rect 83792 39516 83798 39568
rect 84764 39556 84792 39596
rect 85390 39584 85396 39636
rect 85448 39624 85454 39636
rect 86037 39627 86095 39633
rect 86037 39624 86049 39627
rect 85448 39596 86049 39624
rect 85448 39584 85454 39596
rect 86037 39593 86049 39596
rect 86083 39593 86095 39627
rect 86037 39587 86095 39593
rect 85577 39559 85635 39565
rect 85577 39556 85589 39559
rect 84764 39528 85589 39556
rect 77205 39491 77263 39497
rect 77205 39488 77217 39491
rect 76116 39460 77217 39488
rect 77205 39457 77217 39460
rect 77251 39488 77263 39491
rect 78030 39488 78036 39500
rect 77251 39460 78036 39488
rect 77251 39457 77263 39460
rect 77205 39451 77263 39457
rect 78030 39448 78036 39460
rect 78088 39448 78094 39500
rect 79134 39488 79140 39500
rect 79095 39460 79140 39488
rect 79134 39448 79140 39460
rect 79192 39448 79198 39500
rect 79410 39488 79416 39500
rect 79371 39460 79416 39488
rect 79410 39448 79416 39460
rect 79468 39448 79474 39500
rect 80698 39488 80704 39500
rect 80659 39460 80704 39488
rect 80698 39448 80704 39460
rect 80756 39448 80762 39500
rect 84378 39488 84384 39500
rect 84339 39460 84384 39488
rect 84378 39448 84384 39460
rect 84436 39448 84442 39500
rect 84764 39497 84792 39528
rect 85577 39525 85589 39528
rect 85623 39556 85635 39559
rect 85623 39528 85988 39556
rect 85623 39525 85635 39528
rect 85577 39519 85635 39525
rect 85960 39497 85988 39528
rect 84749 39491 84807 39497
rect 84749 39457 84761 39491
rect 84795 39457 84807 39491
rect 84749 39451 84807 39457
rect 84933 39491 84991 39497
rect 84933 39457 84945 39491
rect 84979 39488 84991 39491
rect 85761 39491 85819 39497
rect 85761 39488 85773 39491
rect 84979 39460 85773 39488
rect 84979 39457 84991 39460
rect 84933 39451 84991 39457
rect 85761 39457 85773 39460
rect 85807 39457 85819 39491
rect 85761 39451 85819 39457
rect 85945 39491 86003 39497
rect 85945 39457 85957 39491
rect 85991 39457 86003 39491
rect 85945 39451 86003 39457
rect 75840 39420 75868 39448
rect 77352 39423 77410 39429
rect 77352 39420 77364 39423
rect 75840 39392 77364 39420
rect 77352 39389 77364 39392
rect 77398 39389 77410 39423
rect 77352 39383 77410 39389
rect 77573 39423 77631 39429
rect 77573 39389 77585 39423
rect 77619 39389 77631 39423
rect 77573 39383 77631 39389
rect 77941 39423 77999 39429
rect 77941 39389 77953 39423
rect 77987 39420 77999 39423
rect 79229 39423 79287 39429
rect 79229 39420 79241 39423
rect 77987 39392 79241 39420
rect 77987 39389 77999 39392
rect 77941 39383 77999 39389
rect 79229 39389 79241 39392
rect 79275 39389 79287 39423
rect 84289 39423 84347 39429
rect 84289 39420 84301 39423
rect 79229 39383 79287 39389
rect 83384 39392 84301 39420
rect 76009 39355 76067 39361
rect 76009 39352 76021 39355
rect 75472 39324 76021 39352
rect 76009 39321 76021 39324
rect 76055 39352 76067 39355
rect 76466 39352 76472 39364
rect 76055 39324 76472 39352
rect 76055 39321 76067 39324
rect 76009 39315 76067 39321
rect 76466 39312 76472 39324
rect 76524 39312 76530 39364
rect 77481 39355 77539 39361
rect 77481 39352 77493 39355
rect 76760 39324 77493 39352
rect 70029 39287 70087 39293
rect 70029 39284 70041 39287
rect 68572 39256 70041 39284
rect 70029 39253 70041 39256
rect 70075 39253 70087 39287
rect 70029 39247 70087 39253
rect 76374 39244 76380 39296
rect 76432 39284 76438 39296
rect 76760 39293 76788 39324
rect 77481 39321 77493 39324
rect 77527 39321 77539 39355
rect 77481 39315 77539 39321
rect 76745 39287 76803 39293
rect 76745 39284 76757 39287
rect 76432 39256 76757 39284
rect 76432 39244 76438 39256
rect 76745 39253 76757 39256
rect 76791 39253 76803 39287
rect 76745 39247 76803 39253
rect 77113 39287 77171 39293
rect 77113 39253 77125 39287
rect 77159 39284 77171 39287
rect 77294 39284 77300 39296
rect 77159 39256 77300 39284
rect 77159 39253 77171 39256
rect 77113 39247 77171 39253
rect 77294 39244 77300 39256
rect 77352 39284 77358 39296
rect 77588 39284 77616 39383
rect 77352 39256 77616 39284
rect 77352 39244 77358 39256
rect 82906 39244 82912 39296
rect 82964 39284 82970 39296
rect 83384 39293 83412 39392
rect 84289 39389 84301 39392
rect 84335 39389 84347 39423
rect 84289 39383 84347 39389
rect 84010 39312 84016 39364
rect 84068 39352 84074 39364
rect 84948 39352 84976 39451
rect 84068 39324 84976 39352
rect 84068 39312 84074 39324
rect 83369 39287 83427 39293
rect 83369 39284 83381 39287
rect 82964 39256 83381 39284
rect 82964 39244 82970 39256
rect 83369 39253 83381 39256
rect 83415 39253 83427 39287
rect 83369 39247 83427 39253
rect 1104 39194 111136 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 65686 39194
rect 65738 39142 65750 39194
rect 65802 39142 65814 39194
rect 65866 39142 65878 39194
rect 65930 39142 96406 39194
rect 96458 39142 96470 39194
rect 96522 39142 96534 39194
rect 96586 39142 96598 39194
rect 96650 39142 111136 39194
rect 1104 39120 111136 39142
rect 3786 39040 3792 39092
rect 3844 39080 3850 39092
rect 9766 39080 9772 39092
rect 3844 39052 9772 39080
rect 3844 39040 3850 39052
rect 9766 39040 9772 39052
rect 9824 39040 9830 39092
rect 11514 39040 11520 39092
rect 11572 39080 11578 39092
rect 11701 39083 11759 39089
rect 11701 39080 11713 39083
rect 11572 39052 11713 39080
rect 11572 39040 11578 39052
rect 11701 39049 11713 39052
rect 11747 39080 11759 39083
rect 15473 39083 15531 39089
rect 11747 39052 15240 39080
rect 11747 39049 11759 39052
rect 11701 39043 11759 39049
rect 4062 38972 4068 39024
rect 4120 39012 4126 39024
rect 15010 39012 15016 39024
rect 4120 38984 15016 39012
rect 4120 38972 4126 38984
rect 15010 38972 15016 38984
rect 15068 38972 15074 39024
rect 15212 39012 15240 39052
rect 15473 39049 15485 39083
rect 15519 39080 15531 39083
rect 16666 39080 16672 39092
rect 15519 39052 16672 39080
rect 15519 39049 15531 39052
rect 15473 39043 15531 39049
rect 16666 39040 16672 39052
rect 16724 39040 16730 39092
rect 18141 39083 18199 39089
rect 18141 39049 18153 39083
rect 18187 39080 18199 39083
rect 18187 39052 26924 39080
rect 18187 39049 18199 39052
rect 18141 39043 18199 39049
rect 15841 39015 15899 39021
rect 15841 39012 15853 39015
rect 15212 38984 15853 39012
rect 15841 38981 15853 38984
rect 15887 39012 15899 39015
rect 18156 39012 18184 39043
rect 15887 38984 18184 39012
rect 15887 38981 15899 38984
rect 15841 38975 15899 38981
rect 14642 38944 14648 38956
rect 5736 38916 14648 38944
rect 2590 38836 2596 38888
rect 2648 38876 2654 38888
rect 2685 38879 2743 38885
rect 2685 38876 2697 38879
rect 2648 38848 2697 38876
rect 2648 38836 2654 38848
rect 2685 38845 2697 38848
rect 2731 38845 2743 38879
rect 2685 38839 2743 38845
rect 2961 38879 3019 38885
rect 2961 38845 2973 38879
rect 3007 38876 3019 38879
rect 5258 38876 5264 38888
rect 3007 38848 4108 38876
rect 5219 38848 5264 38876
rect 3007 38845 3019 38848
rect 2961 38839 3019 38845
rect 4080 38808 4108 38848
rect 5258 38836 5264 38848
rect 5316 38836 5322 38888
rect 5736 38885 5764 38916
rect 14642 38904 14648 38916
rect 14700 38904 14706 38956
rect 5721 38879 5779 38885
rect 5721 38845 5733 38879
rect 5767 38845 5779 38879
rect 5721 38839 5779 38845
rect 10781 38879 10839 38885
rect 10781 38845 10793 38879
rect 10827 38845 10839 38879
rect 10962 38876 10968 38888
rect 10923 38848 10968 38876
rect 10781 38839 10839 38845
rect 4080 38780 5304 38808
rect 4154 38700 4160 38752
rect 4212 38740 4218 38752
rect 4249 38743 4307 38749
rect 4249 38740 4261 38743
rect 4212 38712 4261 38740
rect 4212 38700 4218 38712
rect 4249 38709 4261 38712
rect 4295 38709 4307 38743
rect 4430 38740 4436 38752
rect 4391 38712 4436 38740
rect 4249 38703 4307 38709
rect 4430 38700 4436 38712
rect 4488 38700 4494 38752
rect 5276 38749 5304 38780
rect 9766 38768 9772 38820
rect 9824 38808 9830 38820
rect 10321 38811 10379 38817
rect 10321 38808 10333 38811
rect 9824 38780 10333 38808
rect 9824 38768 9830 38780
rect 10321 38777 10333 38780
rect 10367 38777 10379 38811
rect 10796 38808 10824 38839
rect 10962 38836 10968 38848
rect 11020 38836 11026 38888
rect 11238 38836 11244 38888
rect 11296 38876 11302 38888
rect 11333 38879 11391 38885
rect 11333 38876 11345 38879
rect 11296 38848 11345 38876
rect 11296 38836 11302 38848
rect 11333 38845 11345 38848
rect 11379 38845 11391 38879
rect 11514 38876 11520 38888
rect 11475 38848 11520 38876
rect 11333 38839 11391 38845
rect 11514 38836 11520 38848
rect 11572 38836 11578 38888
rect 13262 38836 13268 38888
rect 13320 38876 13326 38888
rect 14415 38879 14473 38885
rect 14415 38876 14427 38879
rect 13320 38848 14427 38876
rect 13320 38836 13326 38848
rect 14415 38845 14427 38848
rect 14461 38845 14473 38879
rect 14415 38839 14473 38845
rect 14553 38879 14611 38885
rect 14553 38845 14565 38879
rect 14599 38876 14611 38879
rect 14826 38876 14832 38888
rect 14599 38848 14832 38876
rect 14599 38845 14611 38848
rect 14553 38839 14611 38845
rect 14826 38836 14832 38848
rect 14884 38836 14890 38888
rect 15010 38876 15016 38888
rect 14971 38848 15016 38876
rect 15010 38836 15016 38848
rect 15068 38836 15074 38888
rect 15197 38879 15255 38885
rect 15197 38845 15209 38879
rect 15243 38845 15255 38879
rect 15197 38839 15255 38845
rect 11793 38811 11851 38817
rect 11793 38808 11805 38811
rect 10796 38780 11805 38808
rect 10321 38771 10379 38777
rect 11793 38777 11805 38780
rect 11839 38777 11851 38811
rect 11793 38771 11851 38777
rect 5261 38743 5319 38749
rect 5261 38709 5273 38743
rect 5307 38709 5319 38743
rect 11808 38740 11836 38771
rect 13998 38768 14004 38820
rect 14056 38808 14062 38820
rect 14093 38811 14151 38817
rect 14093 38808 14105 38811
rect 14056 38780 14105 38808
rect 14056 38768 14062 38780
rect 14093 38777 14105 38780
rect 14139 38777 14151 38811
rect 15212 38808 15240 38839
rect 15856 38808 15884 38975
rect 20438 38972 20444 39024
rect 20496 39012 20502 39024
rect 23842 39012 23848 39024
rect 20496 38984 23848 39012
rect 20496 38972 20502 38984
rect 23842 38972 23848 38984
rect 23900 38972 23906 39024
rect 25958 38972 25964 39024
rect 26016 39021 26022 39024
rect 26016 39015 26065 39021
rect 26016 38981 26019 39015
rect 26053 38981 26065 39015
rect 26016 38975 26065 38981
rect 26145 39015 26203 39021
rect 26145 38981 26157 39015
rect 26191 38981 26203 39015
rect 26145 38975 26203 38981
rect 26016 38972 26022 38975
rect 19334 38904 19340 38956
rect 19392 38944 19398 38956
rect 19705 38947 19763 38953
rect 19705 38944 19717 38947
rect 19392 38916 19717 38944
rect 19392 38904 19398 38916
rect 19705 38913 19717 38916
rect 19751 38913 19763 38947
rect 21174 38944 21180 38956
rect 19705 38907 19763 38913
rect 19812 38916 21180 38944
rect 16577 38879 16635 38885
rect 16577 38845 16589 38879
rect 16623 38876 16635 38879
rect 16666 38876 16672 38888
rect 16623 38848 16672 38876
rect 16623 38845 16635 38848
rect 16577 38839 16635 38845
rect 16666 38836 16672 38848
rect 16724 38876 16730 38888
rect 16942 38876 16948 38888
rect 16724 38848 16948 38876
rect 16724 38836 16730 38848
rect 16942 38836 16948 38848
rect 17000 38836 17006 38888
rect 18046 38876 18052 38888
rect 18007 38848 18052 38876
rect 18046 38836 18052 38848
rect 18104 38836 18110 38888
rect 18966 38836 18972 38888
rect 19024 38876 19030 38888
rect 19429 38879 19487 38885
rect 19429 38876 19441 38879
rect 19024 38848 19441 38876
rect 19024 38836 19030 38848
rect 19429 38845 19441 38848
rect 19475 38876 19487 38879
rect 19812 38876 19840 38916
rect 21174 38904 21180 38916
rect 21232 38904 21238 38956
rect 26160 38888 26188 38975
rect 26234 38904 26240 38956
rect 26292 38944 26298 38956
rect 26896 38944 26924 39052
rect 27430 39040 27436 39092
rect 27488 39080 27494 39092
rect 29730 39080 29736 39092
rect 27488 39052 29736 39080
rect 27488 39040 27494 39052
rect 29730 39040 29736 39052
rect 29788 39040 29794 39092
rect 29822 39040 29828 39092
rect 29880 39080 29886 39092
rect 31386 39080 31392 39092
rect 29880 39052 31392 39080
rect 29880 39040 29886 39052
rect 31386 39040 31392 39052
rect 31444 39040 31450 39092
rect 34606 39040 34612 39092
rect 34664 39080 34670 39092
rect 34664 39052 37872 39080
rect 34664 39040 34670 39052
rect 26970 38972 26976 39024
rect 27028 39012 27034 39024
rect 34698 39012 34704 39024
rect 27028 38984 34704 39012
rect 27028 38972 27034 38984
rect 34698 38972 34704 38984
rect 34756 38972 34762 39024
rect 37642 39012 37648 39024
rect 36648 38984 37648 39012
rect 34790 38944 34796 38956
rect 26292 38916 26337 38944
rect 26896 38916 34796 38944
rect 26292 38904 26298 38916
rect 34790 38904 34796 38916
rect 34848 38904 34854 38956
rect 23661 38879 23719 38885
rect 23661 38876 23673 38879
rect 19475 38848 19840 38876
rect 20824 38848 23673 38876
rect 19475 38845 19487 38848
rect 19429 38839 19487 38845
rect 15212 38780 15884 38808
rect 14093 38771 14151 38777
rect 20824 38752 20852 38848
rect 23661 38845 23673 38848
rect 23707 38845 23719 38879
rect 23842 38876 23848 38888
rect 23803 38848 23848 38876
rect 23661 38839 23719 38845
rect 23842 38836 23848 38848
rect 23900 38836 23906 38888
rect 24394 38876 24400 38888
rect 24355 38848 24400 38876
rect 24394 38836 24400 38848
rect 24452 38836 24458 38888
rect 24581 38879 24639 38885
rect 24581 38845 24593 38879
rect 24627 38876 24639 38879
rect 24762 38876 24768 38888
rect 24627 38848 24768 38876
rect 24627 38845 24639 38848
rect 24581 38839 24639 38845
rect 23477 38811 23535 38817
rect 23477 38777 23489 38811
rect 23523 38808 23535 38811
rect 23566 38808 23572 38820
rect 23523 38780 23572 38808
rect 23523 38777 23535 38780
rect 23477 38771 23535 38777
rect 23566 38768 23572 38780
rect 23624 38808 23630 38820
rect 24596 38808 24624 38839
rect 24762 38836 24768 38848
rect 24820 38836 24826 38888
rect 25222 38876 25228 38888
rect 25183 38848 25228 38876
rect 25222 38836 25228 38848
rect 25280 38836 25286 38888
rect 25774 38836 25780 38888
rect 25832 38876 25838 38888
rect 25869 38879 25927 38885
rect 25869 38876 25881 38879
rect 25832 38848 25881 38876
rect 25832 38836 25838 38848
rect 25869 38845 25881 38848
rect 25915 38845 25927 38879
rect 25869 38839 25927 38845
rect 26142 38836 26148 38888
rect 26200 38836 26206 38888
rect 26786 38836 26792 38888
rect 26844 38876 26850 38888
rect 29454 38876 29460 38888
rect 26844 38848 29460 38876
rect 26844 38836 26850 38848
rect 29454 38836 29460 38848
rect 29512 38836 29518 38888
rect 29638 38876 29644 38888
rect 29551 38848 29644 38876
rect 29638 38836 29644 38848
rect 29696 38876 29702 38888
rect 36648 38885 36676 38984
rect 37642 38972 37648 38984
rect 37700 38972 37706 39024
rect 37734 38944 37740 38956
rect 37695 38916 37740 38944
rect 37734 38904 37740 38916
rect 37792 38904 37798 38956
rect 37844 38944 37872 39052
rect 37918 39040 37924 39092
rect 37976 39080 37982 39092
rect 38197 39083 38255 39089
rect 38197 39080 38209 39083
rect 37976 39052 38209 39080
rect 37976 39040 37982 39052
rect 38197 39049 38209 39052
rect 38243 39080 38255 39083
rect 39482 39080 39488 39092
rect 38243 39052 39488 39080
rect 38243 39049 38255 39052
rect 38197 39043 38255 39049
rect 39482 39040 39488 39052
rect 39540 39080 39546 39092
rect 49326 39080 49332 39092
rect 39540 39052 49332 39080
rect 39540 39040 39546 39052
rect 49326 39040 49332 39052
rect 49384 39040 49390 39092
rect 53374 39040 53380 39092
rect 53432 39080 53438 39092
rect 54205 39083 54263 39089
rect 54205 39080 54217 39083
rect 53432 39052 54217 39080
rect 53432 39040 53438 39052
rect 54205 39049 54217 39052
rect 54251 39080 54263 39083
rect 62114 39080 62120 39092
rect 54251 39052 62120 39080
rect 54251 39049 54263 39052
rect 54205 39043 54263 39049
rect 62114 39040 62120 39052
rect 62172 39040 62178 39092
rect 67634 39080 67640 39092
rect 62224 39052 67640 39080
rect 41049 39015 41107 39021
rect 41049 38981 41061 39015
rect 41095 39012 41107 39015
rect 41095 38984 41828 39012
rect 41095 38981 41107 38984
rect 41049 38975 41107 38981
rect 41138 38944 41144 38956
rect 37844 38916 41144 38944
rect 41138 38904 41144 38916
rect 41196 38944 41202 38956
rect 41196 38916 41276 38944
rect 41196 38904 41202 38916
rect 36449 38879 36507 38885
rect 36449 38876 36461 38879
rect 29696 38848 36461 38876
rect 29696 38836 29702 38848
rect 36449 38845 36461 38848
rect 36495 38845 36507 38879
rect 36449 38839 36507 38845
rect 36633 38879 36691 38885
rect 36633 38845 36645 38879
rect 36679 38845 36691 38879
rect 37090 38876 37096 38888
rect 37051 38848 37096 38876
rect 36633 38839 36691 38845
rect 37090 38836 37096 38848
rect 37148 38836 37154 38888
rect 37185 38879 37243 38885
rect 37185 38845 37197 38879
rect 37231 38876 37243 38879
rect 38470 38876 38476 38888
rect 37231 38848 38476 38876
rect 37231 38845 37243 38848
rect 37185 38839 37243 38845
rect 38470 38836 38476 38848
rect 38528 38836 38534 38888
rect 41248 38876 41276 38916
rect 41417 38879 41475 38885
rect 41417 38876 41429 38879
rect 41248 38848 41429 38876
rect 41417 38845 41429 38848
rect 41463 38876 41475 38879
rect 41509 38879 41567 38885
rect 41509 38876 41521 38879
rect 41463 38848 41521 38876
rect 41463 38845 41475 38848
rect 41417 38839 41475 38845
rect 41509 38845 41521 38848
rect 41555 38845 41567 38879
rect 41509 38839 41567 38845
rect 41598 38836 41604 38888
rect 41656 38876 41662 38888
rect 41693 38879 41751 38885
rect 41693 38876 41705 38879
rect 41656 38848 41705 38876
rect 41656 38836 41662 38848
rect 41693 38845 41705 38848
rect 41739 38845 41751 38879
rect 41800 38876 41828 38984
rect 41874 38972 41880 39024
rect 41932 39012 41938 39024
rect 43349 39015 43407 39021
rect 43349 39012 43361 39015
rect 41932 38984 43361 39012
rect 41932 38972 41938 38984
rect 43349 38981 43361 38984
rect 43395 38981 43407 39015
rect 43530 39012 43536 39024
rect 43491 38984 43536 39012
rect 43349 38975 43407 38981
rect 43530 38972 43536 38984
rect 43588 38972 43594 39024
rect 43622 38972 43628 39024
rect 43680 39012 43686 39024
rect 43855 39015 43913 39021
rect 43855 39012 43867 39015
rect 43680 38984 43867 39012
rect 43680 38972 43686 38984
rect 43855 38981 43867 38984
rect 43901 38981 43913 39015
rect 43990 39012 43996 39024
rect 43951 38984 43996 39012
rect 43855 38975 43913 38981
rect 43990 38972 43996 38984
rect 44048 38972 44054 39024
rect 44361 39015 44419 39021
rect 44361 38981 44373 39015
rect 44407 39012 44419 39015
rect 44542 39012 44548 39024
rect 44407 38984 44548 39012
rect 44407 38981 44419 38984
rect 44361 38975 44419 38981
rect 44542 38972 44548 38984
rect 44600 38972 44606 39024
rect 48866 39012 48872 39024
rect 47504 38984 48872 39012
rect 42702 38944 42708 38956
rect 42663 38916 42708 38944
rect 42702 38904 42708 38916
rect 42760 38904 42766 38956
rect 43073 38947 43131 38953
rect 43073 38913 43085 38947
rect 43119 38944 43131 38947
rect 43162 38944 43168 38956
rect 43119 38916 43168 38944
rect 43119 38913 43131 38916
rect 43073 38907 43131 38913
rect 42153 38879 42211 38885
rect 42153 38876 42165 38879
rect 41800 38848 42165 38876
rect 41693 38839 41751 38845
rect 42153 38845 42165 38848
rect 42199 38845 42211 38879
rect 42153 38839 42211 38845
rect 42242 38836 42248 38888
rect 42300 38876 42306 38888
rect 43088 38876 43116 38907
rect 43162 38904 43168 38916
rect 43220 38904 43226 38956
rect 44085 38947 44143 38953
rect 44085 38913 44097 38947
rect 44131 38944 44143 38947
rect 44266 38944 44272 38956
rect 44131 38916 44272 38944
rect 44131 38913 44143 38916
rect 44085 38907 44143 38913
rect 44266 38904 44272 38916
rect 44324 38904 44330 38956
rect 47394 38944 47400 38956
rect 47355 38916 47400 38944
rect 47394 38904 47400 38916
rect 47452 38904 47458 38956
rect 42300 38848 43116 38876
rect 42300 38836 42306 38848
rect 43530 38836 43536 38888
rect 43588 38876 43594 38888
rect 47504 38885 47532 38984
rect 48866 38972 48872 38984
rect 48924 38972 48930 39024
rect 49053 39015 49111 39021
rect 49053 38981 49065 39015
rect 49099 39012 49111 39015
rect 49142 39012 49148 39024
rect 49099 38984 49148 39012
rect 49099 38981 49111 38984
rect 49053 38975 49111 38981
rect 49142 38972 49148 38984
rect 49200 39012 49206 39024
rect 49200 38984 54432 39012
rect 49200 38972 49206 38984
rect 43717 38879 43775 38885
rect 43717 38876 43729 38879
rect 43588 38848 43729 38876
rect 43588 38836 43594 38848
rect 43717 38845 43729 38848
rect 43763 38845 43775 38879
rect 43717 38839 43775 38845
rect 47489 38879 47547 38885
rect 47489 38845 47501 38879
rect 47535 38845 47547 38879
rect 47489 38839 47547 38845
rect 47578 38836 47584 38888
rect 47636 38876 47642 38888
rect 47949 38879 48007 38885
rect 47949 38876 47961 38879
rect 47636 38848 47961 38876
rect 47636 38836 47642 38848
rect 47949 38845 47961 38848
rect 47995 38845 48007 38879
rect 47949 38839 48007 38845
rect 48038 38836 48044 38888
rect 48096 38876 48102 38888
rect 52641 38879 52699 38885
rect 48096 38848 48141 38876
rect 48096 38836 48102 38848
rect 52641 38845 52653 38879
rect 52687 38845 52699 38879
rect 52641 38839 52699 38845
rect 23624 38780 24624 38808
rect 24949 38811 25007 38817
rect 23624 38768 23630 38780
rect 24949 38777 24961 38811
rect 24995 38808 25007 38811
rect 26050 38808 26056 38820
rect 24995 38780 26056 38808
rect 24995 38777 25007 38780
rect 24949 38771 25007 38777
rect 26050 38768 26056 38780
rect 26108 38768 26114 38820
rect 26602 38808 26608 38820
rect 26563 38780 26608 38808
rect 26602 38768 26608 38780
rect 26660 38768 26666 38820
rect 26694 38768 26700 38820
rect 26752 38808 26758 38820
rect 47854 38808 47860 38820
rect 26752 38780 47860 38808
rect 26752 38768 26758 38780
rect 47854 38768 47860 38780
rect 47912 38768 47918 38820
rect 52546 38768 52552 38820
rect 52604 38808 52610 38820
rect 52656 38808 52684 38839
rect 52822 38836 52828 38888
rect 52880 38876 52886 38888
rect 53282 38876 53288 38888
rect 52880 38848 52925 38876
rect 53243 38848 53288 38876
rect 52880 38836 52886 38848
rect 53282 38836 53288 38848
rect 53340 38836 53346 38888
rect 53374 38836 53380 38888
rect 53432 38876 53438 38888
rect 53432 38848 53477 38876
rect 53432 38836 53438 38848
rect 53558 38808 53564 38820
rect 52604 38780 53564 38808
rect 52604 38768 52610 38780
rect 53558 38768 53564 38780
rect 53616 38808 53622 38820
rect 54297 38811 54355 38817
rect 54297 38808 54309 38811
rect 53616 38780 54309 38808
rect 53616 38768 53622 38780
rect 54297 38777 54309 38780
rect 54343 38777 54355 38811
rect 54297 38771 54355 38777
rect 16574 38740 16580 38752
rect 11808 38712 16580 38740
rect 5261 38703 5319 38709
rect 16574 38700 16580 38712
rect 16632 38700 16638 38752
rect 16761 38743 16819 38749
rect 16761 38709 16773 38743
rect 16807 38740 16819 38743
rect 16850 38740 16856 38752
rect 16807 38712 16856 38740
rect 16807 38709 16819 38712
rect 16761 38703 16819 38709
rect 16850 38700 16856 38712
rect 16908 38700 16914 38752
rect 20806 38740 20812 38752
rect 20767 38712 20812 38740
rect 20806 38700 20812 38712
rect 20864 38700 20870 38752
rect 21174 38740 21180 38752
rect 21135 38712 21180 38740
rect 21174 38700 21180 38712
rect 21232 38700 21238 38752
rect 24394 38700 24400 38752
rect 24452 38740 24458 38752
rect 25406 38740 25412 38752
rect 24452 38712 25412 38740
rect 24452 38700 24458 38712
rect 25406 38700 25412 38712
rect 25464 38740 25470 38752
rect 34054 38740 34060 38752
rect 25464 38712 34060 38740
rect 25464 38700 25470 38712
rect 34054 38700 34060 38712
rect 34112 38700 34118 38752
rect 34146 38700 34152 38752
rect 34204 38740 34210 38752
rect 36906 38740 36912 38752
rect 34204 38712 36912 38740
rect 34204 38700 34210 38712
rect 36906 38700 36912 38712
rect 36964 38700 36970 38752
rect 38013 38743 38071 38749
rect 38013 38709 38025 38743
rect 38059 38740 38071 38743
rect 38470 38740 38476 38752
rect 38059 38712 38476 38740
rect 38059 38709 38071 38712
rect 38013 38703 38071 38709
rect 38470 38700 38476 38712
rect 38528 38700 38534 38752
rect 39574 38700 39580 38752
rect 39632 38740 39638 38752
rect 41049 38743 41107 38749
rect 41049 38740 41061 38743
rect 39632 38712 41061 38740
rect 39632 38700 39638 38712
rect 41049 38709 41061 38712
rect 41095 38740 41107 38743
rect 41141 38743 41199 38749
rect 41141 38740 41153 38743
rect 41095 38712 41153 38740
rect 41095 38709 41107 38712
rect 41049 38703 41107 38709
rect 41141 38709 41153 38712
rect 41187 38709 41199 38743
rect 41141 38703 41199 38709
rect 41690 38700 41696 38752
rect 41748 38740 41754 38752
rect 42518 38740 42524 38752
rect 41748 38712 42524 38740
rect 41748 38700 41754 38712
rect 42518 38700 42524 38712
rect 42576 38700 42582 38752
rect 42886 38700 42892 38752
rect 42944 38740 42950 38752
rect 43254 38740 43260 38752
rect 42944 38712 43260 38740
rect 42944 38700 42950 38712
rect 43254 38700 43260 38712
rect 43312 38700 43318 38752
rect 43349 38743 43407 38749
rect 43349 38709 43361 38743
rect 43395 38740 43407 38743
rect 47213 38743 47271 38749
rect 47213 38740 47225 38743
rect 43395 38712 47225 38740
rect 43395 38709 43407 38712
rect 43349 38703 43407 38709
rect 47213 38709 47225 38712
rect 47259 38740 47271 38743
rect 47578 38740 47584 38752
rect 47259 38712 47584 38740
rect 47259 38709 47271 38712
rect 47213 38703 47271 38709
rect 47578 38700 47584 38712
rect 47636 38700 47642 38752
rect 48130 38700 48136 38752
rect 48188 38740 48194 38752
rect 48406 38740 48412 38752
rect 48188 38712 48412 38740
rect 48188 38700 48194 38712
rect 48406 38700 48412 38712
rect 48464 38700 48470 38752
rect 48498 38700 48504 38752
rect 48556 38740 48562 38752
rect 48556 38712 48601 38740
rect 48556 38700 48562 38712
rect 53742 38700 53748 38752
rect 53800 38740 53806 38752
rect 53837 38743 53895 38749
rect 53837 38740 53849 38743
rect 53800 38712 53849 38740
rect 53800 38700 53806 38712
rect 53837 38709 53849 38712
rect 53883 38709 53895 38743
rect 54404 38740 54432 38984
rect 56226 38972 56232 39024
rect 56284 39012 56290 39024
rect 62224 39012 62252 39052
rect 67634 39040 67640 39052
rect 67692 39040 67698 39092
rect 69017 39083 69075 39089
rect 69017 39049 69029 39083
rect 69063 39080 69075 39083
rect 69106 39080 69112 39092
rect 69063 39052 69112 39080
rect 69063 39049 69075 39052
rect 69017 39043 69075 39049
rect 69106 39040 69112 39052
rect 69164 39040 69170 39092
rect 70946 39080 70952 39092
rect 70859 39052 70952 39080
rect 70946 39040 70952 39052
rect 71004 39080 71010 39092
rect 71004 39052 72556 39080
rect 71004 39040 71010 39052
rect 68738 39012 68744 39024
rect 56284 38984 62252 39012
rect 63604 38984 68744 39012
rect 56284 38972 56290 38984
rect 56134 38904 56140 38956
rect 56192 38944 56198 38956
rect 63604 38944 63632 38984
rect 68738 38972 68744 38984
rect 68796 38972 68802 39024
rect 72528 39012 72556 39052
rect 72602 39040 72608 39092
rect 72660 39080 72666 39092
rect 73982 39080 73988 39092
rect 72660 39052 73988 39080
rect 72660 39040 72666 39052
rect 73982 39040 73988 39052
rect 74040 39040 74046 39092
rect 75178 39080 75184 39092
rect 75139 39052 75184 39080
rect 75178 39040 75184 39052
rect 75236 39040 75242 39092
rect 77205 39083 77263 39089
rect 77205 39049 77217 39083
rect 77251 39080 77263 39083
rect 78950 39080 78956 39092
rect 77251 39052 78956 39080
rect 77251 39049 77263 39052
rect 77205 39043 77263 39049
rect 78950 39040 78956 39052
rect 79008 39040 79014 39092
rect 82722 39080 82728 39092
rect 80164 39052 82728 39080
rect 76837 39015 76895 39021
rect 76837 39012 76849 39015
rect 72528 38984 76849 39012
rect 76837 38981 76849 38984
rect 76883 39012 76895 39015
rect 79778 39012 79784 39024
rect 76883 38984 79784 39012
rect 76883 38981 76895 38984
rect 76837 38975 76895 38981
rect 63770 38944 63776 38956
rect 56192 38916 63632 38944
rect 63731 38916 63776 38944
rect 56192 38904 56198 38916
rect 63770 38904 63776 38916
rect 63828 38904 63834 38956
rect 64046 38904 64052 38956
rect 64104 38944 64110 38956
rect 64506 38944 64512 38956
rect 64104 38916 64512 38944
rect 64104 38904 64110 38916
rect 64506 38904 64512 38916
rect 64564 38944 64570 38956
rect 64693 38947 64751 38953
rect 64693 38944 64705 38947
rect 64564 38916 64705 38944
rect 64564 38904 64570 38916
rect 64693 38913 64705 38916
rect 64739 38913 64751 38947
rect 64693 38907 64751 38913
rect 65518 38904 65524 38956
rect 65576 38944 65582 38956
rect 72329 38947 72387 38953
rect 72329 38944 72341 38947
rect 65576 38916 68784 38944
rect 65576 38904 65582 38916
rect 55674 38876 55680 38888
rect 55635 38848 55680 38876
rect 55674 38836 55680 38848
rect 55732 38836 55738 38888
rect 55766 38836 55772 38888
rect 55824 38876 55830 38888
rect 55824 38848 55869 38876
rect 55824 38836 55830 38848
rect 56042 38836 56048 38888
rect 56100 38876 56106 38888
rect 56100 38848 56145 38876
rect 56100 38836 56106 38848
rect 62298 38836 62304 38888
rect 62356 38876 62362 38888
rect 63218 38876 63224 38888
rect 62356 38848 63224 38876
rect 62356 38836 62362 38848
rect 63218 38836 63224 38848
rect 63276 38836 63282 38888
rect 63405 38879 63463 38885
rect 63405 38845 63417 38879
rect 63451 38876 63463 38879
rect 63678 38876 63684 38888
rect 63451 38848 63684 38876
rect 63451 38845 63463 38848
rect 63405 38839 63463 38845
rect 63678 38836 63684 38848
rect 63736 38876 63742 38888
rect 64601 38879 64659 38885
rect 64601 38876 64613 38879
rect 63736 38848 64613 38876
rect 63736 38836 63742 38848
rect 64601 38845 64613 38848
rect 64647 38876 64659 38879
rect 64782 38876 64788 38888
rect 64647 38848 64788 38876
rect 64647 38845 64659 38848
rect 64601 38839 64659 38845
rect 64782 38836 64788 38848
rect 64840 38836 64846 38888
rect 68554 38876 68560 38888
rect 68515 38848 68560 38876
rect 68554 38836 68560 38848
rect 68612 38836 68618 38888
rect 68756 38876 68784 38916
rect 69400 38916 72341 38944
rect 69400 38876 69428 38916
rect 72329 38913 72341 38916
rect 72375 38944 72387 38947
rect 74905 38947 74963 38953
rect 74905 38944 74917 38947
rect 72375 38916 74917 38944
rect 72375 38913 72387 38916
rect 72329 38907 72387 38913
rect 74905 38913 74917 38916
rect 74951 38944 74963 38947
rect 74951 38916 75684 38944
rect 74951 38913 74963 38916
rect 74905 38907 74963 38913
rect 68756 38848 69428 38876
rect 69661 38879 69719 38885
rect 69661 38845 69673 38879
rect 69707 38845 69719 38879
rect 69661 38839 69719 38845
rect 70765 38879 70823 38885
rect 70765 38845 70777 38879
rect 70811 38876 70823 38879
rect 71406 38876 71412 38888
rect 70811 38848 71412 38876
rect 70811 38845 70823 38848
rect 70765 38839 70823 38845
rect 55858 38768 55864 38820
rect 55916 38808 55922 38820
rect 55916 38780 62068 38808
rect 55916 38768 55922 38780
rect 60826 38740 60832 38752
rect 54404 38712 60832 38740
rect 53837 38703 53895 38709
rect 60826 38700 60832 38712
rect 60884 38700 60890 38752
rect 62040 38740 62068 38780
rect 62114 38768 62120 38820
rect 62172 38808 62178 38820
rect 69474 38808 69480 38820
rect 62172 38780 68738 38808
rect 69435 38780 69480 38808
rect 62172 38768 62178 38780
rect 68710 38752 68738 38780
rect 69474 38768 69480 38780
rect 69532 38808 69538 38820
rect 69676 38808 69704 38839
rect 71406 38836 71412 38848
rect 71464 38836 71470 38888
rect 72237 38879 72295 38885
rect 72237 38845 72249 38879
rect 72283 38876 72295 38879
rect 72602 38876 72608 38888
rect 72283 38848 72608 38876
rect 72283 38845 72295 38848
rect 72237 38839 72295 38845
rect 72602 38836 72608 38848
rect 72660 38836 72666 38888
rect 75656 38885 75684 38916
rect 75730 38904 75736 38956
rect 75788 38944 75794 38956
rect 77570 38944 77576 38956
rect 75788 38916 77576 38944
rect 75788 38904 75794 38916
rect 77570 38904 77576 38916
rect 77628 38904 77634 38956
rect 77680 38953 77708 38984
rect 79778 38972 79784 38984
rect 79836 38972 79842 39024
rect 80057 39015 80115 39021
rect 80057 38981 80069 39015
rect 80103 39012 80115 39015
rect 80164 39012 80192 39052
rect 82722 39040 82728 39052
rect 82780 39040 82786 39092
rect 83458 39080 83464 39092
rect 83419 39052 83464 39080
rect 83458 39040 83464 39052
rect 83516 39040 83522 39092
rect 84378 39040 84384 39092
rect 84436 39080 84442 39092
rect 85298 39080 85304 39092
rect 84436 39052 85304 39080
rect 84436 39040 84442 39052
rect 85298 39040 85304 39052
rect 85356 39080 85362 39092
rect 85485 39083 85543 39089
rect 85485 39080 85497 39083
rect 85356 39052 85497 39080
rect 85356 39040 85362 39052
rect 85485 39049 85497 39052
rect 85531 39049 85543 39083
rect 85485 39043 85543 39049
rect 80103 38984 80192 39012
rect 80103 38981 80115 38984
rect 80057 38975 80115 38981
rect 80238 38972 80244 39024
rect 80296 39012 80302 39024
rect 80977 39015 81035 39021
rect 80977 39012 80989 39015
rect 80296 38984 80989 39012
rect 80296 38972 80302 38984
rect 80977 38981 80989 38984
rect 81023 38981 81035 39015
rect 80977 38975 81035 38981
rect 81084 38984 84148 39012
rect 77665 38947 77723 38953
rect 77665 38913 77677 38947
rect 77711 38913 77723 38947
rect 77665 38907 77723 38913
rect 77864 38916 78352 38944
rect 75365 38879 75423 38885
rect 75365 38845 75377 38879
rect 75411 38845 75423 38879
rect 75365 38839 75423 38845
rect 75641 38879 75699 38885
rect 75641 38845 75653 38879
rect 75687 38876 75699 38879
rect 76374 38876 76380 38888
rect 75687 38848 76380 38876
rect 75687 38845 75699 38848
rect 75641 38839 75699 38845
rect 69532 38780 69704 38808
rect 75380 38808 75408 38839
rect 76374 38836 76380 38848
rect 76432 38836 76438 38888
rect 77754 38876 77760 38888
rect 77715 38848 77760 38876
rect 77754 38836 77760 38848
rect 77812 38836 77818 38888
rect 76098 38808 76104 38820
rect 75380 38780 76104 38808
rect 69532 38768 69538 38780
rect 76098 38768 76104 38780
rect 76156 38768 76162 38820
rect 77018 38768 77024 38820
rect 77076 38808 77082 38820
rect 77864 38808 77892 38916
rect 78324 38885 78352 38916
rect 79594 38904 79600 38956
rect 79652 38944 79658 38956
rect 79928 38947 79986 38953
rect 79928 38944 79940 38947
rect 79652 38916 79940 38944
rect 79652 38904 79658 38916
rect 79928 38913 79940 38916
rect 79974 38944 79986 38947
rect 80146 38947 80204 38953
rect 79974 38913 80008 38944
rect 79928 38907 80008 38913
rect 80146 38913 80158 38947
rect 80192 38944 80204 38947
rect 80256 38944 80284 38972
rect 80192 38916 80284 38944
rect 80192 38913 80204 38916
rect 80146 38907 80204 38913
rect 78125 38879 78183 38885
rect 78125 38845 78137 38879
rect 78171 38845 78183 38879
rect 78125 38839 78183 38845
rect 78309 38879 78367 38885
rect 78309 38845 78321 38879
rect 78355 38876 78367 38879
rect 79980 38876 80008 38907
rect 80330 38904 80336 38956
rect 80388 38944 80394 38956
rect 81084 38944 81112 38984
rect 83734 38944 83740 38956
rect 80388 38916 81112 38944
rect 83695 38916 83740 38944
rect 80388 38904 80394 38916
rect 83734 38904 83740 38916
rect 83792 38944 83798 38956
rect 84120 38953 84148 38984
rect 84105 38947 84163 38953
rect 83792 38916 84056 38944
rect 83792 38904 83798 38916
rect 80793 38879 80851 38885
rect 80793 38876 80805 38879
rect 78355 38848 79916 38876
rect 79980 38848 80805 38876
rect 78355 38845 78367 38848
rect 78309 38839 78367 38845
rect 77076 38780 77892 38808
rect 78141 38808 78169 38839
rect 79778 38808 79784 38820
rect 78141 38780 78260 38808
rect 79739 38780 79784 38808
rect 77076 38768 77082 38780
rect 78232 38752 78260 38780
rect 79778 38768 79784 38780
rect 79836 38768 79842 38820
rect 79888 38808 79916 38848
rect 80793 38845 80805 38848
rect 80839 38845 80851 38879
rect 80793 38839 80851 38845
rect 83642 38836 83648 38888
rect 83700 38885 83706 38888
rect 83700 38876 83708 38885
rect 83921 38879 83979 38885
rect 83700 38848 83745 38876
rect 83700 38839 83708 38848
rect 83921 38845 83933 38879
rect 83967 38845 83979 38879
rect 84028 38876 84056 38916
rect 84105 38913 84117 38947
rect 84151 38913 84163 38947
rect 84105 38907 84163 38913
rect 84473 38879 84531 38885
rect 84473 38876 84485 38879
rect 84028 38848 84485 38876
rect 83921 38839 83979 38845
rect 84473 38845 84485 38848
rect 84519 38876 84531 38879
rect 85206 38876 85212 38888
rect 84519 38848 85212 38876
rect 84519 38845 84531 38848
rect 84473 38839 84531 38845
rect 83700 38836 83706 38839
rect 80238 38808 80244 38820
rect 79888 38780 80244 38808
rect 80238 38768 80244 38780
rect 80296 38768 80302 38820
rect 80609 38811 80667 38817
rect 80609 38808 80621 38811
rect 80348 38780 80621 38808
rect 65978 38740 65984 38752
rect 62040 38712 65984 38740
rect 65978 38700 65984 38712
rect 66036 38700 66042 38752
rect 67266 38700 67272 38752
rect 67324 38740 67330 38752
rect 68462 38740 68468 38752
rect 67324 38712 68468 38740
rect 67324 38700 67330 38712
rect 68462 38700 68468 38712
rect 68520 38700 68526 38752
rect 68710 38712 68744 38752
rect 68738 38700 68744 38712
rect 68796 38740 68802 38752
rect 68796 38712 68889 38740
rect 68796 38700 68802 38712
rect 69750 38700 69756 38752
rect 69808 38740 69814 38752
rect 69845 38743 69903 38749
rect 69845 38740 69857 38743
rect 69808 38712 69857 38740
rect 69808 38700 69814 38712
rect 69845 38709 69857 38712
rect 69891 38740 69903 38743
rect 70302 38740 70308 38752
rect 69891 38712 70308 38740
rect 69891 38709 69903 38712
rect 69845 38703 69903 38709
rect 70302 38700 70308 38712
rect 70360 38700 70366 38752
rect 76282 38700 76288 38752
rect 76340 38740 76346 38752
rect 76650 38740 76656 38752
rect 76340 38712 76656 38740
rect 76340 38700 76346 38712
rect 76650 38700 76656 38712
rect 76708 38740 76714 38752
rect 76929 38743 76987 38749
rect 76929 38740 76941 38743
rect 76708 38712 76941 38740
rect 76708 38700 76714 38712
rect 76929 38709 76941 38712
rect 76975 38740 76987 38743
rect 77570 38740 77576 38752
rect 76975 38712 77576 38740
rect 76975 38709 76987 38712
rect 76929 38703 76987 38709
rect 77570 38700 77576 38712
rect 77628 38700 77634 38752
rect 78214 38700 78220 38752
rect 78272 38700 78278 38752
rect 79796 38740 79824 38768
rect 80348 38740 80376 38780
rect 80609 38777 80621 38780
rect 80655 38777 80667 38811
rect 80609 38771 80667 38777
rect 83458 38768 83464 38820
rect 83516 38808 83522 38820
rect 83936 38808 83964 38839
rect 85206 38836 85212 38848
rect 85264 38836 85270 38888
rect 85390 38876 85396 38888
rect 85351 38848 85396 38876
rect 85390 38836 85396 38848
rect 85448 38836 85454 38888
rect 86497 38879 86555 38885
rect 86497 38876 86509 38879
rect 86420 38848 86509 38876
rect 83516 38780 83964 38808
rect 83516 38768 83522 38780
rect 86420 38752 86448 38848
rect 86497 38845 86509 38848
rect 86543 38845 86555 38879
rect 86770 38876 86776 38888
rect 86731 38848 86776 38876
rect 86497 38839 86555 38845
rect 86770 38836 86776 38848
rect 86828 38836 86834 38888
rect 79796 38712 80376 38740
rect 80425 38743 80483 38749
rect 80425 38709 80437 38743
rect 80471 38740 80483 38743
rect 80514 38740 80520 38752
rect 80471 38712 80520 38740
rect 80471 38709 80483 38712
rect 80425 38703 80483 38709
rect 80514 38700 80520 38712
rect 80572 38700 80578 38752
rect 86402 38740 86408 38752
rect 86363 38712 86408 38740
rect 86402 38700 86408 38712
rect 86460 38700 86466 38752
rect 87874 38740 87880 38752
rect 87835 38712 87880 38740
rect 87874 38700 87880 38712
rect 87932 38700 87938 38752
rect 1104 38650 111136 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 50326 38650
rect 50378 38598 50390 38650
rect 50442 38598 50454 38650
rect 50506 38598 50518 38650
rect 50570 38598 81046 38650
rect 81098 38598 81110 38650
rect 81162 38598 81174 38650
rect 81226 38598 81238 38650
rect 81290 38598 111136 38650
rect 1104 38576 111136 38598
rect 3694 38496 3700 38548
rect 3752 38536 3758 38548
rect 8110 38536 8116 38548
rect 3752 38508 8116 38536
rect 3752 38496 3758 38508
rect 8110 38496 8116 38508
rect 8168 38496 8174 38548
rect 9950 38536 9956 38548
rect 9911 38508 9956 38536
rect 9950 38496 9956 38508
rect 10008 38496 10014 38548
rect 11238 38496 11244 38548
rect 11296 38536 11302 38548
rect 13078 38536 13084 38548
rect 11296 38508 11928 38536
rect 13039 38508 13084 38536
rect 11296 38496 11302 38508
rect 7469 38471 7527 38477
rect 7469 38437 7481 38471
rect 7515 38468 7527 38471
rect 7515 38440 8800 38468
rect 7515 38437 7527 38440
rect 7469 38431 7527 38437
rect 8772 38412 8800 38440
rect 10410 38428 10416 38480
rect 10468 38468 10474 38480
rect 10873 38471 10931 38477
rect 10873 38468 10885 38471
rect 10468 38440 10885 38468
rect 10468 38428 10474 38440
rect 10873 38437 10885 38440
rect 10919 38437 10931 38471
rect 10873 38431 10931 38437
rect 10962 38428 10968 38480
rect 11020 38468 11026 38480
rect 11020 38440 11560 38468
rect 11020 38428 11026 38440
rect 4341 38403 4399 38409
rect 4341 38369 4353 38403
rect 4387 38400 4399 38403
rect 4430 38400 4436 38412
rect 4387 38372 4436 38400
rect 4387 38369 4399 38372
rect 4341 38363 4399 38369
rect 4430 38360 4436 38372
rect 4488 38400 4494 38412
rect 5074 38400 5080 38412
rect 4488 38372 5080 38400
rect 4488 38360 4494 38372
rect 5074 38360 5080 38372
rect 5132 38400 5138 38412
rect 6089 38403 6147 38409
rect 6089 38400 6101 38403
rect 5132 38372 6101 38400
rect 5132 38360 5138 38372
rect 6089 38369 6101 38372
rect 6135 38369 6147 38403
rect 6089 38363 6147 38369
rect 7285 38403 7343 38409
rect 7285 38369 7297 38403
rect 7331 38400 7343 38403
rect 8018 38400 8024 38412
rect 7331 38372 8024 38400
rect 7331 38369 7343 38372
rect 7285 38363 7343 38369
rect 8018 38360 8024 38372
rect 8076 38360 8082 38412
rect 8205 38403 8263 38409
rect 8205 38369 8217 38403
rect 8251 38369 8263 38403
rect 8205 38363 8263 38369
rect 8573 38403 8631 38409
rect 8573 38369 8585 38403
rect 8619 38369 8631 38403
rect 8754 38400 8760 38412
rect 8715 38372 8760 38400
rect 8573 38363 8631 38369
rect 4614 38332 4620 38344
rect 4575 38304 4620 38332
rect 4614 38292 4620 38304
rect 4672 38292 4678 38344
rect 5442 38292 5448 38344
rect 5500 38332 5506 38344
rect 7561 38335 7619 38341
rect 7561 38332 7573 38335
rect 5500 38304 7573 38332
rect 5500 38292 5506 38304
rect 7561 38301 7573 38304
rect 7607 38301 7619 38335
rect 7561 38295 7619 38301
rect 8220 38264 8248 38363
rect 8588 38332 8616 38363
rect 8754 38360 8760 38372
rect 8812 38360 8818 38412
rect 9769 38403 9827 38409
rect 9769 38369 9781 38403
rect 9815 38400 9827 38403
rect 10778 38400 10784 38412
rect 9815 38372 10784 38400
rect 9815 38369 9827 38372
rect 9769 38363 9827 38369
rect 10778 38360 10784 38372
rect 10836 38360 10842 38412
rect 11238 38400 11244 38412
rect 10888 38372 11244 38400
rect 10888 38344 10916 38372
rect 11238 38360 11244 38372
rect 11296 38360 11302 38412
rect 11532 38409 11560 38440
rect 11900 38409 11928 38508
rect 13078 38496 13084 38508
rect 13136 38496 13142 38548
rect 14182 38496 14188 38548
rect 14240 38536 14246 38548
rect 14921 38539 14979 38545
rect 14921 38536 14933 38539
rect 14240 38508 14933 38536
rect 14240 38496 14246 38508
rect 14921 38505 14933 38508
rect 14967 38536 14979 38539
rect 15105 38539 15163 38545
rect 15105 38536 15117 38539
rect 14967 38508 15117 38536
rect 14967 38505 14979 38508
rect 14921 38499 14979 38505
rect 15105 38505 15117 38508
rect 15151 38505 15163 38539
rect 16482 38536 16488 38548
rect 16443 38508 16488 38536
rect 15105 38499 15163 38505
rect 16482 38496 16488 38508
rect 16540 38496 16546 38548
rect 16574 38496 16580 38548
rect 16632 38536 16638 38548
rect 16853 38539 16911 38545
rect 16853 38536 16865 38539
rect 16632 38508 16865 38536
rect 16632 38496 16638 38508
rect 16853 38505 16865 38508
rect 16899 38536 16911 38539
rect 17402 38536 17408 38548
rect 16899 38508 17408 38536
rect 16899 38505 16911 38508
rect 16853 38499 16911 38505
rect 17402 38496 17408 38508
rect 17460 38496 17466 38548
rect 19242 38536 19248 38548
rect 17512 38508 19248 38536
rect 14458 38428 14464 38480
rect 14516 38468 14522 38480
rect 17512 38468 17540 38508
rect 19242 38496 19248 38508
rect 19300 38496 19306 38548
rect 25406 38536 25412 38548
rect 25367 38508 25412 38536
rect 25406 38496 25412 38508
rect 25464 38496 25470 38548
rect 27522 38496 27528 38548
rect 27580 38536 27586 38548
rect 29638 38536 29644 38548
rect 27580 38508 29040 38536
rect 29599 38508 29644 38536
rect 27580 38496 27586 38508
rect 14516 38440 17540 38468
rect 14516 38428 14522 38440
rect 22278 38428 22284 38480
rect 22336 38468 22342 38480
rect 23569 38471 23627 38477
rect 23569 38468 23581 38471
rect 22336 38440 23581 38468
rect 22336 38428 22342 38440
rect 23569 38437 23581 38440
rect 23615 38468 23627 38471
rect 23934 38468 23940 38480
rect 23615 38440 23940 38468
rect 23615 38437 23627 38440
rect 23569 38431 23627 38437
rect 23934 38428 23940 38440
rect 23992 38428 23998 38480
rect 24949 38471 25007 38477
rect 24949 38437 24961 38471
rect 24995 38468 25007 38471
rect 26878 38468 26884 38480
rect 24995 38440 26884 38468
rect 24995 38437 25007 38440
rect 24949 38431 25007 38437
rect 26878 38428 26884 38440
rect 26936 38428 26942 38480
rect 29012 38468 29040 38508
rect 29638 38496 29644 38508
rect 29696 38496 29702 38548
rect 30561 38539 30619 38545
rect 30561 38505 30573 38539
rect 30607 38536 30619 38539
rect 46014 38536 46020 38548
rect 30607 38508 46020 38536
rect 30607 38505 30619 38508
rect 30561 38499 30619 38505
rect 46014 38496 46020 38508
rect 46072 38496 46078 38548
rect 46106 38496 46112 38548
rect 46164 38536 46170 38548
rect 52546 38536 52552 38548
rect 46164 38508 52552 38536
rect 46164 38496 46170 38508
rect 52546 38496 52552 38508
rect 52604 38496 52610 38548
rect 53285 38539 53343 38545
rect 53285 38505 53297 38539
rect 53331 38536 53343 38539
rect 53374 38536 53380 38548
rect 53331 38508 53380 38536
rect 53331 38505 53343 38508
rect 53285 38499 53343 38505
rect 51810 38468 51816 38480
rect 29012 38440 51816 38468
rect 51810 38428 51816 38440
rect 51868 38428 51874 38480
rect 11517 38403 11575 38409
rect 11517 38369 11529 38403
rect 11563 38369 11575 38403
rect 11517 38363 11575 38369
rect 11885 38403 11943 38409
rect 11885 38369 11897 38403
rect 11931 38400 11943 38403
rect 11974 38400 11980 38412
rect 11931 38372 11980 38400
rect 11931 38369 11943 38372
rect 11885 38363 11943 38369
rect 11974 38360 11980 38372
rect 12032 38360 12038 38412
rect 12069 38403 12127 38409
rect 12069 38369 12081 38403
rect 12115 38369 12127 38403
rect 12069 38363 12127 38369
rect 10870 38332 10876 38344
rect 8588 38304 10876 38332
rect 10870 38292 10876 38304
rect 10928 38292 10934 38344
rect 11609 38335 11667 38341
rect 11609 38301 11621 38335
rect 11655 38301 11667 38335
rect 12084 38332 12112 38363
rect 12158 38360 12164 38412
rect 12216 38400 12222 38412
rect 12897 38403 12955 38409
rect 12897 38400 12909 38403
rect 12216 38372 12909 38400
rect 12216 38360 12222 38372
rect 12897 38369 12909 38372
rect 12943 38369 12955 38403
rect 12897 38363 12955 38369
rect 13998 38360 14004 38412
rect 14056 38400 14062 38412
rect 14737 38403 14795 38409
rect 14737 38400 14749 38403
rect 14056 38372 14749 38400
rect 14056 38360 14062 38372
rect 14737 38369 14749 38372
rect 14783 38400 14795 38403
rect 14826 38400 14832 38412
rect 14783 38372 14832 38400
rect 14783 38369 14795 38372
rect 14737 38363 14795 38369
rect 14826 38360 14832 38372
rect 14884 38360 14890 38412
rect 15105 38403 15163 38409
rect 15105 38369 15117 38403
rect 15151 38400 15163 38403
rect 15473 38403 15531 38409
rect 15473 38400 15485 38403
rect 15151 38372 15485 38400
rect 15151 38369 15163 38372
rect 15105 38363 15163 38369
rect 15473 38369 15485 38372
rect 15519 38369 15531 38403
rect 15473 38363 15531 38369
rect 15565 38403 15623 38409
rect 15565 38369 15577 38403
rect 15611 38369 15623 38403
rect 15565 38363 15623 38369
rect 12253 38335 12311 38341
rect 12253 38332 12265 38335
rect 12084 38304 12265 38332
rect 11609 38295 11667 38301
rect 12253 38301 12265 38304
rect 12299 38332 12311 38335
rect 15378 38332 15384 38344
rect 12299 38304 15384 38332
rect 12299 38301 12311 38304
rect 12253 38295 12311 38301
rect 10042 38264 10048 38276
rect 8220 38236 10048 38264
rect 10042 38224 10048 38236
rect 10100 38224 10106 38276
rect 11624 38264 11652 38295
rect 15378 38292 15384 38304
rect 15436 38292 15442 38344
rect 15580 38332 15608 38363
rect 15930 38360 15936 38412
rect 15988 38400 15994 38412
rect 16025 38403 16083 38409
rect 16025 38400 16037 38403
rect 15988 38372 16037 38400
rect 15988 38360 15994 38372
rect 16025 38369 16037 38372
rect 16071 38369 16083 38403
rect 16025 38363 16083 38369
rect 16209 38403 16267 38409
rect 16209 38369 16221 38403
rect 16255 38400 16267 38403
rect 16574 38400 16580 38412
rect 16255 38372 16580 38400
rect 16255 38369 16267 38372
rect 16209 38363 16267 38369
rect 16574 38360 16580 38372
rect 16632 38360 16638 38412
rect 19705 38403 19763 38409
rect 19705 38369 19717 38403
rect 19751 38400 19763 38403
rect 20530 38400 20536 38412
rect 19751 38372 20536 38400
rect 19751 38369 19763 38372
rect 19705 38363 19763 38369
rect 20530 38360 20536 38372
rect 20588 38400 20594 38412
rect 23661 38403 23719 38409
rect 23661 38400 23673 38403
rect 20588 38372 23673 38400
rect 20588 38360 20594 38372
rect 23661 38369 23673 38372
rect 23707 38369 23719 38403
rect 23842 38400 23848 38412
rect 23803 38372 23848 38400
rect 23661 38363 23719 38369
rect 23842 38360 23848 38372
rect 23900 38360 23906 38412
rect 24394 38400 24400 38412
rect 24355 38372 24400 38400
rect 24394 38360 24400 38372
rect 24452 38360 24458 38412
rect 24578 38400 24584 38412
rect 24539 38372 24584 38400
rect 24578 38360 24584 38372
rect 24636 38360 24642 38412
rect 26602 38360 26608 38412
rect 26660 38400 26666 38412
rect 30650 38400 30656 38412
rect 26660 38372 29132 38400
rect 30611 38372 30656 38400
rect 26660 38360 26666 38372
rect 25222 38332 25228 38344
rect 15488 38304 15608 38332
rect 25183 38304 25228 38332
rect 12345 38267 12403 38273
rect 12345 38264 12357 38267
rect 11624 38236 12357 38264
rect 12345 38233 12357 38236
rect 12391 38264 12403 38267
rect 15194 38264 15200 38276
rect 12391 38236 15200 38264
rect 12391 38233 12403 38236
rect 12345 38227 12403 38233
rect 15194 38224 15200 38236
rect 15252 38224 15258 38276
rect 15488 38264 15516 38304
rect 25222 38292 25228 38304
rect 25280 38292 25286 38344
rect 25866 38292 25872 38344
rect 25924 38332 25930 38344
rect 27893 38335 27951 38341
rect 27893 38332 27905 38335
rect 25924 38304 27905 38332
rect 25924 38292 25930 38304
rect 27893 38301 27905 38304
rect 27939 38332 27951 38335
rect 28077 38335 28135 38341
rect 28077 38332 28089 38335
rect 27939 38304 28089 38332
rect 27939 38301 27951 38304
rect 27893 38295 27951 38301
rect 28077 38301 28089 38304
rect 28123 38301 28135 38335
rect 28350 38332 28356 38344
rect 28311 38304 28356 38332
rect 28077 38295 28135 38301
rect 28350 38292 28356 38304
rect 28408 38292 28414 38344
rect 29104 38332 29132 38372
rect 30650 38360 30656 38372
rect 30708 38360 30714 38412
rect 31478 38360 31484 38412
rect 31536 38400 31542 38412
rect 33229 38403 33287 38409
rect 33229 38400 33241 38403
rect 31536 38372 33241 38400
rect 31536 38360 31542 38372
rect 33229 38369 33241 38372
rect 33275 38369 33287 38403
rect 36538 38400 36544 38412
rect 36499 38372 36544 38400
rect 33229 38363 33287 38369
rect 36538 38360 36544 38372
rect 36596 38360 36602 38412
rect 37734 38400 37740 38412
rect 37695 38372 37740 38400
rect 37734 38360 37740 38372
rect 37792 38360 37798 38412
rect 37918 38400 37924 38412
rect 37879 38372 37924 38400
rect 37918 38360 37924 38372
rect 37976 38360 37982 38412
rect 38010 38360 38016 38412
rect 38068 38400 38074 38412
rect 38381 38403 38439 38409
rect 38381 38400 38393 38403
rect 38068 38372 38393 38400
rect 38068 38360 38074 38372
rect 38381 38369 38393 38372
rect 38427 38369 38439 38403
rect 38381 38363 38439 38369
rect 38470 38360 38476 38412
rect 38528 38400 38534 38412
rect 38528 38372 38573 38400
rect 38528 38360 38534 38372
rect 38654 38360 38660 38412
rect 38712 38400 38718 38412
rect 39209 38403 39267 38409
rect 39209 38400 39221 38403
rect 38712 38372 39221 38400
rect 38712 38360 38718 38372
rect 39209 38369 39221 38372
rect 39255 38369 39267 38403
rect 40862 38400 40868 38412
rect 40823 38372 40868 38400
rect 39209 38363 39267 38369
rect 40862 38360 40868 38372
rect 40920 38360 40926 38412
rect 43898 38400 43904 38412
rect 40972 38372 43904 38400
rect 32858 38332 32864 38344
rect 29104 38304 32864 38332
rect 32858 38292 32864 38304
rect 32916 38292 32922 38344
rect 36446 38292 36452 38344
rect 36504 38332 36510 38344
rect 36633 38335 36691 38341
rect 36633 38332 36645 38335
rect 36504 38304 36645 38332
rect 36504 38292 36510 38304
rect 36633 38301 36645 38304
rect 36679 38301 36691 38335
rect 36633 38295 36691 38301
rect 39025 38335 39083 38341
rect 39025 38301 39037 38335
rect 39071 38332 39083 38335
rect 40972 38332 41000 38372
rect 43898 38360 43904 38372
rect 43956 38360 43962 38412
rect 47581 38403 47639 38409
rect 47581 38369 47593 38403
rect 47627 38400 47639 38403
rect 47670 38400 47676 38412
rect 47627 38372 47676 38400
rect 47627 38369 47639 38372
rect 47581 38363 47639 38369
rect 47670 38360 47676 38372
rect 47728 38400 47734 38412
rect 50154 38400 50160 38412
rect 47728 38372 50160 38400
rect 47728 38360 47734 38372
rect 50154 38360 50160 38372
rect 50212 38360 50218 38412
rect 51718 38360 51724 38412
rect 51776 38400 51782 38412
rect 51905 38403 51963 38409
rect 51905 38400 51917 38403
rect 51776 38372 51917 38400
rect 51776 38360 51782 38372
rect 51905 38369 51917 38372
rect 51951 38369 51963 38403
rect 52365 38403 52423 38409
rect 52365 38400 52377 38403
rect 51905 38363 51963 38369
rect 52104 38372 52377 38400
rect 41230 38332 41236 38344
rect 39071 38304 41000 38332
rect 41191 38304 41236 38332
rect 39071 38301 39083 38304
rect 39025 38295 39083 38301
rect 41230 38292 41236 38304
rect 41288 38292 41294 38344
rect 41601 38335 41659 38341
rect 41601 38301 41613 38335
rect 41647 38332 41659 38335
rect 51534 38332 51540 38344
rect 41647 38304 51540 38332
rect 41647 38301 41659 38304
rect 41601 38295 41659 38301
rect 51534 38292 51540 38304
rect 51592 38292 51598 38344
rect 51810 38332 51816 38344
rect 51771 38304 51816 38332
rect 51810 38292 51816 38304
rect 51868 38292 51874 38344
rect 15304 38236 15516 38264
rect 4706 38156 4712 38208
rect 4764 38196 4770 38208
rect 5721 38199 5779 38205
rect 5721 38196 5733 38199
rect 4764 38168 5733 38196
rect 4764 38156 4770 38168
rect 5721 38165 5733 38168
rect 5767 38165 5779 38199
rect 5721 38159 5779 38165
rect 14826 38156 14832 38208
rect 14884 38196 14890 38208
rect 15304 38196 15332 38236
rect 16942 38224 16948 38276
rect 17000 38264 17006 38276
rect 17000 38236 27016 38264
rect 17000 38224 17006 38236
rect 14884 38168 15332 38196
rect 14884 38156 14890 38168
rect 18414 38156 18420 38208
rect 18472 38196 18478 38208
rect 19797 38199 19855 38205
rect 19797 38196 19809 38199
rect 18472 38168 19809 38196
rect 18472 38156 18478 38168
rect 19797 38165 19809 38168
rect 19843 38165 19855 38199
rect 19797 38159 19855 38165
rect 24118 38156 24124 38208
rect 24176 38196 24182 38208
rect 26878 38196 26884 38208
rect 24176 38168 26884 38196
rect 24176 38156 24182 38168
rect 26878 38156 26884 38168
rect 26936 38156 26942 38208
rect 26988 38196 27016 38236
rect 29086 38224 29092 38276
rect 29144 38264 29150 38276
rect 38838 38264 38844 38276
rect 29144 38236 38844 38264
rect 29144 38224 29150 38236
rect 38838 38224 38844 38236
rect 38896 38224 38902 38276
rect 40681 38267 40739 38273
rect 40681 38264 40693 38267
rect 38948 38236 40693 38264
rect 30561 38199 30619 38205
rect 30561 38196 30573 38199
rect 26988 38168 30573 38196
rect 30561 38165 30573 38168
rect 30607 38165 30619 38199
rect 30742 38196 30748 38208
rect 30703 38168 30748 38196
rect 30561 38159 30619 38165
rect 30742 38156 30748 38168
rect 30800 38156 30806 38208
rect 33045 38199 33103 38205
rect 33045 38165 33057 38199
rect 33091 38196 33103 38199
rect 33134 38196 33140 38208
rect 33091 38168 33140 38196
rect 33091 38165 33103 38168
rect 33045 38159 33103 38165
rect 33134 38156 33140 38168
rect 33192 38156 33198 38208
rect 33226 38156 33232 38208
rect 33284 38196 33290 38208
rect 38948 38196 38976 38236
rect 40681 38233 40693 38236
rect 40727 38264 40739 38267
rect 40862 38264 40868 38276
rect 40727 38236 40868 38264
rect 40727 38233 40739 38236
rect 40681 38227 40739 38233
rect 40862 38224 40868 38236
rect 40920 38224 40926 38276
rect 49694 38264 49700 38276
rect 46216 38236 49700 38264
rect 39482 38196 39488 38208
rect 33284 38168 38976 38196
rect 39443 38168 39488 38196
rect 33284 38156 33290 38168
rect 39482 38156 39488 38168
rect 39540 38156 39546 38208
rect 39942 38156 39948 38208
rect 40000 38196 40006 38208
rect 41003 38199 41061 38205
rect 41003 38196 41015 38199
rect 40000 38168 41015 38196
rect 40000 38156 40006 38168
rect 41003 38165 41015 38168
rect 41049 38165 41061 38199
rect 41003 38159 41061 38165
rect 41141 38199 41199 38205
rect 41141 38165 41153 38199
rect 41187 38196 41199 38199
rect 41506 38196 41512 38208
rect 41187 38168 41512 38196
rect 41187 38165 41199 38168
rect 41141 38159 41199 38165
rect 41506 38156 41512 38168
rect 41564 38156 41570 38208
rect 42058 38156 42064 38208
rect 42116 38196 42122 38208
rect 46216 38196 46244 38236
rect 49694 38224 49700 38236
rect 49752 38224 49758 38276
rect 50154 38224 50160 38276
rect 50212 38264 50218 38276
rect 52104 38264 52132 38372
rect 52365 38369 52377 38372
rect 52411 38369 52423 38403
rect 52365 38363 52423 38369
rect 52457 38403 52515 38409
rect 52457 38369 52469 38403
rect 52503 38400 52515 38403
rect 53300 38400 53328 38499
rect 53374 38496 53380 38508
rect 53432 38496 53438 38548
rect 57790 38496 57796 38548
rect 57848 38536 57854 38548
rect 63773 38539 63831 38545
rect 57848 38508 63724 38536
rect 57848 38496 57854 38508
rect 63696 38468 63724 38508
rect 63773 38505 63785 38539
rect 63819 38536 63831 38539
rect 65518 38536 65524 38548
rect 63819 38508 65524 38536
rect 63819 38505 63831 38508
rect 63773 38499 63831 38505
rect 65518 38496 65524 38508
rect 65576 38496 65582 38548
rect 68646 38496 68652 38548
rect 68704 38536 68710 38548
rect 69201 38539 69259 38545
rect 69201 38536 69213 38539
rect 68704 38508 69213 38536
rect 68704 38496 68710 38508
rect 69201 38505 69213 38508
rect 69247 38505 69259 38539
rect 69201 38499 69259 38505
rect 74629 38539 74687 38545
rect 74629 38505 74641 38539
rect 74675 38536 74687 38539
rect 77754 38536 77760 38548
rect 74675 38508 77760 38536
rect 74675 38505 74687 38508
rect 74629 38499 74687 38505
rect 67634 38468 67640 38480
rect 63696 38440 67640 38468
rect 67634 38428 67640 38440
rect 67692 38428 67698 38480
rect 52503 38372 53328 38400
rect 52503 38369 52515 38372
rect 52457 38363 52515 38369
rect 59814 38360 59820 38412
rect 59872 38400 59878 38412
rect 60921 38403 60979 38409
rect 60921 38400 60933 38403
rect 59872 38372 60933 38400
rect 59872 38360 59878 38372
rect 60921 38369 60933 38372
rect 60967 38369 60979 38403
rect 60921 38363 60979 38369
rect 64141 38403 64199 38409
rect 64141 38369 64153 38403
rect 64187 38369 64199 38403
rect 64141 38363 64199 38369
rect 64509 38403 64567 38409
rect 64509 38369 64521 38403
rect 64555 38369 64567 38403
rect 69216 38400 69244 38499
rect 77754 38496 77760 38508
rect 77812 38496 77818 38548
rect 83642 38496 83648 38548
rect 83700 38536 83706 38548
rect 84010 38536 84016 38548
rect 83700 38508 84016 38536
rect 83700 38496 83706 38508
rect 84010 38496 84016 38508
rect 84068 38496 84074 38548
rect 75549 38471 75607 38477
rect 75549 38468 75561 38471
rect 74552 38440 75561 38468
rect 69385 38403 69443 38409
rect 69385 38400 69397 38403
rect 69216 38372 69397 38400
rect 64509 38363 64567 38369
rect 69385 38369 69397 38372
rect 69431 38369 69443 38403
rect 70118 38400 70124 38412
rect 70079 38372 70124 38400
rect 69385 38363 69443 38369
rect 60274 38292 60280 38344
rect 60332 38332 60338 38344
rect 60645 38335 60703 38341
rect 60645 38332 60657 38335
rect 60332 38304 60657 38332
rect 60332 38292 60338 38304
rect 60645 38301 60657 38304
rect 60691 38301 60703 38335
rect 60645 38295 60703 38301
rect 63957 38335 64015 38341
rect 63957 38301 63969 38335
rect 64003 38301 64015 38335
rect 63957 38295 64015 38301
rect 50212 38236 52132 38264
rect 50212 38224 50218 38236
rect 61838 38224 61844 38276
rect 61896 38264 61902 38276
rect 63972 38264 64000 38295
rect 61896 38236 64000 38264
rect 64156 38264 64184 38363
rect 64414 38332 64420 38344
rect 64375 38304 64420 38332
rect 64414 38292 64420 38304
rect 64472 38292 64478 38344
rect 64524 38332 64552 38363
rect 70118 38360 70124 38372
rect 70176 38360 70182 38412
rect 70394 38360 70400 38412
rect 70452 38400 70458 38412
rect 71409 38403 71467 38409
rect 71409 38400 71421 38403
rect 70452 38372 71421 38400
rect 70452 38360 70458 38372
rect 71409 38369 71421 38372
rect 71455 38400 71467 38403
rect 71866 38400 71872 38412
rect 71455 38372 71872 38400
rect 71455 38369 71467 38372
rect 71409 38363 71467 38369
rect 71866 38360 71872 38372
rect 71924 38360 71930 38412
rect 74552 38409 74580 38440
rect 75549 38437 75561 38440
rect 75595 38468 75607 38471
rect 76926 38468 76932 38480
rect 75595 38440 76932 38468
rect 75595 38437 75607 38440
rect 75549 38431 75607 38437
rect 76926 38428 76932 38440
rect 76984 38428 76990 38480
rect 77018 38428 77024 38480
rect 77076 38468 77082 38480
rect 77076 38440 77121 38468
rect 77076 38428 77082 38440
rect 77202 38428 77208 38480
rect 77260 38468 77266 38480
rect 77386 38468 77392 38480
rect 77260 38440 77392 38468
rect 77260 38428 77266 38440
rect 77386 38428 77392 38440
rect 77444 38428 77450 38480
rect 77772 38468 77800 38496
rect 78585 38471 78643 38477
rect 78585 38468 78597 38471
rect 77772 38440 78597 38468
rect 78585 38437 78597 38440
rect 78631 38437 78643 38471
rect 78585 38431 78643 38437
rect 82722 38428 82728 38480
rect 82780 38468 82786 38480
rect 86310 38468 86316 38480
rect 82780 38440 86316 38468
rect 82780 38428 82786 38440
rect 74537 38403 74595 38409
rect 74537 38369 74549 38403
rect 74583 38369 74595 38403
rect 75730 38400 75736 38412
rect 75691 38372 75736 38400
rect 74537 38363 74595 38369
rect 75730 38360 75736 38372
rect 75788 38400 75794 38412
rect 76193 38403 76251 38409
rect 76193 38400 76205 38403
rect 75788 38372 76205 38400
rect 75788 38360 75794 38372
rect 76193 38369 76205 38372
rect 76239 38400 76251 38403
rect 76745 38403 76803 38409
rect 76745 38400 76757 38403
rect 76239 38372 76757 38400
rect 76239 38369 76251 38372
rect 76193 38363 76251 38369
rect 76745 38369 76757 38372
rect 76791 38400 76803 38403
rect 77294 38400 77300 38412
rect 76791 38372 76972 38400
rect 76791 38369 76803 38372
rect 76745 38363 76803 38369
rect 65061 38335 65119 38341
rect 65061 38332 65073 38335
rect 64524 38304 65073 38332
rect 65061 38301 65073 38304
rect 65107 38332 65119 38335
rect 65150 38332 65156 38344
rect 65107 38304 65156 38332
rect 65107 38301 65119 38304
rect 65061 38295 65119 38301
rect 65150 38292 65156 38304
rect 65208 38332 65214 38344
rect 70302 38332 70308 38344
rect 65208 38304 70164 38332
rect 70263 38304 70308 38332
rect 65208 38292 65214 38304
rect 69661 38267 69719 38273
rect 64156 38236 64920 38264
rect 61896 38224 61902 38236
rect 64892 38208 64920 38236
rect 69661 38233 69673 38267
rect 69707 38264 69719 38267
rect 70026 38264 70032 38276
rect 69707 38236 70032 38264
rect 69707 38233 69719 38236
rect 69661 38227 69719 38233
rect 70026 38224 70032 38236
rect 70084 38224 70090 38276
rect 70136 38264 70164 38304
rect 70302 38292 70308 38304
rect 70360 38292 70366 38344
rect 76098 38332 76104 38344
rect 76059 38304 76104 38332
rect 76098 38292 76104 38304
rect 76156 38292 76162 38344
rect 76944 38332 76972 38372
rect 77174 38372 77300 38400
rect 77174 38332 77202 38372
rect 77294 38360 77300 38372
rect 77352 38400 77358 38412
rect 77352 38372 77432 38400
rect 77352 38360 77358 38372
rect 77404 38341 77432 38372
rect 78398 38360 78404 38412
rect 78456 38400 78462 38412
rect 78769 38403 78827 38409
rect 78769 38400 78781 38403
rect 78456 38372 78781 38400
rect 78456 38360 78462 38372
rect 78769 38369 78781 38372
rect 78815 38369 78827 38403
rect 83550 38400 83556 38412
rect 83511 38372 83556 38400
rect 78769 38363 78827 38369
rect 83550 38360 83556 38372
rect 83608 38360 83614 38412
rect 83660 38409 83688 38440
rect 86310 38428 86316 38440
rect 86368 38428 86374 38480
rect 86405 38471 86463 38477
rect 86405 38437 86417 38471
rect 86451 38468 86463 38471
rect 86770 38468 86776 38480
rect 86451 38440 86776 38468
rect 86451 38437 86463 38440
rect 86405 38431 86463 38437
rect 86770 38428 86776 38440
rect 86828 38428 86834 38480
rect 83645 38403 83703 38409
rect 83645 38369 83657 38403
rect 83691 38369 83703 38403
rect 83645 38363 83703 38369
rect 83829 38403 83887 38409
rect 83829 38369 83841 38403
rect 83875 38369 83887 38403
rect 85850 38400 85856 38412
rect 85811 38372 85856 38400
rect 83829 38363 83887 38369
rect 76944 38304 77202 38332
rect 77389 38335 77447 38341
rect 77389 38301 77401 38335
rect 77435 38301 77447 38335
rect 77662 38332 77668 38344
rect 77623 38304 77668 38332
rect 77389 38295 77447 38301
rect 77662 38292 77668 38304
rect 77720 38292 77726 38344
rect 83844 38332 83872 38363
rect 85850 38360 85856 38372
rect 85908 38360 85914 38412
rect 85942 38360 85948 38412
rect 86000 38400 86006 38412
rect 86000 38372 86045 38400
rect 86000 38360 86006 38372
rect 83384 38304 83872 38332
rect 75638 38264 75644 38276
rect 70136 38236 75644 38264
rect 75638 38224 75644 38236
rect 75696 38224 75702 38276
rect 76374 38264 76380 38276
rect 76335 38236 76380 38264
rect 76374 38224 76380 38236
rect 76432 38264 76438 38276
rect 77297 38267 77355 38273
rect 77297 38264 77309 38267
rect 76432 38236 77309 38264
rect 76432 38224 76438 38236
rect 77297 38233 77309 38236
rect 77343 38233 77355 38267
rect 77297 38227 77355 38233
rect 77478 38224 77484 38276
rect 77536 38264 77542 38276
rect 77536 38236 78904 38264
rect 77536 38224 77542 38236
rect 42116 38168 46244 38196
rect 42116 38156 42122 38168
rect 46290 38156 46296 38208
rect 46348 38196 46354 38208
rect 47670 38196 47676 38208
rect 46348 38168 46393 38196
rect 47631 38168 47676 38196
rect 46348 38156 46354 38168
rect 47670 38156 47676 38168
rect 47728 38156 47734 38208
rect 47762 38156 47768 38208
rect 47820 38196 47826 38208
rect 52822 38196 52828 38208
rect 47820 38168 52828 38196
rect 47820 38156 47826 38168
rect 52822 38156 52828 38168
rect 52880 38156 52886 38208
rect 52917 38199 52975 38205
rect 52917 38165 52929 38199
rect 52963 38196 52975 38199
rect 53098 38196 53104 38208
rect 52963 38168 53104 38196
rect 52963 38165 52975 38168
rect 52917 38159 52975 38165
rect 53098 38156 53104 38168
rect 53156 38156 53162 38208
rect 53374 38196 53380 38208
rect 53335 38168 53380 38196
rect 53374 38156 53380 38168
rect 53432 38156 53438 38208
rect 62209 38199 62267 38205
rect 62209 38165 62221 38199
rect 62255 38196 62267 38199
rect 64506 38196 64512 38208
rect 62255 38168 64512 38196
rect 62255 38165 62267 38168
rect 62209 38159 62267 38165
rect 64506 38156 64512 38168
rect 64564 38156 64570 38208
rect 64874 38196 64880 38208
rect 64835 38168 64880 38196
rect 64874 38156 64880 38168
rect 64932 38156 64938 38208
rect 67634 38156 67640 38208
rect 67692 38196 67698 38208
rect 68922 38196 68928 38208
rect 67692 38168 68928 38196
rect 67692 38156 67698 38168
rect 68922 38156 68928 38168
rect 68980 38196 68986 38208
rect 71593 38199 71651 38205
rect 71593 38196 71605 38199
rect 68980 38168 71605 38196
rect 68980 38156 68986 38168
rect 71593 38165 71605 38168
rect 71639 38165 71651 38199
rect 71593 38159 71651 38165
rect 76282 38156 76288 38208
rect 76340 38196 76346 38208
rect 76561 38199 76619 38205
rect 76561 38196 76573 38199
rect 76340 38168 76573 38196
rect 76340 38156 76346 38168
rect 76561 38165 76573 38168
rect 76607 38196 76619 38199
rect 77159 38199 77217 38205
rect 77159 38196 77171 38199
rect 76607 38168 77171 38196
rect 76607 38165 76619 38168
rect 76561 38159 76619 38165
rect 77159 38165 77171 38168
rect 77205 38165 77217 38199
rect 78398 38196 78404 38208
rect 78359 38168 78404 38196
rect 77159 38159 77217 38165
rect 78398 38156 78404 38168
rect 78456 38156 78462 38208
rect 78876 38205 78904 38236
rect 78861 38199 78919 38205
rect 78861 38165 78873 38199
rect 78907 38165 78919 38199
rect 78861 38159 78919 38165
rect 82814 38156 82820 38208
rect 82872 38196 82878 38208
rect 83384 38205 83412 38304
rect 83369 38199 83427 38205
rect 83369 38196 83381 38199
rect 82872 38168 83381 38196
rect 82872 38156 82878 38168
rect 83369 38165 83381 38168
rect 83415 38165 83427 38199
rect 83369 38159 83427 38165
rect 84746 38156 84752 38208
rect 84804 38196 84810 38208
rect 85669 38199 85727 38205
rect 85669 38196 85681 38199
rect 84804 38168 85681 38196
rect 84804 38156 84810 38168
rect 85669 38165 85681 38168
rect 85715 38165 85727 38199
rect 85669 38159 85727 38165
rect 1104 38106 111136 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 65686 38106
rect 65738 38054 65750 38106
rect 65802 38054 65814 38106
rect 65866 38054 65878 38106
rect 65930 38054 96406 38106
rect 96458 38054 96470 38106
rect 96522 38054 96534 38106
rect 96586 38054 96598 38106
rect 96650 38054 111136 38106
rect 1104 38032 111136 38054
rect 3970 37992 3976 38004
rect 3931 37964 3976 37992
rect 3970 37952 3976 37964
rect 4028 37952 4034 38004
rect 6086 37992 6092 38004
rect 6047 37964 6092 37992
rect 6086 37952 6092 37964
rect 6144 37952 6150 38004
rect 9858 37952 9864 38004
rect 9916 37992 9922 38004
rect 12158 37992 12164 38004
rect 9916 37964 12164 37992
rect 9916 37952 9922 37964
rect 12158 37952 12164 37964
rect 12216 37952 12222 38004
rect 14182 37992 14188 38004
rect 14143 37964 14188 37992
rect 14182 37952 14188 37964
rect 14240 37952 14246 38004
rect 14274 37952 14280 38004
rect 14332 37992 14338 38004
rect 14461 37995 14519 38001
rect 14461 37992 14473 37995
rect 14332 37964 14473 37992
rect 14332 37952 14338 37964
rect 14461 37961 14473 37964
rect 14507 37992 14519 37995
rect 16390 37992 16396 38004
rect 14507 37964 16396 37992
rect 14507 37961 14519 37964
rect 14461 37955 14519 37961
rect 16390 37952 16396 37964
rect 16448 37952 16454 38004
rect 16482 37952 16488 38004
rect 16540 37992 16546 38004
rect 20530 37992 20536 38004
rect 16540 37964 20392 37992
rect 20491 37964 20536 37992
rect 16540 37952 16546 37964
rect 3878 37884 3884 37936
rect 3936 37924 3942 37936
rect 3936 37896 11376 37924
rect 3936 37884 3942 37896
rect 2590 37856 2596 37868
rect 2503 37828 2596 37856
rect 2590 37816 2596 37828
rect 2648 37856 2654 37868
rect 4522 37856 4528 37868
rect 2648 37828 4528 37856
rect 2648 37816 2654 37828
rect 4522 37816 4528 37828
rect 4580 37856 4586 37868
rect 5074 37856 5080 37868
rect 4580 37828 5080 37856
rect 4580 37816 4586 37828
rect 5074 37816 5080 37828
rect 5132 37816 5138 37868
rect 5276 37828 6960 37856
rect 5276 37800 5304 37828
rect 2869 37791 2927 37797
rect 2869 37757 2881 37791
rect 2915 37788 2927 37791
rect 5258 37788 5264 37800
rect 2915 37760 4476 37788
rect 5219 37760 5264 37788
rect 2915 37757 2927 37760
rect 2869 37751 2927 37757
rect 4448 37729 4476 37760
rect 5258 37748 5264 37760
rect 5316 37748 5322 37800
rect 5721 37791 5779 37797
rect 5721 37757 5733 37791
rect 5767 37788 5779 37791
rect 6086 37788 6092 37800
rect 5767 37760 6092 37788
rect 5767 37757 5779 37760
rect 5721 37751 5779 37757
rect 6086 37748 6092 37760
rect 6144 37748 6150 37800
rect 6932 37797 6960 37828
rect 10042 37816 10048 37868
rect 10100 37856 10106 37868
rect 10962 37856 10968 37868
rect 10100 37828 10968 37856
rect 10100 37816 10106 37828
rect 6917 37791 6975 37797
rect 6917 37757 6929 37791
rect 6963 37757 6975 37791
rect 6917 37751 6975 37757
rect 7377 37791 7435 37797
rect 7377 37757 7389 37791
rect 7423 37788 7435 37791
rect 10594 37788 10600 37800
rect 7423 37760 10272 37788
rect 10555 37760 10600 37788
rect 7423 37757 7435 37760
rect 7377 37751 7435 37757
rect 4433 37723 4491 37729
rect 4433 37689 4445 37723
rect 4479 37720 4491 37723
rect 5902 37720 5908 37732
rect 4479 37692 5908 37720
rect 4479 37689 4491 37692
rect 4433 37683 4491 37689
rect 5902 37680 5908 37692
rect 5960 37680 5966 37732
rect 10134 37720 10140 37732
rect 10095 37692 10140 37720
rect 10134 37680 10140 37692
rect 10192 37680 10198 37732
rect 10244 37720 10272 37760
rect 10594 37748 10600 37760
rect 10652 37748 10658 37800
rect 10796 37797 10824 37828
rect 10962 37816 10968 37828
rect 11020 37816 11026 37868
rect 11348 37856 11376 37896
rect 11422 37884 11428 37936
rect 11480 37924 11486 37936
rect 18414 37924 18420 37936
rect 11480 37896 18420 37924
rect 11480 37884 11486 37896
rect 18414 37884 18420 37896
rect 18472 37884 18478 37936
rect 20364 37924 20392 37964
rect 20530 37952 20536 37964
rect 20588 37952 20594 38004
rect 20640 37964 36584 37992
rect 20640 37924 20668 37964
rect 20364 37896 20668 37924
rect 20809 37927 20867 37933
rect 20809 37893 20821 37927
rect 20855 37924 20867 37927
rect 21174 37924 21180 37936
rect 20855 37896 21180 37924
rect 20855 37893 20867 37896
rect 20809 37887 20867 37893
rect 21174 37884 21180 37896
rect 21232 37884 21238 37936
rect 23477 37927 23535 37933
rect 23477 37893 23489 37927
rect 23523 37924 23535 37927
rect 29086 37924 29092 37936
rect 23523 37896 29092 37924
rect 23523 37893 23535 37896
rect 23477 37887 23535 37893
rect 29086 37884 29092 37896
rect 29144 37884 29150 37936
rect 30650 37924 30656 37936
rect 30611 37896 30656 37924
rect 30650 37884 30656 37896
rect 30708 37884 30714 37936
rect 31570 37884 31576 37936
rect 31628 37924 31634 37936
rect 31895 37927 31953 37933
rect 31895 37924 31907 37927
rect 31628 37896 31907 37924
rect 31628 37884 31634 37896
rect 31895 37893 31907 37896
rect 31941 37893 31953 37927
rect 31895 37887 31953 37893
rect 32033 37927 32091 37933
rect 32033 37893 32045 37927
rect 32079 37924 32091 37927
rect 32674 37924 32680 37936
rect 32079 37896 32680 37924
rect 32079 37893 32091 37896
rect 32033 37887 32091 37893
rect 32674 37884 32680 37896
rect 32732 37884 32738 37936
rect 33226 37884 33232 37936
rect 33284 37924 33290 37936
rect 34422 37924 34428 37936
rect 33284 37896 34428 37924
rect 33284 37884 33290 37896
rect 34422 37884 34428 37896
rect 34480 37924 34486 37936
rect 35345 37927 35403 37933
rect 35345 37924 35357 37927
rect 34480 37896 35357 37924
rect 34480 37884 34486 37896
rect 35345 37893 35357 37896
rect 35391 37893 35403 37927
rect 36556 37924 36584 37964
rect 36630 37952 36636 38004
rect 36688 37992 36694 38004
rect 47762 37992 47768 38004
rect 36688 37964 47768 37992
rect 36688 37952 36694 37964
rect 47762 37952 47768 37964
rect 47820 37952 47826 38004
rect 51626 37952 51632 38004
rect 51684 37992 51690 38004
rect 51684 37964 53512 37992
rect 51684 37952 51690 37964
rect 42058 37924 42064 37936
rect 36556 37896 42064 37924
rect 35345 37887 35403 37893
rect 14458 37856 14464 37868
rect 11348 37828 14464 37856
rect 14458 37816 14464 37828
rect 14516 37816 14522 37868
rect 15194 37816 15200 37868
rect 15252 37856 15258 37868
rect 17037 37859 17095 37865
rect 15252 37828 16160 37856
rect 15252 37816 15258 37828
rect 10781 37791 10839 37797
rect 10781 37757 10793 37791
rect 10827 37757 10839 37791
rect 10781 37751 10839 37757
rect 10870 37748 10876 37800
rect 10928 37788 10934 37800
rect 11149 37791 11207 37797
rect 11149 37788 11161 37791
rect 10928 37760 11161 37788
rect 10928 37748 10934 37760
rect 11149 37757 11161 37760
rect 11195 37757 11207 37791
rect 11149 37751 11207 37757
rect 11333 37791 11391 37797
rect 11333 37757 11345 37791
rect 11379 37788 11391 37791
rect 12618 37788 12624 37800
rect 11379 37760 12624 37788
rect 11379 37757 11391 37760
rect 11333 37751 11391 37757
rect 12618 37748 12624 37760
rect 12676 37748 12682 37800
rect 14001 37791 14059 37797
rect 14001 37757 14013 37791
rect 14047 37788 14059 37791
rect 14274 37788 14280 37800
rect 14047 37760 14280 37788
rect 14047 37757 14059 37760
rect 14001 37751 14059 37757
rect 14274 37748 14280 37760
rect 14332 37748 14338 37800
rect 15749 37791 15807 37797
rect 15749 37788 15761 37791
rect 15580 37760 15761 37788
rect 15286 37720 15292 37732
rect 10244 37692 15292 37720
rect 15286 37680 15292 37692
rect 15344 37680 15350 37732
rect 15580 37664 15608 37760
rect 15749 37757 15761 37760
rect 15795 37757 15807 37791
rect 15930 37788 15936 37800
rect 15891 37760 15936 37788
rect 15749 37751 15807 37757
rect 15930 37748 15936 37760
rect 15988 37748 15994 37800
rect 16132 37788 16160 37828
rect 17037 37825 17049 37859
rect 17083 37856 17095 37859
rect 26142 37856 26148 37868
rect 17083 37828 25176 37856
rect 17083 37825 17095 37828
rect 17037 37819 17095 37825
rect 16298 37788 16304 37800
rect 16132 37760 16304 37788
rect 16298 37748 16304 37760
rect 16356 37788 16362 37800
rect 16393 37791 16451 37797
rect 16393 37788 16405 37791
rect 16356 37760 16405 37788
rect 16356 37748 16362 37760
rect 16393 37757 16405 37760
rect 16439 37757 16451 37791
rect 16393 37751 16451 37757
rect 16485 37791 16543 37797
rect 16485 37757 16497 37791
rect 16531 37788 16543 37791
rect 16574 37788 16580 37800
rect 16531 37760 16580 37788
rect 16531 37757 16543 37760
rect 16485 37751 16543 37757
rect 16574 37748 16580 37760
rect 16632 37788 16638 37800
rect 16850 37788 16856 37800
rect 16632 37760 16856 37788
rect 16632 37748 16638 37760
rect 16850 37748 16856 37760
rect 16908 37788 16914 37800
rect 17678 37788 17684 37800
rect 16908 37760 17684 37788
rect 16908 37748 16914 37760
rect 17678 37748 17684 37760
rect 17736 37748 17742 37800
rect 18966 37788 18972 37800
rect 18927 37760 18972 37788
rect 18966 37748 18972 37760
rect 19024 37748 19030 37800
rect 19242 37788 19248 37800
rect 19203 37760 19248 37788
rect 19242 37748 19248 37760
rect 19300 37748 19306 37800
rect 25148 37788 25176 37828
rect 25332 37828 26148 37856
rect 25332 37788 25360 37828
rect 26142 37816 26148 37828
rect 26200 37816 26206 37868
rect 27065 37859 27123 37865
rect 27065 37825 27077 37859
rect 27111 37856 27123 37859
rect 29549 37859 29607 37865
rect 29549 37856 29561 37859
rect 27111 37828 29561 37856
rect 27111 37825 27123 37828
rect 27065 37819 27123 37825
rect 29549 37825 29561 37828
rect 29595 37825 29607 37859
rect 32122 37856 32128 37868
rect 32083 37828 32128 37856
rect 29549 37819 29607 37825
rect 32122 37816 32128 37828
rect 32180 37816 32186 37868
rect 35360 37856 35388 37887
rect 42058 37884 42064 37896
rect 42116 37884 42122 37936
rect 45833 37927 45891 37933
rect 45833 37924 45845 37927
rect 42168 37896 45845 37924
rect 35529 37859 35587 37865
rect 35529 37856 35541 37859
rect 35360 37828 35541 37856
rect 35529 37825 35541 37828
rect 35575 37825 35587 37859
rect 35529 37819 35587 37825
rect 35805 37859 35863 37865
rect 35805 37825 35817 37859
rect 35851 37856 35863 37859
rect 35986 37856 35992 37868
rect 35851 37828 35992 37856
rect 35851 37825 35863 37828
rect 35805 37819 35863 37825
rect 35986 37816 35992 37828
rect 36044 37816 36050 37868
rect 36170 37816 36176 37868
rect 36228 37856 36234 37868
rect 38105 37859 38163 37865
rect 38105 37856 38117 37859
rect 36228 37828 38117 37856
rect 36228 37816 36234 37828
rect 38105 37825 38117 37828
rect 38151 37825 38163 37859
rect 38105 37819 38163 37825
rect 41414 37816 41420 37868
rect 41472 37856 41478 37868
rect 42168 37856 42196 37896
rect 45833 37893 45845 37896
rect 45879 37893 45891 37927
rect 45833 37887 45891 37893
rect 41472 37828 42196 37856
rect 45848 37856 45876 37887
rect 46014 37884 46020 37936
rect 46072 37924 46078 37936
rect 47581 37927 47639 37933
rect 46072 37896 47532 37924
rect 46072 37884 46078 37896
rect 46109 37859 46167 37865
rect 46109 37856 46121 37859
rect 45848 37828 46121 37856
rect 41472 37816 41478 37828
rect 46109 37825 46121 37828
rect 46155 37856 46167 37859
rect 47504 37856 47532 37896
rect 47581 37893 47593 37927
rect 47627 37924 47639 37927
rect 49234 37924 49240 37936
rect 47627 37896 49240 37924
rect 47627 37893 47639 37896
rect 47581 37887 47639 37893
rect 49234 37884 49240 37896
rect 49292 37884 49298 37936
rect 53484 37924 53512 37964
rect 53558 37952 53564 38004
rect 53616 37992 53622 38004
rect 54849 37995 54907 38001
rect 54849 37992 54861 37995
rect 53616 37964 54861 37992
rect 53616 37952 53622 37964
rect 54849 37961 54861 37964
rect 54895 37961 54907 37995
rect 54849 37955 54907 37961
rect 56965 37995 57023 38001
rect 56965 37961 56977 37995
rect 57011 37992 57023 37995
rect 57011 37964 57744 37992
rect 57011 37961 57023 37964
rect 56965 37955 57023 37961
rect 57333 37927 57391 37933
rect 57333 37924 57345 37927
rect 53484 37896 57345 37924
rect 57333 37893 57345 37896
rect 57379 37924 57391 37927
rect 57517 37927 57575 37933
rect 57517 37924 57529 37927
rect 57379 37896 57529 37924
rect 57379 37893 57391 37896
rect 57333 37887 57391 37893
rect 57517 37893 57529 37896
rect 57563 37893 57575 37927
rect 57517 37887 57575 37893
rect 51810 37856 51816 37868
rect 46155 37828 46612 37856
rect 47504 37828 51816 37856
rect 46155 37825 46167 37828
rect 46109 37819 46167 37825
rect 25148 37760 25360 37788
rect 25498 37748 25504 37800
rect 25556 37788 25562 37800
rect 25961 37791 26019 37797
rect 25961 37788 25973 37791
rect 25556 37760 25973 37788
rect 25556 37748 25562 37760
rect 25961 37757 25973 37760
rect 26007 37757 26019 37791
rect 25961 37751 26019 37757
rect 26050 37748 26056 37800
rect 26108 37788 26114 37800
rect 26513 37791 26571 37797
rect 26108 37760 26153 37788
rect 26108 37748 26114 37760
rect 26513 37757 26525 37791
rect 26559 37757 26571 37791
rect 26513 37751 26571 37757
rect 26697 37791 26755 37797
rect 26697 37757 26709 37791
rect 26743 37757 26755 37791
rect 26697 37751 26755 37757
rect 25406 37680 25412 37732
rect 25464 37720 25470 37732
rect 26528 37720 26556 37751
rect 25464 37692 26556 37720
rect 26712 37720 26740 37751
rect 26878 37748 26884 37800
rect 26936 37788 26942 37800
rect 29086 37788 29092 37800
rect 26936 37760 29092 37788
rect 26936 37748 26942 37760
rect 29086 37748 29092 37760
rect 29144 37748 29150 37800
rect 29270 37788 29276 37800
rect 29328 37797 29334 37800
rect 29238 37760 29276 37788
rect 29270 37748 29276 37760
rect 29328 37751 29338 37797
rect 30742 37788 30748 37800
rect 29380 37760 30748 37788
rect 29328 37748 29334 37751
rect 27062 37720 27068 37732
rect 26712 37692 27068 37720
rect 25464 37680 25470 37692
rect 27062 37680 27068 37692
rect 27120 37720 27126 37732
rect 29380 37720 29408 37760
rect 30742 37748 30748 37760
rect 30800 37748 30806 37800
rect 32493 37791 32551 37797
rect 32493 37757 32505 37791
rect 32539 37788 32551 37791
rect 36630 37788 36636 37800
rect 32539 37760 36636 37788
rect 32539 37757 32551 37760
rect 32493 37751 32551 37757
rect 36630 37748 36636 37760
rect 36688 37748 36694 37800
rect 37185 37791 37243 37797
rect 37185 37757 37197 37791
rect 37231 37788 37243 37791
rect 38010 37788 38016 37800
rect 37231 37760 38016 37788
rect 37231 37757 37243 37760
rect 37185 37751 37243 37757
rect 38010 37748 38016 37760
rect 38068 37748 38074 37800
rect 40586 37748 40592 37800
rect 40644 37788 40650 37800
rect 41874 37788 41880 37800
rect 40644 37760 41880 37788
rect 40644 37748 40650 37760
rect 41874 37748 41880 37760
rect 41932 37788 41938 37800
rect 41969 37791 42027 37797
rect 41969 37788 41981 37791
rect 41932 37760 41981 37788
rect 41932 37748 41938 37760
rect 41969 37757 41981 37760
rect 42015 37757 42027 37791
rect 41969 37751 42027 37757
rect 42061 37791 42119 37797
rect 42061 37757 42073 37791
rect 42107 37757 42119 37791
rect 42061 37751 42119 37757
rect 42429 37791 42487 37797
rect 42429 37757 42441 37791
rect 42475 37757 42487 37791
rect 42429 37751 42487 37757
rect 42521 37791 42579 37797
rect 42521 37757 42533 37791
rect 42567 37788 42579 37791
rect 42610 37788 42616 37800
rect 42567 37760 42616 37788
rect 42567 37757 42579 37760
rect 42521 37751 42579 37757
rect 30374 37720 30380 37732
rect 27120 37692 29408 37720
rect 30208 37692 30380 37720
rect 27120 37680 27126 37692
rect 4522 37652 4528 37664
rect 4483 37624 4528 37652
rect 4522 37612 4528 37624
rect 4580 37612 4586 37664
rect 4614 37612 4620 37664
rect 4672 37652 4678 37664
rect 5261 37655 5319 37661
rect 5261 37652 5273 37655
rect 4672 37624 5273 37652
rect 4672 37612 4678 37624
rect 5261 37621 5273 37624
rect 5307 37621 5319 37655
rect 6914 37652 6920 37664
rect 6875 37624 6920 37652
rect 5261 37615 5319 37621
rect 6914 37612 6920 37624
rect 6972 37612 6978 37664
rect 15562 37652 15568 37664
rect 15523 37624 15568 37652
rect 15562 37612 15568 37624
rect 15620 37612 15626 37664
rect 16298 37612 16304 37664
rect 16356 37652 16362 37664
rect 17221 37655 17279 37661
rect 17221 37652 17233 37655
rect 16356 37624 17233 37652
rect 16356 37612 16362 37624
rect 17221 37621 17233 37624
rect 17267 37652 17279 37655
rect 23477 37655 23535 37661
rect 23477 37652 23489 37655
rect 17267 37624 23489 37652
rect 17267 37621 17279 37624
rect 17221 37615 17279 37621
rect 23477 37621 23489 37624
rect 23523 37621 23535 37655
rect 25498 37652 25504 37664
rect 25459 37624 25504 37652
rect 23477 37615 23535 37621
rect 25498 37612 25504 37624
rect 25556 37612 25562 37664
rect 25685 37655 25743 37661
rect 25685 37621 25697 37655
rect 25731 37652 25743 37655
rect 26050 37652 26056 37664
rect 25731 37624 26056 37652
rect 25731 37621 25743 37624
rect 25685 37615 25743 37621
rect 26050 37612 26056 37624
rect 26108 37612 26114 37664
rect 26694 37612 26700 37664
rect 26752 37652 26758 37664
rect 30208 37652 30236 37692
rect 30374 37680 30380 37692
rect 30432 37680 30438 37732
rect 31757 37723 31815 37729
rect 31757 37689 31769 37723
rect 31803 37720 31815 37723
rect 33410 37720 33416 37732
rect 31803 37692 33416 37720
rect 31803 37689 31815 37692
rect 31757 37683 31815 37689
rect 33410 37680 33416 37692
rect 33468 37680 33474 37732
rect 36538 37680 36544 37732
rect 36596 37720 36602 37732
rect 41693 37723 41751 37729
rect 41693 37720 41705 37723
rect 36596 37692 41705 37720
rect 36596 37680 36602 37692
rect 41693 37689 41705 37692
rect 41739 37720 41751 37723
rect 42076 37720 42104 37751
rect 41739 37692 42104 37720
rect 41739 37689 41751 37692
rect 41693 37683 41751 37689
rect 26752 37624 30236 37652
rect 26752 37612 26758 37624
rect 30282 37612 30288 37664
rect 30340 37652 30346 37664
rect 31021 37655 31079 37661
rect 31021 37652 31033 37655
rect 30340 37624 31033 37652
rect 30340 37612 30346 37624
rect 31021 37621 31033 37624
rect 31067 37621 31079 37655
rect 31570 37652 31576 37664
rect 31531 37624 31576 37652
rect 31021 37615 31079 37621
rect 31570 37612 31576 37624
rect 31628 37612 31634 37664
rect 38194 37612 38200 37664
rect 38252 37652 38258 37664
rect 41414 37652 41420 37664
rect 38252 37624 41420 37652
rect 38252 37612 38258 37624
rect 41414 37612 41420 37624
rect 41472 37612 41478 37664
rect 41509 37655 41567 37661
rect 41509 37621 41521 37655
rect 41555 37652 41567 37655
rect 41598 37652 41604 37664
rect 41555 37624 41604 37652
rect 41555 37621 41567 37624
rect 41509 37615 41567 37621
rect 41598 37612 41604 37624
rect 41656 37652 41662 37664
rect 42444 37652 42472 37751
rect 42610 37748 42616 37760
rect 42668 37748 42674 37800
rect 46584 37797 46612 37828
rect 51810 37816 51816 37828
rect 51868 37856 51874 37868
rect 53374 37856 53380 37868
rect 51868 37828 53380 37856
rect 51868 37816 51874 37828
rect 53374 37816 53380 37828
rect 53432 37816 53438 37868
rect 54018 37856 54024 37868
rect 53979 37828 54024 37856
rect 54018 37816 54024 37828
rect 54076 37816 54082 37868
rect 46385 37791 46443 37797
rect 46385 37757 46397 37791
rect 46431 37757 46443 37791
rect 46385 37751 46443 37757
rect 46569 37791 46627 37797
rect 46569 37757 46581 37791
rect 46615 37788 46627 37791
rect 47121 37791 47179 37797
rect 47121 37788 47133 37791
rect 46615 37760 47133 37788
rect 46615 37757 46627 37760
rect 46569 37751 46627 37757
rect 47121 37757 47133 37760
rect 47167 37757 47179 37791
rect 47121 37751 47179 37757
rect 47305 37791 47363 37797
rect 47305 37757 47317 37791
rect 47351 37788 47363 37791
rect 47670 37788 47676 37800
rect 47351 37760 47676 37788
rect 47351 37757 47363 37760
rect 47305 37751 47363 37757
rect 43073 37723 43131 37729
rect 43073 37689 43085 37723
rect 43119 37720 43131 37723
rect 44174 37720 44180 37732
rect 43119 37692 44180 37720
rect 43119 37689 43131 37692
rect 43073 37683 43131 37689
rect 44174 37680 44180 37692
rect 44232 37680 44238 37732
rect 46106 37680 46112 37732
rect 46164 37720 46170 37732
rect 46290 37720 46296 37732
rect 46164 37692 46296 37720
rect 46164 37680 46170 37692
rect 46290 37680 46296 37692
rect 46348 37720 46354 37732
rect 46400 37720 46428 37751
rect 46348 37692 46428 37720
rect 47136 37720 47164 37751
rect 47670 37748 47676 37760
rect 47728 37748 47734 37800
rect 48593 37791 48651 37797
rect 48593 37757 48605 37791
rect 48639 37788 48651 37791
rect 48682 37788 48688 37800
rect 48639 37760 48688 37788
rect 48639 37757 48651 37760
rect 48593 37751 48651 37757
rect 48682 37748 48688 37760
rect 48740 37748 48746 37800
rect 51994 37748 52000 37800
rect 52052 37788 52058 37800
rect 52273 37791 52331 37797
rect 52273 37788 52285 37791
rect 52052 37760 52285 37788
rect 52052 37748 52058 37760
rect 52273 37757 52285 37760
rect 52319 37757 52331 37791
rect 52549 37791 52607 37797
rect 52549 37788 52561 37791
rect 52273 37751 52331 37757
rect 52380 37760 52561 37788
rect 51902 37720 51908 37732
rect 47136 37692 51908 37720
rect 46348 37680 46354 37692
rect 51902 37680 51908 37692
rect 51960 37680 51966 37732
rect 52380 37720 52408 37760
rect 52549 37757 52561 37760
rect 52595 37757 52607 37791
rect 52549 37751 52607 37757
rect 52638 37748 52644 37800
rect 52696 37788 52702 37800
rect 53650 37788 53656 37800
rect 52696 37760 53656 37788
rect 52696 37748 52702 37760
rect 53650 37748 53656 37760
rect 53708 37748 53714 37800
rect 53926 37788 53932 37800
rect 53839 37760 53932 37788
rect 53926 37748 53932 37760
rect 53984 37788 53990 37800
rect 54757 37791 54815 37797
rect 54757 37788 54769 37791
rect 53984 37760 54769 37788
rect 53984 37748 53990 37760
rect 54757 37757 54769 37760
rect 54803 37757 54815 37791
rect 57532 37788 57560 37887
rect 57716 37868 57744 37964
rect 58710 37952 58716 38004
rect 58768 37992 58774 38004
rect 58768 37964 61700 37992
rect 58768 37952 58774 37964
rect 57698 37816 57704 37868
rect 57756 37856 57762 37868
rect 58989 37859 59047 37865
rect 57756 37828 57849 37856
rect 57756 37816 57762 37828
rect 58989 37825 59001 37859
rect 59035 37856 59047 37859
rect 60553 37859 60611 37865
rect 60553 37856 60565 37859
rect 59035 37828 60565 37856
rect 59035 37825 59047 37828
rect 58989 37819 59047 37825
rect 60553 37825 60565 37828
rect 60599 37825 60611 37859
rect 61672 37856 61700 37964
rect 61746 37952 61752 38004
rect 61804 37992 61810 38004
rect 61841 37995 61899 38001
rect 61841 37992 61853 37995
rect 61804 37964 61853 37992
rect 61804 37952 61810 37964
rect 61841 37961 61853 37964
rect 61887 37992 61899 37995
rect 64414 37992 64420 38004
rect 61887 37964 64420 37992
rect 61887 37961 61899 37964
rect 61841 37955 61899 37961
rect 64414 37952 64420 37964
rect 64472 37952 64478 38004
rect 65150 37992 65156 38004
rect 65111 37964 65156 37992
rect 65150 37952 65156 37964
rect 65208 37952 65214 38004
rect 69014 37952 69020 38004
rect 69072 37992 69078 38004
rect 69109 37995 69167 38001
rect 69109 37992 69121 37995
rect 69072 37964 69121 37992
rect 69072 37952 69078 37964
rect 69109 37961 69121 37964
rect 69155 37961 69167 37995
rect 69109 37955 69167 37961
rect 70302 37952 70308 38004
rect 70360 37992 70366 38004
rect 72053 37995 72111 38001
rect 72053 37992 72065 37995
rect 70360 37964 72065 37992
rect 70360 37952 70366 37964
rect 72053 37961 72065 37964
rect 72099 37961 72111 37995
rect 72053 37955 72111 37961
rect 76098 37952 76104 38004
rect 76156 37992 76162 38004
rect 77110 37992 77116 38004
rect 76156 37964 77116 37992
rect 76156 37952 76162 37964
rect 77110 37952 77116 37964
rect 77168 37952 77174 38004
rect 83734 37952 83740 38004
rect 83792 37992 83798 38004
rect 83829 37995 83887 38001
rect 83829 37992 83841 37995
rect 83792 37964 83841 37992
rect 83792 37952 83798 37964
rect 83829 37961 83841 37964
rect 83875 37961 83887 37995
rect 83829 37955 83887 37961
rect 86310 37952 86316 38004
rect 86368 37992 86374 38004
rect 86865 37995 86923 38001
rect 86865 37992 86877 37995
rect 86368 37964 86877 37992
rect 86368 37952 86374 37964
rect 86865 37961 86877 37964
rect 86911 37961 86923 37995
rect 86865 37955 86923 37961
rect 65705 37927 65763 37933
rect 65705 37924 65717 37927
rect 64064 37896 65717 37924
rect 64064 37865 64092 37896
rect 65705 37893 65717 37896
rect 65751 37893 65763 37927
rect 65705 37887 65763 37893
rect 64049 37859 64107 37865
rect 64049 37856 64061 37859
rect 61672 37828 64061 37856
rect 60553 37819 60611 37825
rect 64049 37825 64061 37828
rect 64095 37825 64107 37859
rect 64506 37856 64512 37868
rect 64467 37828 64512 37856
rect 64049 37819 64107 37825
rect 64506 37816 64512 37828
rect 64564 37856 64570 37868
rect 75730 37856 75736 37868
rect 64564 37828 65656 37856
rect 64564 37816 64570 37828
rect 57885 37791 57943 37797
rect 57885 37788 57897 37791
rect 57532 37760 57897 37788
rect 54757 37751 54815 37757
rect 57885 37757 57897 37760
rect 57931 37788 57943 37791
rect 58437 37791 58495 37797
rect 58437 37788 58449 37791
rect 57931 37760 58449 37788
rect 57931 37757 57943 37760
rect 57885 37751 57943 37757
rect 58437 37757 58449 37760
rect 58483 37757 58495 37791
rect 58618 37788 58624 37800
rect 58579 37760 58624 37788
rect 58437 37751 58495 37757
rect 58618 37748 58624 37760
rect 58676 37748 58682 37800
rect 60274 37788 60280 37800
rect 60235 37760 60280 37788
rect 60274 37748 60280 37760
rect 60332 37748 60338 37800
rect 61838 37788 61844 37800
rect 60384 37760 61844 37788
rect 58636 37720 58664 37748
rect 60384 37720 60412 37760
rect 61838 37748 61844 37760
rect 61896 37748 61902 37800
rect 64233 37791 64291 37797
rect 64233 37757 64245 37791
rect 64279 37757 64291 37791
rect 64233 37751 64291 37757
rect 64601 37791 64659 37797
rect 64601 37757 64613 37791
rect 64647 37788 64659 37791
rect 65150 37788 65156 37800
rect 64647 37760 65156 37788
rect 64647 37757 64659 37760
rect 64601 37751 64659 37757
rect 52104 37692 52408 37720
rect 53944 37692 54248 37720
rect 58636 37692 60412 37720
rect 52104 37664 52132 37692
rect 41656 37624 42472 37652
rect 43349 37655 43407 37661
rect 41656 37612 41662 37624
rect 43349 37621 43361 37655
rect 43395 37652 43407 37655
rect 43438 37652 43444 37664
rect 43395 37624 43444 37652
rect 43395 37621 43407 37624
rect 43349 37615 43407 37621
rect 43438 37612 43444 37624
rect 43496 37612 43502 37664
rect 47026 37612 47032 37664
rect 47084 37652 47090 37664
rect 48685 37655 48743 37661
rect 48685 37652 48697 37655
rect 47084 37624 48697 37652
rect 47084 37612 47090 37624
rect 48685 37621 48697 37624
rect 48731 37621 48743 37655
rect 52086 37652 52092 37664
rect 52047 37624 52092 37652
rect 48685 37615 48743 37621
rect 52086 37612 52092 37624
rect 52144 37612 52150 37664
rect 52178 37612 52184 37664
rect 52236 37652 52242 37664
rect 53944 37652 53972 37692
rect 52236 37624 53972 37652
rect 54220 37652 54248 37692
rect 62114 37680 62120 37732
rect 62172 37720 62178 37732
rect 63589 37723 63647 37729
rect 63589 37720 63601 37723
rect 62172 37692 63601 37720
rect 62172 37680 62178 37692
rect 63589 37689 63601 37692
rect 63635 37689 63647 37723
rect 64248 37720 64276 37751
rect 65150 37748 65156 37760
rect 65208 37748 65214 37800
rect 65628 37797 65656 37828
rect 65720 37828 75736 37856
rect 65613 37791 65671 37797
rect 65613 37757 65625 37791
rect 65659 37757 65671 37791
rect 65613 37751 65671 37757
rect 64874 37720 64880 37732
rect 64248 37692 64880 37720
rect 63589 37683 63647 37689
rect 64874 37680 64880 37692
rect 64932 37720 64938 37732
rect 64969 37723 65027 37729
rect 64969 37720 64981 37723
rect 64932 37692 64981 37720
rect 64932 37680 64938 37692
rect 64969 37689 64981 37692
rect 65015 37720 65027 37723
rect 65720 37720 65748 37828
rect 75730 37816 75736 37828
rect 75788 37816 75794 37868
rect 78033 37859 78091 37865
rect 78033 37856 78045 37859
rect 75932 37828 78045 37856
rect 69014 37748 69020 37800
rect 69072 37788 69078 37800
rect 69293 37791 69351 37797
rect 69293 37788 69305 37791
rect 69072 37760 69305 37788
rect 69072 37748 69078 37760
rect 69293 37757 69305 37760
rect 69339 37757 69351 37791
rect 69566 37788 69572 37800
rect 69527 37760 69572 37788
rect 69293 37751 69351 37757
rect 69566 37748 69572 37760
rect 69624 37748 69630 37800
rect 71961 37791 72019 37797
rect 71961 37788 71973 37791
rect 71608 37760 71973 37788
rect 65015 37692 65748 37720
rect 65015 37689 65027 37692
rect 64969 37683 65027 37689
rect 56965 37655 57023 37661
rect 56965 37652 56977 37655
rect 54220 37624 56977 37652
rect 52236 37612 52242 37624
rect 56965 37621 56977 37624
rect 57011 37652 57023 37655
rect 57057 37655 57115 37661
rect 57057 37652 57069 37655
rect 57011 37624 57069 37652
rect 57011 37621 57023 37624
rect 56965 37615 57023 37621
rect 57057 37621 57069 37624
rect 57103 37621 57115 37655
rect 57057 37615 57115 37621
rect 57146 37612 57152 37664
rect 57204 37652 57210 37664
rect 67450 37652 67456 37664
rect 57204 37624 67456 37652
rect 57204 37612 57210 37624
rect 67450 37612 67456 37624
rect 67508 37612 67514 37664
rect 70670 37652 70676 37664
rect 70631 37624 70676 37652
rect 70670 37612 70676 37624
rect 70728 37612 70734 37664
rect 71130 37612 71136 37664
rect 71188 37652 71194 37664
rect 71608 37661 71636 37760
rect 71961 37757 71973 37760
rect 72007 37757 72019 37791
rect 75638 37788 75644 37800
rect 75599 37760 75644 37788
rect 71961 37751 72019 37757
rect 75638 37748 75644 37760
rect 75696 37788 75702 37800
rect 75932 37797 75960 37828
rect 78033 37825 78045 37828
rect 78079 37856 78091 37859
rect 78398 37856 78404 37868
rect 78079 37828 78404 37856
rect 78079 37825 78091 37828
rect 78033 37819 78091 37825
rect 78398 37816 78404 37828
rect 78456 37816 78462 37868
rect 80330 37816 80336 37868
rect 80388 37856 80394 37868
rect 84746 37856 84752 37868
rect 80388 37828 84752 37856
rect 80388 37816 80394 37828
rect 84746 37816 84752 37828
rect 84804 37816 84810 37868
rect 85850 37856 85856 37868
rect 85811 37828 85856 37856
rect 85850 37816 85856 37828
rect 85908 37816 85914 37868
rect 87874 37856 87880 37868
rect 86052 37828 87880 37856
rect 75917 37791 75975 37797
rect 75917 37788 75929 37791
rect 75696 37760 75929 37788
rect 75696 37748 75702 37760
rect 75917 37757 75929 37760
rect 75963 37757 75975 37791
rect 75917 37751 75975 37757
rect 76653 37791 76711 37797
rect 76653 37757 76665 37791
rect 76699 37757 76711 37791
rect 76926 37788 76932 37800
rect 76887 37760 76932 37788
rect 76653 37751 76711 37757
rect 71682 37680 71688 37732
rect 71740 37720 71746 37732
rect 71777 37723 71835 37729
rect 71777 37720 71789 37723
rect 71740 37692 71789 37720
rect 71740 37680 71746 37692
rect 71777 37689 71789 37692
rect 71823 37689 71835 37723
rect 71777 37683 71835 37689
rect 71593 37655 71651 37661
rect 71593 37652 71605 37655
rect 71188 37624 71605 37652
rect 71188 37612 71194 37624
rect 71593 37621 71605 37624
rect 71639 37621 71651 37655
rect 71593 37615 71651 37621
rect 76561 37655 76619 37661
rect 76561 37621 76573 37655
rect 76607 37652 76619 37655
rect 76668 37652 76696 37751
rect 76926 37748 76932 37760
rect 76984 37748 76990 37800
rect 82722 37788 82728 37800
rect 82683 37760 82728 37788
rect 82722 37748 82728 37760
rect 82780 37748 82786 37800
rect 83737 37791 83795 37797
rect 83737 37757 83749 37791
rect 83783 37788 83795 37791
rect 84013 37791 84071 37797
rect 84013 37788 84025 37791
rect 83783 37760 84025 37788
rect 83783 37757 83795 37760
rect 83737 37751 83795 37757
rect 84013 37757 84025 37760
rect 84059 37757 84071 37791
rect 84013 37751 84071 37757
rect 82630 37680 82636 37732
rect 82688 37720 82694 37732
rect 83752 37720 83780 37751
rect 82688 37692 83780 37720
rect 84028 37720 84056 37751
rect 85298 37748 85304 37800
rect 85356 37788 85362 37800
rect 86052 37797 86080 37828
rect 87874 37816 87880 37828
rect 87932 37816 87938 37868
rect 85393 37791 85451 37797
rect 85393 37788 85405 37791
rect 85356 37760 85405 37788
rect 85356 37748 85362 37760
rect 85393 37757 85405 37760
rect 85439 37757 85451 37791
rect 85393 37751 85451 37757
rect 85577 37791 85635 37797
rect 85577 37757 85589 37791
rect 85623 37788 85635 37791
rect 86037 37791 86095 37797
rect 86037 37788 86049 37791
rect 85623 37760 86049 37788
rect 85623 37757 85635 37760
rect 85577 37751 85635 37757
rect 86037 37757 86049 37760
rect 86083 37757 86095 37791
rect 86770 37788 86776 37800
rect 86731 37760 86776 37788
rect 86037 37751 86095 37757
rect 85592 37720 85620 37751
rect 86770 37748 86776 37760
rect 86828 37748 86834 37800
rect 84028 37692 85620 37720
rect 82688 37680 82694 37692
rect 77938 37652 77944 37664
rect 76607 37624 77944 37652
rect 76607 37621 76619 37624
rect 76561 37615 76619 37621
rect 77938 37612 77944 37624
rect 77996 37612 78002 37664
rect 80146 37612 80152 37664
rect 80204 37652 80210 37664
rect 82814 37652 82820 37664
rect 80204 37624 82820 37652
rect 80204 37612 80210 37624
rect 82814 37612 82820 37624
rect 82872 37612 82878 37664
rect 1104 37562 111136 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 81046 37562
rect 81098 37510 81110 37562
rect 81162 37510 81174 37562
rect 81226 37510 81238 37562
rect 81290 37510 111136 37562
rect 1104 37488 111136 37510
rect 6733 37451 6791 37457
rect 6733 37448 6745 37451
rect 5000 37420 6745 37448
rect 4798 37272 4804 37324
rect 4856 37312 4862 37324
rect 5000 37321 5028 37420
rect 6733 37417 6745 37420
rect 6779 37417 6791 37451
rect 10042 37448 10048 37460
rect 10003 37420 10048 37448
rect 6733 37411 6791 37417
rect 10042 37408 10048 37420
rect 10100 37408 10106 37460
rect 11057 37451 11115 37457
rect 11057 37448 11069 37451
rect 10152 37420 11069 37448
rect 8294 37340 8300 37392
rect 8352 37380 8358 37392
rect 10152 37380 10180 37420
rect 11057 37417 11069 37420
rect 11103 37417 11115 37451
rect 15562 37448 15568 37460
rect 11057 37411 11115 37417
rect 15028 37420 15568 37448
rect 8352 37352 10180 37380
rect 8352 37340 8358 37352
rect 10962 37340 10968 37392
rect 11020 37380 11026 37392
rect 11020 37352 11652 37380
rect 11020 37340 11026 37352
rect 4985 37315 5043 37321
rect 4985 37312 4997 37315
rect 4856 37284 4997 37312
rect 4856 37272 4862 37284
rect 4985 37281 4997 37284
rect 5031 37281 5043 37315
rect 4985 37275 5043 37281
rect 5261 37315 5319 37321
rect 5261 37281 5273 37315
rect 5307 37312 5319 37315
rect 6914 37312 6920 37324
rect 5307 37284 6920 37312
rect 5307 37281 5319 37284
rect 5261 37275 5319 37281
rect 6914 37272 6920 37284
rect 6972 37272 6978 37324
rect 9858 37312 9864 37324
rect 9819 37284 9864 37312
rect 9858 37272 9864 37284
rect 9916 37272 9922 37324
rect 11422 37312 11428 37324
rect 11383 37284 11428 37312
rect 11422 37272 11428 37284
rect 11480 37272 11486 37324
rect 11624 37321 11652 37352
rect 13538 37340 13544 37392
rect 13596 37380 13602 37392
rect 15028 37389 15056 37420
rect 15013 37383 15071 37389
rect 15013 37380 15025 37383
rect 13596 37352 15025 37380
rect 13596 37340 13602 37352
rect 15013 37349 15025 37352
rect 15059 37349 15071 37383
rect 15013 37343 15071 37349
rect 11609 37315 11667 37321
rect 11609 37281 11621 37315
rect 11655 37281 11667 37315
rect 11974 37312 11980 37324
rect 11935 37284 11980 37312
rect 11609 37275 11667 37281
rect 11974 37272 11980 37284
rect 12032 37272 12038 37324
rect 15304 37321 15332 37420
rect 15562 37408 15568 37420
rect 15620 37408 15626 37460
rect 16482 37448 16488 37460
rect 16443 37420 16488 37448
rect 16482 37408 16488 37420
rect 16540 37408 16546 37460
rect 16574 37408 16580 37460
rect 16632 37448 16638 37460
rect 19889 37451 19947 37457
rect 19889 37448 19901 37451
rect 16632 37420 19901 37448
rect 16632 37408 16638 37420
rect 19889 37417 19901 37420
rect 19935 37417 19947 37451
rect 21082 37448 21088 37460
rect 20995 37420 21088 37448
rect 19889 37411 19947 37417
rect 21082 37408 21088 37420
rect 21140 37448 21146 37460
rect 25406 37448 25412 37460
rect 21140 37420 25412 37448
rect 21140 37408 21146 37420
rect 25406 37408 25412 37420
rect 25464 37408 25470 37460
rect 26050 37448 26056 37460
rect 26011 37420 26056 37448
rect 26050 37408 26056 37420
rect 26108 37408 26114 37460
rect 26142 37408 26148 37460
rect 26200 37448 26206 37460
rect 52086 37448 52092 37460
rect 26200 37420 52092 37448
rect 26200 37408 26206 37420
rect 52086 37408 52092 37420
rect 52144 37408 52150 37460
rect 52822 37408 52828 37460
rect 52880 37448 52886 37460
rect 54297 37451 54355 37457
rect 54297 37448 54309 37451
rect 52880 37420 54309 37448
rect 52880 37408 52886 37420
rect 54297 37417 54309 37420
rect 54343 37417 54355 37451
rect 57054 37448 57060 37460
rect 54297 37411 54355 37417
rect 54956 37420 57060 37448
rect 15378 37340 15384 37392
rect 15436 37380 15442 37392
rect 15436 37352 16252 37380
rect 15436 37340 15442 37352
rect 12161 37315 12219 37321
rect 12161 37281 12173 37315
rect 12207 37312 12219 37315
rect 15289 37315 15347 37321
rect 12207 37284 15240 37312
rect 12207 37281 12219 37284
rect 12161 37275 12219 37281
rect 3510 37204 3516 37256
rect 3568 37244 3574 37256
rect 4890 37244 4896 37256
rect 3568 37216 4896 37244
rect 3568 37204 3574 37216
rect 4890 37204 4896 37216
rect 4948 37204 4954 37256
rect 4062 37136 4068 37188
rect 4120 37176 4126 37188
rect 4706 37176 4712 37188
rect 4120 37148 4712 37176
rect 4120 37136 4126 37148
rect 4706 37136 4712 37148
rect 4764 37136 4770 37188
rect 15212 37176 15240 37284
rect 15289 37281 15301 37315
rect 15335 37281 15347 37315
rect 15470 37312 15476 37324
rect 15431 37284 15476 37312
rect 15289 37275 15347 37281
rect 15470 37272 15476 37284
rect 15528 37312 15534 37324
rect 16224 37321 16252 37352
rect 17770 37340 17776 37392
rect 17828 37380 17834 37392
rect 18785 37383 18843 37389
rect 17828 37352 18552 37380
rect 17828 37340 17834 37352
rect 16025 37315 16083 37321
rect 16025 37312 16037 37315
rect 15528 37284 16037 37312
rect 15528 37272 15534 37284
rect 16025 37281 16037 37284
rect 16071 37281 16083 37315
rect 16025 37275 16083 37281
rect 16209 37315 16267 37321
rect 16209 37281 16221 37315
rect 16255 37312 16267 37315
rect 16853 37315 16911 37321
rect 16853 37312 16865 37315
rect 16255 37284 16865 37312
rect 16255 37281 16267 37284
rect 16209 37275 16267 37281
rect 16853 37281 16865 37284
rect 16899 37312 16911 37315
rect 16942 37312 16948 37324
rect 16899 37284 16948 37312
rect 16899 37281 16911 37284
rect 16853 37275 16911 37281
rect 16942 37272 16948 37284
rect 17000 37272 17006 37324
rect 17678 37312 17684 37324
rect 17591 37284 17684 37312
rect 17678 37272 17684 37284
rect 17736 37312 17742 37324
rect 18233 37315 18291 37321
rect 18233 37312 18245 37315
rect 17736 37284 18245 37312
rect 17736 37272 17742 37284
rect 18233 37281 18245 37284
rect 18279 37281 18291 37315
rect 18414 37312 18420 37324
rect 18375 37284 18420 37312
rect 18233 37275 18291 37281
rect 18414 37272 18420 37284
rect 18472 37272 18478 37324
rect 18524 37312 18552 37352
rect 18785 37349 18797 37383
rect 18831 37380 18843 37383
rect 19242 37380 19248 37392
rect 18831 37352 19248 37380
rect 18831 37349 18843 37352
rect 18785 37343 18843 37349
rect 19242 37340 19248 37352
rect 19300 37340 19306 37392
rect 27801 37383 27859 37389
rect 19352 37352 27568 37380
rect 19352 37312 19380 37352
rect 18524 37284 19380 37312
rect 19797 37315 19855 37321
rect 19797 37281 19809 37315
rect 19843 37312 19855 37315
rect 20806 37312 20812 37324
rect 19843 37284 20812 37312
rect 19843 37281 19855 37284
rect 19797 37275 19855 37281
rect 20806 37272 20812 37284
rect 20864 37272 20870 37324
rect 20898 37272 20904 37324
rect 20956 37312 20962 37324
rect 21269 37315 21327 37321
rect 21269 37312 21281 37315
rect 20956 37284 21281 37312
rect 20956 37272 20962 37284
rect 21269 37281 21281 37284
rect 21315 37312 21327 37315
rect 21818 37312 21824 37324
rect 21315 37284 21824 37312
rect 21315 37281 21327 37284
rect 21269 37275 21327 37281
rect 21818 37272 21824 37284
rect 21876 37272 21882 37324
rect 25225 37315 25283 37321
rect 25225 37312 25237 37315
rect 25056 37284 25237 37312
rect 17497 37247 17555 37253
rect 17497 37244 17509 37247
rect 17328 37216 17509 37244
rect 16482 37176 16488 37188
rect 15212 37148 16488 37176
rect 16482 37136 16488 37148
rect 16540 37136 16546 37188
rect 6362 37108 6368 37120
rect 6323 37080 6368 37108
rect 6362 37068 6368 37080
rect 6420 37068 6426 37120
rect 14918 37068 14924 37120
rect 14976 37108 14982 37120
rect 17328 37117 17356 37216
rect 17497 37213 17509 37216
rect 17543 37213 17555 37247
rect 17497 37207 17555 37213
rect 24762 37136 24768 37188
rect 24820 37176 24826 37188
rect 25056 37185 25084 37284
rect 25225 37281 25237 37284
rect 25271 37281 25283 37315
rect 26237 37315 26295 37321
rect 26237 37312 26249 37315
rect 25225 37275 25283 37281
rect 25424 37284 26249 37312
rect 25424 37185 25452 37284
rect 26237 37281 26249 37284
rect 26283 37312 26295 37315
rect 26694 37312 26700 37324
rect 26283 37284 26700 37312
rect 26283 37281 26295 37284
rect 26237 37275 26295 37281
rect 26694 37272 26700 37284
rect 26752 37272 26758 37324
rect 27246 37312 27252 37324
rect 27207 37284 27252 37312
rect 27246 37272 27252 37284
rect 27304 37272 27310 37324
rect 27430 37312 27436 37324
rect 27391 37284 27436 37312
rect 27430 37272 27436 37284
rect 27488 37272 27494 37324
rect 27540 37312 27568 37352
rect 27801 37349 27813 37383
rect 27847 37380 27859 37383
rect 28350 37380 28356 37392
rect 27847 37352 28356 37380
rect 27847 37349 27859 37352
rect 27801 37343 27859 37349
rect 28350 37340 28356 37352
rect 28408 37340 28414 37392
rect 28994 37340 29000 37392
rect 29052 37380 29058 37392
rect 29825 37383 29883 37389
rect 29825 37380 29837 37383
rect 29052 37352 29837 37380
rect 29052 37340 29058 37352
rect 29825 37349 29837 37352
rect 29871 37349 29883 37383
rect 29825 37343 29883 37349
rect 30374 37340 30380 37392
rect 30432 37380 30438 37392
rect 36817 37383 36875 37389
rect 30432 37352 35296 37380
rect 30432 37340 30438 37352
rect 29641 37315 29699 37321
rect 29641 37312 29653 37315
rect 27540 37284 29653 37312
rect 29641 37281 29653 37284
rect 29687 37312 29699 37315
rect 29972 37315 30030 37321
rect 29972 37312 29984 37315
rect 29687 37284 29984 37312
rect 29687 37281 29699 37284
rect 29641 37275 29699 37281
rect 29972 37281 29984 37284
rect 30018 37281 30030 37315
rect 29972 37275 30030 37281
rect 30164 37315 30222 37321
rect 30164 37281 30176 37315
rect 30210 37312 30222 37315
rect 30834 37312 30840 37324
rect 30210 37284 30840 37312
rect 30210 37281 30222 37284
rect 30164 37275 30222 37281
rect 30834 37272 30840 37284
rect 30892 37272 30898 37324
rect 31662 37312 31668 37324
rect 31623 37284 31668 37312
rect 31662 37272 31668 37284
rect 31720 37312 31726 37324
rect 31757 37315 31815 37321
rect 31757 37312 31769 37315
rect 31720 37284 31769 37312
rect 31720 37272 31726 37284
rect 31757 37281 31769 37284
rect 31803 37281 31815 37315
rect 31757 37275 31815 37281
rect 34422 37272 34428 37324
rect 34480 37312 34486 37324
rect 34977 37315 35035 37321
rect 34977 37312 34989 37315
rect 34480 37284 34989 37312
rect 34480 37272 34486 37284
rect 34977 37281 34989 37284
rect 35023 37312 35035 37315
rect 35161 37315 35219 37321
rect 35161 37312 35173 37315
rect 35023 37284 35173 37312
rect 35023 37281 35035 37284
rect 34977 37275 35035 37281
rect 35161 37281 35173 37284
rect 35207 37281 35219 37315
rect 35268 37312 35296 37352
rect 36817 37349 36829 37383
rect 36863 37380 36875 37383
rect 37090 37380 37096 37392
rect 36863 37352 37096 37380
rect 36863 37349 36875 37352
rect 36817 37343 36875 37349
rect 37090 37340 37096 37352
rect 37148 37340 37154 37392
rect 39758 37340 39764 37392
rect 39816 37380 39822 37392
rect 40221 37383 40279 37389
rect 40221 37380 40233 37383
rect 39816 37352 40233 37380
rect 39816 37340 39822 37352
rect 40221 37349 40233 37352
rect 40267 37380 40279 37383
rect 41969 37383 42027 37389
rect 41969 37380 41981 37383
rect 40267 37352 40448 37380
rect 40267 37349 40279 37352
rect 40221 37343 40279 37349
rect 38194 37312 38200 37324
rect 35268 37284 38200 37312
rect 35161 37275 35219 37281
rect 38194 37272 38200 37284
rect 38252 37272 38258 37324
rect 38286 37272 38292 37324
rect 38344 37312 38350 37324
rect 40420 37321 40448 37352
rect 41156 37352 41981 37380
rect 40037 37315 40095 37321
rect 40037 37312 40049 37315
rect 38344 37284 40049 37312
rect 38344 37272 38350 37284
rect 40037 37281 40049 37284
rect 40083 37312 40095 37315
rect 40405 37315 40463 37321
rect 40083 37284 40356 37312
rect 40083 37281 40095 37284
rect 40037 37275 40095 37281
rect 26050 37204 26056 37256
rect 26108 37244 26114 37256
rect 26513 37247 26571 37253
rect 26513 37244 26525 37247
rect 26108 37216 26525 37244
rect 26108 37204 26114 37216
rect 26513 37213 26525 37216
rect 26559 37213 26571 37247
rect 35434 37244 35440 37256
rect 26513 37207 26571 37213
rect 27632 37216 35204 37244
rect 35395 37216 35440 37244
rect 25041 37179 25099 37185
rect 25041 37176 25053 37179
rect 24820 37148 25053 37176
rect 24820 37136 24826 37148
rect 25041 37145 25053 37148
rect 25087 37145 25099 37179
rect 25041 37139 25099 37145
rect 25409 37179 25467 37185
rect 25409 37145 25421 37179
rect 25455 37145 25467 37179
rect 25409 37139 25467 37145
rect 17313 37111 17371 37117
rect 17313 37108 17325 37111
rect 14976 37080 17325 37108
rect 14976 37068 14982 37080
rect 17313 37077 17325 37080
rect 17359 37077 17371 37111
rect 17313 37071 17371 37077
rect 21358 37068 21364 37120
rect 21416 37108 21422 37120
rect 27632 37108 27660 37216
rect 30101 37179 30159 37185
rect 30101 37145 30113 37179
rect 30147 37176 30159 37179
rect 30558 37176 30564 37188
rect 30147 37148 30564 37176
rect 30147 37145 30159 37148
rect 30101 37139 30159 37145
rect 30558 37136 30564 37148
rect 30616 37136 30622 37188
rect 30466 37108 30472 37120
rect 21416 37080 27660 37108
rect 30427 37080 30472 37108
rect 21416 37068 21422 37080
rect 30466 37068 30472 37080
rect 30524 37068 30530 37120
rect 31478 37108 31484 37120
rect 31439 37080 31484 37108
rect 31478 37068 31484 37080
rect 31536 37068 31542 37120
rect 34606 37068 34612 37120
rect 34664 37108 34670 37120
rect 34701 37111 34759 37117
rect 34701 37108 34713 37111
rect 34664 37080 34713 37108
rect 34664 37068 34670 37080
rect 34701 37077 34713 37080
rect 34747 37077 34759 37111
rect 35176 37108 35204 37216
rect 35434 37204 35440 37216
rect 35492 37204 35498 37256
rect 40328 37244 40356 37284
rect 40405 37281 40417 37315
rect 40451 37281 40463 37315
rect 40586 37312 40592 37324
rect 40547 37284 40592 37312
rect 40405 37275 40463 37281
rect 40586 37272 40592 37284
rect 40644 37272 40650 37324
rect 41156 37321 41184 37352
rect 41969 37349 41981 37352
rect 42015 37380 42027 37383
rect 42610 37380 42616 37392
rect 42015 37352 42616 37380
rect 42015 37349 42027 37352
rect 41969 37343 42027 37349
rect 42610 37340 42616 37352
rect 42668 37340 42674 37392
rect 47949 37383 48007 37389
rect 47949 37349 47961 37383
rect 47995 37380 48007 37383
rect 48682 37380 48688 37392
rect 47995 37352 48688 37380
rect 47995 37349 48007 37352
rect 47949 37343 48007 37349
rect 48682 37340 48688 37352
rect 48740 37340 48746 37392
rect 49694 37380 49700 37392
rect 49655 37352 49700 37380
rect 49694 37340 49700 37352
rect 49752 37380 49758 37392
rect 51537 37383 51595 37389
rect 49752 37352 50016 37380
rect 49752 37340 49758 37352
rect 41049 37315 41107 37321
rect 41049 37312 41061 37315
rect 40696 37284 41061 37312
rect 40696 37244 40724 37284
rect 41049 37281 41061 37284
rect 41095 37281 41107 37315
rect 41049 37275 41107 37281
rect 41141 37315 41199 37321
rect 41141 37281 41153 37315
rect 41187 37281 41199 37315
rect 41141 37275 41199 37281
rect 41874 37272 41880 37324
rect 41932 37312 41938 37324
rect 43346 37312 43352 37324
rect 41932 37284 43352 37312
rect 41932 37272 41938 37284
rect 43346 37272 43352 37284
rect 43404 37272 43410 37324
rect 46293 37315 46351 37321
rect 46293 37281 46305 37315
rect 46339 37312 46351 37315
rect 46569 37315 46627 37321
rect 46339 37284 46520 37312
rect 46339 37281 46351 37284
rect 46293 37275 46351 37281
rect 40328 37216 40724 37244
rect 46492 37244 46520 37284
rect 46569 37281 46581 37315
rect 46615 37312 46627 37315
rect 47210 37312 47216 37324
rect 46615 37284 47216 37312
rect 46615 37281 46627 37284
rect 46569 37275 46627 37281
rect 47210 37272 47216 37284
rect 47268 37272 47274 37324
rect 48041 37315 48099 37321
rect 48041 37312 48053 37315
rect 47320 37284 48053 37312
rect 47320 37244 47348 37284
rect 48041 37281 48053 37284
rect 48087 37312 48099 37315
rect 49881 37315 49939 37321
rect 49881 37312 49893 37315
rect 48087 37284 49893 37312
rect 48087 37281 48099 37284
rect 48041 37275 48099 37281
rect 49881 37281 49893 37284
rect 49927 37281 49939 37315
rect 49988 37312 50016 37352
rect 51537 37349 51549 37383
rect 51583 37380 51595 37383
rect 51718 37380 51724 37392
rect 51583 37352 51724 37380
rect 51583 37349 51595 37352
rect 51537 37343 51595 37349
rect 51718 37340 51724 37352
rect 51776 37380 51782 37392
rect 54312 37380 54340 37411
rect 51776 37352 53420 37380
rect 54312 37352 54708 37380
rect 51776 37340 51782 37352
rect 50157 37315 50215 37321
rect 50157 37312 50169 37315
rect 49988 37284 50169 37312
rect 49881 37275 49939 37281
rect 50157 37281 50169 37284
rect 50203 37281 50215 37315
rect 50982 37312 50988 37324
rect 50157 37275 50215 37281
rect 50264 37284 50988 37312
rect 46492 37216 47348 37244
rect 49896 37244 49924 37275
rect 50264 37244 50292 37284
rect 50982 37272 50988 37284
rect 51040 37312 51046 37324
rect 51629 37315 51687 37321
rect 51629 37312 51641 37315
rect 51040 37284 51641 37312
rect 51040 37272 51046 37284
rect 51629 37281 51641 37284
rect 51675 37312 51687 37315
rect 51994 37312 52000 37324
rect 51675 37284 52000 37312
rect 51675 37281 51687 37284
rect 51629 37275 51687 37281
rect 51994 37272 52000 37284
rect 52052 37272 52058 37324
rect 53006 37312 53012 37324
rect 52967 37284 53012 37312
rect 53006 37272 53012 37284
rect 53064 37272 53070 37324
rect 53098 37272 53104 37324
rect 53156 37312 53162 37324
rect 53392 37321 53420 37352
rect 53377 37315 53435 37321
rect 53156 37284 53201 37312
rect 53156 37272 53162 37284
rect 53377 37281 53389 37315
rect 53423 37281 53435 37315
rect 53377 37275 53435 37281
rect 53466 37272 53472 37324
rect 53524 37312 53530 37324
rect 53524 37284 53569 37312
rect 53524 37272 53530 37284
rect 53650 37272 53656 37324
rect 53708 37312 53714 37324
rect 54573 37315 54631 37321
rect 54573 37312 54585 37315
rect 53708 37284 54585 37312
rect 53708 37272 53714 37284
rect 54573 37281 54585 37284
rect 54619 37281 54631 37315
rect 54680 37312 54708 37352
rect 54956 37321 54984 37420
rect 57054 37408 57060 37420
rect 57112 37408 57118 37460
rect 57238 37448 57244 37460
rect 57199 37420 57244 37448
rect 57238 37408 57244 37420
rect 57296 37448 57302 37460
rect 57425 37451 57483 37457
rect 57425 37448 57437 37451
rect 57296 37420 57437 37448
rect 57296 37408 57302 37420
rect 57425 37417 57437 37420
rect 57471 37417 57483 37451
rect 57698 37448 57704 37460
rect 57659 37420 57704 37448
rect 57425 37411 57483 37417
rect 54803 37315 54861 37321
rect 54803 37312 54815 37315
rect 54680 37284 54815 37312
rect 54573 37275 54631 37281
rect 54803 37281 54815 37284
rect 54849 37281 54861 37315
rect 54803 37275 54861 37281
rect 54912 37315 54984 37321
rect 54912 37281 54924 37315
rect 54958 37284 54984 37315
rect 55306 37312 55312 37324
rect 55267 37284 55312 37312
rect 54958 37281 54970 37284
rect 54912 37275 54970 37281
rect 55306 37272 55312 37284
rect 55364 37272 55370 37324
rect 57440 37312 57468 37411
rect 57698 37408 57704 37420
rect 57756 37408 57762 37460
rect 57790 37408 57796 37460
rect 57848 37448 57854 37460
rect 60550 37448 60556 37460
rect 57848 37420 60556 37448
rect 57848 37408 57854 37420
rect 60550 37408 60556 37420
rect 60608 37408 60614 37460
rect 61838 37448 61844 37460
rect 61799 37420 61844 37448
rect 61838 37408 61844 37420
rect 61896 37408 61902 37460
rect 63037 37451 63095 37457
rect 63037 37417 63049 37451
rect 63083 37448 63095 37451
rect 64782 37448 64788 37460
rect 63083 37420 64788 37448
rect 63083 37417 63095 37420
rect 63037 37411 63095 37417
rect 64782 37408 64788 37420
rect 64840 37408 64846 37460
rect 67174 37448 67180 37460
rect 67135 37420 67180 37448
rect 67174 37408 67180 37420
rect 67232 37408 67238 37460
rect 67361 37451 67419 37457
rect 67361 37417 67373 37451
rect 67407 37448 67419 37451
rect 82630 37448 82636 37460
rect 67407 37420 82636 37448
rect 67407 37417 67419 37420
rect 67361 37411 67419 37417
rect 64046 37380 64052 37392
rect 63604 37352 64052 37380
rect 63604 37324 63632 37352
rect 64046 37340 64052 37352
rect 64104 37340 64110 37392
rect 67192 37380 67220 37408
rect 66456 37352 67220 37380
rect 66456 37324 66484 37352
rect 57977 37315 58035 37321
rect 57977 37312 57989 37315
rect 57440 37284 57989 37312
rect 57977 37281 57989 37284
rect 58023 37312 58035 37315
rect 58529 37315 58587 37321
rect 58529 37312 58541 37315
rect 58023 37284 58541 37312
rect 58023 37281 58035 37284
rect 57977 37275 58035 37281
rect 58529 37281 58541 37284
rect 58575 37281 58587 37315
rect 58710 37312 58716 37324
rect 58671 37284 58716 37312
rect 58529 37275 58587 37281
rect 58710 37272 58716 37284
rect 58768 37272 58774 37324
rect 61746 37312 61752 37324
rect 60660 37284 60780 37312
rect 61707 37284 61752 37312
rect 49896 37216 50292 37244
rect 50338 37204 50344 37256
rect 50396 37244 50402 37256
rect 50396 37216 53512 37244
rect 50396 37204 50402 37216
rect 53484 37176 53512 37216
rect 57698 37204 57704 37256
rect 57756 37244 57762 37256
rect 57793 37247 57851 37253
rect 57793 37244 57805 37247
rect 57756 37216 57805 37244
rect 57756 37204 57762 37216
rect 57793 37213 57805 37216
rect 57839 37213 57851 37247
rect 57793 37207 57851 37213
rect 59081 37247 59139 37253
rect 59081 37213 59093 37247
rect 59127 37244 59139 37247
rect 59814 37244 59820 37256
rect 59127 37216 59820 37244
rect 59127 37213 59139 37216
rect 59081 37207 59139 37213
rect 59814 37204 59820 37216
rect 59872 37204 59878 37256
rect 60660 37176 60688 37284
rect 60752 37244 60780 37284
rect 61746 37272 61752 37284
rect 61804 37272 61810 37324
rect 62574 37312 62580 37324
rect 62535 37284 62580 37312
rect 62574 37272 62580 37284
rect 62632 37312 62638 37324
rect 63221 37315 63279 37321
rect 63221 37312 63233 37315
rect 62632 37284 63233 37312
rect 62632 37272 62638 37284
rect 63221 37281 63233 37284
rect 63267 37281 63279 37315
rect 63221 37275 63279 37281
rect 63405 37315 63463 37321
rect 63405 37281 63417 37315
rect 63451 37312 63463 37315
rect 63586 37312 63592 37324
rect 63451 37284 63592 37312
rect 63451 37281 63463 37284
rect 63405 37275 63463 37281
rect 63586 37272 63592 37284
rect 63644 37272 63650 37324
rect 63678 37272 63684 37324
rect 63736 37312 63742 37324
rect 63773 37315 63831 37321
rect 63773 37312 63785 37315
rect 63736 37284 63785 37312
rect 63736 37272 63742 37284
rect 63773 37281 63785 37284
rect 63819 37281 63831 37315
rect 63773 37275 63831 37281
rect 63957 37315 64015 37321
rect 63957 37281 63969 37315
rect 64003 37312 64015 37315
rect 64322 37312 64328 37324
rect 64003 37284 64328 37312
rect 64003 37281 64015 37284
rect 63957 37275 64015 37281
rect 64322 37272 64328 37284
rect 64380 37272 64386 37324
rect 66254 37312 66260 37324
rect 66215 37284 66260 37312
rect 66254 37272 66260 37284
rect 66312 37272 66318 37324
rect 66438 37312 66444 37324
rect 66351 37284 66444 37312
rect 66438 37272 66444 37284
rect 66496 37272 66502 37324
rect 66622 37272 66628 37324
rect 66680 37312 66686 37324
rect 66809 37315 66867 37321
rect 66809 37312 66821 37315
rect 66680 37284 66821 37312
rect 66680 37272 66686 37284
rect 66809 37281 66821 37284
rect 66855 37312 66867 37315
rect 67376 37312 67404 37411
rect 82630 37408 82636 37420
rect 82688 37408 82694 37460
rect 82722 37408 82728 37460
rect 82780 37448 82786 37460
rect 84473 37451 84531 37457
rect 84473 37448 84485 37451
rect 82780 37420 84485 37448
rect 82780 37408 82786 37420
rect 84473 37417 84485 37420
rect 84519 37417 84531 37451
rect 84473 37411 84531 37417
rect 69477 37383 69535 37389
rect 69477 37349 69489 37383
rect 69523 37380 69535 37383
rect 69566 37380 69572 37392
rect 69523 37352 69572 37380
rect 69523 37349 69535 37352
rect 69477 37343 69535 37349
rect 69566 37340 69572 37352
rect 69624 37340 69630 37392
rect 71130 37380 71136 37392
rect 69676 37352 71136 37380
rect 66855 37284 67404 37312
rect 66855 37281 66867 37284
rect 66809 37275 66867 37281
rect 67450 37272 67456 37324
rect 67508 37312 67514 37324
rect 69106 37312 69112 37324
rect 67508 37284 69112 37312
rect 67508 37272 67514 37284
rect 69106 37272 69112 37284
rect 69164 37312 69170 37324
rect 69676 37312 69704 37352
rect 71130 37340 71136 37352
rect 71188 37380 71194 37392
rect 71188 37352 72004 37380
rect 71188 37340 71194 37352
rect 70026 37312 70032 37324
rect 69164 37284 69704 37312
rect 69987 37284 70032 37312
rect 69164 37272 69170 37284
rect 70026 37272 70032 37284
rect 70084 37272 70090 37324
rect 70118 37272 70124 37324
rect 70176 37321 70182 37324
rect 70176 37315 70225 37321
rect 70176 37281 70179 37315
rect 70213 37281 70225 37315
rect 70302 37312 70308 37324
rect 70263 37284 70308 37312
rect 70176 37275 70225 37281
rect 70176 37272 70182 37275
rect 70302 37272 70308 37284
rect 70360 37272 70366 37324
rect 71682 37312 71688 37324
rect 71643 37284 71688 37312
rect 71682 37272 71688 37284
rect 71740 37272 71746 37324
rect 71976 37321 72004 37352
rect 76926 37340 76932 37392
rect 76984 37380 76990 37392
rect 77757 37383 77815 37389
rect 77757 37380 77769 37383
rect 76984 37352 77769 37380
rect 76984 37340 76990 37352
rect 77757 37349 77769 37352
rect 77803 37349 77815 37383
rect 80330 37380 80336 37392
rect 77757 37343 77815 37349
rect 77864 37352 80336 37380
rect 71961 37315 72019 37321
rect 71961 37281 71973 37315
rect 72007 37281 72019 37315
rect 71961 37275 72019 37281
rect 72050 37272 72056 37324
rect 72108 37312 72114 37324
rect 75273 37315 75331 37321
rect 75273 37312 75285 37315
rect 72108 37284 75285 37312
rect 72108 37272 72114 37284
rect 75273 37281 75285 37284
rect 75319 37281 75331 37315
rect 77202 37312 77208 37324
rect 77163 37284 77208 37312
rect 75273 37275 75331 37281
rect 77202 37272 77208 37284
rect 77260 37272 77266 37324
rect 77338 37315 77396 37321
rect 77338 37281 77350 37315
rect 77384 37312 77396 37315
rect 77478 37312 77484 37324
rect 77384 37284 77484 37312
rect 77384 37281 77396 37284
rect 77338 37275 77396 37281
rect 77478 37272 77484 37284
rect 77536 37272 77542 37324
rect 66162 37244 66168 37256
rect 60752 37216 66168 37244
rect 66162 37204 66168 37216
rect 66220 37204 66226 37256
rect 66714 37244 66720 37256
rect 66675 37216 66720 37244
rect 66714 37204 66720 37216
rect 66772 37204 66778 37256
rect 75178 37244 75184 37256
rect 66824 37216 75184 37244
rect 66824 37176 66852 37216
rect 75178 37204 75184 37216
rect 75236 37204 75242 37256
rect 77021 37247 77079 37253
rect 77021 37213 77033 37247
rect 77067 37244 77079 37247
rect 77864 37244 77892 37352
rect 80330 37340 80336 37352
rect 80388 37340 80394 37392
rect 83182 37380 83188 37392
rect 81544 37352 83188 37380
rect 78585 37315 78643 37321
rect 78585 37281 78597 37315
rect 78631 37312 78643 37315
rect 78674 37312 78680 37324
rect 78631 37284 78680 37312
rect 78631 37281 78643 37284
rect 78585 37275 78643 37281
rect 78674 37272 78680 37284
rect 78732 37272 78738 37324
rect 81544 37321 81572 37352
rect 83182 37340 83188 37352
rect 83240 37340 83246 37392
rect 86402 37380 86408 37392
rect 84672 37352 86408 37380
rect 81529 37315 81587 37321
rect 78784 37284 81480 37312
rect 77067 37216 77892 37244
rect 77067 37213 77079 37216
rect 77021 37207 77079 37213
rect 36096 37148 46336 37176
rect 53484 37148 60688 37176
rect 62868 37148 66852 37176
rect 36096 37108 36124 37148
rect 35176 37080 36124 37108
rect 34701 37071 34759 37077
rect 40862 37068 40868 37120
rect 40920 37108 40926 37120
rect 41601 37111 41659 37117
rect 41601 37108 41613 37111
rect 40920 37080 41613 37108
rect 40920 37068 40926 37080
rect 41601 37077 41613 37080
rect 41647 37077 41659 37111
rect 41601 37071 41659 37077
rect 46017 37111 46075 37117
rect 46017 37077 46029 37111
rect 46063 37108 46075 37111
rect 46106 37108 46112 37120
rect 46063 37080 46112 37108
rect 46063 37077 46075 37080
rect 46017 37071 46075 37077
rect 46106 37068 46112 37080
rect 46164 37068 46170 37120
rect 46308 37108 46336 37148
rect 50982 37108 50988 37120
rect 46308 37080 50988 37108
rect 50982 37068 50988 37080
rect 51040 37068 51046 37120
rect 52454 37108 52460 37120
rect 52415 37080 52460 37108
rect 52454 37068 52460 37080
rect 52512 37068 52518 37120
rect 54386 37068 54392 37120
rect 54444 37108 54450 37120
rect 54711 37111 54769 37117
rect 54711 37108 54723 37111
rect 54444 37080 54723 37108
rect 54444 37068 54450 37080
rect 54711 37077 54723 37080
rect 54757 37077 54769 37111
rect 54711 37071 54769 37077
rect 54846 37068 54852 37120
rect 54904 37108 54910 37120
rect 62868 37108 62896 37148
rect 69934 37136 69940 37188
rect 69992 37176 69998 37188
rect 71501 37179 71559 37185
rect 71501 37176 71513 37179
rect 69992 37148 71513 37176
rect 69992 37136 69998 37148
rect 71501 37145 71513 37148
rect 71547 37145 71559 37179
rect 71501 37139 71559 37145
rect 75457 37179 75515 37185
rect 75457 37145 75469 37179
rect 75503 37176 75515 37179
rect 77036 37176 77064 37207
rect 77938 37204 77944 37256
rect 77996 37244 78002 37256
rect 78784 37244 78812 37284
rect 77996 37216 78812 37244
rect 77996 37204 78002 37216
rect 75503 37148 77064 37176
rect 81452 37176 81480 37284
rect 81529 37281 81541 37315
rect 81575 37281 81587 37315
rect 81529 37275 81587 37281
rect 81621 37315 81679 37321
rect 81621 37281 81633 37315
rect 81667 37312 81679 37315
rect 83369 37315 83427 37321
rect 83369 37312 83381 37315
rect 81667 37284 83381 37312
rect 81667 37281 81679 37284
rect 81621 37275 81679 37281
rect 83369 37281 83381 37284
rect 83415 37281 83427 37315
rect 84672 37312 84700 37352
rect 86402 37340 86408 37352
rect 86460 37380 86466 37392
rect 86862 37380 86868 37392
rect 86460 37352 86868 37380
rect 86460 37340 86466 37352
rect 86862 37340 86868 37352
rect 86920 37340 86926 37392
rect 83369 37275 83427 37281
rect 83476 37284 84700 37312
rect 83093 37247 83151 37253
rect 83093 37213 83105 37247
rect 83139 37244 83151 37247
rect 83476 37244 83504 37284
rect 84746 37272 84752 37324
rect 84804 37312 84810 37324
rect 84804 37284 85896 37312
rect 84804 37272 84810 37284
rect 83139 37216 83504 37244
rect 83139 37213 83151 37216
rect 83093 37207 83151 37213
rect 82909 37179 82967 37185
rect 82909 37176 82921 37179
rect 81452 37148 82921 37176
rect 75503 37145 75515 37148
rect 75457 37139 75515 37145
rect 82909 37145 82921 37148
rect 82955 37176 82967 37179
rect 83108 37176 83136 37207
rect 82955 37148 83136 37176
rect 85868 37176 85896 37284
rect 85942 37272 85948 37324
rect 86000 37312 86006 37324
rect 86129 37315 86187 37321
rect 86129 37312 86141 37315
rect 86000 37284 86141 37312
rect 86000 37272 86006 37284
rect 86129 37281 86141 37284
rect 86175 37281 86187 37315
rect 86129 37275 86187 37281
rect 86218 37272 86224 37324
rect 86276 37312 86282 37324
rect 86681 37315 86739 37321
rect 86276 37284 86321 37312
rect 86276 37272 86282 37284
rect 86681 37281 86693 37315
rect 86727 37312 86739 37315
rect 87414 37312 87420 37324
rect 86727 37284 87420 37312
rect 86727 37281 86739 37284
rect 86681 37275 86739 37281
rect 87414 37272 87420 37284
rect 87472 37272 87478 37324
rect 85945 37179 86003 37185
rect 85945 37176 85957 37179
rect 85868 37148 85957 37176
rect 82955 37145 82967 37148
rect 82909 37139 82967 37145
rect 85945 37145 85957 37148
rect 85991 37145 86003 37179
rect 85945 37139 86003 37145
rect 54904 37080 62896 37108
rect 54904 37068 54910 37080
rect 65978 37068 65984 37120
rect 66036 37108 66042 37120
rect 66073 37111 66131 37117
rect 66073 37108 66085 37111
rect 66036 37080 66085 37108
rect 66036 37068 66042 37080
rect 66073 37077 66085 37080
rect 66119 37077 66131 37111
rect 66073 37071 66131 37077
rect 66162 37068 66168 37120
rect 66220 37108 66226 37120
rect 67726 37108 67732 37120
rect 66220 37080 67732 37108
rect 66220 37068 66226 37080
rect 67726 37068 67732 37080
rect 67784 37068 67790 37120
rect 68646 37068 68652 37120
rect 68704 37108 68710 37120
rect 70670 37108 70676 37120
rect 68704 37080 70676 37108
rect 68704 37068 68710 37080
rect 70670 37068 70676 37080
rect 70728 37068 70734 37120
rect 77018 37068 77024 37120
rect 77076 37108 77082 37120
rect 78677 37111 78735 37117
rect 78677 37108 78689 37111
rect 77076 37080 78689 37108
rect 77076 37068 77082 37080
rect 78677 37077 78689 37080
rect 78723 37077 78735 37111
rect 78677 37071 78735 37077
rect 80422 37068 80428 37120
rect 80480 37108 80486 37120
rect 83550 37108 83556 37120
rect 80480 37080 83556 37108
rect 80480 37068 80486 37080
rect 83550 37068 83556 37080
rect 83608 37068 83614 37120
rect 1104 37018 111136 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 65686 37018
rect 65738 36966 65750 37018
rect 65802 36966 65814 37018
rect 65866 36966 65878 37018
rect 65930 36966 96406 37018
rect 96458 36966 96470 37018
rect 96522 36966 96534 37018
rect 96586 36966 96598 37018
rect 96650 36966 111136 37018
rect 1104 36944 111136 36966
rect 10870 36864 10876 36916
rect 10928 36904 10934 36916
rect 10965 36907 11023 36913
rect 10965 36904 10977 36907
rect 10928 36876 10977 36904
rect 10928 36864 10934 36876
rect 10965 36873 10977 36876
rect 11011 36873 11023 36907
rect 10965 36867 11023 36873
rect 18230 36864 18236 36916
rect 18288 36904 18294 36916
rect 18325 36907 18383 36913
rect 18325 36904 18337 36907
rect 18288 36876 18337 36904
rect 18288 36864 18294 36876
rect 18325 36873 18337 36876
rect 18371 36873 18383 36907
rect 26602 36904 26608 36916
rect 18325 36867 18383 36873
rect 18432 36876 26608 36904
rect 5534 36796 5540 36848
rect 5592 36836 5598 36848
rect 18432 36836 18460 36876
rect 26602 36864 26608 36876
rect 26660 36864 26666 36916
rect 30466 36864 30472 36916
rect 30524 36904 30530 36916
rect 41322 36904 41328 36916
rect 30524 36876 41328 36904
rect 30524 36864 30530 36876
rect 41322 36864 41328 36876
rect 41380 36864 41386 36916
rect 41506 36904 41512 36916
rect 41467 36876 41512 36904
rect 41506 36864 41512 36876
rect 41564 36864 41570 36916
rect 43990 36864 43996 36916
rect 44048 36904 44054 36916
rect 44637 36907 44695 36913
rect 44637 36904 44649 36907
rect 44048 36876 44649 36904
rect 44048 36864 44054 36876
rect 44637 36873 44649 36876
rect 44683 36873 44695 36907
rect 44637 36867 44695 36873
rect 46842 36864 46848 36916
rect 46900 36904 46906 36916
rect 51626 36904 51632 36916
rect 46900 36876 51632 36904
rect 46900 36864 46906 36876
rect 51626 36864 51632 36876
rect 51684 36864 51690 36916
rect 51810 36904 51816 36916
rect 51771 36876 51816 36904
rect 51810 36864 51816 36876
rect 51868 36864 51874 36916
rect 53101 36907 53159 36913
rect 53101 36873 53113 36907
rect 53147 36904 53159 36907
rect 54386 36904 54392 36916
rect 53147 36876 54392 36904
rect 53147 36873 53159 36876
rect 53101 36867 53159 36873
rect 54386 36864 54392 36876
rect 54444 36864 54450 36916
rect 54478 36864 54484 36916
rect 54536 36904 54542 36916
rect 60642 36904 60648 36916
rect 54536 36876 60648 36904
rect 54536 36864 54542 36876
rect 60642 36864 60648 36876
rect 60700 36864 60706 36916
rect 60734 36864 60740 36916
rect 60792 36904 60798 36916
rect 61197 36907 61255 36913
rect 60792 36876 61148 36904
rect 60792 36864 60798 36876
rect 5592 36808 18460 36836
rect 18785 36839 18843 36845
rect 5592 36796 5598 36808
rect 18785 36805 18797 36839
rect 18831 36836 18843 36839
rect 21358 36836 21364 36848
rect 18831 36808 21364 36836
rect 18831 36805 18843 36808
rect 18785 36799 18843 36805
rect 15470 36768 15476 36780
rect 15304 36740 15476 36768
rect 5258 36700 5264 36712
rect 5219 36672 5264 36700
rect 5258 36660 5264 36672
rect 5316 36660 5322 36712
rect 5629 36703 5687 36709
rect 5629 36669 5641 36703
rect 5675 36700 5687 36703
rect 8846 36700 8852 36712
rect 5675 36672 8852 36700
rect 5675 36669 5687 36672
rect 5629 36663 5687 36669
rect 8846 36660 8852 36672
rect 8904 36660 8910 36712
rect 10778 36700 10784 36712
rect 10739 36672 10784 36700
rect 10778 36660 10784 36672
rect 10836 36660 10842 36712
rect 15304 36709 15332 36740
rect 15470 36728 15476 36740
rect 15528 36728 15534 36780
rect 18049 36771 18107 36777
rect 18049 36737 18061 36771
rect 18095 36768 18107 36771
rect 18414 36768 18420 36780
rect 18095 36740 18420 36768
rect 18095 36737 18107 36740
rect 18049 36731 18107 36737
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 15105 36703 15163 36709
rect 15105 36700 15117 36703
rect 14936 36672 15117 36700
rect 14936 36576 14964 36672
rect 15105 36669 15117 36672
rect 15151 36669 15163 36703
rect 15105 36663 15163 36669
rect 15289 36703 15347 36709
rect 15289 36669 15301 36703
rect 15335 36669 15347 36703
rect 15289 36663 15347 36669
rect 15841 36703 15899 36709
rect 15841 36669 15853 36703
rect 15887 36669 15899 36703
rect 15841 36663 15899 36669
rect 16025 36703 16083 36709
rect 16025 36669 16037 36703
rect 16071 36700 16083 36703
rect 16482 36700 16488 36712
rect 16071 36672 16488 36700
rect 16071 36669 16083 36672
rect 16025 36663 16083 36669
rect 15304 36632 15332 36663
rect 15856 36632 15884 36663
rect 16482 36660 16488 36672
rect 16540 36660 16546 36712
rect 17218 36660 17224 36712
rect 17276 36700 17282 36712
rect 18141 36703 18199 36709
rect 18141 36700 18153 36703
rect 17276 36672 18153 36700
rect 17276 36660 17282 36672
rect 18141 36669 18153 36672
rect 18187 36700 18199 36703
rect 18800 36700 18828 36799
rect 21358 36796 21364 36808
rect 21416 36796 21422 36848
rect 25406 36796 25412 36848
rect 25464 36836 25470 36848
rect 25464 36808 25728 36836
rect 25464 36796 25470 36808
rect 19429 36771 19487 36777
rect 19429 36737 19441 36771
rect 19475 36768 19487 36771
rect 19475 36740 19840 36768
rect 19475 36737 19487 36740
rect 19429 36731 19487 36737
rect 19812 36709 19840 36740
rect 18187 36672 18828 36700
rect 19705 36703 19763 36709
rect 18187 36669 18199 36672
rect 18141 36663 18199 36669
rect 19705 36669 19717 36703
rect 19751 36669 19763 36703
rect 19705 36663 19763 36669
rect 19797 36703 19855 36709
rect 19797 36669 19809 36703
rect 19843 36700 19855 36703
rect 19886 36700 19892 36712
rect 19843 36672 19892 36700
rect 19843 36669 19855 36672
rect 19797 36663 19855 36669
rect 15304 36604 15884 36632
rect 19720 36632 19748 36663
rect 19886 36660 19892 36672
rect 19944 36660 19950 36712
rect 20162 36700 20168 36712
rect 20123 36672 20168 36700
rect 20162 36660 20168 36672
rect 20220 36660 20226 36712
rect 20257 36703 20315 36709
rect 20257 36669 20269 36703
rect 20303 36700 20315 36703
rect 21082 36700 21088 36712
rect 20303 36672 21088 36700
rect 20303 36669 20315 36672
rect 20257 36663 20315 36669
rect 20272 36632 20300 36663
rect 21082 36660 21088 36672
rect 21140 36660 21146 36712
rect 21726 36700 21732 36712
rect 21687 36672 21732 36700
rect 21726 36660 21732 36672
rect 21784 36660 21790 36712
rect 25406 36660 25412 36712
rect 25464 36709 25470 36712
rect 25464 36703 25513 36709
rect 25464 36669 25467 36703
rect 25501 36669 25513 36703
rect 25590 36700 25596 36712
rect 25551 36672 25596 36700
rect 25464 36663 25513 36669
rect 25464 36660 25470 36663
rect 25590 36660 25596 36672
rect 25648 36660 25654 36712
rect 25700 36700 25728 36808
rect 33134 36796 33140 36848
rect 33192 36836 33198 36848
rect 34425 36839 34483 36845
rect 34425 36836 34437 36839
rect 33192 36808 34437 36836
rect 33192 36796 33198 36808
rect 34425 36805 34437 36808
rect 34471 36836 34483 36839
rect 34517 36839 34575 36845
rect 34517 36836 34529 36839
rect 34471 36808 34529 36836
rect 34471 36805 34483 36808
rect 34425 36799 34483 36805
rect 34517 36805 34529 36808
rect 34563 36836 34575 36839
rect 35986 36836 35992 36848
rect 34563 36808 35112 36836
rect 35947 36808 35992 36836
rect 34563 36805 34575 36808
rect 34517 36799 34575 36805
rect 27154 36728 27160 36780
rect 27212 36768 27218 36780
rect 27430 36768 27436 36780
rect 27212 36740 27436 36768
rect 27212 36728 27218 36740
rect 27430 36728 27436 36740
rect 27488 36728 27494 36780
rect 34606 36728 34612 36780
rect 34664 36768 34670 36780
rect 34885 36771 34943 36777
rect 34885 36768 34897 36771
rect 34664 36740 34897 36768
rect 34664 36728 34670 36740
rect 34885 36737 34897 36740
rect 34931 36737 34943 36771
rect 34885 36731 34943 36737
rect 35084 36709 35112 36808
rect 35986 36796 35992 36808
rect 36044 36796 36050 36848
rect 39758 36796 39764 36848
rect 39816 36836 39822 36848
rect 41141 36839 41199 36845
rect 41141 36836 41153 36839
rect 39816 36808 41153 36836
rect 39816 36796 39822 36808
rect 41141 36805 41153 36808
rect 41187 36805 41199 36839
rect 41141 36799 41199 36805
rect 41414 36796 41420 36848
rect 41472 36836 41478 36848
rect 44453 36839 44511 36845
rect 41472 36808 44404 36836
rect 41472 36796 41478 36808
rect 39482 36728 39488 36780
rect 39540 36768 39546 36780
rect 41012 36771 41070 36777
rect 41012 36768 41024 36771
rect 39540 36740 41024 36768
rect 39540 36728 39546 36740
rect 41012 36737 41024 36740
rect 41058 36737 41070 36771
rect 41012 36731 41070 36737
rect 41233 36771 41291 36777
rect 41233 36737 41245 36771
rect 41279 36768 41291 36771
rect 41690 36768 41696 36780
rect 41279 36740 41696 36768
rect 41279 36737 41291 36740
rect 41233 36731 41291 36737
rect 41690 36728 41696 36740
rect 41748 36728 41754 36780
rect 44376 36768 44404 36808
rect 44453 36805 44465 36839
rect 44499 36836 44511 36839
rect 46934 36836 46940 36848
rect 44499 36808 46940 36836
rect 44499 36805 44511 36808
rect 44453 36799 44511 36805
rect 46934 36796 46940 36808
rect 46992 36796 46998 36848
rect 47210 36836 47216 36848
rect 47171 36808 47216 36836
rect 47210 36796 47216 36808
rect 47268 36796 47274 36848
rect 47302 36796 47308 36848
rect 47360 36836 47366 36848
rect 50706 36836 50712 36848
rect 47360 36808 50712 36836
rect 47360 36796 47366 36808
rect 50706 36796 50712 36808
rect 50764 36796 50770 36848
rect 53466 36796 53472 36848
rect 53524 36836 53530 36848
rect 61120 36836 61148 36876
rect 61197 36873 61209 36907
rect 61243 36904 61255 36907
rect 70946 36904 70952 36916
rect 61243 36876 70952 36904
rect 61243 36873 61255 36876
rect 61197 36867 61255 36873
rect 70946 36864 70952 36876
rect 71004 36864 71010 36916
rect 71130 36904 71136 36916
rect 71091 36876 71136 36904
rect 71130 36864 71136 36876
rect 71188 36864 71194 36916
rect 77018 36904 77024 36916
rect 71424 36876 77024 36904
rect 71424 36836 71452 36876
rect 77018 36864 77024 36876
rect 77076 36864 77082 36916
rect 82906 36904 82912 36916
rect 82867 36876 82912 36904
rect 82906 36864 82912 36876
rect 82964 36864 82970 36916
rect 83182 36864 83188 36916
rect 83240 36904 83246 36916
rect 83277 36907 83335 36913
rect 83277 36904 83289 36907
rect 83240 36876 83289 36904
rect 83240 36864 83246 36876
rect 83277 36873 83289 36876
rect 83323 36873 83335 36907
rect 83918 36904 83924 36916
rect 83277 36867 83335 36873
rect 83384 36876 83924 36904
rect 53524 36808 54248 36836
rect 61120 36808 71452 36836
rect 53524 36796 53530 36808
rect 45557 36771 45615 36777
rect 45557 36768 45569 36771
rect 44376 36740 45569 36768
rect 45557 36737 45569 36740
rect 45603 36768 45615 36771
rect 45741 36771 45799 36777
rect 45741 36768 45753 36771
rect 45603 36740 45753 36768
rect 45603 36737 45615 36740
rect 45557 36731 45615 36737
rect 45741 36737 45753 36740
rect 45787 36768 45799 36771
rect 48869 36771 48927 36777
rect 45787 36740 46336 36768
rect 45787 36737 45799 36740
rect 45741 36731 45799 36737
rect 26053 36703 26111 36709
rect 26053 36700 26065 36703
rect 25700 36672 26065 36700
rect 26053 36669 26065 36672
rect 26099 36669 26111 36703
rect 26053 36663 26111 36669
rect 26237 36703 26295 36709
rect 26237 36669 26249 36703
rect 26283 36700 26295 36703
rect 26789 36703 26847 36709
rect 26789 36700 26801 36703
rect 26283 36672 26801 36700
rect 26283 36669 26295 36672
rect 26237 36663 26295 36669
rect 26789 36669 26801 36672
rect 26835 36700 26847 36703
rect 35069 36703 35127 36709
rect 26835 36672 35020 36700
rect 26835 36669 26847 36672
rect 26789 36663 26847 36669
rect 19720 36604 20300 36632
rect 20364 36604 21588 36632
rect 5166 36564 5172 36576
rect 5127 36536 5172 36564
rect 5166 36524 5172 36536
rect 5224 36524 5230 36576
rect 14918 36564 14924 36576
rect 14879 36536 14924 36564
rect 14918 36524 14924 36536
rect 14976 36524 14982 36576
rect 16301 36567 16359 36573
rect 16301 36533 16313 36567
rect 16347 36564 16359 36567
rect 19334 36564 19340 36576
rect 16347 36536 19340 36564
rect 16347 36533 16359 36536
rect 16301 36527 16359 36533
rect 19334 36524 19340 36536
rect 19392 36524 19398 36576
rect 20162 36524 20168 36576
rect 20220 36564 20226 36576
rect 20364 36564 20392 36604
rect 21560 36576 21588 36604
rect 24854 36592 24860 36644
rect 24912 36632 24918 36644
rect 26252 36632 26280 36663
rect 24912 36604 26280 36632
rect 26605 36635 26663 36641
rect 24912 36592 24918 36604
rect 26605 36601 26617 36635
rect 26651 36632 26663 36635
rect 32398 36632 32404 36644
rect 26651 36604 32404 36632
rect 26651 36601 26663 36604
rect 26605 36595 26663 36601
rect 32398 36592 32404 36604
rect 32456 36592 32462 36644
rect 20714 36564 20720 36576
rect 20220 36536 20392 36564
rect 20675 36536 20720 36564
rect 20220 36524 20226 36536
rect 20714 36524 20720 36536
rect 20772 36524 20778 36576
rect 21542 36524 21548 36576
rect 21600 36564 21606 36576
rect 21821 36567 21879 36573
rect 21821 36564 21833 36567
rect 21600 36536 21833 36564
rect 21600 36524 21606 36536
rect 21821 36533 21833 36536
rect 21867 36533 21879 36567
rect 21821 36527 21879 36533
rect 25225 36567 25283 36573
rect 25225 36533 25237 36567
rect 25271 36564 25283 36567
rect 25406 36564 25412 36576
rect 25271 36536 25412 36564
rect 25271 36533 25283 36536
rect 25225 36527 25283 36533
rect 25406 36524 25412 36536
rect 25464 36564 25470 36576
rect 25590 36564 25596 36576
rect 25464 36536 25596 36564
rect 25464 36524 25470 36536
rect 25590 36524 25596 36536
rect 25648 36524 25654 36576
rect 34992 36564 35020 36672
rect 35069 36669 35081 36703
rect 35115 36700 35127 36703
rect 35618 36700 35624 36712
rect 35115 36672 35624 36700
rect 35115 36669 35127 36672
rect 35069 36663 35127 36669
rect 35618 36660 35624 36672
rect 35676 36660 35682 36712
rect 35802 36700 35808 36712
rect 35763 36672 35808 36700
rect 35802 36660 35808 36672
rect 35860 36660 35866 36712
rect 35986 36660 35992 36712
rect 36044 36700 36050 36712
rect 41322 36700 41328 36712
rect 36044 36672 41328 36700
rect 36044 36660 36050 36672
rect 41322 36660 41328 36672
rect 41380 36660 41386 36712
rect 42429 36703 42487 36709
rect 42429 36700 42441 36703
rect 41432 36672 42441 36700
rect 40862 36592 40868 36644
rect 40920 36632 40926 36644
rect 40920 36604 40965 36632
rect 40920 36592 40926 36604
rect 36538 36564 36544 36576
rect 34992 36536 36544 36564
rect 36538 36524 36544 36536
rect 36596 36524 36602 36576
rect 36630 36524 36636 36576
rect 36688 36564 36694 36576
rect 41432 36564 41460 36672
rect 42429 36669 42441 36672
rect 42475 36700 42487 36703
rect 43990 36700 43996 36712
rect 42475 36672 43996 36700
rect 42475 36669 42487 36672
rect 42429 36663 42487 36669
rect 43990 36660 43996 36672
rect 44048 36660 44054 36712
rect 44174 36700 44180 36712
rect 44135 36672 44180 36700
rect 44174 36660 44180 36672
rect 44232 36660 44238 36712
rect 44542 36709 44548 36712
rect 44324 36703 44382 36709
rect 44324 36669 44336 36703
rect 44370 36669 44382 36703
rect 44324 36663 44382 36669
rect 44516 36703 44548 36709
rect 44516 36669 44528 36703
rect 44516 36663 44548 36669
rect 44339 36632 44367 36663
rect 44542 36660 44548 36663
rect 44600 36660 44606 36712
rect 46106 36700 46112 36712
rect 46067 36672 46112 36700
rect 46106 36660 46112 36672
rect 46164 36660 46170 36712
rect 46308 36709 46336 36740
rect 48869 36737 48881 36771
rect 48915 36768 48927 36771
rect 49234 36768 49240 36780
rect 48915 36740 49240 36768
rect 48915 36737 48927 36740
rect 48869 36731 48927 36737
rect 49234 36728 49240 36740
rect 49292 36728 49298 36780
rect 53742 36768 53748 36780
rect 53703 36740 53748 36768
rect 53742 36728 53748 36740
rect 53800 36728 53806 36780
rect 54113 36771 54171 36777
rect 54113 36737 54125 36771
rect 54159 36768 54171 36771
rect 54220 36768 54248 36808
rect 71498 36796 71504 36848
rect 71556 36836 71562 36848
rect 72881 36839 72939 36845
rect 72881 36836 72893 36839
rect 71556 36808 72893 36836
rect 71556 36796 71562 36808
rect 72881 36805 72893 36808
rect 72927 36805 72939 36839
rect 72881 36799 72939 36805
rect 75178 36796 75184 36848
rect 75236 36836 75242 36848
rect 80146 36836 80152 36848
rect 75236 36808 80152 36836
rect 75236 36796 75242 36808
rect 80146 36796 80152 36808
rect 80204 36796 80210 36848
rect 82924 36836 82952 36864
rect 83384 36836 83412 36876
rect 83918 36864 83924 36876
rect 83976 36864 83982 36916
rect 86954 36904 86960 36916
rect 86915 36876 86960 36904
rect 86954 36864 86960 36876
rect 87012 36864 87018 36916
rect 82924 36808 83412 36836
rect 54159 36740 54248 36768
rect 54159 36737 54171 36740
rect 54113 36731 54171 36737
rect 54294 36728 54300 36780
rect 54352 36768 54358 36780
rect 61197 36771 61255 36777
rect 61197 36768 61209 36771
rect 54352 36740 61209 36768
rect 54352 36728 54358 36740
rect 61197 36737 61209 36740
rect 61243 36737 61255 36771
rect 65061 36771 65119 36777
rect 65061 36768 65073 36771
rect 61197 36731 61255 36737
rect 61304 36740 65073 36768
rect 46293 36703 46351 36709
rect 46293 36669 46305 36703
rect 46339 36700 46351 36703
rect 46842 36700 46848 36712
rect 46339 36672 46848 36700
rect 46339 36669 46351 36672
rect 46293 36663 46351 36669
rect 46842 36660 46848 36672
rect 46900 36660 46906 36712
rect 47026 36700 47032 36712
rect 46987 36672 47032 36700
rect 47026 36660 47032 36672
rect 47084 36660 47090 36712
rect 48406 36660 48412 36712
rect 48464 36700 48470 36712
rect 48685 36703 48743 36709
rect 48685 36700 48697 36703
rect 48464 36672 48697 36700
rect 48464 36660 48470 36672
rect 48685 36669 48697 36672
rect 48731 36700 48743 36703
rect 48961 36703 49019 36709
rect 48961 36700 48973 36703
rect 48731 36672 48973 36700
rect 48731 36669 48743 36672
rect 48685 36663 48743 36669
rect 48961 36669 48973 36672
rect 49007 36669 49019 36703
rect 48961 36663 49019 36669
rect 49145 36703 49203 36709
rect 49145 36669 49157 36703
rect 49191 36669 49203 36703
rect 49252 36700 49280 36728
rect 49605 36703 49663 36709
rect 49605 36700 49617 36703
rect 49252 36672 49617 36700
rect 49145 36663 49203 36669
rect 49605 36669 49617 36672
rect 49651 36669 49663 36703
rect 49605 36663 49663 36669
rect 49160 36632 49188 36663
rect 49694 36660 49700 36712
rect 49752 36700 49758 36712
rect 50709 36703 50767 36709
rect 50709 36700 50721 36703
rect 49752 36672 50721 36700
rect 49752 36660 49758 36672
rect 50709 36669 50721 36672
rect 50755 36700 50767 36703
rect 50798 36700 50804 36712
rect 50755 36672 50804 36700
rect 50755 36669 50767 36672
rect 50709 36663 50767 36669
rect 50798 36660 50804 36672
rect 50856 36660 50862 36712
rect 51718 36700 51724 36712
rect 51679 36672 51724 36700
rect 51718 36660 51724 36672
rect 51776 36660 51782 36712
rect 53650 36700 53656 36712
rect 53611 36672 53656 36700
rect 53650 36660 53656 36672
rect 53708 36660 53714 36712
rect 53926 36660 53932 36712
rect 53984 36700 53990 36712
rect 54021 36703 54079 36709
rect 54021 36700 54033 36703
rect 53984 36672 54033 36700
rect 53984 36660 53990 36672
rect 54021 36669 54033 36672
rect 54067 36669 54079 36703
rect 54021 36663 54079 36669
rect 54202 36660 54208 36712
rect 54260 36700 54266 36712
rect 61102 36700 61108 36712
rect 54260 36672 61108 36700
rect 54260 36660 54266 36672
rect 61102 36660 61108 36672
rect 61160 36660 61166 36712
rect 61304 36709 61332 36740
rect 65061 36737 65073 36740
rect 65107 36737 65119 36771
rect 66622 36768 66628 36780
rect 65061 36731 65119 36737
rect 66088 36740 66628 36768
rect 61289 36703 61347 36709
rect 61289 36669 61301 36703
rect 61335 36669 61347 36703
rect 61289 36663 61347 36669
rect 61381 36703 61439 36709
rect 61381 36669 61393 36703
rect 61427 36669 61439 36703
rect 61381 36663 61439 36669
rect 61565 36703 61623 36709
rect 61565 36669 61577 36703
rect 61611 36700 61623 36703
rect 63037 36703 63095 36709
rect 63037 36700 63049 36703
rect 61611 36672 63049 36700
rect 61611 36669 61623 36672
rect 61565 36663 61623 36669
rect 63037 36669 63049 36672
rect 63083 36669 63095 36703
rect 63037 36663 63095 36669
rect 63497 36703 63555 36709
rect 63497 36669 63509 36703
rect 63543 36669 63555 36703
rect 63497 36663 63555 36669
rect 50525 36635 50583 36641
rect 50525 36632 50537 36635
rect 44339 36604 48728 36632
rect 49160 36604 50537 36632
rect 36688 36536 41460 36564
rect 36688 36524 36694 36536
rect 41506 36524 41512 36576
rect 41564 36564 41570 36576
rect 42518 36564 42524 36576
rect 41564 36536 42524 36564
rect 41564 36524 41570 36536
rect 42518 36524 42524 36536
rect 42576 36524 42582 36576
rect 48700 36564 48728 36604
rect 50525 36601 50537 36604
rect 50571 36632 50583 36635
rect 54846 36632 54852 36644
rect 50571 36604 54852 36632
rect 50571 36601 50583 36604
rect 50525 36595 50583 36601
rect 54846 36592 54852 36604
rect 54904 36592 54910 36644
rect 61396 36632 61424 36663
rect 62114 36632 62120 36644
rect 61396 36604 62120 36632
rect 62114 36592 62120 36604
rect 62172 36592 62178 36644
rect 50157 36567 50215 36573
rect 50157 36564 50169 36567
rect 48700 36536 50169 36564
rect 50157 36533 50169 36536
rect 50203 36533 50215 36567
rect 50157 36527 50215 36533
rect 51626 36524 51632 36576
rect 51684 36564 51690 36576
rect 55030 36564 55036 36576
rect 51684 36536 55036 36564
rect 51684 36524 51690 36536
rect 55030 36524 55036 36536
rect 55088 36524 55094 36576
rect 56594 36524 56600 36576
rect 56652 36564 56658 36576
rect 61749 36567 61807 36573
rect 61749 36564 61761 36567
rect 56652 36536 61761 36564
rect 56652 36524 56658 36536
rect 61749 36533 61761 36536
rect 61795 36533 61807 36567
rect 63512 36564 63540 36663
rect 63586 36660 63592 36712
rect 63644 36700 63650 36712
rect 63681 36703 63739 36709
rect 63681 36700 63693 36703
rect 63644 36672 63693 36700
rect 63644 36660 63650 36672
rect 63681 36669 63693 36672
rect 63727 36669 63739 36703
rect 63681 36663 63739 36669
rect 63770 36660 63776 36712
rect 63828 36700 63834 36712
rect 64049 36703 64107 36709
rect 64049 36700 64061 36703
rect 63828 36672 64061 36700
rect 63828 36660 63834 36672
rect 64049 36669 64061 36672
rect 64095 36669 64107 36703
rect 64049 36663 64107 36669
rect 64233 36703 64291 36709
rect 64233 36669 64245 36703
rect 64279 36700 64291 36703
rect 64506 36700 64512 36712
rect 64279 36672 64512 36700
rect 64279 36669 64291 36672
rect 64233 36663 64291 36669
rect 64506 36660 64512 36672
rect 64564 36660 64570 36712
rect 65426 36660 65432 36712
rect 65484 36700 65490 36712
rect 66088 36709 66116 36740
rect 66622 36728 66628 36740
rect 66680 36728 66686 36780
rect 71130 36728 71136 36780
rect 71188 36768 71194 36780
rect 71372 36771 71430 36777
rect 71372 36768 71384 36771
rect 71188 36740 71384 36768
rect 71188 36728 71194 36740
rect 71372 36737 71384 36740
rect 71418 36737 71430 36771
rect 71590 36768 71596 36780
rect 71551 36740 71596 36768
rect 71372 36731 71430 36737
rect 71590 36728 71596 36740
rect 71648 36728 71654 36780
rect 71958 36728 71964 36780
rect 72016 36768 72022 36780
rect 72016 36740 82032 36768
rect 72016 36728 72022 36740
rect 65521 36703 65579 36709
rect 65521 36700 65533 36703
rect 65484 36672 65533 36700
rect 65484 36660 65490 36672
rect 65521 36669 65533 36672
rect 65567 36669 65579 36703
rect 65521 36663 65579 36669
rect 65705 36703 65763 36709
rect 65705 36669 65717 36703
rect 65751 36669 65763 36703
rect 65705 36663 65763 36669
rect 66073 36703 66131 36709
rect 66073 36669 66085 36703
rect 66119 36669 66131 36703
rect 66073 36663 66131 36669
rect 65720 36632 65748 36663
rect 66162 36660 66168 36712
rect 66220 36700 66226 36712
rect 66438 36700 66444 36712
rect 66220 36672 66265 36700
rect 66399 36672 66444 36700
rect 66220 36660 66226 36672
rect 66438 36660 66444 36672
rect 66496 36660 66502 36712
rect 68646 36700 68652 36712
rect 68607 36672 68652 36700
rect 68646 36660 68652 36672
rect 68704 36700 68710 36712
rect 68925 36703 68983 36709
rect 68925 36700 68937 36703
rect 68704 36672 68937 36700
rect 68704 36660 68710 36672
rect 68925 36669 68937 36672
rect 68971 36669 68983 36703
rect 69750 36700 69756 36712
rect 69711 36672 69756 36700
rect 68925 36663 68983 36669
rect 69750 36660 69756 36672
rect 69808 36660 69814 36712
rect 69934 36700 69940 36712
rect 69895 36672 69940 36700
rect 69934 36660 69940 36672
rect 69992 36660 69998 36712
rect 71608 36700 71636 36728
rect 72053 36703 72111 36709
rect 72053 36700 72065 36703
rect 71608 36672 72065 36700
rect 72053 36669 72065 36672
rect 72099 36700 72111 36703
rect 72602 36700 72608 36712
rect 72099 36672 72608 36700
rect 72099 36669 72111 36672
rect 72053 36663 72111 36669
rect 72602 36660 72608 36672
rect 72660 36660 72666 36712
rect 72786 36700 72792 36712
rect 72747 36672 72792 36700
rect 72786 36660 72792 36672
rect 72844 36660 72850 36712
rect 76834 36660 76840 36712
rect 76892 36700 76898 36712
rect 76929 36703 76987 36709
rect 76929 36700 76941 36703
rect 76892 36672 76941 36700
rect 76892 36660 76898 36672
rect 76929 36669 76941 36672
rect 76975 36700 76987 36703
rect 77297 36703 77355 36709
rect 77297 36700 77309 36703
rect 76975 36672 77309 36700
rect 76975 36669 76987 36672
rect 76929 36663 76987 36669
rect 77297 36669 77309 36672
rect 77343 36669 77355 36703
rect 77297 36663 77355 36669
rect 77849 36703 77907 36709
rect 77849 36669 77861 36703
rect 77895 36669 77907 36703
rect 78214 36700 78220 36712
rect 78175 36672 78220 36700
rect 77849 36663 77907 36669
rect 66456 36632 66484 36660
rect 65720 36604 66484 36632
rect 68741 36635 68799 36641
rect 68741 36601 68753 36635
rect 68787 36632 68799 36635
rect 69845 36635 69903 36641
rect 68787 36604 69796 36632
rect 68787 36601 68799 36604
rect 68741 36595 68799 36601
rect 64417 36567 64475 36573
rect 64417 36564 64429 36567
rect 63512 36536 64429 36564
rect 61749 36527 61807 36533
rect 64417 36533 64429 36536
rect 64463 36564 64475 36567
rect 64598 36564 64604 36576
rect 64463 36536 64604 36564
rect 64463 36533 64475 36536
rect 64417 36527 64475 36533
rect 64598 36524 64604 36536
rect 64656 36524 64662 36576
rect 69768 36564 69796 36604
rect 69845 36601 69857 36635
rect 69891 36632 69903 36635
rect 70302 36632 70308 36644
rect 69891 36604 70308 36632
rect 69891 36601 69903 36604
rect 69845 36595 69903 36601
rect 70302 36592 70308 36604
rect 70360 36592 70366 36644
rect 70397 36635 70455 36641
rect 70397 36601 70409 36635
rect 70443 36632 70455 36635
rect 70578 36632 70584 36644
rect 70443 36604 70584 36632
rect 70443 36601 70455 36604
rect 70397 36595 70455 36601
rect 70578 36592 70584 36604
rect 70636 36592 70642 36644
rect 71225 36635 71283 36641
rect 71225 36632 71237 36635
rect 70780 36604 71237 36632
rect 70118 36564 70124 36576
rect 69768 36536 70124 36564
rect 70118 36524 70124 36536
rect 70176 36564 70182 36576
rect 70780 36564 70808 36604
rect 71225 36601 71237 36604
rect 71271 36601 71283 36635
rect 71225 36595 71283 36601
rect 71961 36635 72019 36641
rect 71961 36601 71973 36635
rect 72007 36632 72019 36635
rect 74442 36632 74448 36644
rect 72007 36604 74448 36632
rect 72007 36601 72019 36604
rect 71961 36595 72019 36601
rect 74442 36592 74448 36604
rect 74500 36592 74506 36644
rect 77864 36632 77892 36663
rect 78214 36660 78220 36672
rect 78272 36660 78278 36712
rect 77220 36604 77892 36632
rect 82004 36632 82032 36740
rect 83550 36728 83556 36780
rect 83608 36768 83614 36780
rect 84289 36771 84347 36777
rect 84289 36768 84301 36771
rect 83608 36740 84301 36768
rect 83608 36728 83614 36740
rect 84289 36737 84301 36740
rect 84335 36737 84347 36771
rect 85942 36768 85948 36780
rect 85903 36740 85948 36768
rect 84289 36731 84347 36737
rect 85942 36728 85948 36740
rect 86000 36728 86006 36780
rect 86972 36768 87000 36864
rect 87141 36771 87199 36777
rect 87141 36768 87153 36771
rect 86972 36740 87153 36768
rect 87141 36737 87153 36740
rect 87187 36737 87199 36771
rect 87414 36768 87420 36780
rect 87375 36740 87420 36768
rect 87141 36731 87199 36737
rect 87414 36728 87420 36740
rect 87472 36728 87478 36780
rect 82170 36700 82176 36712
rect 82131 36672 82176 36700
rect 82170 36660 82176 36672
rect 82228 36660 82234 36712
rect 82265 36703 82323 36709
rect 82265 36669 82277 36703
rect 82311 36700 82323 36703
rect 83829 36703 83887 36709
rect 83829 36700 83841 36703
rect 82311 36672 83841 36700
rect 82311 36669 82323 36672
rect 82265 36663 82323 36669
rect 83829 36669 83841 36672
rect 83875 36669 83887 36703
rect 83829 36663 83887 36669
rect 83844 36632 83872 36663
rect 83918 36660 83924 36712
rect 83976 36700 83982 36712
rect 84194 36700 84200 36712
rect 83976 36672 84021 36700
rect 84155 36672 84200 36700
rect 83976 36660 83982 36672
rect 84194 36660 84200 36672
rect 84252 36660 84258 36712
rect 85577 36703 85635 36709
rect 85577 36669 85589 36703
rect 85623 36700 85635 36703
rect 86037 36703 86095 36709
rect 86037 36700 86049 36703
rect 85623 36672 86049 36700
rect 85623 36669 85635 36672
rect 85577 36663 85635 36669
rect 86037 36669 86049 36672
rect 86083 36700 86095 36703
rect 86954 36700 86960 36712
rect 86083 36672 86960 36700
rect 86083 36669 86095 36672
rect 86037 36663 86095 36669
rect 85393 36635 85451 36641
rect 85393 36632 85405 36635
rect 82004 36604 83780 36632
rect 83844 36604 85405 36632
rect 77220 36576 77248 36604
rect 77202 36564 77208 36576
rect 70176 36536 70808 36564
rect 77163 36536 77208 36564
rect 70176 36524 70182 36536
rect 77202 36524 77208 36536
rect 77260 36524 77266 36576
rect 77389 36567 77447 36573
rect 77389 36533 77401 36567
rect 77435 36564 77447 36567
rect 77846 36564 77852 36576
rect 77435 36536 77852 36564
rect 77435 36533 77447 36536
rect 77389 36527 77447 36533
rect 77846 36524 77852 36536
rect 77904 36524 77910 36576
rect 82998 36564 83004 36576
rect 82959 36536 83004 36564
rect 82998 36524 83004 36536
rect 83056 36524 83062 36576
rect 83752 36564 83780 36604
rect 85393 36601 85405 36604
rect 85439 36601 85451 36635
rect 85393 36595 85451 36601
rect 85592 36564 85620 36663
rect 86954 36660 86960 36672
rect 87012 36660 87018 36712
rect 86770 36592 86776 36644
rect 86828 36632 86834 36644
rect 86828 36604 87092 36632
rect 86828 36592 86834 36604
rect 83752 36536 85620 36564
rect 87064 36564 87092 36604
rect 88521 36567 88579 36573
rect 88521 36564 88533 36567
rect 87064 36536 88533 36564
rect 88521 36533 88533 36536
rect 88567 36533 88579 36567
rect 88521 36527 88579 36533
rect 1104 36474 111136 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 81046 36474
rect 81098 36422 81110 36474
rect 81162 36422 81174 36474
rect 81226 36422 81238 36474
rect 81290 36422 111136 36474
rect 1104 36400 111136 36422
rect 4982 36360 4988 36372
rect 4943 36332 4988 36360
rect 4982 36320 4988 36332
rect 5040 36320 5046 36372
rect 15470 36360 15476 36372
rect 15431 36332 15476 36360
rect 15470 36320 15476 36332
rect 15528 36320 15534 36372
rect 17218 36360 17224 36372
rect 17179 36332 17224 36360
rect 17218 36320 17224 36332
rect 17276 36320 17282 36372
rect 25409 36363 25467 36369
rect 25409 36329 25421 36363
rect 25455 36329 25467 36363
rect 26602 36360 26608 36372
rect 26563 36332 26608 36360
rect 25409 36323 25467 36329
rect 9858 36252 9864 36304
rect 9916 36292 9922 36304
rect 10594 36292 10600 36304
rect 9916 36264 10600 36292
rect 9916 36252 9922 36264
rect 10594 36252 10600 36264
rect 10652 36252 10658 36304
rect 11333 36295 11391 36301
rect 11333 36261 11345 36295
rect 11379 36292 11391 36295
rect 16758 36292 16764 36304
rect 11379 36264 16764 36292
rect 11379 36261 11391 36264
rect 11333 36255 11391 36261
rect 5169 36227 5227 36233
rect 5169 36193 5181 36227
rect 5215 36193 5227 36227
rect 5350 36224 5356 36236
rect 5311 36196 5356 36224
rect 5169 36187 5227 36193
rect 5184 36156 5212 36187
rect 5350 36184 5356 36196
rect 5408 36184 5414 36236
rect 6457 36227 6515 36233
rect 6457 36193 6469 36227
rect 6503 36224 6515 36227
rect 8202 36224 8208 36236
rect 6503 36196 8208 36224
rect 6503 36193 6515 36196
rect 6457 36187 6515 36193
rect 8202 36184 8208 36196
rect 8260 36184 8266 36236
rect 10781 36227 10839 36233
rect 10781 36193 10793 36227
rect 10827 36224 10839 36227
rect 11348 36224 11376 36255
rect 16758 36252 16764 36264
rect 16816 36252 16822 36304
rect 10827 36196 11376 36224
rect 15289 36227 15347 36233
rect 10827 36193 10839 36196
rect 10781 36187 10839 36193
rect 15289 36193 15301 36227
rect 15335 36193 15347 36227
rect 16482 36224 16488 36236
rect 16443 36196 16488 36224
rect 15289 36187 15347 36193
rect 5258 36156 5264 36168
rect 5171 36128 5264 36156
rect 5258 36116 5264 36128
rect 5316 36156 5322 36168
rect 11054 36156 11060 36168
rect 5316 36128 6684 36156
rect 11015 36128 11060 36156
rect 5316 36116 5322 36128
rect 6656 36097 6684 36128
rect 11054 36116 11060 36128
rect 11112 36116 11118 36168
rect 15304 36156 15332 36187
rect 16482 36184 16488 36196
rect 16540 36184 16546 36236
rect 16577 36227 16635 36233
rect 16577 36193 16589 36227
rect 16623 36224 16635 36227
rect 17236 36224 17264 36320
rect 25424 36292 25452 36323
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 33686 36360 33692 36372
rect 27080 36332 33692 36360
rect 25498 36292 25504 36304
rect 25411 36264 25504 36292
rect 25498 36252 25504 36264
rect 25556 36292 25562 36304
rect 27080 36292 27108 36332
rect 33686 36320 33692 36332
rect 33744 36320 33750 36372
rect 35434 36320 35440 36372
rect 35492 36360 35498 36372
rect 35805 36363 35863 36369
rect 35805 36360 35817 36363
rect 35492 36332 35817 36360
rect 35492 36320 35498 36332
rect 35805 36329 35817 36332
rect 35851 36329 35863 36363
rect 35805 36323 35863 36329
rect 36538 36320 36544 36372
rect 36596 36360 36602 36372
rect 41322 36360 41328 36372
rect 36596 36332 41328 36360
rect 36596 36320 36602 36332
rect 41322 36320 41328 36332
rect 41380 36320 41386 36372
rect 41690 36360 41696 36372
rect 41651 36332 41696 36360
rect 41690 36320 41696 36332
rect 41748 36320 41754 36372
rect 41782 36320 41788 36372
rect 41840 36360 41846 36372
rect 42245 36363 42303 36369
rect 42245 36360 42257 36363
rect 41840 36332 42257 36360
rect 41840 36320 41846 36332
rect 42245 36329 42257 36332
rect 42291 36360 42303 36363
rect 44542 36360 44548 36372
rect 42291 36332 43484 36360
rect 44503 36332 44548 36360
rect 42291 36329 42303 36332
rect 42245 36323 42303 36329
rect 32214 36292 32220 36304
rect 25556 36264 27108 36292
rect 27172 36264 32220 36292
rect 25556 36252 25562 36264
rect 24854 36224 24860 36236
rect 16623 36196 17264 36224
rect 17328 36196 24860 36224
rect 16623 36193 16635 36196
rect 16577 36187 16635 36193
rect 16393 36159 16451 36165
rect 16393 36156 16405 36159
rect 15304 36128 16405 36156
rect 16393 36125 16405 36128
rect 16439 36125 16451 36159
rect 16393 36119 16451 36125
rect 16758 36116 16764 36168
rect 16816 36156 16822 36168
rect 17328 36156 17356 36196
rect 24854 36184 24860 36196
rect 24912 36184 24918 36236
rect 24946 36184 24952 36236
rect 25004 36224 25010 36236
rect 25133 36227 25191 36233
rect 25133 36224 25145 36227
rect 25004 36196 25145 36224
rect 25004 36184 25010 36196
rect 25133 36193 25145 36196
rect 25179 36224 25191 36227
rect 25225 36227 25283 36233
rect 25225 36224 25237 36227
rect 25179 36196 25237 36224
rect 25179 36193 25191 36196
rect 25133 36187 25191 36193
rect 25225 36193 25237 36196
rect 25271 36193 25283 36227
rect 26142 36224 26148 36236
rect 26055 36196 26148 36224
rect 25225 36187 25283 36193
rect 26142 36184 26148 36196
rect 26200 36224 26206 36236
rect 27172 36233 27200 36264
rect 32214 36252 32220 36264
rect 32272 36252 32278 36304
rect 33781 36295 33839 36301
rect 33781 36261 33793 36295
rect 33827 36292 33839 36295
rect 36630 36292 36636 36304
rect 33827 36264 36636 36292
rect 33827 36261 33839 36264
rect 33781 36255 33839 36261
rect 36630 36252 36636 36264
rect 36688 36252 36694 36304
rect 43456 36292 43484 36332
rect 44542 36320 44548 36332
rect 44600 36320 44606 36372
rect 45097 36363 45155 36369
rect 45097 36329 45109 36363
rect 45143 36360 45155 36363
rect 49970 36360 49976 36372
rect 45143 36332 49976 36360
rect 45143 36329 45155 36332
rect 45097 36323 45155 36329
rect 39500 36264 41184 36292
rect 43456 36264 44128 36292
rect 27157 36227 27215 36233
rect 27157 36224 27169 36227
rect 26200 36196 27169 36224
rect 26200 36184 26206 36196
rect 27157 36193 27169 36196
rect 27203 36193 27215 36227
rect 27157 36187 27215 36193
rect 27525 36227 27583 36233
rect 27525 36193 27537 36227
rect 27571 36193 27583 36227
rect 27525 36187 27583 36193
rect 30101 36227 30159 36233
rect 30101 36193 30113 36227
rect 30147 36224 30159 36227
rect 31478 36224 31484 36236
rect 30147 36196 31484 36224
rect 30147 36193 30159 36196
rect 30101 36187 30159 36193
rect 20990 36156 20996 36168
rect 16816 36128 17356 36156
rect 20951 36128 20996 36156
rect 16816 36116 16822 36128
rect 20990 36116 20996 36128
rect 21048 36116 21054 36168
rect 21266 36156 21272 36168
rect 21227 36128 21272 36156
rect 21266 36116 21272 36128
rect 21324 36116 21330 36168
rect 27062 36156 27068 36168
rect 27023 36128 27068 36156
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 27430 36156 27436 36168
rect 27391 36128 27436 36156
rect 27430 36116 27436 36128
rect 27488 36116 27494 36168
rect 27540 36100 27568 36187
rect 31478 36184 31484 36196
rect 31536 36184 31542 36236
rect 32398 36224 32404 36236
rect 32359 36196 32404 36224
rect 32398 36184 32404 36196
rect 32456 36184 32462 36236
rect 34146 36224 34152 36236
rect 34059 36196 34152 36224
rect 34146 36184 34152 36196
rect 34204 36224 34210 36236
rect 34333 36227 34391 36233
rect 34333 36224 34345 36227
rect 34204 36196 34345 36224
rect 34204 36184 34210 36196
rect 34333 36193 34345 36196
rect 34379 36224 34391 36227
rect 34793 36227 34851 36233
rect 34793 36224 34805 36227
rect 34379 36196 34805 36224
rect 34379 36193 34391 36196
rect 34333 36187 34391 36193
rect 34793 36193 34805 36196
rect 34839 36224 34851 36227
rect 35342 36224 35348 36236
rect 34839 36196 35348 36224
rect 34839 36193 34851 36196
rect 34793 36187 34851 36193
rect 35342 36184 35348 36196
rect 35400 36184 35406 36236
rect 35529 36227 35587 36233
rect 35529 36193 35541 36227
rect 35575 36224 35587 36227
rect 35986 36224 35992 36236
rect 35575 36196 35992 36224
rect 35575 36193 35587 36196
rect 35529 36187 35587 36193
rect 35986 36184 35992 36196
rect 36044 36224 36050 36236
rect 36446 36224 36452 36236
rect 36044 36196 36452 36224
rect 36044 36184 36050 36196
rect 36446 36184 36452 36196
rect 36504 36184 36510 36236
rect 39114 36184 39120 36236
rect 39172 36224 39178 36236
rect 39500 36233 39528 36264
rect 39485 36227 39543 36233
rect 39485 36224 39497 36227
rect 39172 36196 39497 36224
rect 39172 36184 39178 36196
rect 39485 36193 39497 36196
rect 39531 36193 39543 36227
rect 40678 36224 40684 36236
rect 40639 36196 40684 36224
rect 39485 36187 39543 36193
rect 40678 36184 40684 36196
rect 40736 36184 40742 36236
rect 41156 36233 41184 36264
rect 41141 36227 41199 36233
rect 41141 36193 41153 36227
rect 41187 36193 41199 36227
rect 41141 36187 41199 36193
rect 41233 36227 41291 36233
rect 41233 36193 41245 36227
rect 41279 36224 41291 36227
rect 41782 36224 41788 36236
rect 41279 36196 41788 36224
rect 41279 36193 41291 36196
rect 41233 36187 41291 36193
rect 41782 36184 41788 36196
rect 41840 36184 41846 36236
rect 42061 36227 42119 36233
rect 42061 36193 42073 36227
rect 42107 36224 42119 36227
rect 42242 36224 42248 36236
rect 42107 36196 42248 36224
rect 42107 36193 42119 36196
rect 42061 36187 42119 36193
rect 42242 36184 42248 36196
rect 42300 36224 42306 36236
rect 43530 36224 43536 36236
rect 42300 36196 43536 36224
rect 42300 36184 42306 36196
rect 43530 36184 43536 36196
rect 43588 36184 43594 36236
rect 43625 36227 43683 36233
rect 43625 36193 43637 36227
rect 43671 36224 43683 36227
rect 43714 36224 43720 36236
rect 43671 36196 43720 36224
rect 43671 36193 43683 36196
rect 43625 36187 43683 36193
rect 30282 36156 30288 36168
rect 29932 36128 30288 36156
rect 6641 36091 6699 36097
rect 6641 36057 6653 36091
rect 6687 36057 6699 36091
rect 22741 36091 22799 36097
rect 22741 36088 22753 36091
rect 6641 36051 6699 36057
rect 22112 36060 22753 36088
rect 16393 36023 16451 36029
rect 16393 35989 16405 36023
rect 16439 36020 16451 36023
rect 16482 36020 16488 36032
rect 16439 35992 16488 36020
rect 16439 35989 16451 35992
rect 16393 35983 16451 35989
rect 16482 35980 16488 35992
rect 16540 35980 16546 36032
rect 16758 36020 16764 36032
rect 16719 35992 16764 36020
rect 16758 35980 16764 35992
rect 16816 35980 16822 36032
rect 20990 35980 20996 36032
rect 21048 36020 21054 36032
rect 22002 36020 22008 36032
rect 21048 35992 22008 36020
rect 21048 35980 21054 35992
rect 22002 35980 22008 35992
rect 22060 36020 22066 36032
rect 22112 36020 22140 36060
rect 22741 36057 22753 36060
rect 22787 36057 22799 36091
rect 22741 36051 22799 36057
rect 25314 36048 25320 36100
rect 25372 36088 25378 36100
rect 25866 36088 25872 36100
rect 25372 36060 25872 36088
rect 25372 36048 25378 36060
rect 25866 36048 25872 36060
rect 25924 36048 25930 36100
rect 27522 36088 27528 36100
rect 26252 36060 27528 36088
rect 26252 36032 26280 36060
rect 27522 36048 27528 36060
rect 27580 36048 27586 36100
rect 29178 36048 29184 36100
rect 29236 36088 29242 36100
rect 29932 36097 29960 36128
rect 30282 36116 30288 36128
rect 30340 36156 30346 36168
rect 31941 36159 31999 36165
rect 31941 36156 31953 36159
rect 30340 36128 31953 36156
rect 30340 36116 30346 36128
rect 31941 36125 31953 36128
rect 31987 36156 31999 36159
rect 32125 36159 32183 36165
rect 32125 36156 32137 36159
rect 31987 36128 32137 36156
rect 31987 36125 31999 36128
rect 31941 36119 31999 36125
rect 32125 36125 32137 36128
rect 32171 36125 32183 36159
rect 32125 36119 32183 36125
rect 34609 36159 34667 36165
rect 34609 36125 34621 36159
rect 34655 36125 34667 36159
rect 34609 36119 34667 36125
rect 29917 36091 29975 36097
rect 29917 36088 29929 36091
rect 29236 36060 29929 36088
rect 29236 36048 29242 36060
rect 29917 36057 29929 36060
rect 29963 36057 29975 36091
rect 29917 36051 29975 36057
rect 34624 36032 34652 36119
rect 35894 36116 35900 36168
rect 35952 36156 35958 36168
rect 37550 36156 37556 36168
rect 35952 36128 37556 36156
rect 35952 36116 35958 36128
rect 37550 36116 37556 36128
rect 37608 36116 37614 36168
rect 40218 36116 40224 36168
rect 40276 36156 40282 36168
rect 40497 36159 40555 36165
rect 40497 36156 40509 36159
rect 40276 36128 40509 36156
rect 40276 36116 40282 36128
rect 40497 36125 40509 36128
rect 40543 36125 40555 36159
rect 40497 36119 40555 36125
rect 43165 36159 43223 36165
rect 43165 36125 43177 36159
rect 43211 36156 43223 36159
rect 43640 36156 43668 36187
rect 43714 36184 43720 36196
rect 43772 36184 43778 36236
rect 43990 36224 43996 36236
rect 43951 36196 43996 36224
rect 43990 36184 43996 36196
rect 44048 36184 44054 36236
rect 44100 36233 44128 36264
rect 44085 36227 44143 36233
rect 44085 36193 44097 36227
rect 44131 36224 44143 36227
rect 45112 36224 45140 36323
rect 49970 36320 49976 36332
rect 50028 36320 50034 36372
rect 51629 36363 51687 36369
rect 51629 36360 51641 36363
rect 50080 36332 51641 36360
rect 46584 36264 46796 36292
rect 46014 36224 46020 36236
rect 44131 36196 45140 36224
rect 45975 36196 46020 36224
rect 44131 36193 44143 36196
rect 44085 36187 44143 36193
rect 46014 36184 46020 36196
rect 46072 36184 46078 36236
rect 44910 36156 44916 36168
rect 43211 36128 43668 36156
rect 44823 36128 44916 36156
rect 43211 36125 43223 36128
rect 43165 36119 43223 36125
rect 44910 36116 44916 36128
rect 44968 36156 44974 36168
rect 45557 36159 45615 36165
rect 45557 36156 45569 36159
rect 44968 36128 45569 36156
rect 44968 36116 44974 36128
rect 45557 36125 45569 36128
rect 45603 36125 45615 36159
rect 45830 36156 45836 36168
rect 45791 36128 45836 36156
rect 45557 36119 45615 36125
rect 45830 36116 45836 36128
rect 45888 36156 45894 36168
rect 46584 36156 46612 36264
rect 46661 36227 46719 36233
rect 46661 36193 46673 36227
rect 46707 36193 46719 36227
rect 46768 36224 46796 36264
rect 46934 36252 46940 36304
rect 46992 36292 46998 36304
rect 46992 36264 50016 36292
rect 46992 36252 46998 36264
rect 47029 36227 47087 36233
rect 47029 36224 47041 36227
rect 46768 36196 47041 36224
rect 46661 36187 46719 36193
rect 47029 36193 47041 36196
rect 47075 36193 47087 36227
rect 47029 36187 47087 36193
rect 47213 36227 47271 36233
rect 47213 36193 47225 36227
rect 47259 36224 47271 36227
rect 47670 36224 47676 36236
rect 47259 36196 47676 36224
rect 47259 36193 47271 36196
rect 47213 36187 47271 36193
rect 45888 36128 46612 36156
rect 45888 36116 45894 36128
rect 35250 36048 35256 36100
rect 35308 36088 35314 36100
rect 45649 36091 45707 36097
rect 45649 36088 45661 36091
rect 35308 36060 45661 36088
rect 35308 36048 35314 36060
rect 45649 36057 45661 36060
rect 45695 36088 45707 36091
rect 46676 36088 46704 36187
rect 46753 36159 46811 36165
rect 46753 36125 46765 36159
rect 46799 36156 46811 36159
rect 46934 36156 46940 36168
rect 46799 36128 46940 36156
rect 46799 36125 46811 36128
rect 46753 36119 46811 36125
rect 46934 36116 46940 36128
rect 46992 36116 46998 36168
rect 47044 36156 47072 36187
rect 47670 36184 47676 36196
rect 47728 36184 47734 36236
rect 49050 36184 49056 36236
rect 49108 36224 49114 36236
rect 49513 36227 49571 36233
rect 49513 36224 49525 36227
rect 49108 36196 49525 36224
rect 49108 36184 49114 36196
rect 49513 36193 49525 36196
rect 49559 36224 49571 36227
rect 49881 36227 49939 36233
rect 49881 36224 49893 36227
rect 49559 36196 49893 36224
rect 49559 36193 49571 36196
rect 49513 36187 49571 36193
rect 49881 36193 49893 36196
rect 49927 36193 49939 36227
rect 49881 36187 49939 36193
rect 49786 36156 49792 36168
rect 47044 36128 49792 36156
rect 49786 36116 49792 36128
rect 49844 36116 49850 36168
rect 49988 36088 50016 36264
rect 50080 36233 50108 36332
rect 51629 36329 51641 36332
rect 51675 36360 51687 36363
rect 54478 36360 54484 36372
rect 51675 36332 54484 36360
rect 51675 36329 51687 36332
rect 51629 36323 51687 36329
rect 54478 36320 54484 36332
rect 54536 36320 54542 36372
rect 61102 36320 61108 36372
rect 61160 36360 61166 36372
rect 68646 36360 68652 36372
rect 61160 36332 68652 36360
rect 61160 36320 61166 36332
rect 68646 36320 68652 36332
rect 68704 36320 68710 36372
rect 72786 36320 72792 36372
rect 72844 36360 72850 36372
rect 73617 36363 73675 36369
rect 73617 36360 73629 36363
rect 72844 36332 73629 36360
rect 72844 36320 72850 36332
rect 73617 36329 73629 36332
rect 73663 36329 73675 36363
rect 73617 36323 73675 36329
rect 77205 36363 77263 36369
rect 77205 36329 77217 36363
rect 77251 36360 77263 36363
rect 77938 36360 77944 36372
rect 77251 36332 77944 36360
rect 77251 36329 77263 36332
rect 77205 36323 77263 36329
rect 51166 36292 51172 36304
rect 50632 36264 51172 36292
rect 50065 36227 50123 36233
rect 50065 36193 50077 36227
rect 50111 36193 50123 36227
rect 50065 36187 50123 36193
rect 50154 36184 50160 36236
rect 50212 36224 50218 36236
rect 50632 36233 50660 36264
rect 51166 36252 51172 36264
rect 51224 36252 51230 36304
rect 51534 36252 51540 36304
rect 51592 36292 51598 36304
rect 52089 36295 52147 36301
rect 52089 36292 52101 36295
rect 51592 36264 52101 36292
rect 51592 36252 51598 36264
rect 52089 36261 52101 36264
rect 52135 36261 52147 36295
rect 52454 36292 52460 36304
rect 52089 36255 52147 36261
rect 52288 36264 52460 36292
rect 50525 36227 50583 36233
rect 50525 36224 50537 36227
rect 50212 36196 50537 36224
rect 50212 36184 50218 36196
rect 50525 36193 50537 36196
rect 50571 36193 50583 36227
rect 50525 36187 50583 36193
rect 50617 36227 50675 36233
rect 50617 36193 50629 36227
rect 50663 36193 50675 36227
rect 50617 36187 50675 36193
rect 50706 36184 50712 36236
rect 50764 36224 50770 36236
rect 52288 36233 52316 36264
rect 52454 36252 52460 36264
rect 52512 36252 52518 36304
rect 58618 36292 58624 36304
rect 57348 36264 58624 36292
rect 51813 36227 51871 36233
rect 51813 36224 51825 36227
rect 50764 36196 51825 36224
rect 50764 36184 50770 36196
rect 51813 36193 51825 36196
rect 51859 36224 51871 36227
rect 51905 36227 51963 36233
rect 51905 36224 51917 36227
rect 51859 36196 51917 36224
rect 51859 36193 51871 36196
rect 51813 36187 51871 36193
rect 51905 36193 51917 36196
rect 51951 36193 51963 36227
rect 51905 36187 51963 36193
rect 52236 36227 52316 36233
rect 52236 36193 52248 36227
rect 52282 36196 52316 36227
rect 54294 36224 54300 36236
rect 52380 36196 54300 36224
rect 52282 36193 52294 36196
rect 52236 36187 52294 36193
rect 51166 36116 51172 36168
rect 51224 36156 51230 36168
rect 51353 36159 51411 36165
rect 51353 36156 51365 36159
rect 51224 36128 51365 36156
rect 51224 36116 51230 36128
rect 51353 36125 51365 36128
rect 51399 36125 51411 36159
rect 52380 36156 52408 36196
rect 54294 36184 54300 36196
rect 54352 36184 54358 36236
rect 57348 36233 57376 36264
rect 58618 36252 58624 36264
rect 58676 36252 58682 36304
rect 64782 36252 64788 36304
rect 64840 36292 64846 36304
rect 69937 36295 69995 36301
rect 64840 36264 66116 36292
rect 64840 36252 64846 36264
rect 57333 36227 57391 36233
rect 57333 36193 57345 36227
rect 57379 36193 57391 36227
rect 57333 36187 57391 36193
rect 57517 36227 57575 36233
rect 57517 36193 57529 36227
rect 57563 36193 57575 36227
rect 57885 36227 57943 36233
rect 57885 36224 57897 36227
rect 57517 36187 57575 36193
rect 57624 36196 57897 36224
rect 51353 36119 51411 36125
rect 51460 36128 52408 36156
rect 52457 36159 52515 36165
rect 50985 36091 51043 36097
rect 50985 36088 50997 36091
rect 45695 36060 49832 36088
rect 49988 36060 50997 36088
rect 45695 36057 45707 36060
rect 45649 36051 45707 36057
rect 22060 35992 22140 36020
rect 22557 36023 22615 36029
rect 22060 35980 22066 35992
rect 22557 35989 22569 36023
rect 22603 36020 22615 36023
rect 23658 36020 23664 36032
rect 22603 35992 23664 36020
rect 22603 35989 22615 35992
rect 22557 35983 22615 35989
rect 23658 35980 23664 35992
rect 23716 35980 23722 36032
rect 26234 36020 26240 36032
rect 26195 35992 26240 36020
rect 26234 35980 26240 35992
rect 26292 35980 26298 36032
rect 27154 35980 27160 36032
rect 27212 36020 27218 36032
rect 27430 36020 27436 36032
rect 27212 35992 27436 36020
rect 27212 35980 27218 35992
rect 27430 35980 27436 35992
rect 27488 35980 27494 36032
rect 34517 36023 34575 36029
rect 34517 35989 34529 36023
rect 34563 36020 34575 36023
rect 34606 36020 34612 36032
rect 34563 35992 34612 36020
rect 34563 35989 34575 35992
rect 34517 35983 34575 35989
rect 34606 35980 34612 35992
rect 34664 35980 34670 36032
rect 38746 35980 38752 36032
rect 38804 36020 38810 36032
rect 39574 36020 39580 36032
rect 38804 35992 39580 36020
rect 38804 35980 38810 35992
rect 39574 35980 39580 35992
rect 39632 35980 39638 36032
rect 39853 36023 39911 36029
rect 39853 35989 39865 36023
rect 39899 36020 39911 36023
rect 39942 36020 39948 36032
rect 39899 35992 39948 36020
rect 39899 35989 39911 35992
rect 39853 35983 39911 35989
rect 39942 35980 39948 35992
rect 40000 35980 40006 36032
rect 40218 35980 40224 36032
rect 40276 36020 40282 36032
rect 40313 36023 40371 36029
rect 40313 36020 40325 36023
rect 40276 35992 40325 36020
rect 40276 35980 40282 35992
rect 40313 35989 40325 35992
rect 40359 35989 40371 36023
rect 40313 35983 40371 35989
rect 45557 36023 45615 36029
rect 45557 35989 45569 36023
rect 45603 36020 45615 36023
rect 49142 36020 49148 36032
rect 45603 35992 49148 36020
rect 45603 35989 45615 35992
rect 45557 35983 45615 35989
rect 49142 35980 49148 35992
rect 49200 35980 49206 36032
rect 49510 35980 49516 36032
rect 49568 36020 49574 36032
rect 49697 36023 49755 36029
rect 49697 36020 49709 36023
rect 49568 35992 49709 36020
rect 49568 35980 49574 35992
rect 49697 35989 49709 35992
rect 49743 35989 49755 36023
rect 49804 36020 49832 36060
rect 50985 36057 50997 36060
rect 51031 36057 51043 36091
rect 50985 36051 51043 36057
rect 51258 36048 51264 36100
rect 51316 36088 51322 36100
rect 51460 36088 51488 36128
rect 52457 36125 52469 36159
rect 52503 36156 52515 36159
rect 56594 36156 56600 36168
rect 52503 36128 56600 36156
rect 52503 36125 52515 36128
rect 52457 36119 52515 36125
rect 56594 36116 56600 36128
rect 56652 36116 56658 36168
rect 56870 36156 56876 36168
rect 56831 36128 56876 36156
rect 56870 36116 56876 36128
rect 56928 36116 56934 36168
rect 51316 36060 51488 36088
rect 51813 36091 51871 36097
rect 51316 36048 51322 36060
rect 51813 36057 51825 36091
rect 51859 36088 51871 36091
rect 52365 36091 52423 36097
rect 52365 36088 52377 36091
rect 51859 36060 52377 36088
rect 51859 36057 51871 36060
rect 51813 36051 51871 36057
rect 52365 36057 52377 36060
rect 52411 36057 52423 36091
rect 54846 36088 54852 36100
rect 52365 36051 52423 36057
rect 52656 36060 54852 36088
rect 52656 36020 52684 36060
rect 54846 36048 54852 36060
rect 54904 36088 54910 36100
rect 55950 36088 55956 36100
rect 54904 36060 55956 36088
rect 54904 36048 54910 36060
rect 55950 36048 55956 36060
rect 56008 36088 56014 36100
rect 56505 36091 56563 36097
rect 56505 36088 56517 36091
rect 56008 36060 56517 36088
rect 56008 36048 56014 36060
rect 56505 36057 56517 36060
rect 56551 36088 56563 36091
rect 57532 36088 57560 36187
rect 56551 36060 57560 36088
rect 56551 36057 56563 36060
rect 56505 36051 56563 36057
rect 49804 35992 52684 36020
rect 52733 36023 52791 36029
rect 49697 35983 49755 35989
rect 52733 35989 52745 36023
rect 52779 36020 52791 36023
rect 53282 36020 53288 36032
rect 52779 35992 53288 36020
rect 52779 35989 52791 35992
rect 52733 35983 52791 35989
rect 53282 35980 53288 35992
rect 53340 35980 53346 36032
rect 55030 35980 55036 36032
rect 55088 36020 55094 36032
rect 56689 36023 56747 36029
rect 56689 36020 56701 36023
rect 55088 35992 56701 36020
rect 55088 35980 55094 35992
rect 56689 35989 56701 35992
rect 56735 36020 56747 36023
rect 57624 36020 57652 36196
rect 57885 36193 57897 36196
rect 57931 36193 57943 36227
rect 57885 36187 57943 36193
rect 58069 36227 58127 36233
rect 58069 36193 58081 36227
rect 58115 36224 58127 36227
rect 58710 36224 58716 36236
rect 58115 36196 58716 36224
rect 58115 36193 58127 36196
rect 58069 36187 58127 36193
rect 58710 36184 58716 36196
rect 58768 36184 58774 36236
rect 62206 36184 62212 36236
rect 62264 36224 62270 36236
rect 62669 36227 62727 36233
rect 62669 36224 62681 36227
rect 62264 36196 62681 36224
rect 62264 36184 62270 36196
rect 62669 36193 62681 36196
rect 62715 36193 62727 36227
rect 62669 36187 62727 36193
rect 65797 36227 65855 36233
rect 65797 36193 65809 36227
rect 65843 36224 65855 36227
rect 65978 36224 65984 36236
rect 65843 36196 65984 36224
rect 65843 36193 65855 36196
rect 65797 36187 65855 36193
rect 65978 36184 65984 36196
rect 66036 36184 66042 36236
rect 66088 36233 66116 36264
rect 69937 36261 69949 36295
rect 69983 36292 69995 36295
rect 71498 36292 71504 36304
rect 69983 36264 71504 36292
rect 69983 36261 69995 36264
rect 69937 36255 69995 36261
rect 71498 36252 71504 36264
rect 71556 36252 71562 36304
rect 77312 36236 77340 36332
rect 77938 36320 77944 36332
rect 77996 36320 78002 36372
rect 78674 36360 78680 36372
rect 78635 36332 78680 36360
rect 78674 36320 78680 36332
rect 78732 36320 78738 36372
rect 82170 36320 82176 36372
rect 82228 36360 82234 36372
rect 84197 36363 84255 36369
rect 84197 36360 84209 36363
rect 82228 36332 84209 36360
rect 82228 36320 82234 36332
rect 84197 36329 84209 36332
rect 84243 36329 84255 36363
rect 86954 36360 86960 36372
rect 86915 36332 86960 36360
rect 84197 36323 84255 36329
rect 79781 36295 79839 36301
rect 79781 36261 79793 36295
rect 79827 36292 79839 36295
rect 81342 36292 81348 36304
rect 79827 36264 81348 36292
rect 79827 36261 79839 36264
rect 79781 36255 79839 36261
rect 81342 36252 81348 36264
rect 81400 36252 81406 36304
rect 83550 36252 83556 36304
rect 83608 36292 83614 36304
rect 83921 36295 83979 36301
rect 83921 36292 83933 36295
rect 83608 36264 83933 36292
rect 83608 36252 83614 36264
rect 83921 36261 83933 36264
rect 83967 36261 83979 36295
rect 84212 36292 84240 36323
rect 86954 36320 86960 36332
rect 87012 36320 87018 36372
rect 85393 36295 85451 36301
rect 85393 36292 85405 36295
rect 84212 36264 85405 36292
rect 83921 36255 83979 36261
rect 85393 36261 85405 36264
rect 85439 36261 85451 36295
rect 85393 36255 85451 36261
rect 85945 36295 86003 36301
rect 85945 36261 85957 36295
rect 85991 36292 86003 36295
rect 86218 36292 86224 36304
rect 85991 36264 86224 36292
rect 85991 36261 86003 36264
rect 85945 36255 86003 36261
rect 86218 36252 86224 36264
rect 86276 36252 86282 36304
rect 66073 36227 66131 36233
rect 66073 36193 66085 36227
rect 66119 36193 66131 36227
rect 66073 36187 66131 36193
rect 69566 36184 69572 36236
rect 69624 36224 69630 36236
rect 70121 36227 70179 36233
rect 70121 36224 70133 36227
rect 69624 36196 70133 36224
rect 69624 36184 69630 36196
rect 70121 36193 70133 36196
rect 70167 36193 70179 36227
rect 70121 36187 70179 36193
rect 70489 36227 70547 36233
rect 70489 36193 70501 36227
rect 70535 36224 70547 36227
rect 71682 36224 71688 36236
rect 70535 36196 71688 36224
rect 70535 36193 70547 36196
rect 70489 36187 70547 36193
rect 62114 36116 62120 36168
rect 62172 36156 62178 36168
rect 62393 36159 62451 36165
rect 62393 36156 62405 36159
rect 62172 36128 62405 36156
rect 62172 36116 62178 36128
rect 62393 36125 62405 36128
rect 62439 36125 62451 36159
rect 62393 36119 62451 36125
rect 65518 36116 65524 36168
rect 65576 36156 65582 36168
rect 65889 36159 65947 36165
rect 65889 36156 65901 36159
rect 65576 36128 65901 36156
rect 65576 36116 65582 36128
rect 65889 36125 65901 36128
rect 65935 36125 65947 36159
rect 65889 36119 65947 36125
rect 66257 36159 66315 36165
rect 66257 36125 66269 36159
rect 66303 36125 66315 36159
rect 70136 36156 70164 36187
rect 71682 36184 71688 36196
rect 71740 36184 71746 36236
rect 72145 36227 72203 36233
rect 72145 36193 72157 36227
rect 72191 36224 72203 36227
rect 72237 36227 72295 36233
rect 72237 36224 72249 36227
rect 72191 36196 72249 36224
rect 72191 36193 72203 36196
rect 72145 36187 72203 36193
rect 72237 36193 72249 36196
rect 72283 36224 72295 36227
rect 77294 36224 77300 36236
rect 72283 36196 77300 36224
rect 72283 36193 72295 36196
rect 72237 36187 72295 36193
rect 70581 36159 70639 36165
rect 70581 36156 70593 36159
rect 70136 36128 70593 36156
rect 66257 36119 66315 36125
rect 70581 36125 70593 36128
rect 70627 36156 70639 36159
rect 71590 36156 71596 36168
rect 70627 36128 71596 36156
rect 70627 36125 70639 36128
rect 70581 36119 70639 36125
rect 60550 36048 60556 36100
rect 60608 36088 60614 36100
rect 66272 36088 66300 36119
rect 71590 36116 71596 36128
rect 71648 36116 71654 36168
rect 60608 36060 62344 36088
rect 60608 36048 60614 36060
rect 62206 36020 62212 36032
rect 56735 35992 57652 36020
rect 62167 35992 62212 36020
rect 56735 35989 56747 35992
rect 56689 35983 56747 35989
rect 62206 35980 62212 35992
rect 62264 35980 62270 36032
rect 62316 36020 62344 36060
rect 63328 36060 66300 36088
rect 63328 36020 63356 36060
rect 62316 35992 63356 36020
rect 63957 36023 64015 36029
rect 63957 35989 63969 36023
rect 64003 36020 64015 36023
rect 64506 36020 64512 36032
rect 64003 35992 64512 36020
rect 64003 35989 64015 35992
rect 63957 35983 64015 35989
rect 64506 35980 64512 35992
rect 64564 35980 64570 36032
rect 69014 35980 69020 36032
rect 69072 36020 69078 36032
rect 70118 36020 70124 36032
rect 69072 35992 70124 36020
rect 69072 35980 69078 35992
rect 70118 35980 70124 35992
rect 70176 36020 70182 36032
rect 72160 36020 72188 36187
rect 77294 36184 77300 36196
rect 77352 36184 77358 36236
rect 79962 36224 79968 36236
rect 79923 36196 79968 36224
rect 79962 36184 79968 36196
rect 80020 36184 80026 36236
rect 82814 36224 82820 36236
rect 82775 36196 82820 36224
rect 82814 36184 82820 36196
rect 82872 36224 82878 36236
rect 83185 36227 83243 36233
rect 83185 36224 83197 36227
rect 82872 36196 83197 36224
rect 82872 36184 82878 36196
rect 83185 36193 83197 36196
rect 83231 36193 83243 36227
rect 84105 36227 84163 36233
rect 84105 36224 84117 36227
rect 83185 36187 83243 36193
rect 83752 36196 84117 36224
rect 72510 36156 72516 36168
rect 72471 36128 72516 36156
rect 72510 36116 72516 36128
rect 72568 36116 72574 36168
rect 77570 36156 77576 36168
rect 77531 36128 77576 36156
rect 77570 36116 77576 36128
rect 77628 36116 77634 36168
rect 79686 36048 79692 36100
rect 79744 36088 79750 36100
rect 82998 36088 83004 36100
rect 79744 36060 83004 36088
rect 79744 36048 79750 36060
rect 82998 36048 83004 36060
rect 83056 36088 83062 36100
rect 83752 36097 83780 36196
rect 84105 36193 84117 36196
rect 84151 36224 84163 36227
rect 84194 36224 84200 36236
rect 84151 36196 84200 36224
rect 84151 36193 84163 36196
rect 84105 36187 84163 36193
rect 84194 36184 84200 36196
rect 84252 36184 84258 36236
rect 85577 36227 85635 36233
rect 85577 36193 85589 36227
rect 85623 36224 85635 36227
rect 86310 36224 86316 36236
rect 85623 36196 86316 36224
rect 85623 36193 85635 36196
rect 85577 36187 85635 36193
rect 86310 36184 86316 36196
rect 86368 36184 86374 36236
rect 86770 36224 86776 36236
rect 86731 36196 86776 36224
rect 86770 36184 86776 36196
rect 86828 36184 86834 36236
rect 83737 36091 83795 36097
rect 83737 36088 83749 36091
rect 83056 36060 83749 36088
rect 83056 36048 83062 36060
rect 83737 36057 83749 36060
rect 83783 36057 83795 36091
rect 83737 36051 83795 36057
rect 70176 35992 72188 36020
rect 70176 35980 70182 35992
rect 78214 35980 78220 36032
rect 78272 36020 78278 36032
rect 80057 36023 80115 36029
rect 80057 36020 80069 36023
rect 78272 35992 80069 36020
rect 78272 35980 78278 35992
rect 80057 35989 80069 35992
rect 80103 36020 80115 36023
rect 80238 36020 80244 36032
rect 80103 35992 80244 36020
rect 80103 35989 80115 35992
rect 80057 35983 80115 35989
rect 80238 35980 80244 35992
rect 80296 35980 80302 36032
rect 1104 35930 111136 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 65686 35930
rect 65738 35878 65750 35930
rect 65802 35878 65814 35930
rect 65866 35878 65878 35930
rect 65930 35878 96406 35930
rect 96458 35878 96470 35930
rect 96522 35878 96534 35930
rect 96586 35878 96598 35930
rect 96650 35878 111136 35930
rect 1104 35856 111136 35878
rect 4062 35776 4068 35828
rect 4120 35816 4126 35828
rect 6362 35816 6368 35828
rect 4120 35788 6368 35816
rect 4120 35776 4126 35788
rect 6362 35776 6368 35788
rect 6420 35776 6426 35828
rect 16025 35819 16083 35825
rect 16025 35785 16037 35819
rect 16071 35816 16083 35819
rect 26142 35816 26148 35828
rect 16071 35788 26148 35816
rect 16071 35785 16083 35788
rect 16025 35779 16083 35785
rect 26142 35776 26148 35788
rect 26200 35776 26206 35828
rect 27157 35819 27215 35825
rect 27157 35785 27169 35819
rect 27203 35816 27215 35819
rect 30834 35816 30840 35828
rect 27203 35788 30840 35816
rect 27203 35785 27215 35788
rect 27157 35779 27215 35785
rect 21726 35748 21732 35760
rect 21687 35720 21732 35748
rect 21726 35708 21732 35720
rect 21784 35708 21790 35760
rect 22462 35708 22468 35760
rect 22520 35748 22526 35760
rect 27172 35748 27200 35779
rect 30834 35776 30840 35788
rect 30892 35776 30898 35828
rect 30926 35776 30932 35828
rect 30984 35816 30990 35828
rect 31021 35819 31079 35825
rect 31021 35816 31033 35819
rect 30984 35788 31033 35816
rect 30984 35776 30990 35788
rect 31021 35785 31033 35788
rect 31067 35816 31079 35819
rect 31662 35816 31668 35828
rect 31067 35788 31668 35816
rect 31067 35785 31079 35788
rect 31021 35779 31079 35785
rect 31662 35776 31668 35788
rect 31720 35816 31726 35828
rect 32214 35816 32220 35828
rect 31720 35788 32220 35816
rect 31720 35776 31726 35788
rect 32214 35776 32220 35788
rect 32272 35776 32278 35828
rect 32306 35776 32312 35828
rect 32364 35816 32370 35828
rect 34425 35819 34483 35825
rect 34425 35816 34437 35819
rect 32364 35788 34437 35816
rect 32364 35776 32370 35788
rect 34425 35785 34437 35788
rect 34471 35816 34483 35819
rect 35250 35816 35256 35828
rect 34471 35788 35256 35816
rect 34471 35785 34483 35788
rect 34425 35779 34483 35785
rect 35250 35776 35256 35788
rect 35308 35776 35314 35828
rect 35342 35776 35348 35828
rect 35400 35816 35406 35828
rect 38378 35816 38384 35828
rect 35400 35788 38384 35816
rect 35400 35776 35406 35788
rect 38378 35776 38384 35788
rect 38436 35776 38442 35828
rect 38470 35776 38476 35828
rect 38528 35816 38534 35828
rect 39669 35819 39727 35825
rect 39669 35816 39681 35819
rect 38528 35788 39681 35816
rect 38528 35776 38534 35788
rect 39669 35785 39681 35788
rect 39715 35816 39727 35819
rect 40770 35816 40776 35828
rect 39715 35788 40776 35816
rect 39715 35785 39727 35788
rect 39669 35779 39727 35785
rect 40770 35776 40776 35788
rect 40828 35776 40834 35828
rect 40862 35776 40868 35828
rect 40920 35816 40926 35828
rect 40920 35788 46244 35816
rect 40920 35776 40926 35788
rect 22520 35720 27200 35748
rect 22520 35708 22526 35720
rect 3881 35683 3939 35689
rect 3881 35649 3893 35683
rect 3927 35680 3939 35683
rect 5166 35680 5172 35692
rect 3927 35652 5172 35680
rect 3927 35649 3939 35652
rect 3881 35643 3939 35649
rect 5166 35640 5172 35652
rect 5224 35640 5230 35692
rect 5626 35640 5632 35692
rect 5684 35680 5690 35692
rect 14918 35680 14924 35692
rect 5684 35652 14924 35680
rect 5684 35640 5690 35652
rect 14918 35640 14924 35652
rect 14976 35640 14982 35692
rect 20625 35683 20683 35689
rect 20625 35649 20637 35683
rect 20671 35680 20683 35683
rect 20714 35680 20720 35692
rect 20671 35652 20720 35680
rect 20671 35649 20683 35652
rect 20625 35643 20683 35649
rect 20714 35640 20720 35652
rect 20772 35640 20778 35692
rect 3605 35615 3663 35621
rect 3605 35581 3617 35615
rect 3651 35612 3663 35615
rect 3694 35612 3700 35624
rect 3651 35584 3700 35612
rect 3651 35581 3663 35584
rect 3605 35575 3663 35581
rect 3694 35572 3700 35584
rect 3752 35572 3758 35624
rect 6270 35572 6276 35624
rect 6328 35612 6334 35624
rect 6825 35615 6883 35621
rect 6825 35612 6837 35615
rect 6328 35584 6837 35612
rect 6328 35572 6334 35584
rect 6825 35581 6837 35584
rect 6871 35581 6883 35615
rect 6825 35575 6883 35581
rect 7377 35615 7435 35621
rect 7377 35581 7389 35615
rect 7423 35612 7435 35615
rect 10134 35612 10140 35624
rect 7423 35584 10140 35612
rect 7423 35581 7435 35584
rect 7377 35575 7435 35581
rect 10134 35572 10140 35584
rect 10192 35572 10198 35624
rect 10873 35615 10931 35621
rect 10873 35581 10885 35615
rect 10919 35581 10931 35615
rect 10873 35575 10931 35581
rect 4798 35504 4804 35556
rect 4856 35544 4862 35556
rect 5353 35547 5411 35553
rect 5353 35544 5365 35547
rect 4856 35516 5365 35544
rect 4856 35504 4862 35516
rect 5353 35513 5365 35516
rect 5399 35513 5411 35547
rect 10318 35544 10324 35556
rect 10279 35516 10324 35544
rect 5353 35507 5411 35513
rect 10318 35504 10324 35516
rect 10376 35504 10382 35556
rect 4154 35436 4160 35488
rect 4212 35476 4218 35488
rect 4985 35479 5043 35485
rect 4985 35476 4997 35479
rect 4212 35448 4997 35476
rect 4212 35436 4218 35448
rect 4985 35445 4997 35448
rect 5031 35445 5043 35479
rect 4985 35439 5043 35445
rect 6086 35436 6092 35488
rect 6144 35476 6150 35488
rect 6917 35479 6975 35485
rect 6917 35476 6929 35479
rect 6144 35448 6929 35476
rect 6144 35436 6150 35448
rect 6917 35445 6929 35448
rect 6963 35445 6975 35479
rect 10226 35476 10232 35488
rect 10187 35448 10232 35476
rect 6917 35439 6975 35445
rect 10226 35436 10232 35448
rect 10284 35476 10290 35488
rect 10888 35476 10916 35575
rect 10962 35572 10968 35624
rect 11020 35612 11026 35624
rect 11149 35615 11207 35621
rect 11149 35612 11161 35615
rect 11020 35584 11161 35612
rect 11020 35572 11026 35584
rect 11149 35581 11161 35584
rect 11195 35581 11207 35615
rect 11149 35575 11207 35581
rect 11333 35615 11391 35621
rect 11333 35581 11345 35615
rect 11379 35612 11391 35615
rect 13357 35615 13415 35621
rect 11379 35584 11560 35612
rect 11379 35581 11391 35584
rect 11333 35575 11391 35581
rect 11532 35488 11560 35584
rect 13357 35581 13369 35615
rect 13403 35581 13415 35615
rect 13630 35612 13636 35624
rect 13591 35584 13636 35612
rect 13357 35575 13415 35581
rect 11514 35476 11520 35488
rect 10284 35448 10916 35476
rect 11475 35448 11520 35476
rect 10284 35436 10290 35448
rect 11514 35436 11520 35448
rect 11572 35436 11578 35488
rect 13265 35479 13323 35485
rect 13265 35445 13277 35479
rect 13311 35476 13323 35479
rect 13372 35476 13400 35575
rect 13630 35572 13636 35584
rect 13688 35572 13694 35624
rect 14550 35572 14556 35624
rect 14608 35612 14614 35624
rect 15749 35615 15807 35621
rect 15749 35612 15761 35615
rect 14608 35584 15761 35612
rect 14608 35572 14614 35584
rect 15749 35581 15761 35584
rect 15795 35612 15807 35615
rect 15841 35615 15899 35621
rect 15841 35612 15853 35615
rect 15795 35584 15853 35612
rect 15795 35581 15807 35584
rect 15749 35575 15807 35581
rect 15841 35581 15853 35584
rect 15887 35581 15899 35615
rect 15841 35575 15899 35581
rect 20349 35615 20407 35621
rect 20349 35581 20361 35615
rect 20395 35612 20407 35615
rect 20990 35612 20996 35624
rect 20395 35584 20996 35612
rect 20395 35581 20407 35584
rect 20349 35575 20407 35581
rect 20990 35572 20996 35584
rect 21048 35572 21054 35624
rect 22922 35612 22928 35624
rect 21284 35584 22928 35612
rect 15010 35544 15016 35556
rect 14923 35516 15016 35544
rect 15010 35504 15016 35516
rect 15068 35544 15074 35556
rect 15068 35516 16252 35544
rect 15068 35504 15074 35516
rect 13446 35476 13452 35488
rect 13311 35448 13452 35476
rect 13311 35445 13323 35448
rect 13265 35439 13323 35445
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 16224 35476 16252 35516
rect 21284 35476 21312 35584
rect 22922 35572 22928 35584
rect 22980 35572 22986 35624
rect 25406 35612 25412 35624
rect 25367 35584 25412 35612
rect 25406 35572 25412 35584
rect 25464 35612 25470 35624
rect 25593 35615 25651 35621
rect 25593 35612 25605 35615
rect 25464 35584 25605 35612
rect 25464 35572 25470 35584
rect 25593 35581 25605 35584
rect 25639 35581 25651 35615
rect 25593 35575 25651 35581
rect 25777 35615 25835 35621
rect 25777 35581 25789 35615
rect 25823 35612 25835 35615
rect 25976 35612 26004 35720
rect 27522 35708 27528 35760
rect 27580 35748 27586 35760
rect 31386 35748 31392 35760
rect 27580 35720 31392 35748
rect 27580 35708 27586 35720
rect 31386 35708 31392 35720
rect 31444 35708 31450 35760
rect 31496 35720 31800 35748
rect 30558 35680 30564 35692
rect 29288 35652 29592 35680
rect 30519 35652 30564 35680
rect 26237 35615 26295 35621
rect 26237 35612 26249 35615
rect 25823 35584 25912 35612
rect 25976 35584 26249 35612
rect 25823 35581 25835 35584
rect 25777 35575 25835 35581
rect 21358 35504 21364 35556
rect 21416 35544 21422 35556
rect 25884 35544 25912 35584
rect 26237 35581 26249 35584
rect 26283 35581 26295 35615
rect 26237 35575 26295 35581
rect 26329 35615 26387 35621
rect 26329 35581 26341 35615
rect 26375 35612 26387 35615
rect 27246 35612 27252 35624
rect 26375 35584 27252 35612
rect 26375 35581 26387 35584
rect 26329 35575 26387 35581
rect 26344 35544 26372 35575
rect 27246 35572 27252 35584
rect 27304 35572 27310 35624
rect 28626 35572 28632 35624
rect 28684 35612 28690 35624
rect 29288 35621 29316 35652
rect 29273 35615 29331 35621
rect 29273 35612 29285 35615
rect 28684 35584 29285 35612
rect 28684 35572 28690 35584
rect 29273 35581 29285 35584
rect 29319 35581 29331 35615
rect 29454 35612 29460 35624
rect 29415 35584 29460 35612
rect 29273 35575 29331 35581
rect 29454 35572 29460 35584
rect 29512 35572 29518 35624
rect 29564 35612 29592 35652
rect 30558 35640 30564 35652
rect 30616 35640 30622 35692
rect 30837 35683 30895 35689
rect 30837 35649 30849 35683
rect 30883 35680 30895 35683
rect 30926 35680 30932 35692
rect 30883 35652 30932 35680
rect 30883 35649 30895 35652
rect 30837 35643 30895 35649
rect 29917 35615 29975 35621
rect 29917 35612 29929 35615
rect 29564 35584 29929 35612
rect 29917 35581 29929 35584
rect 29963 35581 29975 35615
rect 29917 35575 29975 35581
rect 30006 35572 30012 35624
rect 30064 35612 30070 35624
rect 30852 35612 30880 35643
rect 30926 35640 30932 35652
rect 30984 35640 30990 35692
rect 30064 35584 30880 35612
rect 30064 35572 30070 35584
rect 31018 35572 31024 35624
rect 31076 35612 31082 35624
rect 31496 35621 31524 35720
rect 31481 35615 31539 35621
rect 31481 35612 31493 35615
rect 31076 35584 31493 35612
rect 31076 35572 31082 35584
rect 31481 35581 31493 35584
rect 31527 35581 31539 35615
rect 31481 35575 31539 35581
rect 31570 35572 31576 35624
rect 31628 35621 31634 35624
rect 31628 35615 31677 35621
rect 31628 35581 31631 35615
rect 31665 35581 31677 35615
rect 31772 35612 31800 35720
rect 32674 35708 32680 35760
rect 32732 35748 32738 35760
rect 33045 35751 33103 35757
rect 32732 35720 32777 35748
rect 32732 35708 32738 35720
rect 33045 35717 33057 35751
rect 33091 35748 33103 35751
rect 33229 35751 33287 35757
rect 33229 35748 33241 35751
rect 33091 35720 33241 35748
rect 33091 35717 33103 35720
rect 33045 35711 33103 35717
rect 33229 35717 33241 35720
rect 33275 35748 33287 35751
rect 41322 35748 41328 35760
rect 33275 35720 41328 35748
rect 33275 35717 33287 35720
rect 33229 35711 33287 35717
rect 32125 35615 32183 35621
rect 32125 35612 32137 35615
rect 31772 35584 32137 35612
rect 31628 35575 31677 35581
rect 32125 35581 32137 35584
rect 32171 35581 32183 35615
rect 32125 35575 32183 35581
rect 31628 35572 31634 35575
rect 32214 35572 32220 35624
rect 32272 35612 32278 35624
rect 33060 35612 33088 35711
rect 41322 35708 41328 35720
rect 41380 35708 41386 35760
rect 41966 35708 41972 35760
rect 42024 35748 42030 35760
rect 42981 35751 43039 35757
rect 42981 35748 42993 35751
rect 42024 35720 42993 35748
rect 42024 35708 42030 35720
rect 42981 35717 42993 35720
rect 43027 35717 43039 35751
rect 46216 35748 46244 35788
rect 48958 35776 48964 35828
rect 49016 35816 49022 35828
rect 49694 35816 49700 35828
rect 49016 35788 49700 35816
rect 49016 35776 49022 35788
rect 49694 35776 49700 35788
rect 49752 35776 49758 35828
rect 50798 35776 50804 35828
rect 50856 35816 50862 35828
rect 51077 35819 51135 35825
rect 51077 35816 51089 35819
rect 50856 35788 51089 35816
rect 50856 35776 50862 35788
rect 51077 35785 51089 35788
rect 51123 35785 51135 35819
rect 52365 35819 52423 35825
rect 51077 35779 51135 35785
rect 51883 35788 52316 35816
rect 51883 35748 51911 35788
rect 51994 35748 52000 35760
rect 46216 35720 51911 35748
rect 51955 35720 52000 35748
rect 42981 35711 43039 35717
rect 51994 35708 52000 35720
rect 52052 35708 52058 35760
rect 52288 35748 52316 35788
rect 52365 35785 52377 35819
rect 52411 35816 52423 35819
rect 53650 35816 53656 35828
rect 52411 35788 53656 35816
rect 52411 35785 52423 35788
rect 52365 35779 52423 35785
rect 53650 35776 53656 35788
rect 53708 35776 53714 35828
rect 54846 35816 54852 35828
rect 54807 35788 54852 35816
rect 54846 35776 54852 35788
rect 54904 35776 54910 35828
rect 55030 35816 55036 35828
rect 54991 35788 55036 35816
rect 55030 35776 55036 35788
rect 55088 35776 55094 35828
rect 55674 35776 55680 35828
rect 55732 35816 55738 35828
rect 58250 35816 58256 35828
rect 55732 35788 58256 35816
rect 55732 35776 55738 35788
rect 58250 35776 58256 35788
rect 58308 35776 58314 35828
rect 63681 35819 63739 35825
rect 58452 35788 63632 35816
rect 56781 35751 56839 35757
rect 56781 35748 56793 35751
rect 52288 35720 56793 35748
rect 56781 35717 56793 35720
rect 56827 35748 56839 35751
rect 56965 35751 57023 35757
rect 56965 35748 56977 35751
rect 56827 35720 56977 35748
rect 56827 35717 56839 35720
rect 56781 35711 56839 35717
rect 56965 35717 56977 35720
rect 57011 35748 57023 35751
rect 57011 35720 57560 35748
rect 57011 35717 57023 35720
rect 56965 35711 57023 35717
rect 35621 35683 35679 35689
rect 35621 35649 35633 35683
rect 35667 35680 35679 35683
rect 35710 35680 35716 35692
rect 35667 35652 35716 35680
rect 35667 35649 35679 35652
rect 35621 35643 35679 35649
rect 35710 35640 35716 35652
rect 35768 35640 35774 35692
rect 35805 35683 35863 35689
rect 35805 35649 35817 35683
rect 35851 35680 35863 35683
rect 35986 35680 35992 35692
rect 35851 35652 35992 35680
rect 35851 35649 35863 35652
rect 35805 35643 35863 35649
rect 35986 35640 35992 35652
rect 36044 35640 36050 35692
rect 38562 35680 38568 35692
rect 36188 35652 38568 35680
rect 32272 35584 33088 35612
rect 35529 35615 35587 35621
rect 32272 35572 32278 35584
rect 35529 35581 35541 35615
rect 35575 35612 35587 35615
rect 35897 35615 35955 35621
rect 35575 35584 35664 35612
rect 35575 35581 35587 35584
rect 35529 35575 35587 35581
rect 21416 35516 26372 35544
rect 26881 35547 26939 35553
rect 21416 35504 21422 35516
rect 26881 35513 26893 35547
rect 26927 35544 26939 35547
rect 33410 35544 33416 35556
rect 26927 35516 33416 35544
rect 26927 35513 26939 35516
rect 26881 35507 26939 35513
rect 33410 35504 33416 35516
rect 33468 35504 33474 35556
rect 33502 35504 33508 35556
rect 33560 35544 33566 35556
rect 34885 35547 34943 35553
rect 34885 35544 34897 35547
rect 33560 35516 34897 35544
rect 33560 35504 33566 35516
rect 34885 35513 34897 35516
rect 34931 35513 34943 35547
rect 34885 35507 34943 35513
rect 35250 35504 35256 35556
rect 35308 35544 35314 35556
rect 35636 35544 35664 35584
rect 35897 35581 35909 35615
rect 35943 35612 35955 35615
rect 36188 35612 36216 35652
rect 38562 35640 38568 35652
rect 38620 35640 38626 35692
rect 39482 35680 39488 35692
rect 39443 35652 39488 35680
rect 39482 35640 39488 35652
rect 39540 35640 39546 35692
rect 40313 35683 40371 35689
rect 40313 35649 40325 35683
rect 40359 35680 40371 35683
rect 41785 35683 41843 35689
rect 40359 35652 40908 35680
rect 40359 35649 40371 35652
rect 40313 35643 40371 35649
rect 38197 35615 38255 35621
rect 38197 35612 38209 35615
rect 35943 35584 36216 35612
rect 37844 35584 38209 35612
rect 35943 35581 35955 35584
rect 35897 35575 35955 35581
rect 35308 35516 35664 35544
rect 35308 35504 35314 35516
rect 16224 35448 21312 35476
rect 22002 35436 22008 35488
rect 22060 35476 22066 35488
rect 22097 35479 22155 35485
rect 22097 35476 22109 35479
rect 22060 35448 22109 35476
rect 22060 35436 22066 35448
rect 22097 35445 22109 35448
rect 22143 35476 22155 35479
rect 26510 35476 26516 35488
rect 22143 35448 26516 35476
rect 22143 35445 22155 35448
rect 22097 35439 22155 35445
rect 26510 35436 26516 35448
rect 26568 35436 26574 35488
rect 28626 35436 28632 35488
rect 28684 35476 28690 35488
rect 28813 35479 28871 35485
rect 28813 35476 28825 35479
rect 28684 35448 28825 35476
rect 28684 35436 28690 35448
rect 28813 35445 28825 35448
rect 28859 35476 28871 35479
rect 28997 35479 29055 35485
rect 28997 35476 29009 35479
rect 28859 35448 29009 35476
rect 28859 35445 28871 35448
rect 28813 35439 28871 35445
rect 28997 35445 29009 35448
rect 29043 35445 29055 35479
rect 28997 35439 29055 35445
rect 29454 35436 29460 35488
rect 29512 35476 29518 35488
rect 30006 35476 30012 35488
rect 29512 35448 30012 35476
rect 29512 35436 29518 35448
rect 30006 35436 30012 35448
rect 30064 35436 30070 35488
rect 31018 35436 31024 35488
rect 31076 35476 31082 35488
rect 31113 35479 31171 35485
rect 31113 35476 31125 35479
rect 31076 35448 31125 35476
rect 31076 35436 31082 35448
rect 31113 35445 31125 35448
rect 31159 35476 31171 35479
rect 31297 35479 31355 35485
rect 31297 35476 31309 35479
rect 31159 35448 31309 35476
rect 31159 35445 31171 35448
rect 31113 35439 31171 35445
rect 31297 35445 31309 35448
rect 31343 35445 31355 35479
rect 31297 35439 31355 35445
rect 31386 35436 31392 35488
rect 31444 35476 31450 35488
rect 34609 35479 34667 35485
rect 34609 35476 34621 35479
rect 31444 35448 34621 35476
rect 31444 35436 31450 35448
rect 34609 35445 34621 35448
rect 34655 35476 34667 35479
rect 35912 35476 35940 35575
rect 37844 35488 37872 35584
rect 38197 35581 38209 35584
rect 38243 35581 38255 35615
rect 38197 35575 38255 35581
rect 38381 35615 38439 35621
rect 38381 35581 38393 35615
rect 38427 35581 38439 35615
rect 38381 35575 38439 35581
rect 38396 35544 38424 35575
rect 38470 35572 38476 35624
rect 38528 35612 38534 35624
rect 38841 35615 38899 35621
rect 38841 35612 38853 35615
rect 38528 35584 38853 35612
rect 38528 35572 38534 35584
rect 38841 35581 38853 35584
rect 38887 35581 38899 35615
rect 38841 35575 38899 35581
rect 38933 35615 38991 35621
rect 38933 35581 38945 35615
rect 38979 35612 38991 35615
rect 39853 35615 39911 35621
rect 39853 35612 39865 35615
rect 38979 35584 39865 35612
rect 38979 35581 38991 35584
rect 38933 35575 38991 35581
rect 39853 35581 39865 35584
rect 39899 35612 39911 35615
rect 40635 35615 40693 35621
rect 40635 35612 40647 35615
rect 39899 35584 40647 35612
rect 39899 35581 39911 35584
rect 39853 35575 39911 35581
rect 40635 35581 40647 35584
rect 40681 35581 40693 35615
rect 40770 35612 40776 35624
rect 40731 35584 40776 35612
rect 40635 35575 40693 35581
rect 39942 35544 39948 35556
rect 38396 35516 39948 35544
rect 39942 35504 39948 35516
rect 40000 35504 40006 35556
rect 37826 35476 37832 35488
rect 34655 35448 35940 35476
rect 37787 35448 37832 35476
rect 34655 35445 34667 35448
rect 34609 35439 34667 35445
rect 37826 35436 37832 35448
rect 37884 35436 37890 35488
rect 38010 35476 38016 35488
rect 37971 35448 38016 35476
rect 38010 35436 38016 35448
rect 38068 35476 38074 35488
rect 38378 35476 38384 35488
rect 38068 35448 38384 35476
rect 38068 35436 38074 35448
rect 38378 35436 38384 35448
rect 38436 35436 38442 35488
rect 38470 35436 38476 35488
rect 38528 35476 38534 35488
rect 40129 35479 40187 35485
rect 40129 35476 40141 35479
rect 38528 35448 40141 35476
rect 38528 35436 38534 35448
rect 40129 35445 40141 35448
rect 40175 35476 40187 35479
rect 40313 35479 40371 35485
rect 40313 35476 40325 35479
rect 40175 35448 40325 35476
rect 40175 35445 40187 35448
rect 40129 35439 40187 35445
rect 40313 35445 40325 35448
rect 40359 35445 40371 35479
rect 40650 35476 40678 35575
rect 40770 35572 40776 35584
rect 40828 35572 40834 35624
rect 40880 35612 40908 35652
rect 41785 35649 41797 35683
rect 41831 35680 41843 35683
rect 42852 35683 42910 35689
rect 42852 35680 42864 35683
rect 41831 35652 42864 35680
rect 41831 35649 41843 35652
rect 41785 35643 41843 35649
rect 42852 35649 42864 35652
rect 42898 35649 42910 35683
rect 42852 35643 42910 35649
rect 43073 35683 43131 35689
rect 43073 35649 43085 35683
rect 43119 35680 43131 35683
rect 43622 35680 43628 35692
rect 43119 35652 43628 35680
rect 43119 35649 43131 35652
rect 43073 35643 43131 35649
rect 43622 35640 43628 35652
rect 43680 35640 43686 35692
rect 49050 35640 49056 35692
rect 49108 35680 49114 35692
rect 50709 35683 50767 35689
rect 49108 35652 49832 35680
rect 49108 35640 49114 35652
rect 41141 35615 41199 35621
rect 41141 35612 41153 35615
rect 40880 35584 41153 35612
rect 41141 35581 41153 35584
rect 41187 35581 41199 35615
rect 41141 35575 41199 35581
rect 41230 35572 41236 35624
rect 41288 35612 41294 35624
rect 42061 35615 42119 35621
rect 42061 35612 42073 35615
rect 41288 35584 42073 35612
rect 41288 35572 41294 35584
rect 42061 35581 42073 35584
rect 42107 35612 42119 35615
rect 42107 35584 49096 35612
rect 42107 35581 42119 35584
rect 42061 35575 42119 35581
rect 42702 35544 42708 35556
rect 42663 35516 42708 35544
rect 42702 35504 42708 35516
rect 42760 35504 42766 35556
rect 48958 35544 48964 35556
rect 42812 35516 48964 35544
rect 42245 35479 42303 35485
rect 42245 35476 42257 35479
rect 40650 35448 42257 35476
rect 40313 35439 40371 35445
rect 42245 35445 42257 35448
rect 42291 35476 42303 35479
rect 42812 35476 42840 35516
rect 48958 35504 48964 35516
rect 49016 35504 49022 35556
rect 49068 35544 49096 35584
rect 49418 35572 49424 35624
rect 49476 35612 49482 35624
rect 49605 35615 49663 35621
rect 49476 35584 49521 35612
rect 49476 35572 49482 35584
rect 49605 35581 49617 35615
rect 49651 35612 49663 35615
rect 49694 35612 49700 35624
rect 49651 35584 49700 35612
rect 49651 35581 49663 35584
rect 49605 35575 49663 35581
rect 49694 35572 49700 35584
rect 49752 35572 49758 35624
rect 49804 35612 49832 35652
rect 50709 35649 50721 35683
rect 50755 35680 50767 35683
rect 51868 35683 51926 35689
rect 51868 35680 51880 35683
rect 50755 35652 51880 35680
rect 50755 35649 50767 35652
rect 50709 35643 50767 35649
rect 51868 35649 51880 35652
rect 51914 35649 51926 35683
rect 51868 35643 51926 35649
rect 52089 35683 52147 35689
rect 52089 35649 52101 35683
rect 52135 35680 52147 35683
rect 53190 35680 53196 35692
rect 52135 35652 53196 35680
rect 52135 35649 52147 35652
rect 52089 35643 52147 35649
rect 53190 35640 53196 35652
rect 53248 35640 53254 35692
rect 57149 35683 57207 35689
rect 57149 35680 57161 35683
rect 53392 35652 57161 35680
rect 50065 35615 50123 35621
rect 50065 35612 50077 35615
rect 49804 35584 50077 35612
rect 50065 35581 50077 35584
rect 50111 35581 50123 35615
rect 50065 35575 50123 35581
rect 50157 35615 50215 35621
rect 50157 35581 50169 35615
rect 50203 35581 50215 35615
rect 50157 35575 50215 35581
rect 50172 35544 50200 35575
rect 51442 35572 51448 35624
rect 51500 35612 51506 35624
rect 53006 35612 53012 35624
rect 51500 35584 53012 35612
rect 51500 35572 51506 35584
rect 53006 35572 53012 35584
rect 53064 35572 53070 35624
rect 53282 35612 53288 35624
rect 53243 35584 53288 35612
rect 53282 35572 53288 35584
rect 53340 35572 53346 35624
rect 50893 35547 50951 35553
rect 50893 35544 50905 35547
rect 49068 35516 50905 35544
rect 50893 35513 50905 35516
rect 50939 35513 50951 35547
rect 50893 35507 50951 35513
rect 43346 35476 43352 35488
rect 42291 35448 42840 35476
rect 43307 35448 43352 35476
rect 42291 35445 42303 35448
rect 42245 35439 42303 35445
rect 43346 35436 43352 35448
rect 43404 35436 43410 35488
rect 49050 35476 49056 35488
rect 49011 35448 49056 35476
rect 49050 35436 49056 35448
rect 49108 35436 49114 35488
rect 49234 35476 49240 35488
rect 49195 35448 49240 35476
rect 49234 35436 49240 35448
rect 49292 35436 49298 35488
rect 49510 35436 49516 35488
rect 49568 35476 49574 35488
rect 50154 35476 50160 35488
rect 49568 35448 50160 35476
rect 49568 35436 49574 35448
rect 50154 35436 50160 35448
rect 50212 35436 50218 35488
rect 50908 35476 50936 35507
rect 50982 35504 50988 35556
rect 51040 35544 51046 35556
rect 51721 35547 51779 35553
rect 51721 35544 51733 35547
rect 51040 35516 51733 35544
rect 51040 35504 51046 35516
rect 51721 35513 51733 35516
rect 51767 35513 51779 35547
rect 53392 35544 53420 35652
rect 57149 35649 57161 35652
rect 57195 35649 57207 35683
rect 57149 35643 57207 35649
rect 55030 35572 55036 35624
rect 55088 35612 55094 35624
rect 55088 35584 55628 35612
rect 55088 35572 55094 35584
rect 55214 35544 55220 35556
rect 51721 35507 51779 35513
rect 53300 35516 53420 35544
rect 55175 35516 55220 35544
rect 53300 35476 53328 35516
rect 55214 35504 55220 35516
rect 55272 35504 55278 35556
rect 55600 35544 55628 35584
rect 55674 35572 55680 35624
rect 55732 35612 55738 35624
rect 55861 35615 55919 35621
rect 55732 35584 55777 35612
rect 55732 35572 55738 35584
rect 55861 35581 55873 35615
rect 55907 35612 55919 35615
rect 55950 35612 55956 35624
rect 55907 35584 55956 35612
rect 55907 35581 55919 35584
rect 55861 35575 55919 35581
rect 55950 35572 55956 35584
rect 56008 35572 56014 35624
rect 56229 35615 56287 35621
rect 56229 35581 56241 35615
rect 56275 35581 56287 35615
rect 56229 35575 56287 35581
rect 56413 35615 56471 35621
rect 56413 35581 56425 35615
rect 56459 35581 56471 35615
rect 56594 35612 56600 35624
rect 56555 35584 56600 35612
rect 56413 35575 56471 35581
rect 56244 35544 56272 35575
rect 55600 35516 56272 35544
rect 56428 35544 56456 35575
rect 56594 35572 56600 35584
rect 56652 35612 56658 35624
rect 57532 35621 57560 35720
rect 57333 35615 57391 35621
rect 57333 35612 57345 35615
rect 56652 35584 57345 35612
rect 56652 35572 56658 35584
rect 57333 35581 57345 35584
rect 57379 35581 57391 35615
rect 57333 35575 57391 35581
rect 57517 35615 57575 35621
rect 57517 35581 57529 35615
rect 57563 35612 57575 35615
rect 58069 35615 58127 35621
rect 58069 35612 58081 35615
rect 57563 35584 58081 35612
rect 57563 35581 57575 35584
rect 57517 35575 57575 35581
rect 58069 35581 58081 35584
rect 58115 35581 58127 35615
rect 58069 35575 58127 35581
rect 58253 35615 58311 35621
rect 58253 35581 58265 35615
rect 58299 35612 58311 35615
rect 58452 35612 58480 35788
rect 59538 35708 59544 35760
rect 59596 35748 59602 35760
rect 60274 35748 60280 35760
rect 59596 35720 60280 35748
rect 59596 35708 59602 35720
rect 60274 35708 60280 35720
rect 60332 35748 60338 35760
rect 62114 35748 62120 35760
rect 60332 35720 62120 35748
rect 60332 35708 60338 35720
rect 62114 35708 62120 35720
rect 62172 35748 62178 35760
rect 62942 35748 62948 35760
rect 62172 35720 62948 35748
rect 62172 35708 62178 35720
rect 62942 35708 62948 35720
rect 63000 35708 63006 35760
rect 63604 35748 63632 35788
rect 63681 35785 63693 35819
rect 63727 35816 63739 35819
rect 63727 35788 74396 35816
rect 63727 35785 63739 35788
rect 63681 35779 63739 35785
rect 63770 35748 63776 35760
rect 63604 35720 63776 35748
rect 63770 35708 63776 35720
rect 63828 35708 63834 35760
rect 68922 35708 68928 35760
rect 68980 35748 68986 35760
rect 69753 35751 69811 35757
rect 69753 35748 69765 35751
rect 68980 35720 69765 35748
rect 68980 35708 68986 35720
rect 69753 35717 69765 35720
rect 69799 35717 69811 35751
rect 70118 35748 70124 35760
rect 70079 35720 70124 35748
rect 69753 35711 69811 35717
rect 70118 35708 70124 35720
rect 70176 35708 70182 35760
rect 71314 35708 71320 35760
rect 71372 35748 71378 35760
rect 71685 35751 71743 35757
rect 71685 35748 71697 35751
rect 71372 35720 71697 35748
rect 71372 35708 71378 35720
rect 71685 35717 71697 35720
rect 71731 35717 71743 35751
rect 74368 35748 74396 35788
rect 74442 35776 74448 35828
rect 74500 35816 74506 35828
rect 79413 35819 79471 35825
rect 79413 35816 79425 35819
rect 74500 35788 79425 35816
rect 74500 35776 74506 35788
rect 79413 35785 79425 35788
rect 79459 35816 79471 35819
rect 79597 35819 79655 35825
rect 79597 35816 79609 35819
rect 79459 35788 79609 35816
rect 79459 35785 79471 35788
rect 79413 35779 79471 35785
rect 79597 35785 79609 35788
rect 79643 35785 79655 35819
rect 80057 35819 80115 35825
rect 80057 35816 80069 35819
rect 79597 35779 79655 35785
rect 79704 35788 80069 35816
rect 77113 35751 77171 35757
rect 77113 35748 77125 35751
rect 74368 35720 77125 35748
rect 71685 35711 71743 35717
rect 77113 35717 77125 35720
rect 77159 35748 77171 35751
rect 77202 35748 77208 35760
rect 77159 35720 77208 35748
rect 77159 35717 77171 35720
rect 77113 35711 77171 35717
rect 77202 35708 77208 35720
rect 77260 35748 77266 35760
rect 79137 35751 79195 35757
rect 77260 35720 78352 35748
rect 77260 35708 77266 35720
rect 77297 35683 77355 35689
rect 58299 35584 58480 35612
rect 58544 35652 75224 35680
rect 58299 35581 58311 35584
rect 58253 35575 58311 35581
rect 58268 35544 58296 35575
rect 56428 35516 58296 35544
rect 58342 35504 58348 35556
rect 58400 35544 58406 35556
rect 58544 35544 58572 35652
rect 62942 35572 62948 35624
rect 63000 35612 63006 35624
rect 63773 35615 63831 35621
rect 63773 35612 63785 35615
rect 63000 35584 63785 35612
rect 63000 35572 63006 35584
rect 63773 35581 63785 35584
rect 63819 35581 63831 35615
rect 64049 35615 64107 35621
rect 64049 35612 64061 35615
rect 63773 35575 63831 35581
rect 63880 35584 64061 35612
rect 58400 35516 58572 35544
rect 58621 35547 58679 35553
rect 58400 35504 58406 35516
rect 58621 35513 58633 35547
rect 58667 35544 58679 35547
rect 63880 35544 63908 35584
rect 64049 35581 64061 35584
rect 64095 35581 64107 35615
rect 64049 35575 64107 35581
rect 65429 35615 65487 35621
rect 65429 35581 65441 35615
rect 65475 35612 65487 35615
rect 66162 35612 66168 35624
rect 65475 35584 66168 35612
rect 65475 35581 65487 35584
rect 65429 35575 65487 35581
rect 66162 35572 66168 35584
rect 66220 35612 66226 35624
rect 66257 35615 66315 35621
rect 66257 35612 66269 35615
rect 66220 35584 66269 35612
rect 66220 35572 66226 35584
rect 66257 35581 66269 35584
rect 66303 35581 66315 35615
rect 68922 35612 68928 35624
rect 68883 35584 68928 35612
rect 66257 35575 66315 35581
rect 68922 35572 68928 35584
rect 68980 35572 68986 35624
rect 69014 35572 69020 35624
rect 69072 35612 69078 35624
rect 69477 35615 69535 35621
rect 69072 35584 69117 35612
rect 69072 35572 69078 35584
rect 69477 35581 69489 35615
rect 69523 35612 69535 35615
rect 70118 35612 70124 35624
rect 69523 35584 70124 35612
rect 69523 35581 69535 35584
rect 69477 35575 69535 35581
rect 70118 35572 70124 35584
rect 70176 35572 70182 35624
rect 70210 35572 70216 35624
rect 70268 35612 70274 35624
rect 70305 35615 70363 35621
rect 70305 35612 70317 35615
rect 70268 35584 70317 35612
rect 70268 35572 70274 35584
rect 70305 35581 70317 35584
rect 70351 35581 70363 35615
rect 70578 35612 70584 35624
rect 70539 35584 70584 35612
rect 70305 35575 70363 35581
rect 70578 35572 70584 35584
rect 70636 35572 70642 35624
rect 70670 35572 70676 35624
rect 70728 35612 70734 35624
rect 72786 35612 72792 35624
rect 70728 35584 71268 35612
rect 72747 35584 72792 35612
rect 70728 35572 70734 35584
rect 58667 35516 63908 35544
rect 69032 35544 69060 35572
rect 69566 35544 69572 35556
rect 69032 35516 69572 35544
rect 58667 35513 58679 35516
rect 58621 35507 58679 35513
rect 69566 35504 69572 35516
rect 69624 35504 69630 35556
rect 71240 35544 71268 35584
rect 72786 35572 72792 35584
rect 72844 35572 72850 35624
rect 75196 35612 75224 35652
rect 77297 35649 77309 35683
rect 77343 35680 77355 35683
rect 77570 35680 77576 35692
rect 77343 35652 77576 35680
rect 77343 35649 77355 35652
rect 77297 35643 77355 35649
rect 77570 35640 77576 35652
rect 77628 35640 77634 35692
rect 77846 35680 77852 35692
rect 77807 35652 77852 35680
rect 77846 35640 77852 35652
rect 77904 35640 77910 35692
rect 78324 35689 78352 35720
rect 79137 35717 79149 35751
rect 79183 35748 79195 35751
rect 79704 35748 79732 35788
rect 80057 35785 80069 35788
rect 80103 35785 80115 35819
rect 80422 35816 80428 35828
rect 80383 35788 80428 35816
rect 80057 35779 80115 35785
rect 80422 35776 80428 35788
rect 80480 35776 80486 35828
rect 82814 35776 82820 35828
rect 82872 35816 82878 35828
rect 86037 35819 86095 35825
rect 86037 35816 86049 35819
rect 82872 35788 86049 35816
rect 82872 35776 82878 35788
rect 82357 35751 82415 35757
rect 82357 35748 82369 35751
rect 79183 35720 79732 35748
rect 79796 35720 82369 35748
rect 79183 35717 79195 35720
rect 79137 35711 79195 35717
rect 78309 35683 78367 35689
rect 77956 35652 78260 35680
rect 77956 35612 77984 35652
rect 78122 35612 78128 35624
rect 75196 35584 77984 35612
rect 78083 35584 78128 35612
rect 78122 35572 78128 35584
rect 78180 35572 78186 35624
rect 78232 35612 78260 35652
rect 78309 35649 78321 35683
rect 78355 35649 78367 35683
rect 79796 35680 79824 35720
rect 82357 35717 82369 35720
rect 82403 35748 82415 35751
rect 83090 35748 83096 35760
rect 82403 35720 83096 35748
rect 82403 35717 82415 35720
rect 82357 35711 82415 35717
rect 83090 35708 83096 35720
rect 83148 35748 83154 35760
rect 83148 35720 84332 35748
rect 83148 35708 83154 35720
rect 79962 35689 79968 35692
rect 78309 35643 78367 35649
rect 78416 35652 79824 35680
rect 79928 35683 79968 35689
rect 78416 35612 78444 35652
rect 79928 35649 79940 35683
rect 79928 35643 79968 35649
rect 79962 35640 79968 35643
rect 80020 35640 80026 35692
rect 80146 35680 80152 35692
rect 80107 35652 80152 35680
rect 80146 35640 80152 35652
rect 80204 35640 80210 35692
rect 82817 35683 82875 35689
rect 82817 35649 82829 35683
rect 82863 35680 82875 35683
rect 82906 35680 82912 35692
rect 82863 35652 82912 35680
rect 82863 35649 82875 35652
rect 82817 35643 82875 35649
rect 82906 35640 82912 35652
rect 82964 35640 82970 35692
rect 83277 35683 83335 35689
rect 83277 35649 83289 35683
rect 83323 35680 83335 35683
rect 84194 35680 84200 35692
rect 83323 35652 84200 35680
rect 83323 35649 83335 35652
rect 83277 35643 83335 35649
rect 84194 35640 84200 35652
rect 84252 35640 84258 35692
rect 78232 35584 78444 35612
rect 79597 35615 79655 35621
rect 79597 35581 79609 35615
rect 79643 35612 79655 35615
rect 79781 35615 79839 35621
rect 79781 35612 79793 35615
rect 79643 35584 79793 35612
rect 79643 35581 79655 35584
rect 79597 35575 79655 35581
rect 79781 35581 79793 35584
rect 79827 35612 79839 35615
rect 82173 35615 82231 35621
rect 79827 35584 81848 35612
rect 79827 35581 79839 35584
rect 79781 35575 79839 35581
rect 79686 35544 79692 35556
rect 71240 35516 79692 35544
rect 79686 35504 79692 35516
rect 79744 35504 79750 35556
rect 81820 35544 81848 35584
rect 82173 35581 82185 35615
rect 82219 35612 82231 35615
rect 82722 35612 82728 35624
rect 82219 35584 82728 35612
rect 82219 35581 82231 35584
rect 82173 35575 82231 35581
rect 82722 35572 82728 35584
rect 82780 35572 82786 35624
rect 82924 35612 82952 35640
rect 83918 35612 83924 35624
rect 82924 35584 83780 35612
rect 83879 35584 83924 35612
rect 82909 35547 82967 35553
rect 82909 35544 82921 35547
rect 81820 35516 82921 35544
rect 82909 35513 82921 35516
rect 82955 35544 82967 35547
rect 82998 35544 83004 35556
rect 82955 35516 83004 35544
rect 82955 35513 82967 35516
rect 82909 35507 82967 35513
rect 82998 35504 83004 35516
rect 83056 35504 83062 35556
rect 83752 35544 83780 35584
rect 83918 35572 83924 35584
rect 83976 35572 83982 35624
rect 84304 35621 84332 35720
rect 84013 35615 84071 35621
rect 84013 35581 84025 35615
rect 84059 35581 84071 35615
rect 84013 35575 84071 35581
rect 84289 35615 84347 35621
rect 84289 35581 84301 35615
rect 84335 35581 84347 35615
rect 84289 35575 84347 35581
rect 84028 35544 84056 35575
rect 84378 35572 84384 35624
rect 84436 35612 84442 35624
rect 85592 35621 85620 35788
rect 86037 35785 86049 35788
rect 86083 35816 86095 35819
rect 86494 35816 86500 35828
rect 86083 35788 86500 35816
rect 86083 35785 86095 35788
rect 86037 35779 86095 35785
rect 86494 35776 86500 35788
rect 86552 35776 86558 35828
rect 86862 35776 86868 35828
rect 86920 35816 86926 35828
rect 86957 35819 87015 35825
rect 86957 35816 86969 35819
rect 86920 35788 86969 35816
rect 86920 35776 86926 35788
rect 86957 35785 86969 35788
rect 87003 35785 87015 35819
rect 86957 35779 87015 35785
rect 85577 35615 85635 35621
rect 84436 35584 84481 35612
rect 84436 35572 84442 35584
rect 85577 35581 85589 35615
rect 85623 35581 85635 35615
rect 85577 35575 85635 35581
rect 86862 35572 86868 35624
rect 86920 35612 86926 35624
rect 87141 35615 87199 35621
rect 87141 35612 87153 35615
rect 86920 35584 87153 35612
rect 86920 35572 86926 35584
rect 87141 35581 87153 35584
rect 87187 35581 87199 35615
rect 87141 35575 87199 35581
rect 87417 35615 87475 35621
rect 87417 35581 87429 35615
rect 87463 35612 87475 35615
rect 88334 35612 88340 35624
rect 87463 35584 88340 35612
rect 87463 35581 87475 35584
rect 87417 35575 87475 35581
rect 88334 35572 88340 35584
rect 88392 35572 88398 35624
rect 85393 35547 85451 35553
rect 85393 35544 85405 35547
rect 83752 35516 84056 35544
rect 84580 35516 85405 35544
rect 50908 35448 53328 35476
rect 53377 35479 53435 35485
rect 53377 35445 53389 35479
rect 53423 35476 53435 35479
rect 53834 35476 53840 35488
rect 53423 35448 53840 35476
rect 53423 35445 53435 35448
rect 53377 35439 53435 35445
rect 53834 35436 53840 35448
rect 53892 35436 53898 35488
rect 57149 35479 57207 35485
rect 57149 35445 57161 35479
rect 57195 35476 57207 35479
rect 63681 35479 63739 35485
rect 63681 35476 63693 35479
rect 57195 35448 63693 35476
rect 57195 35445 57207 35448
rect 57149 35439 57207 35445
rect 63681 35445 63693 35448
rect 63727 35445 63739 35479
rect 63681 35439 63739 35445
rect 63770 35436 63776 35488
rect 63828 35476 63834 35488
rect 65426 35476 65432 35488
rect 63828 35448 65432 35476
rect 63828 35436 63834 35448
rect 65426 35436 65432 35448
rect 65484 35476 65490 35488
rect 66349 35479 66407 35485
rect 66349 35476 66361 35479
rect 65484 35448 66361 35476
rect 65484 35436 65490 35448
rect 66349 35445 66361 35448
rect 66395 35445 66407 35479
rect 66349 35439 66407 35445
rect 69842 35436 69848 35488
rect 69900 35476 69906 35488
rect 70854 35476 70860 35488
rect 69900 35448 70860 35476
rect 69900 35436 69906 35448
rect 70854 35436 70860 35448
rect 70912 35476 70918 35488
rect 72973 35479 73031 35485
rect 72973 35476 72985 35479
rect 70912 35448 72985 35476
rect 70912 35436 70918 35448
rect 72973 35445 72985 35448
rect 73019 35445 73031 35479
rect 72973 35439 73031 35445
rect 77018 35436 77024 35488
rect 77076 35476 77082 35488
rect 79137 35479 79195 35485
rect 79137 35476 79149 35479
rect 77076 35448 79149 35476
rect 77076 35436 77082 35448
rect 79137 35445 79149 35448
rect 79183 35476 79195 35479
rect 79229 35479 79287 35485
rect 79229 35476 79241 35479
rect 79183 35448 79241 35476
rect 79183 35445 79195 35448
rect 79137 35439 79195 35445
rect 79229 35445 79241 35448
rect 79275 35445 79287 35479
rect 79229 35439 79287 35445
rect 80146 35436 80152 35488
rect 80204 35476 80210 35488
rect 80701 35479 80759 35485
rect 80701 35476 80713 35479
rect 80204 35448 80713 35476
rect 80204 35436 80210 35448
rect 80701 35445 80713 35448
rect 80747 35476 80759 35479
rect 82633 35479 82691 35485
rect 82633 35476 82645 35479
rect 80747 35448 82645 35476
rect 80747 35445 80759 35448
rect 80701 35439 80759 35445
rect 82633 35445 82645 35448
rect 82679 35476 82691 35479
rect 82722 35476 82728 35488
rect 82679 35448 82728 35476
rect 82679 35445 82691 35448
rect 82633 35439 82691 35445
rect 82722 35436 82728 35448
rect 82780 35436 82786 35488
rect 83918 35436 83924 35488
rect 83976 35476 83982 35488
rect 84580 35476 84608 35516
rect 85393 35513 85405 35516
rect 85439 35513 85451 35547
rect 85393 35507 85451 35513
rect 83976 35448 84608 35476
rect 83976 35436 83982 35448
rect 85022 35436 85028 35488
rect 85080 35476 85086 35488
rect 85669 35479 85727 35485
rect 85669 35476 85681 35479
rect 85080 35448 85681 35476
rect 85080 35436 85086 35448
rect 85669 35445 85681 35448
rect 85715 35445 85727 35479
rect 85669 35439 85727 35445
rect 88242 35436 88248 35488
rect 88300 35476 88306 35488
rect 88521 35479 88579 35485
rect 88521 35476 88533 35479
rect 88300 35448 88533 35476
rect 88300 35436 88306 35448
rect 88521 35445 88533 35448
rect 88567 35445 88579 35479
rect 88521 35439 88579 35445
rect 1104 35386 111136 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 81046 35386
rect 81098 35334 81110 35386
rect 81162 35334 81174 35386
rect 81226 35334 81238 35386
rect 81290 35334 111136 35386
rect 1104 35312 111136 35334
rect 4706 35272 4712 35284
rect 4667 35244 4712 35272
rect 4706 35232 4712 35244
rect 4764 35232 4770 35284
rect 11517 35275 11575 35281
rect 11517 35241 11529 35275
rect 11563 35272 11575 35275
rect 12342 35272 12348 35284
rect 11563 35244 12348 35272
rect 11563 35241 11575 35244
rect 11517 35235 11575 35241
rect 9766 35204 9772 35216
rect 4724 35176 5396 35204
rect 4724 35145 4752 35176
rect 5368 35148 5396 35176
rect 6564 35176 9772 35204
rect 4709 35139 4767 35145
rect 4709 35105 4721 35139
rect 4755 35105 4767 35139
rect 4709 35099 4767 35105
rect 4985 35139 5043 35145
rect 4985 35105 4997 35139
rect 5031 35105 5043 35139
rect 4985 35099 5043 35105
rect 5000 35068 5028 35099
rect 5350 35096 5356 35148
rect 5408 35136 5414 35148
rect 6270 35136 6276 35148
rect 5408 35108 6276 35136
rect 5408 35096 5414 35108
rect 6270 35096 6276 35108
rect 6328 35096 6334 35148
rect 6564 35145 6592 35176
rect 9766 35164 9772 35176
rect 9824 35164 9830 35216
rect 11054 35204 11060 35216
rect 10244 35176 11060 35204
rect 6549 35139 6607 35145
rect 6549 35105 6561 35139
rect 6595 35105 6607 35139
rect 8294 35136 8300 35148
rect 6549 35099 6607 35105
rect 6656 35108 8300 35136
rect 6656 35068 6684 35108
rect 8294 35096 8300 35108
rect 8352 35096 8358 35148
rect 10244 35145 10272 35176
rect 11054 35164 11060 35176
rect 11112 35164 11118 35216
rect 9677 35139 9735 35145
rect 9677 35105 9689 35139
rect 9723 35105 9735 35139
rect 9677 35099 9735 35105
rect 10229 35139 10287 35145
rect 10229 35105 10241 35139
rect 10275 35105 10287 35139
rect 10229 35099 10287 35105
rect 5000 35040 6684 35068
rect 6733 35071 6791 35077
rect 6733 35037 6745 35071
rect 6779 35037 6791 35071
rect 6733 35031 6791 35037
rect 2866 34960 2872 35012
rect 2924 35000 2930 35012
rect 6748 35000 6776 35031
rect 8202 35028 8208 35080
rect 8260 35068 8266 35080
rect 9692 35068 9720 35099
rect 10318 35096 10324 35148
rect 10376 35136 10382 35148
rect 11624 35145 11652 35244
rect 12342 35232 12348 35244
rect 12400 35272 12406 35284
rect 15657 35275 15715 35281
rect 15657 35272 15669 35275
rect 12400 35244 15669 35272
rect 12400 35232 12406 35244
rect 10505 35139 10563 35145
rect 10505 35136 10517 35139
rect 10376 35108 10517 35136
rect 10376 35096 10382 35108
rect 10505 35105 10517 35108
rect 10551 35105 10563 35139
rect 10505 35099 10563 35105
rect 11609 35139 11667 35145
rect 11609 35105 11621 35139
rect 11655 35105 11667 35139
rect 11609 35099 11667 35105
rect 13817 35139 13875 35145
rect 13817 35105 13829 35139
rect 13863 35136 13875 35139
rect 14185 35139 14243 35145
rect 14185 35136 14197 35139
rect 13863 35108 14197 35136
rect 13863 35105 13875 35108
rect 13817 35099 13875 35105
rect 14185 35105 14197 35108
rect 14231 35136 14243 35139
rect 15010 35136 15016 35148
rect 14231 35108 15016 35136
rect 14231 35105 14243 35108
rect 14185 35099 14243 35105
rect 15010 35096 15016 35108
rect 15068 35096 15074 35148
rect 15304 35145 15332 35244
rect 15657 35241 15669 35244
rect 15703 35241 15715 35275
rect 15657 35235 15715 35241
rect 21085 35275 21143 35281
rect 21085 35241 21097 35275
rect 21131 35272 21143 35275
rect 21358 35272 21364 35284
rect 21131 35244 21364 35272
rect 21131 35241 21143 35244
rect 21085 35235 21143 35241
rect 21358 35232 21364 35244
rect 21416 35232 21422 35284
rect 22741 35275 22799 35281
rect 22741 35241 22753 35275
rect 22787 35272 22799 35275
rect 32766 35272 32772 35284
rect 22787 35244 26280 35272
rect 22787 35241 22799 35244
rect 22741 35235 22799 35241
rect 22462 35204 22468 35216
rect 15396 35176 22468 35204
rect 15289 35139 15347 35145
rect 15289 35105 15301 35139
rect 15335 35105 15347 35139
rect 15289 35099 15347 35105
rect 8260 35040 9720 35068
rect 8260 35028 8266 35040
rect 11514 35028 11520 35080
rect 11572 35068 11578 35080
rect 15396 35068 15424 35176
rect 22462 35164 22468 35176
rect 22520 35164 22526 35216
rect 26252 35213 26280 35244
rect 27264 35244 32772 35272
rect 26237 35207 26295 35213
rect 26237 35173 26249 35207
rect 26283 35204 26295 35207
rect 27264 35204 27292 35244
rect 32766 35232 32772 35244
rect 32824 35232 32830 35284
rect 41230 35272 41236 35284
rect 32968 35244 41236 35272
rect 26283 35176 27292 35204
rect 26283 35173 26295 35176
rect 26237 35167 26295 35173
rect 16390 35136 16396 35148
rect 16351 35108 16396 35136
rect 16390 35096 16396 35108
rect 16448 35136 16454 35148
rect 16761 35139 16819 35145
rect 16761 35136 16773 35139
rect 16448 35108 16773 35136
rect 16448 35096 16454 35108
rect 16761 35105 16773 35108
rect 16807 35105 16819 35139
rect 20901 35139 20959 35145
rect 20901 35136 20913 35139
rect 16761 35099 16819 35105
rect 18708 35108 20913 35136
rect 11572 35040 15424 35068
rect 11572 35028 11578 35040
rect 16482 35028 16488 35080
rect 16540 35068 16546 35080
rect 18708 35068 18736 35108
rect 20901 35105 20913 35108
rect 20947 35136 20959 35139
rect 21726 35136 21732 35148
rect 20947 35108 21732 35136
rect 20947 35105 20959 35108
rect 20901 35099 20959 35105
rect 21726 35096 21732 35108
rect 21784 35096 21790 35148
rect 21818 35096 21824 35148
rect 21876 35136 21882 35148
rect 22373 35139 22431 35145
rect 22373 35136 22385 35139
rect 21876 35108 22385 35136
rect 21876 35096 21882 35108
rect 22373 35105 22385 35108
rect 22419 35136 22431 35139
rect 22557 35139 22615 35145
rect 22557 35136 22569 35139
rect 22419 35108 22569 35136
rect 22419 35105 22431 35108
rect 22373 35099 22431 35105
rect 22557 35105 22569 35108
rect 22603 35105 22615 35139
rect 23658 35136 23664 35148
rect 23619 35108 23664 35136
rect 22557 35099 22615 35105
rect 23658 35096 23664 35108
rect 23716 35096 23722 35148
rect 25130 35096 25136 35148
rect 25188 35136 25194 35148
rect 25188 35108 26648 35136
rect 25188 35096 25194 35108
rect 16540 35040 18736 35068
rect 16540 35028 16546 35040
rect 20714 35028 20720 35080
rect 20772 35068 20778 35080
rect 22002 35068 22008 35080
rect 20772 35040 22008 35068
rect 20772 35028 20778 35040
rect 22002 35028 22008 35040
rect 22060 35068 22066 35080
rect 23753 35071 23811 35077
rect 23753 35068 23765 35071
rect 22060 35040 23765 35068
rect 22060 35028 22066 35040
rect 23753 35037 23765 35040
rect 23799 35037 23811 35071
rect 26513 35071 26571 35077
rect 26513 35068 26525 35071
rect 23753 35031 23811 35037
rect 26344 35040 26525 35068
rect 2924 34972 6776 35000
rect 2924 34960 2930 34972
rect 9122 34960 9128 35012
rect 9180 35000 9186 35012
rect 9769 35003 9827 35009
rect 9769 35000 9781 35003
rect 9180 34972 9781 35000
rect 9180 34960 9186 34972
rect 9769 34969 9781 34972
rect 9815 34969 9827 35003
rect 9769 34963 9827 34969
rect 10962 34960 10968 35012
rect 11020 35000 11026 35012
rect 11793 35003 11851 35009
rect 11793 35000 11805 35003
rect 11020 34972 11805 35000
rect 11020 34960 11026 34972
rect 11793 34969 11805 34972
rect 11839 34969 11851 35003
rect 11793 34963 11851 34969
rect 15473 35003 15531 35009
rect 15473 34969 15485 35003
rect 15519 35000 15531 35003
rect 26234 35000 26240 35012
rect 15519 34972 26240 35000
rect 15519 34969 15531 34972
rect 15473 34963 15531 34969
rect 26234 34960 26240 34972
rect 26292 34960 26298 35012
rect 13906 34932 13912 34944
rect 13867 34904 13912 34932
rect 13906 34892 13912 34904
rect 13964 34892 13970 34944
rect 16574 34932 16580 34944
rect 16535 34904 16580 34932
rect 16574 34892 16580 34904
rect 16632 34892 16638 34944
rect 25866 34892 25872 34944
rect 25924 34932 25930 34944
rect 25961 34935 26019 34941
rect 25961 34932 25973 34935
rect 25924 34904 25973 34932
rect 25924 34892 25930 34904
rect 25961 34901 25973 34904
rect 26007 34932 26019 34935
rect 26344 34932 26372 35040
rect 26513 35037 26525 35040
rect 26559 35037 26571 35071
rect 26620 35068 26648 35108
rect 26694 35096 26700 35148
rect 26752 35136 26758 35148
rect 27264 35145 27292 35176
rect 27890 35164 27896 35216
rect 27948 35204 27954 35216
rect 32861 35207 32919 35213
rect 32861 35204 32873 35207
rect 27948 35176 32873 35204
rect 27948 35164 27954 35176
rect 32861 35173 32873 35176
rect 32907 35173 32919 35207
rect 32861 35167 32919 35173
rect 27157 35139 27215 35145
rect 27157 35136 27169 35139
rect 26752 35108 26797 35136
rect 26896 35108 27169 35136
rect 26752 35096 26758 35108
rect 26896 35068 26924 35108
rect 27157 35105 27169 35108
rect 27203 35105 27215 35139
rect 27157 35099 27215 35105
rect 27249 35139 27307 35145
rect 27249 35105 27261 35139
rect 27295 35105 27307 35139
rect 27249 35099 27307 35105
rect 28166 35096 28172 35148
rect 28224 35136 28230 35148
rect 28805 35139 28863 35145
rect 28805 35136 28817 35139
rect 28224 35108 28817 35136
rect 28224 35096 28230 35108
rect 28805 35105 28817 35108
rect 28851 35105 28863 35139
rect 28805 35099 28863 35105
rect 28902 35096 28908 35148
rect 28960 35136 28966 35148
rect 30374 35136 30380 35148
rect 28960 35108 29005 35136
rect 30335 35108 30380 35136
rect 28960 35096 28966 35108
rect 30374 35096 30380 35108
rect 30432 35096 30438 35148
rect 30469 35139 30527 35145
rect 30469 35105 30481 35139
rect 30515 35136 30527 35139
rect 32968 35136 32996 35244
rect 41230 35232 41236 35244
rect 41288 35232 41294 35284
rect 41322 35232 41328 35284
rect 41380 35272 41386 35284
rect 61286 35272 61292 35284
rect 41380 35244 61292 35272
rect 41380 35232 41386 35244
rect 61286 35232 61292 35244
rect 61344 35232 61350 35284
rect 70578 35272 70584 35284
rect 61488 35244 70584 35272
rect 34793 35207 34851 35213
rect 34793 35173 34805 35207
rect 34839 35204 34851 35207
rect 39114 35204 39120 35216
rect 34839 35176 39120 35204
rect 34839 35173 34851 35176
rect 34793 35167 34851 35173
rect 39114 35164 39120 35176
rect 39172 35164 39178 35216
rect 39945 35207 40003 35213
rect 39945 35204 39957 35207
rect 39224 35176 39957 35204
rect 30515 35108 32996 35136
rect 33045 35139 33103 35145
rect 30515 35105 30527 35108
rect 30469 35099 30527 35105
rect 33045 35105 33057 35139
rect 33091 35136 33103 35139
rect 33137 35139 33195 35145
rect 33137 35136 33149 35139
rect 33091 35108 33149 35136
rect 33091 35105 33103 35108
rect 33045 35099 33103 35105
rect 33137 35105 33149 35108
rect 33183 35136 33195 35139
rect 33226 35136 33232 35148
rect 33183 35108 33232 35136
rect 33183 35105 33195 35108
rect 33137 35099 33195 35105
rect 27798 35068 27804 35080
rect 26620 35040 26924 35068
rect 27759 35040 27804 35068
rect 26513 35031 26571 35037
rect 26007 34904 26372 34932
rect 26896 34932 26924 35040
rect 27798 35028 27804 35040
rect 27856 35028 27862 35080
rect 28077 34935 28135 34941
rect 28077 34932 28089 34935
rect 26896 34904 28089 34932
rect 26007 34901 26019 34904
rect 25961 34895 26019 34901
rect 28077 34901 28089 34904
rect 28123 34932 28135 34935
rect 30484 34932 30512 35099
rect 33226 35096 33232 35108
rect 33284 35096 33290 35148
rect 33410 35136 33416 35148
rect 33371 35108 33416 35136
rect 33410 35096 33416 35108
rect 33468 35096 33474 35148
rect 39224 35145 39252 35176
rect 39945 35173 39957 35176
rect 39991 35204 40003 35207
rect 39991 35176 41092 35204
rect 39991 35173 40003 35176
rect 39945 35167 40003 35173
rect 38657 35139 38715 35145
rect 38657 35105 38669 35139
rect 38703 35105 38715 35139
rect 38657 35099 38715 35105
rect 39209 35139 39267 35145
rect 39209 35105 39221 35139
rect 39255 35105 39267 35139
rect 39390 35136 39396 35148
rect 39351 35108 39396 35136
rect 39209 35099 39267 35105
rect 38102 35028 38108 35080
rect 38160 35068 38166 35080
rect 38470 35068 38476 35080
rect 38160 35040 38476 35068
rect 38160 35028 38166 35040
rect 38470 35028 38476 35040
rect 38528 35028 38534 35080
rect 35618 34960 35624 35012
rect 35676 35000 35682 35012
rect 38562 35000 38568 35012
rect 35676 34972 38568 35000
rect 35676 34960 35682 34972
rect 38562 34960 38568 34972
rect 38620 34960 38626 35012
rect 38672 35000 38700 35099
rect 39390 35096 39396 35108
rect 39448 35136 39454 35148
rect 40880 35145 40908 35176
rect 40681 35139 40739 35145
rect 40681 35136 40693 35139
rect 39448 35108 40693 35136
rect 39448 35096 39454 35108
rect 40681 35105 40693 35108
rect 40727 35105 40739 35139
rect 40681 35099 40739 35105
rect 40865 35139 40923 35145
rect 40865 35105 40877 35139
rect 40911 35105 40923 35139
rect 40865 35099 40923 35105
rect 39758 35068 39764 35080
rect 39719 35040 39764 35068
rect 39758 35028 39764 35040
rect 39816 35028 39822 35080
rect 40218 35028 40224 35080
rect 40276 35068 40282 35080
rect 40497 35071 40555 35077
rect 40497 35068 40509 35071
rect 40276 35040 40509 35068
rect 40276 35028 40282 35040
rect 40497 35037 40509 35040
rect 40543 35068 40555 35071
rect 40954 35068 40960 35080
rect 40543 35040 40960 35068
rect 40543 35037 40555 35040
rect 40497 35031 40555 35037
rect 40954 35028 40960 35040
rect 41012 35028 41018 35080
rect 40129 35003 40187 35009
rect 40129 35000 40141 35003
rect 38672 34972 40141 35000
rect 40129 34969 40141 34972
rect 40175 35000 40187 35003
rect 40862 35000 40868 35012
rect 40175 34972 40868 35000
rect 40175 34969 40187 34972
rect 40129 34963 40187 34969
rect 40862 34960 40868 34972
rect 40920 34960 40926 35012
rect 41064 35000 41092 35176
rect 41506 35164 41512 35216
rect 41564 35204 41570 35216
rect 41966 35204 41972 35216
rect 41564 35176 41644 35204
rect 41927 35176 41972 35204
rect 41564 35164 41570 35176
rect 41230 35096 41236 35148
rect 41288 35136 41294 35148
rect 41325 35139 41383 35145
rect 41325 35136 41337 35139
rect 41288 35108 41337 35136
rect 41288 35096 41294 35108
rect 41325 35105 41337 35108
rect 41371 35105 41383 35139
rect 41325 35099 41383 35105
rect 41414 35096 41420 35148
rect 41472 35136 41478 35148
rect 41616 35136 41644 35176
rect 41966 35164 41972 35176
rect 42024 35164 42030 35216
rect 43714 35204 43720 35216
rect 42076 35176 43720 35204
rect 42076 35136 42104 35176
rect 43714 35164 43720 35176
rect 43772 35204 43778 35216
rect 49605 35207 49663 35213
rect 49605 35204 49617 35207
rect 43772 35176 49617 35204
rect 43772 35164 43778 35176
rect 49605 35173 49617 35176
rect 49651 35204 49663 35207
rect 50985 35207 51043 35213
rect 49651 35176 50384 35204
rect 49651 35173 49663 35176
rect 49605 35167 49663 35173
rect 42242 35136 42248 35148
rect 41472 35108 41517 35136
rect 41616 35108 42104 35136
rect 42203 35108 42248 35136
rect 41472 35096 41478 35108
rect 42242 35096 42248 35108
rect 42300 35096 42306 35148
rect 42429 35139 42487 35145
rect 42429 35105 42441 35139
rect 42475 35136 42487 35139
rect 49878 35136 49884 35148
rect 42475 35108 49884 35136
rect 42475 35105 42487 35108
rect 42429 35099 42487 35105
rect 42444 35000 42472 35099
rect 49878 35096 49884 35108
rect 49936 35096 49942 35148
rect 50356 35145 50384 35176
rect 50985 35173 50997 35207
rect 51031 35204 51043 35207
rect 51994 35204 52000 35216
rect 51031 35176 52000 35204
rect 51031 35173 51043 35176
rect 50985 35167 51043 35173
rect 51994 35164 52000 35176
rect 52052 35164 52058 35216
rect 53190 35204 53196 35216
rect 53151 35176 53196 35204
rect 53190 35164 53196 35176
rect 53248 35164 53254 35216
rect 56134 35204 56140 35216
rect 53576 35176 56140 35204
rect 50341 35139 50399 35145
rect 50341 35105 50353 35139
rect 50387 35105 50399 35139
rect 50341 35099 50399 35105
rect 50430 35096 50436 35148
rect 50488 35136 50494 35148
rect 50488 35108 50533 35136
rect 50488 35096 50494 35108
rect 51166 35096 51172 35148
rect 51224 35136 51230 35148
rect 51445 35139 51503 35145
rect 51445 35136 51457 35139
rect 51224 35108 51457 35136
rect 51224 35096 51230 35108
rect 51445 35105 51457 35108
rect 51491 35136 51503 35139
rect 51810 35136 51816 35148
rect 51491 35108 51816 35136
rect 51491 35105 51503 35108
rect 51445 35099 51503 35105
rect 51810 35096 51816 35108
rect 51868 35096 51874 35148
rect 52086 35136 52092 35148
rect 52047 35108 52092 35136
rect 52086 35096 52092 35108
rect 52144 35096 52150 35148
rect 52549 35139 52607 35145
rect 52549 35136 52561 35139
rect 52196 35108 52561 35136
rect 42518 35028 42524 35080
rect 42576 35068 42582 35080
rect 49418 35068 49424 35080
rect 42576 35040 49424 35068
rect 42576 35028 42582 35040
rect 49418 35028 49424 35040
rect 49476 35028 49482 35080
rect 49694 35068 49700 35080
rect 49655 35040 49700 35068
rect 49694 35028 49700 35040
rect 49752 35028 49758 35080
rect 51718 35028 51724 35080
rect 51776 35068 51782 35080
rect 51905 35071 51963 35077
rect 51905 35068 51917 35071
rect 51776 35040 51917 35068
rect 51776 35028 51782 35040
rect 51905 35037 51917 35040
rect 51951 35068 51963 35071
rect 52196 35068 52224 35108
rect 52549 35105 52561 35108
rect 52595 35105 52607 35139
rect 52549 35099 52607 35105
rect 52638 35096 52644 35148
rect 52696 35136 52702 35148
rect 53576 35145 53604 35176
rect 56134 35164 56140 35176
rect 56192 35164 56198 35216
rect 57054 35164 57060 35216
rect 57112 35204 57118 35216
rect 58342 35204 58348 35216
rect 57112 35176 58348 35204
rect 57112 35164 57118 35176
rect 58342 35164 58348 35176
rect 58400 35164 58406 35216
rect 58437 35207 58495 35213
rect 58437 35173 58449 35207
rect 58483 35204 58495 35207
rect 58483 35176 58756 35204
rect 58483 35173 58495 35176
rect 58437 35167 58495 35173
rect 58728 35148 58756 35176
rect 58802 35164 58808 35216
rect 58860 35204 58866 35216
rect 61488 35204 61516 35244
rect 70578 35232 70584 35244
rect 70636 35232 70642 35284
rect 70673 35275 70731 35281
rect 70673 35241 70685 35275
rect 70719 35272 70731 35275
rect 70854 35272 70860 35284
rect 70719 35244 70860 35272
rect 70719 35241 70731 35244
rect 70673 35235 70731 35241
rect 70854 35232 70860 35244
rect 70912 35232 70918 35284
rect 82814 35272 82820 35284
rect 72344 35244 82820 35272
rect 58860 35176 61516 35204
rect 58860 35164 58866 35176
rect 63034 35164 63040 35216
rect 63092 35204 63098 35216
rect 72344 35204 72372 35244
rect 82814 35232 82820 35244
rect 82872 35232 82878 35284
rect 82998 35272 83004 35284
rect 82959 35244 83004 35272
rect 82998 35232 83004 35244
rect 83056 35232 83062 35284
rect 83090 35232 83096 35284
rect 83148 35272 83154 35284
rect 83185 35275 83243 35281
rect 83185 35272 83197 35275
rect 83148 35244 83197 35272
rect 83148 35232 83154 35244
rect 83185 35241 83197 35244
rect 83231 35241 83243 35275
rect 83185 35235 83243 35241
rect 83274 35232 83280 35284
rect 83332 35272 83338 35284
rect 86494 35272 86500 35284
rect 83332 35244 85068 35272
rect 86455 35244 86500 35272
rect 83332 35232 83338 35244
rect 63092 35176 72372 35204
rect 72421 35207 72479 35213
rect 63092 35164 63098 35176
rect 72421 35173 72433 35207
rect 72467 35204 72479 35207
rect 72510 35204 72516 35216
rect 72467 35176 72516 35204
rect 72467 35173 72479 35176
rect 72421 35167 72479 35173
rect 72510 35164 72516 35176
rect 72568 35164 72574 35216
rect 80054 35204 80060 35216
rect 72620 35176 80060 35204
rect 53561 35139 53619 35145
rect 53561 35136 53573 35139
rect 52696 35108 53573 35136
rect 52696 35096 52702 35108
rect 53561 35105 53573 35108
rect 53607 35105 53619 35139
rect 53561 35099 53619 35105
rect 55769 35139 55827 35145
rect 55769 35105 55781 35139
rect 55815 35136 55827 35139
rect 58710 35136 58716 35148
rect 55815 35108 58572 35136
rect 58671 35108 58716 35136
rect 55815 35105 55827 35108
rect 55769 35099 55827 35105
rect 55950 35068 55956 35080
rect 51951 35040 52224 35068
rect 53392 35040 55956 35068
rect 51951 35037 51963 35040
rect 51905 35031 51963 35037
rect 41064 34972 42472 35000
rect 43346 34960 43352 35012
rect 43404 35000 43410 35012
rect 51442 35000 51448 35012
rect 43404 34972 51448 35000
rect 43404 34960 43410 34972
rect 51442 34960 51448 34972
rect 51500 34960 51506 35012
rect 28123 34904 30512 34932
rect 32861 34935 32919 34941
rect 28123 34901 28135 34904
rect 28077 34895 28135 34901
rect 32861 34901 32873 34935
rect 32907 34932 32919 34935
rect 38102 34932 38108 34944
rect 32907 34904 38108 34932
rect 32907 34901 32919 34904
rect 32861 34895 32919 34901
rect 38102 34892 38108 34904
rect 38160 34892 38166 34944
rect 38286 34932 38292 34944
rect 38247 34904 38292 34932
rect 38286 34892 38292 34904
rect 38344 34932 38350 34944
rect 39390 34932 39396 34944
rect 38344 34904 39396 34932
rect 38344 34892 38350 34904
rect 39390 34892 39396 34904
rect 39448 34932 39454 34944
rect 40313 34935 40371 34941
rect 40313 34932 40325 34935
rect 39448 34904 40325 34932
rect 39448 34892 39454 34904
rect 40313 34901 40325 34904
rect 40359 34901 40371 34935
rect 40313 34895 40371 34901
rect 40402 34892 40408 34944
rect 40460 34932 40466 34944
rect 48866 34932 48872 34944
rect 40460 34904 48872 34932
rect 40460 34892 40466 34904
rect 48866 34892 48872 34904
rect 48924 34892 48930 34944
rect 49326 34932 49332 34944
rect 49287 34904 49332 34932
rect 49326 34892 49332 34904
rect 49384 34932 49390 34944
rect 49510 34932 49516 34944
rect 49384 34904 49516 34932
rect 49384 34892 49390 34904
rect 49510 34892 49516 34904
rect 49568 34932 49574 34944
rect 49694 34932 49700 34944
rect 49568 34904 49700 34932
rect 49568 34892 49574 34904
rect 49694 34892 49700 34904
rect 49752 34892 49758 34944
rect 49878 34892 49884 34944
rect 49936 34932 49942 34944
rect 51166 34932 51172 34944
rect 49936 34904 51172 34932
rect 49936 34892 49942 34904
rect 51166 34892 51172 34904
rect 51224 34892 51230 34944
rect 51258 34892 51264 34944
rect 51316 34932 51322 34944
rect 51534 34932 51540 34944
rect 51316 34904 51361 34932
rect 51495 34904 51540 34932
rect 51316 34892 51322 34904
rect 51534 34892 51540 34904
rect 51592 34932 51598 34944
rect 51718 34932 51724 34944
rect 51592 34904 51724 34932
rect 51592 34892 51598 34904
rect 51718 34892 51724 34904
rect 51776 34892 51782 34944
rect 51810 34892 51816 34944
rect 51868 34932 51874 34944
rect 53392 34932 53420 35040
rect 55950 35028 55956 35040
rect 56008 35028 56014 35080
rect 56042 35028 56048 35080
rect 56100 35068 56106 35080
rect 56318 35068 56324 35080
rect 56100 35040 56145 35068
rect 56279 35040 56324 35068
rect 56100 35028 56106 35040
rect 56318 35028 56324 35040
rect 56376 35028 56382 35080
rect 56410 35028 56416 35080
rect 56468 35068 56474 35080
rect 58434 35068 58440 35080
rect 56468 35040 58440 35068
rect 56468 35028 56474 35040
rect 58434 35028 58440 35040
rect 58492 35028 58498 35080
rect 58544 35068 58572 35108
rect 58710 35096 58716 35108
rect 58768 35096 58774 35148
rect 62022 35136 62028 35148
rect 61983 35108 62028 35136
rect 62022 35096 62028 35108
rect 62080 35096 62086 35148
rect 64506 35136 64512 35148
rect 64467 35108 64512 35136
rect 64506 35096 64512 35108
rect 64564 35096 64570 35148
rect 65521 35139 65579 35145
rect 65521 35105 65533 35139
rect 65567 35136 65579 35139
rect 65797 35139 65855 35145
rect 65797 35136 65809 35139
rect 65567 35108 65809 35136
rect 65567 35105 65579 35108
rect 65521 35099 65579 35105
rect 65797 35105 65809 35108
rect 65843 35136 65855 35139
rect 66714 35136 66720 35148
rect 65843 35108 66720 35136
rect 65843 35105 65855 35108
rect 65797 35099 65855 35105
rect 66714 35096 66720 35108
rect 66772 35096 66778 35148
rect 68925 35139 68983 35145
rect 68925 35105 68937 35139
rect 68971 35136 68983 35139
rect 69290 35136 69296 35148
rect 68971 35108 69296 35136
rect 68971 35105 68983 35108
rect 68925 35099 68983 35105
rect 69290 35096 69296 35108
rect 69348 35096 69354 35148
rect 69842 35096 69848 35148
rect 69900 35136 69906 35148
rect 69937 35139 69995 35145
rect 69937 35136 69949 35139
rect 69900 35108 69949 35136
rect 69900 35096 69906 35108
rect 69937 35105 69949 35108
rect 69983 35105 69995 35139
rect 69937 35099 69995 35105
rect 70026 35096 70032 35148
rect 70084 35136 70090 35148
rect 70121 35139 70179 35145
rect 70121 35136 70133 35139
rect 70084 35108 70133 35136
rect 70084 35096 70090 35108
rect 70121 35105 70133 35108
rect 70167 35136 70179 35139
rect 70765 35139 70823 35145
rect 70765 35136 70777 35139
rect 70167 35108 70777 35136
rect 70167 35105 70179 35108
rect 70121 35099 70179 35105
rect 70765 35105 70777 35108
rect 70811 35136 70823 35139
rect 71406 35136 71412 35148
rect 70811 35108 71412 35136
rect 70811 35105 70823 35108
rect 70765 35099 70823 35105
rect 71406 35096 71412 35108
rect 71464 35096 71470 35148
rect 71682 35096 71688 35148
rect 71740 35136 71746 35148
rect 71869 35139 71927 35145
rect 71869 35136 71881 35139
rect 71740 35108 71881 35136
rect 71740 35096 71746 35108
rect 71869 35105 71881 35108
rect 71915 35105 71927 35139
rect 71869 35099 71927 35105
rect 71961 35139 72019 35145
rect 71961 35105 71973 35139
rect 72007 35105 72019 35139
rect 71961 35099 72019 35105
rect 59630 35068 59636 35080
rect 58544 35040 59636 35068
rect 53466 34960 53472 35012
rect 53524 35000 53530 35012
rect 58544 35009 58572 35040
rect 59630 35028 59636 35040
rect 59688 35028 59694 35080
rect 62298 35028 62304 35080
rect 62356 35068 62362 35080
rect 69860 35068 69888 35096
rect 62356 35040 62401 35068
rect 63328 35040 69888 35068
rect 70489 35071 70547 35077
rect 62356 35028 62362 35040
rect 58529 35003 58587 35009
rect 53524 34972 55720 35000
rect 53524 34960 53530 34972
rect 55582 34932 55588 34944
rect 51868 34904 53420 34932
rect 55543 34904 55588 34932
rect 51868 34892 51874 34904
rect 55582 34892 55588 34904
rect 55640 34892 55646 34944
rect 55692 34932 55720 34972
rect 56980 34972 57560 35000
rect 56980 34932 57008 34972
rect 57422 34932 57428 34944
rect 55692 34904 57008 34932
rect 57383 34904 57428 34932
rect 57422 34892 57428 34904
rect 57480 34892 57486 34944
rect 57532 34932 57560 34972
rect 58529 34969 58541 35003
rect 58575 34969 58587 35003
rect 62022 35000 62028 35012
rect 58529 34963 58587 34969
rect 58636 34972 62028 35000
rect 58636 34932 58664 34972
rect 62022 34960 62028 34972
rect 62080 34960 62086 35012
rect 58802 34932 58808 34944
rect 57532 34904 58664 34932
rect 58763 34904 58808 34932
rect 58802 34892 58808 34904
rect 58860 34892 58866 34944
rect 58894 34892 58900 34944
rect 58952 34932 58958 34944
rect 58989 34935 59047 34941
rect 58989 34932 59001 34935
rect 58952 34904 59001 34932
rect 58952 34892 58958 34904
rect 58989 34901 59001 34904
rect 59035 34901 59047 34935
rect 58989 34895 59047 34901
rect 59078 34892 59084 34944
rect 59136 34932 59142 34944
rect 59173 34935 59231 34941
rect 59173 34932 59185 34935
rect 59136 34904 59185 34932
rect 59136 34892 59142 34904
rect 59173 34901 59185 34904
rect 59219 34901 59231 34935
rect 59173 34895 59231 34901
rect 59449 34935 59507 34941
rect 59449 34901 59461 34935
rect 59495 34932 59507 34935
rect 59722 34932 59728 34944
rect 59495 34904 59728 34932
rect 59495 34901 59507 34904
rect 59449 34895 59507 34901
rect 59722 34892 59728 34904
rect 59780 34892 59786 34944
rect 61286 34892 61292 34944
rect 61344 34932 61350 34944
rect 63328 34932 63356 35040
rect 70489 35037 70501 35071
rect 70535 35037 70547 35071
rect 70489 35031 70547 35037
rect 63589 35003 63647 35009
rect 63589 34969 63601 35003
rect 63635 35000 63647 35003
rect 65521 35003 65579 35009
rect 65521 35000 65533 35003
rect 63635 34972 65533 35000
rect 63635 34969 63647 34972
rect 63589 34963 63647 34969
rect 65521 34969 65533 34972
rect 65567 34969 65579 35003
rect 65521 34963 65579 34969
rect 69017 35003 69075 35009
rect 69017 34969 69029 35003
rect 69063 35000 69075 35003
rect 69106 35000 69112 35012
rect 69063 34972 69112 35000
rect 69063 34969 69075 34972
rect 69017 34963 69075 34969
rect 69106 34960 69112 34972
rect 69164 34960 69170 35012
rect 64598 34932 64604 34944
rect 61344 34904 63356 34932
rect 64559 34904 64604 34932
rect 61344 34892 61350 34904
rect 64598 34892 64604 34904
rect 64656 34892 64662 34944
rect 64690 34892 64696 34944
rect 64748 34932 64754 34944
rect 65889 34935 65947 34941
rect 65889 34932 65901 34935
rect 64748 34904 65901 34932
rect 64748 34892 64754 34904
rect 65889 34901 65901 34904
rect 65935 34932 65947 34935
rect 66254 34932 66260 34944
rect 65935 34904 66260 34932
rect 65935 34901 65947 34904
rect 65889 34895 65947 34901
rect 66254 34892 66260 34904
rect 66312 34892 66318 34944
rect 70504 34932 70532 35031
rect 71590 35028 71596 35080
rect 71648 35068 71654 35080
rect 71976 35068 72004 35099
rect 72234 35096 72240 35148
rect 72292 35136 72298 35148
rect 72620 35136 72648 35176
rect 80054 35164 80060 35176
rect 80112 35164 80118 35216
rect 80238 35204 80244 35216
rect 80199 35176 80244 35204
rect 80238 35164 80244 35176
rect 80296 35164 80302 35216
rect 83016 35204 83044 35232
rect 83369 35207 83427 35213
rect 83369 35204 83381 35207
rect 83016 35176 83381 35204
rect 83369 35173 83381 35176
rect 83415 35204 83427 35207
rect 84378 35204 84384 35216
rect 83415 35176 84384 35204
rect 83415 35173 83427 35176
rect 83369 35167 83427 35173
rect 84378 35164 84384 35176
rect 84436 35164 84442 35216
rect 84930 35204 84936 35216
rect 84891 35176 84936 35204
rect 84930 35164 84936 35176
rect 84988 35164 84994 35216
rect 85040 35204 85068 35244
rect 86494 35232 86500 35244
rect 86552 35232 86558 35284
rect 88337 35207 88395 35213
rect 88337 35204 88349 35207
rect 85040 35176 88349 35204
rect 88337 35173 88349 35176
rect 88383 35173 88395 35207
rect 88337 35167 88395 35173
rect 72292 35108 72648 35136
rect 75917 35139 75975 35145
rect 72292 35096 72298 35108
rect 75917 35105 75929 35139
rect 75963 35105 75975 35139
rect 77018 35136 77024 35148
rect 76979 35108 77024 35136
rect 75917 35099 75975 35105
rect 71648 35040 72004 35068
rect 71648 35028 71654 35040
rect 72142 35028 72148 35080
rect 72200 35068 72206 35080
rect 75932 35068 75960 35099
rect 77018 35096 77024 35108
rect 77076 35136 77082 35148
rect 77389 35139 77447 35145
rect 77389 35136 77401 35139
rect 77076 35108 77401 35136
rect 77076 35096 77082 35108
rect 77389 35105 77401 35108
rect 77435 35105 77447 35139
rect 78582 35136 78588 35148
rect 78543 35108 78588 35136
rect 77389 35099 77447 35105
rect 78582 35096 78588 35108
rect 78640 35096 78646 35148
rect 78950 35096 78956 35148
rect 79008 35136 79014 35148
rect 79045 35139 79103 35145
rect 79045 35136 79057 35139
rect 79008 35108 79057 35136
rect 79008 35096 79014 35108
rect 79045 35105 79057 35108
rect 79091 35105 79103 35139
rect 80146 35136 80152 35148
rect 80107 35108 80152 35136
rect 79045 35099 79103 35105
rect 80146 35096 80152 35108
rect 80204 35096 80210 35148
rect 80333 35139 80391 35145
rect 80333 35105 80345 35139
rect 80379 35105 80391 35139
rect 80333 35099 80391 35105
rect 76193 35071 76251 35077
rect 76193 35068 76205 35071
rect 72200 35040 76205 35068
rect 72200 35028 72206 35040
rect 76193 35037 76205 35040
rect 76239 35068 76251 35071
rect 77754 35068 77760 35080
rect 76239 35040 77760 35068
rect 76239 35037 76251 35040
rect 76193 35031 76251 35037
rect 77754 35028 77760 35040
rect 77812 35028 77818 35080
rect 78861 35071 78919 35077
rect 78861 35037 78873 35071
rect 78907 35068 78919 35071
rect 80348 35068 80376 35099
rect 83090 35096 83096 35148
rect 83148 35136 83154 35148
rect 83553 35139 83611 35145
rect 83553 35136 83565 35139
rect 83148 35108 83565 35136
rect 83148 35096 83154 35108
rect 83553 35105 83565 35108
rect 83599 35105 83611 35139
rect 84746 35136 84752 35148
rect 84707 35108 84752 35136
rect 83553 35099 83611 35105
rect 84746 35096 84752 35108
rect 84804 35096 84810 35148
rect 85022 35136 85028 35148
rect 84983 35108 85028 35136
rect 85022 35096 85028 35108
rect 85080 35096 85086 35148
rect 86313 35139 86371 35145
rect 86313 35136 86325 35139
rect 85224 35108 86325 35136
rect 78907 35040 80376 35068
rect 78907 35037 78919 35040
rect 78861 35031 78919 35037
rect 82170 35028 82176 35080
rect 82228 35068 82234 35080
rect 85224 35068 85252 35108
rect 86313 35105 86325 35108
rect 86359 35136 86371 35139
rect 86862 35136 86868 35148
rect 86359 35108 86868 35136
rect 86359 35105 86371 35108
rect 86313 35099 86371 35105
rect 86862 35096 86868 35108
rect 86920 35096 86926 35148
rect 86957 35139 87015 35145
rect 86957 35105 86969 35139
rect 87003 35136 87015 35139
rect 87322 35136 87328 35148
rect 87003 35108 87328 35136
rect 87003 35105 87015 35108
rect 86957 35099 87015 35105
rect 87322 35096 87328 35108
rect 87380 35096 87386 35148
rect 88242 35136 88248 35148
rect 88203 35108 88248 35136
rect 88242 35096 88248 35108
rect 88300 35096 88306 35148
rect 85482 35068 85488 35080
rect 82228 35040 85252 35068
rect 85443 35040 85488 35068
rect 82228 35028 82234 35040
rect 85482 35028 85488 35040
rect 85540 35028 85546 35080
rect 87141 35071 87199 35077
rect 87141 35037 87153 35071
rect 87187 35068 87199 35071
rect 87230 35068 87236 35080
rect 87187 35040 87236 35068
rect 87187 35037 87199 35040
rect 87141 35031 87199 35037
rect 87230 35028 87236 35040
rect 87288 35028 87294 35080
rect 78309 35003 78367 35009
rect 78309 35000 78321 35003
rect 76024 34972 78321 35000
rect 76024 34944 76052 34972
rect 78309 34969 78321 34972
rect 78355 35000 78367 35003
rect 78674 35000 78680 35012
rect 78355 34972 78680 35000
rect 78355 34969 78367 34972
rect 78309 34963 78367 34969
rect 78674 34960 78680 34972
rect 78732 34960 78738 35012
rect 84194 34960 84200 35012
rect 84252 35000 84258 35012
rect 88242 35000 88248 35012
rect 84252 34972 88248 35000
rect 84252 34960 84258 34972
rect 88242 34960 88248 34972
rect 88300 34960 88306 35012
rect 71590 34932 71596 34944
rect 70504 34904 71596 34932
rect 71590 34892 71596 34904
rect 71648 34892 71654 34944
rect 71685 34935 71743 34941
rect 71685 34901 71697 34935
rect 71731 34932 71743 34935
rect 71866 34932 71872 34944
rect 71731 34904 71872 34932
rect 71731 34901 71743 34904
rect 71685 34895 71743 34901
rect 71866 34892 71872 34904
rect 71924 34892 71930 34944
rect 76006 34932 76012 34944
rect 75967 34904 76012 34932
rect 76006 34892 76012 34904
rect 76064 34892 76070 34944
rect 77202 34932 77208 34944
rect 77163 34904 77208 34932
rect 77202 34892 77208 34904
rect 77260 34892 77266 34944
rect 80514 34932 80520 34944
rect 80475 34904 80520 34932
rect 80514 34892 80520 34904
rect 80572 34892 80578 34944
rect 83274 34892 83280 34944
rect 83332 34932 83338 34944
rect 83645 34935 83703 34941
rect 83645 34932 83657 34935
rect 83332 34904 83657 34932
rect 83332 34892 83338 34904
rect 83645 34901 83657 34904
rect 83691 34901 83703 34935
rect 85942 34932 85948 34944
rect 85903 34904 85948 34932
rect 83645 34895 83703 34901
rect 85942 34892 85948 34904
rect 86000 34892 86006 34944
rect 86126 34932 86132 34944
rect 86087 34904 86132 34932
rect 86126 34892 86132 34904
rect 86184 34892 86190 34944
rect 86678 34932 86684 34944
rect 86639 34904 86684 34932
rect 86678 34892 86684 34904
rect 86736 34892 86742 34944
rect 87325 34935 87383 34941
rect 87325 34901 87337 34935
rect 87371 34932 87383 34935
rect 87506 34932 87512 34944
rect 87371 34904 87512 34932
rect 87371 34901 87383 34904
rect 87325 34895 87383 34901
rect 87506 34892 87512 34904
rect 87564 34892 87570 34944
rect 1104 34842 111136 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 65686 34842
rect 65738 34790 65750 34842
rect 65802 34790 65814 34842
rect 65866 34790 65878 34842
rect 65930 34790 96406 34842
rect 96458 34790 96470 34842
rect 96522 34790 96534 34842
rect 96586 34790 96598 34842
rect 96650 34790 111136 34842
rect 1104 34768 111136 34790
rect 9401 34731 9459 34737
rect 9401 34697 9413 34731
rect 9447 34728 9459 34731
rect 11885 34731 11943 34737
rect 9447 34700 10640 34728
rect 9447 34697 9459 34700
rect 9401 34691 9459 34697
rect 10612 34672 10640 34700
rect 11885 34697 11897 34731
rect 11931 34728 11943 34731
rect 25130 34728 25136 34740
rect 11931 34700 25136 34728
rect 11931 34697 11943 34700
rect 11885 34691 11943 34697
rect 10410 34660 10416 34672
rect 6748 34632 10416 34660
rect 2869 34595 2927 34601
rect 2869 34561 2881 34595
rect 2915 34592 2927 34595
rect 4982 34592 4988 34604
rect 2915 34564 4988 34592
rect 2915 34561 2927 34564
rect 2869 34555 2927 34561
rect 4982 34552 4988 34564
rect 5040 34552 5046 34604
rect 5626 34592 5632 34604
rect 5587 34564 5632 34592
rect 5626 34552 5632 34564
rect 5684 34552 5690 34604
rect 2593 34527 2651 34533
rect 2593 34493 2605 34527
rect 2639 34524 2651 34527
rect 3694 34524 3700 34536
rect 2639 34496 3700 34524
rect 2639 34493 2651 34496
rect 2593 34487 2651 34493
rect 3694 34484 3700 34496
rect 3752 34524 3758 34536
rect 4433 34527 4491 34533
rect 4433 34524 4445 34527
rect 3752 34496 4445 34524
rect 3752 34484 3758 34496
rect 4433 34493 4445 34496
rect 4479 34524 4491 34527
rect 4798 34524 4804 34536
rect 4479 34496 4804 34524
rect 4479 34493 4491 34496
rect 4433 34487 4491 34493
rect 4798 34484 4804 34496
rect 4856 34484 4862 34536
rect 5350 34524 5356 34536
rect 5311 34496 5356 34524
rect 5350 34484 5356 34496
rect 5408 34484 5414 34536
rect 5537 34527 5595 34533
rect 5537 34493 5549 34527
rect 5583 34524 5595 34527
rect 6748 34524 6776 34632
rect 10410 34620 10416 34632
rect 10468 34620 10474 34672
rect 10594 34620 10600 34672
rect 10652 34660 10658 34672
rect 11900 34660 11928 34691
rect 25130 34688 25136 34700
rect 25188 34688 25194 34740
rect 25498 34728 25504 34740
rect 25459 34700 25504 34728
rect 25498 34688 25504 34700
rect 25556 34728 25562 34740
rect 25866 34728 25872 34740
rect 25556 34700 25872 34728
rect 25556 34688 25562 34700
rect 25866 34688 25872 34700
rect 25924 34688 25930 34740
rect 28920 34700 30236 34728
rect 10652 34632 11008 34660
rect 10652 34620 10658 34632
rect 9677 34595 9735 34601
rect 9677 34592 9689 34595
rect 9232 34564 9689 34592
rect 9232 34533 9260 34564
rect 9677 34561 9689 34564
rect 9723 34592 9735 34595
rect 9858 34592 9864 34604
rect 9723 34564 9864 34592
rect 9723 34561 9735 34564
rect 9677 34555 9735 34561
rect 9858 34552 9864 34564
rect 9916 34592 9922 34604
rect 9916 34564 10916 34592
rect 9916 34552 9922 34564
rect 5583 34496 6776 34524
rect 9217 34527 9275 34533
rect 5583 34493 5595 34496
rect 5537 34487 5595 34493
rect 9217 34493 9229 34527
rect 9263 34493 9275 34527
rect 9217 34487 9275 34493
rect 9398 34484 9404 34536
rect 9456 34524 9462 34536
rect 10321 34527 10379 34533
rect 10321 34524 10333 34527
rect 9456 34496 10333 34524
rect 9456 34484 9462 34496
rect 10321 34493 10333 34496
rect 10367 34493 10379 34527
rect 10321 34487 10379 34493
rect 10888 34456 10916 34564
rect 10980 34533 11008 34632
rect 11072 34632 11928 34660
rect 15565 34663 15623 34669
rect 11072 34601 11100 34632
rect 15565 34629 15577 34663
rect 15611 34660 15623 34663
rect 15746 34660 15752 34672
rect 15611 34632 15752 34660
rect 15611 34629 15623 34632
rect 15565 34623 15623 34629
rect 15746 34620 15752 34632
rect 15804 34620 15810 34672
rect 22373 34663 22431 34669
rect 17236 34632 22324 34660
rect 11057 34595 11115 34601
rect 11057 34561 11069 34595
rect 11103 34561 11115 34595
rect 11701 34595 11759 34601
rect 11701 34592 11713 34595
rect 11057 34555 11115 34561
rect 11532 34564 11713 34592
rect 10965 34527 11023 34533
rect 10965 34493 10977 34527
rect 11011 34493 11023 34527
rect 10965 34487 11023 34493
rect 11146 34484 11152 34536
rect 11204 34524 11210 34536
rect 11532 34533 11560 34564
rect 11701 34561 11713 34564
rect 11747 34592 11759 34595
rect 17236 34592 17264 34632
rect 11747 34564 17264 34592
rect 22296 34592 22324 34632
rect 22373 34629 22385 34663
rect 22419 34660 22431 34663
rect 25225 34663 25283 34669
rect 25225 34660 25237 34663
rect 22419 34632 25237 34660
rect 22419 34629 22431 34632
rect 22373 34623 22431 34629
rect 25225 34629 25237 34632
rect 25271 34660 25283 34663
rect 26418 34660 26424 34672
rect 25271 34632 26424 34660
rect 25271 34629 25283 34632
rect 25225 34623 25283 34629
rect 26418 34620 26424 34632
rect 26476 34620 26482 34672
rect 26970 34620 26976 34672
rect 27028 34660 27034 34672
rect 28920 34660 28948 34700
rect 27028 34632 28948 34660
rect 30208 34660 30236 34700
rect 30374 34688 30380 34740
rect 30432 34728 30438 34740
rect 30653 34731 30711 34737
rect 30653 34728 30665 34731
rect 30432 34700 30665 34728
rect 30432 34688 30438 34700
rect 30653 34697 30665 34700
rect 30699 34697 30711 34731
rect 30653 34691 30711 34697
rect 30742 34688 30748 34740
rect 30800 34728 30806 34740
rect 37826 34728 37832 34740
rect 30800 34700 37832 34728
rect 30800 34688 30806 34700
rect 37826 34688 37832 34700
rect 37884 34688 37890 34740
rect 38562 34688 38568 34740
rect 38620 34728 38626 34740
rect 39298 34728 39304 34740
rect 38620 34700 39304 34728
rect 38620 34688 38626 34700
rect 39298 34688 39304 34700
rect 39356 34688 39362 34740
rect 39393 34731 39451 34737
rect 39393 34697 39405 34731
rect 39439 34728 39451 34731
rect 42702 34728 42708 34740
rect 39439 34700 42708 34728
rect 39439 34697 39451 34700
rect 39393 34691 39451 34697
rect 42702 34688 42708 34700
rect 42760 34688 42766 34740
rect 43622 34728 43628 34740
rect 43583 34700 43628 34728
rect 43622 34688 43628 34700
rect 43680 34688 43686 34740
rect 46750 34688 46756 34740
rect 46808 34728 46814 34740
rect 46845 34731 46903 34737
rect 46845 34728 46857 34731
rect 46808 34700 46857 34728
rect 46808 34688 46814 34700
rect 46845 34697 46857 34700
rect 46891 34697 46903 34731
rect 48406 34728 48412 34740
rect 48367 34700 48412 34728
rect 46845 34691 46903 34697
rect 48406 34688 48412 34700
rect 48464 34688 48470 34740
rect 48866 34688 48872 34740
rect 48924 34728 48930 34740
rect 48924 34700 49924 34728
rect 48924 34688 48930 34700
rect 38013 34663 38071 34669
rect 38013 34660 38025 34663
rect 30208 34632 38025 34660
rect 27028 34620 27034 34632
rect 38013 34629 38025 34632
rect 38059 34660 38071 34663
rect 38378 34660 38384 34672
rect 38059 34632 38240 34660
rect 38059 34629 38071 34632
rect 38013 34623 38071 34629
rect 22296 34564 26004 34592
rect 11747 34561 11759 34564
rect 11701 34555 11759 34561
rect 11333 34527 11391 34533
rect 11333 34524 11345 34527
rect 11204 34496 11345 34524
rect 11204 34484 11210 34496
rect 11333 34493 11345 34496
rect 11379 34493 11391 34527
rect 11333 34487 11391 34493
rect 11517 34527 11575 34533
rect 11517 34493 11529 34527
rect 11563 34493 11575 34527
rect 11517 34487 11575 34493
rect 11624 34496 13216 34524
rect 11624 34456 11652 34496
rect 10888 34428 11652 34456
rect 13188 34456 13216 34496
rect 13446 34484 13452 34536
rect 13504 34524 13510 34536
rect 13817 34527 13875 34533
rect 13817 34524 13829 34527
rect 13504 34496 13829 34524
rect 13504 34484 13510 34496
rect 13817 34493 13829 34496
rect 13863 34524 13875 34527
rect 14001 34527 14059 34533
rect 14001 34524 14013 34527
rect 13863 34496 14013 34524
rect 13863 34493 13875 34496
rect 13817 34487 13875 34493
rect 14001 34493 14013 34496
rect 14047 34493 14059 34527
rect 14274 34524 14280 34536
rect 14235 34496 14280 34524
rect 14001 34487 14059 34493
rect 14274 34484 14280 34496
rect 14332 34484 14338 34536
rect 19889 34527 19947 34533
rect 19889 34493 19901 34527
rect 19935 34524 19947 34527
rect 19978 34524 19984 34536
rect 19935 34496 19984 34524
rect 19935 34493 19947 34496
rect 19889 34487 19947 34493
rect 19978 34484 19984 34496
rect 20036 34484 20042 34536
rect 20165 34527 20223 34533
rect 20165 34493 20177 34527
rect 20211 34493 20223 34527
rect 20622 34524 20628 34536
rect 20583 34496 20628 34524
rect 20165 34487 20223 34493
rect 20180 34456 20208 34487
rect 20622 34484 20628 34496
rect 20680 34484 20686 34536
rect 20717 34527 20775 34533
rect 20717 34493 20729 34527
rect 20763 34524 20775 34527
rect 21358 34524 21364 34536
rect 20763 34496 21364 34524
rect 20763 34493 20775 34496
rect 20717 34487 20775 34493
rect 20732 34456 20760 34487
rect 21358 34484 21364 34496
rect 21416 34484 21422 34536
rect 21726 34484 21732 34536
rect 21784 34524 21790 34536
rect 22189 34527 22247 34533
rect 22189 34524 22201 34527
rect 21784 34496 22201 34524
rect 21784 34484 21790 34496
rect 22189 34493 22201 34496
rect 22235 34493 22247 34527
rect 25731 34527 25789 34533
rect 25731 34524 25743 34527
rect 22189 34487 22247 34493
rect 25056 34496 25743 34524
rect 21266 34456 21272 34468
rect 13188 34428 13860 34456
rect 20180 34428 20760 34456
rect 21227 34428 21272 34456
rect 3970 34388 3976 34400
rect 3931 34360 3976 34388
rect 3970 34348 3976 34360
rect 4028 34348 4034 34400
rect 13832 34388 13860 34428
rect 21266 34416 21272 34428
rect 21324 34416 21330 34468
rect 14550 34388 14556 34400
rect 13832 34360 14556 34388
rect 14550 34348 14556 34360
rect 14608 34348 14614 34400
rect 19334 34348 19340 34400
rect 19392 34388 19398 34400
rect 20254 34388 20260 34400
rect 19392 34360 20260 34388
rect 19392 34348 19398 34360
rect 20254 34348 20260 34360
rect 20312 34388 20318 34400
rect 21818 34388 21824 34400
rect 20312 34360 21824 34388
rect 20312 34348 20318 34360
rect 21818 34348 21824 34360
rect 21876 34348 21882 34400
rect 24670 34348 24676 34400
rect 24728 34388 24734 34400
rect 25056 34397 25084 34496
rect 25731 34493 25743 34496
rect 25777 34493 25789 34527
rect 25866 34524 25872 34536
rect 25827 34496 25872 34524
rect 25731 34487 25789 34493
rect 25866 34484 25872 34496
rect 25924 34484 25930 34536
rect 25976 34524 26004 34564
rect 27338 34552 27344 34604
rect 27396 34592 27402 34604
rect 30742 34592 30748 34604
rect 27396 34564 30748 34592
rect 27396 34552 27402 34564
rect 30742 34552 30748 34564
rect 30800 34552 30806 34604
rect 30834 34552 30840 34604
rect 30892 34592 30898 34604
rect 38212 34601 38240 34632
rect 38304 34632 38384 34660
rect 38197 34595 38255 34601
rect 30892 34564 38148 34592
rect 30892 34552 30898 34564
rect 26237 34527 26295 34533
rect 26237 34524 26249 34527
rect 25976 34496 26249 34524
rect 26237 34493 26249 34496
rect 26283 34493 26295 34527
rect 26237 34487 26295 34493
rect 26329 34527 26387 34533
rect 26329 34493 26341 34527
rect 26375 34524 26387 34527
rect 26418 34524 26424 34536
rect 26375 34496 26424 34524
rect 26375 34493 26387 34496
rect 26329 34487 26387 34493
rect 26252 34456 26280 34487
rect 26418 34484 26424 34496
rect 26476 34524 26482 34536
rect 26476 34496 29132 34524
rect 26476 34484 26482 34496
rect 27065 34459 27123 34465
rect 27065 34456 27077 34459
rect 26252 34428 27077 34456
rect 27065 34425 27077 34428
rect 27111 34456 27123 34459
rect 28902 34456 28908 34468
rect 27111 34428 28908 34456
rect 27111 34425 27123 34428
rect 27065 34419 27123 34425
rect 28902 34416 28908 34428
rect 28960 34416 28966 34468
rect 25041 34391 25099 34397
rect 25041 34388 25053 34391
rect 24728 34360 25053 34388
rect 24728 34348 24734 34360
rect 25041 34357 25053 34360
rect 25087 34357 25099 34391
rect 26786 34388 26792 34400
rect 26747 34360 26792 34388
rect 25041 34351 25099 34357
rect 26786 34348 26792 34360
rect 26844 34348 26850 34400
rect 29104 34388 29132 34496
rect 29178 34484 29184 34536
rect 29236 34524 29242 34536
rect 29280 34527 29338 34533
rect 29280 34524 29292 34527
rect 29236 34496 29292 34524
rect 29236 34484 29242 34496
rect 29280 34493 29292 34496
rect 29326 34493 29338 34527
rect 29546 34524 29552 34536
rect 29507 34496 29552 34524
rect 29280 34487 29338 34493
rect 29546 34484 29552 34496
rect 29604 34484 29610 34536
rect 34146 34524 34152 34536
rect 30208 34496 34152 34524
rect 30208 34388 30236 34496
rect 34146 34484 34152 34496
rect 34204 34484 34210 34536
rect 38120 34524 38148 34564
rect 38197 34561 38209 34595
rect 38243 34561 38255 34595
rect 38197 34555 38255 34561
rect 38304 34524 38332 34632
rect 38378 34620 38384 34632
rect 38436 34620 38442 34672
rect 39945 34663 40003 34669
rect 39945 34660 39957 34663
rect 38488 34632 39957 34660
rect 38120 34496 38332 34524
rect 38381 34527 38439 34533
rect 38381 34493 38393 34527
rect 38427 34524 38439 34527
rect 38488 34524 38516 34632
rect 39945 34629 39957 34632
rect 39991 34660 40003 34663
rect 40402 34660 40408 34672
rect 39991 34632 40408 34660
rect 39991 34629 40003 34632
rect 39945 34623 40003 34629
rect 40402 34620 40408 34632
rect 40460 34620 40466 34672
rect 49786 34660 49792 34672
rect 40512 34632 49792 34660
rect 39390 34552 39396 34604
rect 39448 34592 39454 34604
rect 40512 34592 40540 34632
rect 49786 34620 49792 34632
rect 49844 34620 49850 34672
rect 49896 34660 49924 34700
rect 50246 34688 50252 34740
rect 50304 34728 50310 34740
rect 50304 34700 50349 34728
rect 50304 34688 50310 34700
rect 52086 34688 52092 34740
rect 52144 34728 52150 34740
rect 53190 34728 53196 34740
rect 52144 34700 53196 34728
rect 52144 34688 52150 34700
rect 53190 34688 53196 34700
rect 53248 34688 53254 34740
rect 56137 34731 56195 34737
rect 53583 34700 54524 34728
rect 50433 34663 50491 34669
rect 50433 34660 50445 34663
rect 49896 34632 50445 34660
rect 50433 34629 50445 34632
rect 50479 34660 50491 34663
rect 50479 34632 51028 34660
rect 50479 34629 50491 34632
rect 50433 34623 50491 34629
rect 46658 34592 46664 34604
rect 39448 34564 40540 34592
rect 42444 34564 42748 34592
rect 46619 34564 46664 34592
rect 39448 34552 39454 34564
rect 38427 34496 38516 34524
rect 38427 34493 38439 34496
rect 38381 34487 38439 34493
rect 38562 34484 38568 34536
rect 38620 34524 38626 34536
rect 38841 34527 38899 34533
rect 38841 34524 38853 34527
rect 38620 34496 38853 34524
rect 38620 34484 38626 34496
rect 38841 34493 38853 34496
rect 38887 34493 38899 34527
rect 38841 34487 38899 34493
rect 38933 34527 38991 34533
rect 38933 34493 38945 34527
rect 38979 34524 38991 34527
rect 39761 34527 39819 34533
rect 39761 34524 39773 34527
rect 38979 34496 39773 34524
rect 38979 34493 38991 34496
rect 38933 34487 38991 34493
rect 39761 34493 39773 34496
rect 39807 34524 39819 34527
rect 39942 34524 39948 34536
rect 39807 34496 39948 34524
rect 39807 34493 39819 34496
rect 39761 34487 39819 34493
rect 39942 34484 39948 34496
rect 40000 34484 40006 34536
rect 42058 34524 42064 34536
rect 42019 34496 42064 34524
rect 42058 34484 42064 34496
rect 42116 34524 42122 34536
rect 42444 34533 42472 34564
rect 42245 34527 42303 34533
rect 42245 34524 42257 34527
rect 42116 34496 42257 34524
rect 42116 34484 42122 34496
rect 42245 34493 42257 34496
rect 42291 34524 42303 34527
rect 42429 34527 42487 34533
rect 42429 34524 42441 34527
rect 42291 34496 42441 34524
rect 42291 34493 42303 34496
rect 42245 34487 42303 34493
rect 42429 34493 42441 34496
rect 42475 34493 42487 34527
rect 42429 34487 42487 34493
rect 42613 34527 42671 34533
rect 42613 34493 42625 34527
rect 42659 34493 42671 34527
rect 42720 34524 42748 34564
rect 46658 34552 46664 34564
rect 46716 34592 46722 34604
rect 48958 34592 48964 34604
rect 46716 34564 47072 34592
rect 46716 34552 46722 34564
rect 47044 34533 47072 34564
rect 47136 34564 48964 34592
rect 43073 34527 43131 34533
rect 43073 34524 43085 34527
rect 42720 34496 43085 34524
rect 42613 34487 42671 34493
rect 43073 34493 43085 34496
rect 43119 34493 43131 34527
rect 43073 34487 43131 34493
rect 43165 34527 43223 34533
rect 43165 34493 43177 34527
rect 43211 34524 43223 34527
rect 43993 34527 44051 34533
rect 43993 34524 44005 34527
rect 43211 34496 44005 34524
rect 43211 34493 43223 34496
rect 43165 34487 43223 34493
rect 43993 34493 44005 34496
rect 44039 34524 44051 34527
rect 44177 34527 44235 34533
rect 44177 34524 44189 34527
rect 44039 34496 44189 34524
rect 44039 34493 44051 34496
rect 43993 34487 44051 34493
rect 44177 34493 44189 34496
rect 44223 34524 44235 34527
rect 47029 34527 47087 34533
rect 44223 34496 46980 34524
rect 44223 34493 44235 34496
rect 44177 34487 44235 34493
rect 30282 34416 30288 34468
rect 30340 34456 30346 34468
rect 42628 34456 42656 34487
rect 43180 34456 43208 34487
rect 30340 34428 40172 34456
rect 42628 34428 43208 34456
rect 46952 34456 46980 34496
rect 47029 34493 47041 34527
rect 47075 34493 47087 34527
rect 47029 34487 47087 34493
rect 47136 34456 47164 34564
rect 48958 34552 48964 34564
rect 49016 34552 49022 34604
rect 51000 34592 51028 34632
rect 53583 34592 53611 34700
rect 54496 34660 54524 34700
rect 56137 34697 56149 34731
rect 56183 34728 56195 34731
rect 56318 34728 56324 34740
rect 56183 34700 56324 34728
rect 56183 34697 56195 34700
rect 56137 34691 56195 34697
rect 56318 34688 56324 34700
rect 56376 34688 56382 34740
rect 57422 34688 57428 34740
rect 57480 34728 57486 34740
rect 58805 34731 58863 34737
rect 58805 34728 58817 34731
rect 57480 34700 58817 34728
rect 57480 34688 57486 34700
rect 58805 34697 58817 34700
rect 58851 34697 58863 34731
rect 58805 34691 58863 34697
rect 62022 34688 62028 34740
rect 62080 34728 62086 34740
rect 71406 34728 71412 34740
rect 62080 34700 71268 34728
rect 71367 34700 71412 34728
rect 62080 34688 62086 34700
rect 61930 34660 61936 34672
rect 54496 34632 60136 34660
rect 61891 34632 61936 34660
rect 53834 34592 53840 34604
rect 51000 34564 53611 34592
rect 53795 34564 53840 34592
rect 53834 34552 53840 34564
rect 53892 34552 53898 34604
rect 56778 34592 56784 34604
rect 56739 34564 56784 34592
rect 56778 34552 56784 34564
rect 56836 34592 56842 34604
rect 56965 34595 57023 34601
rect 56965 34592 56977 34595
rect 56836 34564 56977 34592
rect 56836 34552 56842 34564
rect 56965 34561 56977 34564
rect 57011 34592 57023 34595
rect 58618 34592 58624 34604
rect 57011 34564 57560 34592
rect 58579 34564 58624 34592
rect 57011 34561 57023 34564
rect 56965 34555 57023 34561
rect 48685 34527 48743 34533
rect 48685 34524 48697 34527
rect 46952 34428 47164 34456
rect 48516 34496 48697 34524
rect 30340 34416 30346 34428
rect 29104 34360 30236 34388
rect 30374 34348 30380 34400
rect 30432 34388 30438 34400
rect 31021 34391 31079 34397
rect 31021 34388 31033 34391
rect 30432 34360 31033 34388
rect 30432 34348 30438 34360
rect 31021 34357 31033 34360
rect 31067 34357 31079 34391
rect 31021 34351 31079 34357
rect 37826 34348 37832 34400
rect 37884 34388 37890 34400
rect 38562 34388 38568 34400
rect 37884 34360 38568 34388
rect 37884 34348 37890 34360
rect 38562 34348 38568 34360
rect 38620 34348 38626 34400
rect 40144 34388 40172 34428
rect 48516 34400 48544 34496
rect 48685 34493 48697 34496
rect 48731 34493 48743 34527
rect 48866 34524 48872 34536
rect 48827 34496 48872 34524
rect 48685 34487 48743 34493
rect 48866 34484 48872 34496
rect 48924 34484 48930 34536
rect 49418 34484 49424 34536
rect 49476 34524 49482 34536
rect 49605 34527 49663 34533
rect 49476 34496 49521 34524
rect 49476 34484 49482 34496
rect 49605 34493 49617 34527
rect 49651 34493 49663 34527
rect 49605 34487 49663 34493
rect 49620 34456 49648 34487
rect 50614 34484 50620 34536
rect 50672 34484 50678 34536
rect 53561 34527 53619 34533
rect 53561 34493 53573 34527
rect 53607 34493 53619 34527
rect 53561 34487 53619 34493
rect 49436 34428 49648 34456
rect 49973 34459 50031 34465
rect 48314 34388 48320 34400
rect 40144 34360 48320 34388
rect 48314 34348 48320 34360
rect 48372 34348 48378 34400
rect 48498 34388 48504 34400
rect 48459 34360 48504 34388
rect 48498 34348 48504 34360
rect 48556 34348 48562 34400
rect 48590 34348 48596 34400
rect 48648 34388 48654 34400
rect 49436 34388 49464 34428
rect 49973 34425 49985 34459
rect 50019 34456 50031 34459
rect 50632 34456 50660 34484
rect 50019 34428 50660 34456
rect 50019 34425 50031 34428
rect 49973 34419 50031 34425
rect 48648 34360 49464 34388
rect 53576 34388 53604 34487
rect 55306 34484 55312 34536
rect 55364 34524 55370 34536
rect 56045 34527 56103 34533
rect 56045 34524 56057 34527
rect 55364 34496 56057 34524
rect 55364 34484 55370 34496
rect 56045 34493 56057 34496
rect 56091 34493 56103 34527
rect 56045 34487 56103 34493
rect 56134 34484 56140 34536
rect 56192 34524 56198 34536
rect 56594 34524 56600 34536
rect 56192 34496 56456 34524
rect 56555 34496 56600 34524
rect 56192 34484 56198 34496
rect 55401 34459 55459 34465
rect 55401 34456 55413 34459
rect 54496 34428 55413 34456
rect 53926 34388 53932 34400
rect 53576 34360 53932 34388
rect 48648 34348 48654 34360
rect 53926 34348 53932 34360
rect 53984 34388 53990 34400
rect 54496 34388 54524 34428
rect 55401 34425 55413 34428
rect 55447 34456 55459 34459
rect 55582 34456 55588 34468
rect 55447 34428 55588 34456
rect 55447 34425 55459 34428
rect 55401 34419 55459 34425
rect 55582 34416 55588 34428
rect 55640 34416 55646 34468
rect 55122 34388 55128 34400
rect 53984 34360 54524 34388
rect 55083 34360 55128 34388
rect 53984 34348 53990 34360
rect 55122 34348 55128 34360
rect 55180 34348 55186 34400
rect 56428 34388 56456 34496
rect 56594 34484 56600 34496
rect 56652 34524 56658 34536
rect 57532 34533 57560 34564
rect 58618 34552 58624 34564
rect 58676 34552 58682 34604
rect 59446 34552 59452 34604
rect 59504 34592 59510 34604
rect 60001 34595 60059 34601
rect 60001 34592 60013 34595
rect 59504 34564 60013 34592
rect 59504 34552 59510 34564
rect 60001 34561 60013 34564
rect 60047 34561 60059 34595
rect 60108 34592 60136 34632
rect 61930 34620 61936 34632
rect 61988 34660 61994 34672
rect 62574 34660 62580 34672
rect 61988 34632 62580 34660
rect 61988 34620 61994 34632
rect 62574 34620 62580 34632
rect 62632 34620 62638 34672
rect 64322 34660 64328 34672
rect 64283 34632 64328 34660
rect 64322 34620 64328 34632
rect 64380 34620 64386 34672
rect 69934 34660 69940 34672
rect 69895 34632 69940 34660
rect 69934 34620 69940 34632
rect 69992 34620 69998 34672
rect 71240 34660 71268 34700
rect 71406 34688 71412 34700
rect 71464 34728 71470 34740
rect 72329 34731 72387 34737
rect 72329 34728 72341 34731
rect 71464 34700 72341 34728
rect 71464 34688 71470 34700
rect 72329 34697 72341 34700
rect 72375 34697 72387 34731
rect 72602 34728 72608 34740
rect 72563 34700 72608 34728
rect 72329 34691 72387 34697
rect 72234 34660 72240 34672
rect 71240 34632 72240 34660
rect 72234 34620 72240 34632
rect 72292 34620 72298 34672
rect 72142 34592 72148 34604
rect 60108 34564 72148 34592
rect 60001 34555 60059 34561
rect 72142 34552 72148 34564
rect 72200 34552 72206 34604
rect 57333 34527 57391 34533
rect 57333 34524 57345 34527
rect 56652 34496 57345 34524
rect 56652 34484 56658 34496
rect 57333 34493 57345 34496
rect 57379 34493 57391 34527
rect 57333 34487 57391 34493
rect 57517 34527 57575 34533
rect 57517 34493 57529 34527
rect 57563 34524 57575 34527
rect 58069 34527 58127 34533
rect 58069 34524 58081 34527
rect 57563 34496 58081 34524
rect 57563 34493 57575 34496
rect 57517 34487 57575 34493
rect 58069 34493 58081 34496
rect 58115 34493 58127 34527
rect 58250 34524 58256 34536
rect 58211 34496 58256 34524
rect 58069 34487 58127 34493
rect 58250 34484 58256 34496
rect 58308 34524 58314 34536
rect 58986 34524 58992 34536
rect 58308 34496 58848 34524
rect 58947 34496 58992 34524
rect 58308 34484 58314 34496
rect 58820 34456 58848 34496
rect 58986 34484 58992 34496
rect 59044 34484 59050 34536
rect 59170 34524 59176 34536
rect 59131 34496 59176 34524
rect 59170 34484 59176 34496
rect 59228 34484 59234 34536
rect 59354 34524 59360 34536
rect 59315 34496 59360 34524
rect 59354 34484 59360 34496
rect 59412 34484 59418 34536
rect 59630 34484 59636 34536
rect 59688 34524 59694 34536
rect 59725 34527 59783 34533
rect 59725 34524 59737 34527
rect 59688 34496 59737 34524
rect 59688 34484 59694 34496
rect 59725 34493 59737 34496
rect 59771 34493 59783 34527
rect 61746 34524 61752 34536
rect 59725 34487 59783 34493
rect 60016 34496 61752 34524
rect 60016 34456 60044 34496
rect 61746 34484 61752 34496
rect 61804 34484 61810 34536
rect 61841 34527 61899 34533
rect 61841 34493 61853 34527
rect 61887 34524 61899 34527
rect 62942 34524 62948 34536
rect 61887 34496 62528 34524
rect 62903 34496 62948 34524
rect 61887 34493 61899 34496
rect 61841 34487 61899 34493
rect 58820 34428 60044 34456
rect 59538 34388 59544 34400
rect 56428 34360 59544 34388
rect 59538 34348 59544 34360
rect 59596 34348 59602 34400
rect 59630 34348 59636 34400
rect 59688 34388 59694 34400
rect 59817 34391 59875 34397
rect 59817 34388 59829 34391
rect 59688 34360 59829 34388
rect 59688 34348 59694 34360
rect 59817 34357 59829 34360
rect 59863 34357 59875 34391
rect 62500 34388 62528 34496
rect 62942 34484 62948 34496
rect 63000 34484 63006 34536
rect 63221 34527 63279 34533
rect 63221 34524 63233 34527
rect 63052 34496 63233 34524
rect 62666 34456 62672 34468
rect 62627 34428 62672 34456
rect 62666 34416 62672 34428
rect 62724 34456 62730 34468
rect 63052 34456 63080 34496
rect 63221 34493 63233 34496
rect 63267 34493 63279 34527
rect 64322 34524 64328 34536
rect 63221 34487 63279 34493
rect 63880 34496 64328 34524
rect 62724 34428 63080 34456
rect 62724 34416 62730 34428
rect 63880 34388 63908 34496
rect 64322 34484 64328 34496
rect 64380 34484 64386 34536
rect 69934 34484 69940 34536
rect 69992 34524 69998 34536
rect 70029 34527 70087 34533
rect 70029 34524 70041 34527
rect 69992 34496 70041 34524
rect 69992 34484 69998 34496
rect 70029 34493 70041 34496
rect 70075 34493 70087 34527
rect 70029 34487 70087 34493
rect 70118 34484 70124 34536
rect 70176 34524 70182 34536
rect 70305 34527 70363 34533
rect 70305 34524 70317 34527
rect 70176 34496 70317 34524
rect 70176 34484 70182 34496
rect 70305 34493 70317 34496
rect 70351 34493 70363 34527
rect 72344 34524 72372 34691
rect 72602 34688 72608 34700
rect 72660 34688 72666 34740
rect 76285 34731 76343 34737
rect 76285 34697 76297 34731
rect 76331 34728 76343 34731
rect 77294 34728 77300 34740
rect 76331 34700 77300 34728
rect 76331 34697 76343 34700
rect 76285 34691 76343 34697
rect 76392 34601 76420 34700
rect 77294 34688 77300 34700
rect 77352 34688 77358 34740
rect 77754 34728 77760 34740
rect 77715 34700 77760 34728
rect 77754 34688 77760 34700
rect 77812 34688 77818 34740
rect 79962 34688 79968 34740
rect 80020 34728 80026 34740
rect 80057 34731 80115 34737
rect 80057 34728 80069 34731
rect 80020 34700 80069 34728
rect 80020 34688 80026 34700
rect 80057 34697 80069 34700
rect 80103 34697 80115 34731
rect 80057 34691 80115 34697
rect 81253 34731 81311 34737
rect 81253 34697 81265 34731
rect 81299 34728 81311 34731
rect 83918 34728 83924 34740
rect 81299 34700 83924 34728
rect 81299 34697 81311 34700
rect 81253 34691 81311 34697
rect 83918 34688 83924 34700
rect 83976 34688 83982 34740
rect 85669 34731 85727 34737
rect 85669 34697 85681 34731
rect 85715 34728 85727 34731
rect 85758 34728 85764 34740
rect 85715 34700 85764 34728
rect 85715 34697 85727 34700
rect 85669 34691 85727 34697
rect 85758 34688 85764 34700
rect 85816 34728 85822 34740
rect 86770 34728 86776 34740
rect 85816 34700 86776 34728
rect 85816 34688 85822 34700
rect 86770 34688 86776 34700
rect 86828 34688 86834 34740
rect 86862 34688 86868 34740
rect 86920 34728 86926 34740
rect 87141 34731 87199 34737
rect 87141 34728 87153 34731
rect 86920 34700 87153 34728
rect 86920 34688 86926 34700
rect 87141 34697 87153 34700
rect 87187 34697 87199 34731
rect 88334 34728 88340 34740
rect 88295 34700 88340 34728
rect 87141 34691 87199 34697
rect 88334 34688 88340 34700
rect 88392 34688 88398 34740
rect 79597 34663 79655 34669
rect 79597 34629 79609 34663
rect 79643 34660 79655 34663
rect 80425 34663 80483 34669
rect 80425 34660 80437 34663
rect 79643 34632 80437 34660
rect 79643 34629 79655 34632
rect 79597 34623 79655 34629
rect 80425 34629 80437 34632
rect 80471 34629 80483 34663
rect 80425 34623 80483 34629
rect 87046 34620 87052 34672
rect 87104 34660 87110 34672
rect 87693 34663 87751 34669
rect 87693 34660 87705 34663
rect 87104 34632 87705 34660
rect 87104 34620 87110 34632
rect 87693 34629 87705 34632
rect 87739 34629 87751 34663
rect 87693 34623 87751 34629
rect 76377 34595 76435 34601
rect 76377 34561 76389 34595
rect 76423 34561 76435 34595
rect 76377 34555 76435 34561
rect 76653 34595 76711 34601
rect 76653 34561 76665 34595
rect 76699 34592 76711 34595
rect 80514 34592 80520 34604
rect 76699 34564 80520 34592
rect 76699 34561 76711 34564
rect 76653 34555 76711 34561
rect 80514 34552 80520 34564
rect 80572 34552 80578 34604
rect 82265 34595 82323 34601
rect 82265 34592 82277 34595
rect 81084 34564 82277 34592
rect 72513 34527 72571 34533
rect 72513 34524 72525 34527
rect 72344 34496 72525 34524
rect 70305 34487 70363 34493
rect 72513 34493 72525 34496
rect 72559 34493 72571 34527
rect 72513 34487 72571 34493
rect 78950 34484 78956 34536
rect 79008 34524 79014 34536
rect 79597 34527 79655 34533
rect 79597 34524 79609 34527
rect 79008 34496 79609 34524
rect 79008 34484 79014 34496
rect 79597 34493 79609 34496
rect 79643 34524 79655 34527
rect 79781 34527 79839 34533
rect 79781 34524 79793 34527
rect 79643 34496 79793 34524
rect 79643 34493 79655 34496
rect 79597 34487 79655 34493
rect 79781 34493 79793 34496
rect 79827 34493 79839 34527
rect 79781 34487 79839 34493
rect 79965 34527 80023 34533
rect 79965 34493 79977 34527
rect 80011 34524 80023 34527
rect 81084 34524 81112 34564
rect 82265 34561 82277 34564
rect 82311 34592 82323 34595
rect 82311 34564 83412 34592
rect 82311 34561 82323 34564
rect 82265 34555 82323 34561
rect 80011 34496 81112 34524
rect 81161 34527 81219 34533
rect 80011 34493 80023 34496
rect 79965 34487 80023 34493
rect 81161 34493 81173 34527
rect 81207 34524 81219 34527
rect 81342 34524 81348 34536
rect 81207 34496 81348 34524
rect 81207 34493 81219 34496
rect 81161 34487 81219 34493
rect 81342 34484 81348 34496
rect 81400 34524 81406 34536
rect 82170 34524 82176 34536
rect 81400 34496 82032 34524
rect 82131 34496 82176 34524
rect 81400 34484 81406 34496
rect 82004 34456 82032 34496
rect 82170 34484 82176 34496
rect 82228 34484 82234 34536
rect 83185 34527 83243 34533
rect 83185 34524 83197 34527
rect 82280 34496 83197 34524
rect 82280 34456 82308 34496
rect 83185 34493 83197 34496
rect 83231 34524 83243 34527
rect 83274 34524 83280 34536
rect 83231 34496 83280 34524
rect 83231 34493 83243 34496
rect 83185 34487 83243 34493
rect 83274 34484 83280 34496
rect 83332 34484 83338 34536
rect 83384 34533 83412 34564
rect 85482 34552 85488 34604
rect 85540 34592 85546 34604
rect 86037 34595 86095 34601
rect 86037 34592 86049 34595
rect 85540 34564 86049 34592
rect 85540 34552 85546 34564
rect 86037 34561 86049 34564
rect 86083 34561 86095 34595
rect 86037 34555 86095 34561
rect 87414 34552 87420 34604
rect 87472 34592 87478 34604
rect 88061 34595 88119 34601
rect 88061 34592 88073 34595
rect 87472 34564 88073 34592
rect 87472 34552 87478 34564
rect 88061 34561 88073 34564
rect 88107 34561 88119 34595
rect 88061 34555 88119 34561
rect 83369 34527 83427 34533
rect 83369 34493 83381 34527
rect 83415 34493 83427 34527
rect 85758 34524 85764 34536
rect 85719 34496 85764 34524
rect 83369 34487 83427 34493
rect 85758 34484 85764 34496
rect 85816 34484 85822 34536
rect 86954 34484 86960 34536
rect 87012 34524 87018 34536
rect 87509 34527 87567 34533
rect 87509 34524 87521 34527
rect 87012 34496 87521 34524
rect 87012 34484 87018 34496
rect 87509 34493 87521 34496
rect 87555 34493 87567 34527
rect 87874 34524 87880 34536
rect 87835 34496 87880 34524
rect 87509 34487 87567 34493
rect 87874 34484 87880 34496
rect 87932 34484 87938 34536
rect 88242 34524 88248 34536
rect 88203 34496 88248 34524
rect 88242 34484 88248 34496
rect 88300 34484 88306 34536
rect 82004 34428 82308 34456
rect 62500 34360 63908 34388
rect 59817 34351 59875 34357
rect 78582 34348 78588 34400
rect 78640 34388 78646 34400
rect 83461 34391 83519 34397
rect 83461 34388 83473 34391
rect 78640 34360 83473 34388
rect 78640 34348 78646 34360
rect 83461 34357 83473 34360
rect 83507 34388 83519 34391
rect 84930 34388 84936 34400
rect 83507 34360 84936 34388
rect 83507 34357 83519 34360
rect 83461 34351 83519 34357
rect 84930 34348 84936 34360
rect 84988 34348 84994 34400
rect 1104 34298 111136 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 81046 34298
rect 81098 34246 81110 34298
rect 81162 34246 81174 34298
rect 81226 34246 81238 34298
rect 81290 34246 111136 34298
rect 1104 34224 111136 34246
rect 4062 34144 4068 34196
rect 4120 34184 4126 34196
rect 13538 34184 13544 34196
rect 4120 34156 13544 34184
rect 4120 34144 4126 34156
rect 13538 34144 13544 34156
rect 13596 34144 13602 34196
rect 15381 34187 15439 34193
rect 15381 34184 15393 34187
rect 13648 34156 15393 34184
rect 5350 34116 5356 34128
rect 5092 34088 5356 34116
rect 5092 34057 5120 34088
rect 5350 34076 5356 34088
rect 5408 34076 5414 34128
rect 13648 34116 13676 34156
rect 15381 34153 15393 34156
rect 15427 34153 15439 34187
rect 15381 34147 15439 34153
rect 15657 34187 15715 34193
rect 15657 34153 15669 34187
rect 15703 34184 15715 34187
rect 15746 34184 15752 34196
rect 15703 34156 15752 34184
rect 15703 34153 15715 34156
rect 15657 34147 15715 34153
rect 14274 34116 14280 34128
rect 10704 34088 13676 34116
rect 14235 34088 14280 34116
rect 5077 34051 5135 34057
rect 5077 34017 5089 34051
rect 5123 34017 5135 34051
rect 5077 34011 5135 34017
rect 5261 34051 5319 34057
rect 5261 34017 5273 34051
rect 5307 34048 5319 34051
rect 5442 34048 5448 34060
rect 5307 34020 5448 34048
rect 5307 34017 5319 34020
rect 5261 34011 5319 34017
rect 5442 34008 5448 34020
rect 5500 34008 5506 34060
rect 10505 34051 10563 34057
rect 5552 34020 10364 34048
rect 3694 33940 3700 33992
rect 3752 33980 3758 33992
rect 5353 33983 5411 33989
rect 5353 33980 5365 33983
rect 3752 33952 5365 33980
rect 3752 33940 3758 33952
rect 5353 33949 5365 33952
rect 5399 33949 5411 33983
rect 5353 33943 5411 33949
rect 5442 33872 5448 33924
rect 5500 33912 5506 33924
rect 5552 33912 5580 34020
rect 9030 33940 9036 33992
rect 9088 33980 9094 33992
rect 9677 33983 9735 33989
rect 9677 33980 9689 33983
rect 9088 33952 9689 33980
rect 9088 33940 9094 33952
rect 9677 33949 9689 33952
rect 9723 33949 9735 33983
rect 10226 33980 10232 33992
rect 10139 33952 10232 33980
rect 9677 33943 9735 33949
rect 10226 33940 10232 33952
rect 10284 33940 10290 33992
rect 5500 33884 5580 33912
rect 5500 33872 5506 33884
rect 9490 33844 9496 33856
rect 9451 33816 9496 33844
rect 9490 33804 9496 33816
rect 9548 33844 9554 33856
rect 10244 33844 10272 33940
rect 10336 33912 10364 34020
rect 10505 34017 10517 34051
rect 10551 34048 10563 34051
rect 10594 34048 10600 34060
rect 10551 34020 10600 34048
rect 10551 34017 10563 34020
rect 10505 34011 10563 34017
rect 10594 34008 10600 34020
rect 10652 34008 10658 34060
rect 10704 34057 10732 34088
rect 10689 34051 10747 34057
rect 10689 34017 10701 34051
rect 10735 34017 10747 34051
rect 13170 34048 13176 34060
rect 13131 34020 13176 34048
rect 10689 34011 10747 34017
rect 13170 34008 13176 34020
rect 13228 34008 13234 34060
rect 13648 34057 13676 34088
rect 14274 34076 14280 34088
rect 14332 34076 14338 34128
rect 13633 34051 13691 34057
rect 13633 34017 13645 34051
rect 13679 34017 13691 34051
rect 13633 34011 13691 34017
rect 13725 34051 13783 34057
rect 13725 34017 13737 34051
rect 13771 34048 13783 34051
rect 15289 34051 15347 34057
rect 13771 34020 15240 34048
rect 13771 34017 13783 34020
rect 13725 34011 13783 34017
rect 12802 33940 12808 33992
rect 12860 33980 12866 33992
rect 12989 33983 13047 33989
rect 12989 33980 13001 33983
rect 12860 33952 13001 33980
rect 12860 33940 12866 33952
rect 12989 33949 13001 33952
rect 13035 33949 13047 33983
rect 15212 33980 15240 34020
rect 15289 34017 15301 34051
rect 15335 34048 15347 34051
rect 15672 34048 15700 34147
rect 15746 34144 15752 34156
rect 15804 34144 15810 34196
rect 21100 34156 21680 34184
rect 21100 34116 21128 34156
rect 15335 34020 15700 34048
rect 18708 34088 21128 34116
rect 15335 34017 15347 34020
rect 15289 34011 15347 34017
rect 18708 33992 18736 34088
rect 18874 34008 18880 34060
rect 18932 34048 18938 34060
rect 19429 34051 19487 34057
rect 19429 34048 19441 34051
rect 18932 34020 19441 34048
rect 18932 34008 18938 34020
rect 19429 34017 19441 34020
rect 19475 34048 19487 34051
rect 19475 34020 19656 34048
rect 19475 34017 19487 34020
rect 19429 34011 19487 34017
rect 18690 33980 18696 33992
rect 15212 33952 18696 33980
rect 12989 33943 13047 33949
rect 18690 33940 18696 33952
rect 18748 33940 18754 33992
rect 18785 33983 18843 33989
rect 18785 33949 18797 33983
rect 18831 33949 18843 33983
rect 18785 33943 18843 33949
rect 19521 33983 19579 33989
rect 19521 33949 19533 33983
rect 19567 33949 19579 33983
rect 19628 33980 19656 34020
rect 19702 34008 19708 34060
rect 19760 34048 19766 34060
rect 19797 34051 19855 34057
rect 19797 34048 19809 34051
rect 19760 34020 19809 34048
rect 19760 34008 19766 34020
rect 19797 34017 19809 34020
rect 19843 34017 19855 34051
rect 19797 34011 19855 34017
rect 19981 34051 20039 34057
rect 19981 34017 19993 34051
rect 20027 34048 20039 34051
rect 20162 34048 20168 34060
rect 20027 34020 20168 34048
rect 20027 34017 20039 34020
rect 19981 34011 20039 34017
rect 20162 34008 20168 34020
rect 20220 34008 20226 34060
rect 21100 34057 21128 34088
rect 21085 34051 21143 34057
rect 20272 34020 21036 34048
rect 20272 33980 20300 34020
rect 19628 33952 20300 33980
rect 19521 33943 19579 33949
rect 18800 33912 18828 33943
rect 10336 33884 18828 33912
rect 19536 33912 19564 33943
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 20901 33983 20959 33989
rect 20901 33980 20913 33983
rect 20680 33952 20913 33980
rect 20680 33940 20686 33952
rect 20901 33949 20913 33952
rect 20947 33949 20959 33983
rect 21008 33980 21036 34020
rect 21085 34017 21097 34051
rect 21131 34017 21143 34051
rect 21542 34048 21548 34060
rect 21085 34011 21143 34017
rect 21192 34020 21548 34048
rect 21192 33980 21220 34020
rect 21542 34008 21548 34020
rect 21600 34008 21606 34060
rect 21652 34057 21680 34156
rect 21818 34144 21824 34196
rect 21876 34184 21882 34196
rect 30282 34184 30288 34196
rect 21876 34156 30288 34184
rect 21876 34144 21882 34156
rect 30282 34144 30288 34156
rect 30340 34144 30346 34196
rect 51534 34184 51540 34196
rect 30392 34156 51540 34184
rect 28166 34116 28172 34128
rect 28127 34088 28172 34116
rect 28166 34076 28172 34088
rect 28224 34076 28230 34128
rect 28350 34076 28356 34128
rect 28408 34116 28414 34128
rect 30392 34116 30420 34156
rect 51534 34144 51540 34156
rect 51592 34144 51598 34196
rect 56597 34187 56655 34193
rect 56597 34153 56609 34187
rect 56643 34184 56655 34187
rect 62666 34184 62672 34196
rect 56643 34156 62672 34184
rect 56643 34153 56655 34156
rect 56597 34147 56655 34153
rect 62666 34144 62672 34156
rect 62724 34144 62730 34196
rect 42058 34116 42064 34128
rect 28408 34088 30420 34116
rect 30484 34088 42064 34116
rect 28408 34076 28414 34088
rect 21637 34051 21695 34057
rect 21637 34017 21649 34051
rect 21683 34017 21695 34051
rect 21637 34011 21695 34017
rect 21821 34051 21879 34057
rect 21821 34017 21833 34051
rect 21867 34048 21879 34051
rect 22465 34051 22523 34057
rect 22465 34048 22477 34051
rect 21867 34020 22477 34048
rect 21867 34017 21879 34020
rect 21821 34011 21879 34017
rect 21008 33952 21220 33980
rect 20901 33943 20959 33949
rect 20257 33915 20315 33921
rect 20257 33912 20269 33915
rect 19536 33884 20269 33912
rect 20257 33881 20269 33884
rect 20303 33912 20315 33915
rect 22020 33912 22048 34020
rect 22465 34017 22477 34020
rect 22511 34048 22523 34051
rect 26786 34048 26792 34060
rect 22511 34020 26648 34048
rect 26747 34020 26792 34048
rect 22511 34017 22523 34020
rect 22465 34011 22523 34017
rect 26510 33980 26516 33992
rect 26471 33952 26516 33980
rect 26510 33940 26516 33952
rect 26568 33940 26574 33992
rect 26620 33980 26648 34020
rect 26786 34008 26792 34020
rect 26844 34008 26850 34060
rect 27982 34008 27988 34060
rect 28040 34048 28046 34060
rect 30484 34048 30512 34088
rect 42058 34076 42064 34088
rect 42116 34076 42122 34128
rect 28040 34020 30512 34048
rect 30561 34051 30619 34057
rect 28040 34008 28046 34020
rect 30561 34017 30573 34051
rect 30607 34048 30619 34051
rect 70026 34048 70032 34060
rect 30607 34020 70032 34048
rect 30607 34017 30619 34020
rect 30561 34011 30619 34017
rect 70026 34008 70032 34020
rect 70084 34008 70090 34060
rect 29365 33983 29423 33989
rect 29365 33980 29377 33983
rect 26620 33952 29377 33980
rect 29365 33949 29377 33952
rect 29411 33949 29423 33983
rect 29365 33943 29423 33949
rect 31680 33952 42196 33980
rect 31680 33912 31708 33952
rect 20303 33884 22048 33912
rect 27448 33884 31708 33912
rect 42168 33912 42196 33952
rect 56597 33915 56655 33921
rect 56597 33912 56609 33915
rect 42168 33884 56609 33912
rect 20303 33881 20315 33884
rect 20257 33875 20315 33881
rect 12802 33844 12808 33856
rect 9548 33816 10272 33844
rect 12763 33816 12808 33844
rect 9548 33804 9554 33816
rect 12802 33804 12808 33816
rect 12860 33804 12866 33856
rect 20162 33844 20168 33856
rect 20123 33816 20168 33844
rect 20162 33804 20168 33816
rect 20220 33804 20226 33856
rect 20622 33844 20628 33856
rect 20583 33816 20628 33844
rect 20622 33804 20628 33816
rect 20680 33804 20686 33856
rect 22097 33847 22155 33853
rect 22097 33813 22109 33847
rect 22143 33844 22155 33847
rect 27448 33844 27476 33884
rect 56597 33881 56609 33884
rect 56643 33881 56655 33915
rect 56597 33875 56655 33881
rect 22143 33816 27476 33844
rect 22143 33813 22155 33816
rect 22097 33807 22155 33813
rect 28258 33804 28264 33856
rect 28316 33844 28322 33856
rect 29178 33844 29184 33856
rect 28316 33816 29184 33844
rect 28316 33804 28322 33816
rect 29178 33804 29184 33816
rect 29236 33804 29242 33856
rect 1104 33754 29256 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 29256 33754
rect 1104 33680 29256 33702
rect 5261 33643 5319 33649
rect 5261 33609 5273 33643
rect 5307 33640 5319 33643
rect 5350 33640 5356 33652
rect 5307 33612 5356 33640
rect 5307 33609 5319 33612
rect 5261 33603 5319 33609
rect 5350 33600 5356 33612
rect 5408 33600 5414 33652
rect 13630 33640 13636 33652
rect 13591 33612 13636 33640
rect 13630 33600 13636 33612
rect 13688 33600 13694 33652
rect 14550 33640 14556 33652
rect 14511 33612 14556 33640
rect 14550 33600 14556 33612
rect 14608 33600 14614 33652
rect 18690 33600 18696 33652
rect 18748 33640 18754 33652
rect 19061 33643 19119 33649
rect 19061 33640 19073 33643
rect 18748 33612 19073 33640
rect 18748 33600 18754 33612
rect 19061 33609 19073 33612
rect 19107 33609 19119 33643
rect 19334 33640 19340 33652
rect 19295 33612 19340 33640
rect 19061 33603 19119 33609
rect 19334 33600 19340 33612
rect 19392 33600 19398 33652
rect 20162 33600 20168 33652
rect 20220 33640 20226 33652
rect 21545 33643 21603 33649
rect 21545 33640 21557 33643
rect 20220 33612 21557 33640
rect 20220 33600 20226 33612
rect 12452 33544 13584 33572
rect 2869 33507 2927 33513
rect 2869 33473 2881 33507
rect 2915 33504 2927 33507
rect 4706 33504 4712 33516
rect 2915 33476 4712 33504
rect 2915 33473 2927 33476
rect 2869 33467 2927 33473
rect 4706 33464 4712 33476
rect 4764 33464 4770 33516
rect 9030 33504 9036 33516
rect 8991 33476 9036 33504
rect 9030 33464 9036 33476
rect 9088 33464 9094 33516
rect 10873 33507 10931 33513
rect 10873 33504 10885 33507
rect 9140 33476 10885 33504
rect 2593 33439 2651 33445
rect 2593 33405 2605 33439
rect 2639 33436 2651 33439
rect 2639 33408 4292 33436
rect 2639 33405 2651 33408
rect 2593 33399 2651 33405
rect 4264 33368 4292 33408
rect 4338 33396 4344 33448
rect 4396 33436 4402 33448
rect 5077 33439 5135 33445
rect 5077 33436 5089 33439
rect 4396 33408 5089 33436
rect 4396 33396 4402 33408
rect 5077 33405 5089 33408
rect 5123 33436 5135 33439
rect 8202 33436 8208 33448
rect 5123 33408 8208 33436
rect 5123 33405 5135 33408
rect 5077 33399 5135 33405
rect 8202 33396 8208 33408
rect 8260 33396 8266 33448
rect 8757 33439 8815 33445
rect 8757 33405 8769 33439
rect 8803 33436 8815 33439
rect 9140 33436 9168 33476
rect 10873 33473 10885 33476
rect 10919 33473 10931 33507
rect 10873 33467 10931 33473
rect 8803 33408 9168 33436
rect 10597 33439 10655 33445
rect 8803 33405 8815 33408
rect 8757 33399 8815 33405
rect 10597 33405 10609 33439
rect 10643 33436 10655 33439
rect 12452 33436 12480 33544
rect 10643 33408 12480 33436
rect 10643 33405 10655 33408
rect 10597 33399 10655 33405
rect 12526 33396 12532 33448
rect 12584 33445 12590 33448
rect 12584 33439 12633 33445
rect 12584 33405 12587 33439
rect 12621 33405 12633 33439
rect 12584 33399 12633 33405
rect 12713 33439 12771 33445
rect 12713 33405 12725 33439
rect 12759 33436 12771 33439
rect 12802 33436 12808 33448
rect 12759 33408 12808 33436
rect 12759 33405 12771 33408
rect 12713 33399 12771 33405
rect 12584 33396 12590 33399
rect 10413 33371 10471 33377
rect 4264 33340 4476 33368
rect 4154 33300 4160 33312
rect 4115 33272 4160 33300
rect 4154 33260 4160 33272
rect 4212 33260 4218 33312
rect 4448 33309 4476 33340
rect 10413 33337 10425 33371
rect 10459 33368 10471 33371
rect 10870 33368 10876 33380
rect 10459 33340 10876 33368
rect 10459 33337 10471 33340
rect 10413 33331 10471 33337
rect 10870 33328 10876 33340
rect 10928 33328 10934 33380
rect 4433 33303 4491 33309
rect 4433 33269 4445 33303
rect 4479 33300 4491 33303
rect 4614 33300 4620 33312
rect 4479 33272 4620 33300
rect 4479 33269 4491 33272
rect 4433 33263 4491 33269
rect 4614 33260 4620 33272
rect 4672 33300 4678 33312
rect 4890 33300 4896 33312
rect 4672 33272 4896 33300
rect 4672 33260 4678 33272
rect 4890 33260 4896 33272
rect 4948 33260 4954 33312
rect 8113 33303 8171 33309
rect 8113 33269 8125 33303
rect 8159 33300 8171 33303
rect 8294 33300 8300 33312
rect 8159 33272 8300 33300
rect 8159 33269 8171 33272
rect 8113 33263 8171 33269
rect 8294 33260 8300 33272
rect 8352 33260 8358 33312
rect 10962 33260 10968 33312
rect 11020 33300 11026 33312
rect 12161 33303 12219 33309
rect 12161 33300 12173 33303
rect 11020 33272 12173 33300
rect 11020 33260 11026 33272
rect 12161 33269 12173 33272
rect 12207 33300 12219 33303
rect 12728 33300 12756 33399
rect 12802 33396 12808 33408
rect 12860 33396 12866 33448
rect 13173 33439 13231 33445
rect 13173 33405 13185 33439
rect 13219 33405 13231 33439
rect 13173 33399 13231 33405
rect 13357 33439 13415 33445
rect 13357 33405 13369 33439
rect 13403 33436 13415 33439
rect 13556 33436 13584 33544
rect 13906 33436 13912 33448
rect 13403 33408 13912 33436
rect 13403 33405 13415 33408
rect 13357 33399 13415 33405
rect 13188 33368 13216 33399
rect 13906 33396 13912 33408
rect 13964 33396 13970 33448
rect 14550 33396 14556 33448
rect 14608 33436 14614 33448
rect 14645 33439 14703 33445
rect 14645 33436 14657 33439
rect 14608 33408 14657 33436
rect 14608 33396 14614 33408
rect 14645 33405 14657 33408
rect 14691 33405 14703 33439
rect 14645 33399 14703 33405
rect 18877 33439 18935 33445
rect 18877 33405 18889 33439
rect 18923 33436 18935 33439
rect 19334 33436 19340 33448
rect 18923 33408 19340 33436
rect 18923 33405 18935 33408
rect 18877 33399 18935 33405
rect 19334 33396 19340 33408
rect 19392 33396 19398 33448
rect 19981 33439 20039 33445
rect 19981 33405 19993 33439
rect 20027 33405 20039 33439
rect 19981 33399 20039 33405
rect 14734 33368 14740 33380
rect 13188 33340 14740 33368
rect 14734 33328 14740 33340
rect 14792 33328 14798 33380
rect 19996 33368 20024 33399
rect 20070 33396 20076 33448
rect 20128 33436 20134 33448
rect 20165 33439 20223 33445
rect 20165 33436 20177 33439
rect 20128 33408 20177 33436
rect 20128 33396 20134 33408
rect 20165 33405 20177 33408
rect 20211 33436 20223 33439
rect 20717 33439 20775 33445
rect 20717 33436 20729 33439
rect 20211 33408 20729 33436
rect 20211 33405 20223 33408
rect 20165 33399 20223 33405
rect 20717 33405 20729 33408
rect 20763 33405 20775 33439
rect 20717 33399 20775 33405
rect 20901 33439 20959 33445
rect 20901 33405 20913 33439
rect 20947 33436 20959 33439
rect 21100 33436 21128 33612
rect 21545 33609 21557 33612
rect 21591 33640 21603 33643
rect 26050 33640 26056 33652
rect 21591 33612 26056 33640
rect 21591 33609 21603 33612
rect 21545 33603 21603 33609
rect 26050 33600 26056 33612
rect 26108 33600 26114 33652
rect 26694 33600 26700 33652
rect 26752 33640 26758 33652
rect 27246 33640 27252 33652
rect 26752 33612 27252 33640
rect 26752 33600 26758 33612
rect 27246 33600 27252 33612
rect 27304 33640 27310 33652
rect 28258 33640 28264 33652
rect 27304 33612 28264 33640
rect 27304 33600 27310 33612
rect 28258 33600 28264 33612
rect 28316 33600 28322 33652
rect 29365 33643 29423 33649
rect 29365 33609 29377 33643
rect 29411 33640 29423 33643
rect 61930 33640 61936 33652
rect 29411 33612 61936 33640
rect 29411 33609 29423 33612
rect 29365 33603 29423 33609
rect 61930 33600 61936 33612
rect 61988 33600 61994 33652
rect 21177 33575 21235 33581
rect 21177 33541 21189 33575
rect 21223 33572 21235 33575
rect 62206 33572 62212 33584
rect 21223 33544 62212 33572
rect 21223 33541 21235 33544
rect 21177 33535 21235 33541
rect 62206 33532 62212 33544
rect 62264 33532 62270 33584
rect 25038 33504 25044 33516
rect 24872 33476 25044 33504
rect 20947 33408 21128 33436
rect 20947 33405 20959 33408
rect 20901 33399 20959 33405
rect 24394 33396 24400 33448
rect 24452 33436 24458 33448
rect 24872 33445 24900 33476
rect 25038 33464 25044 33476
rect 25096 33464 25102 33516
rect 25958 33504 25964 33516
rect 25919 33476 25964 33504
rect 25958 33464 25964 33476
rect 26016 33464 26022 33516
rect 26050 33464 26056 33516
rect 26108 33504 26114 33516
rect 64598 33504 64604 33516
rect 26108 33476 64604 33504
rect 26108 33464 26114 33476
rect 64598 33464 64604 33476
rect 64656 33464 64662 33516
rect 24857 33439 24915 33445
rect 24857 33436 24869 33439
rect 24452 33408 24869 33436
rect 24452 33396 24458 33408
rect 24857 33405 24869 33408
rect 24903 33405 24915 33439
rect 24857 33399 24915 33405
rect 24949 33439 25007 33445
rect 24949 33405 24961 33439
rect 24995 33436 25007 33439
rect 25222 33436 25228 33448
rect 24995 33408 25228 33436
rect 24995 33405 25007 33408
rect 24949 33399 25007 33405
rect 25222 33396 25228 33408
rect 25280 33396 25286 33448
rect 25317 33439 25375 33445
rect 25317 33405 25329 33439
rect 25363 33405 25375 33439
rect 25317 33399 25375 33405
rect 25409 33439 25467 33445
rect 25409 33405 25421 33439
rect 25455 33405 25467 33439
rect 25409 33399 25467 33405
rect 20622 33368 20628 33380
rect 19996 33340 20628 33368
rect 14826 33300 14832 33312
rect 12207 33272 12756 33300
rect 14787 33272 14832 33300
rect 12207 33269 12219 33272
rect 12161 33263 12219 33269
rect 14826 33260 14832 33272
rect 14884 33260 14890 33312
rect 19334 33260 19340 33312
rect 19392 33300 19398 33312
rect 19797 33303 19855 33309
rect 19797 33300 19809 33303
rect 19392 33272 19809 33300
rect 19392 33260 19398 33272
rect 19797 33269 19809 33272
rect 19843 33300 19855 33303
rect 19996 33300 20024 33340
rect 20622 33328 20628 33340
rect 20680 33328 20686 33380
rect 25332 33368 25360 33399
rect 24504 33340 25360 33368
rect 25424 33368 25452 33399
rect 25866 33396 25872 33448
rect 25924 33436 25930 33448
rect 30561 33439 30619 33445
rect 30561 33436 30573 33439
rect 25924 33408 30573 33436
rect 25924 33396 25930 33408
rect 30561 33405 30573 33408
rect 30607 33405 30619 33439
rect 30561 33399 30619 33405
rect 26050 33368 26056 33380
rect 25424 33340 26056 33368
rect 19843 33272 20024 33300
rect 19843 33269 19855 33272
rect 19797 33263 19855 33269
rect 23566 33260 23572 33312
rect 23624 33300 23630 33312
rect 24504 33309 24532 33340
rect 26050 33328 26056 33340
rect 26108 33368 26114 33380
rect 26421 33371 26479 33377
rect 26421 33368 26433 33371
rect 26108 33340 26433 33368
rect 26108 33328 26114 33340
rect 26421 33337 26433 33340
rect 26467 33368 26479 33371
rect 69290 33368 69296 33380
rect 26467 33340 69296 33368
rect 26467 33337 26479 33340
rect 26421 33331 26479 33337
rect 69290 33328 69296 33340
rect 69348 33328 69354 33380
rect 24489 33303 24547 33309
rect 24489 33300 24501 33303
rect 23624 33272 24501 33300
rect 23624 33260 23630 33272
rect 24489 33269 24501 33272
rect 24535 33269 24547 33303
rect 24489 33263 24547 33269
rect 25038 33260 25044 33312
rect 25096 33300 25102 33312
rect 25774 33300 25780 33312
rect 25096 33272 25780 33300
rect 25096 33260 25102 33272
rect 25774 33260 25780 33272
rect 25832 33300 25838 33312
rect 26237 33303 26295 33309
rect 26237 33300 26249 33303
rect 25832 33272 26249 33300
rect 25832 33260 25838 33272
rect 26237 33269 26249 33272
rect 26283 33300 26295 33303
rect 76006 33300 76012 33312
rect 26283 33272 76012 33300
rect 26283 33269 26295 33272
rect 26237 33263 26295 33269
rect 76006 33260 76012 33272
rect 76064 33260 76070 33312
rect 1104 33210 29256 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 29256 33210
rect 1104 33136 29256 33158
rect 3234 33056 3240 33108
rect 3292 33096 3298 33108
rect 13998 33096 14004 33108
rect 3292 33068 14004 33096
rect 3292 33056 3298 33068
rect 13998 33056 14004 33068
rect 14056 33056 14062 33108
rect 16666 33056 16672 33108
rect 16724 33096 16730 33108
rect 20993 33099 21051 33105
rect 20993 33096 21005 33099
rect 16724 33068 21005 33096
rect 16724 33056 16730 33068
rect 20993 33065 21005 33068
rect 21039 33065 21051 33099
rect 25774 33096 25780 33108
rect 25735 33068 25780 33096
rect 20993 33059 21051 33065
rect 25774 33056 25780 33068
rect 25832 33056 25838 33108
rect 25958 33056 25964 33108
rect 26016 33096 26022 33108
rect 34606 33096 34612 33108
rect 26016 33068 34612 33096
rect 26016 33056 26022 33068
rect 34606 33056 34612 33068
rect 34664 33056 34670 33108
rect 9398 33028 9404 33040
rect 7484 33000 9404 33028
rect 4338 32960 4344 32972
rect 4299 32932 4344 32960
rect 4338 32920 4344 32932
rect 4396 32920 4402 32972
rect 4617 32963 4675 32969
rect 4617 32929 4629 32963
rect 4663 32960 4675 32963
rect 7484 32960 7512 33000
rect 9398 32988 9404 33000
rect 9456 32988 9462 33040
rect 12894 33028 12900 33040
rect 12544 33000 12900 33028
rect 8202 32960 8208 32972
rect 4663 32932 7512 32960
rect 8163 32932 8208 32960
rect 4663 32929 4675 32932
rect 4617 32923 4675 32929
rect 8202 32920 8208 32932
rect 8260 32920 8266 32972
rect 12544 32969 12572 33000
rect 12894 32988 12900 33000
rect 12952 33028 12958 33040
rect 12989 33031 13047 33037
rect 12989 33028 13001 33031
rect 12952 33000 13001 33028
rect 12952 32988 12958 33000
rect 12989 32997 13001 33000
rect 13035 33028 13047 33031
rect 13354 33028 13360 33040
rect 13035 33000 13360 33028
rect 13035 32997 13047 33000
rect 12989 32991 13047 32997
rect 13354 32988 13360 33000
rect 13412 33028 13418 33040
rect 13412 33000 14412 33028
rect 13412 32988 13418 33000
rect 12529 32963 12587 32969
rect 12529 32929 12541 32963
rect 12575 32929 12587 32963
rect 12529 32923 12587 32929
rect 13449 32963 13507 32969
rect 13449 32929 13461 32963
rect 13495 32960 13507 32963
rect 13725 32963 13783 32969
rect 13725 32960 13737 32963
rect 13495 32932 13737 32960
rect 13495 32929 13507 32932
rect 13449 32923 13507 32929
rect 13725 32929 13737 32932
rect 13771 32929 13783 32963
rect 14384 32960 14412 33000
rect 17218 32988 17224 33040
rect 17276 33028 17282 33040
rect 55122 33028 55128 33040
rect 17276 33000 55128 33028
rect 17276 32988 17282 33000
rect 55122 32988 55128 33000
rect 55180 32988 55186 33040
rect 18509 32963 18567 32969
rect 14384 32932 18460 32960
rect 13725 32923 13783 32929
rect 4801 32895 4859 32901
rect 4801 32861 4813 32895
rect 4847 32892 4859 32895
rect 5350 32892 5356 32904
rect 4847 32864 5356 32892
rect 4847 32861 4859 32864
rect 4801 32855 4859 32861
rect 5350 32852 5356 32864
rect 5408 32852 5414 32904
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32861 5779 32895
rect 5994 32892 6000 32904
rect 5955 32864 6000 32892
rect 5721 32855 5779 32861
rect 4890 32716 4896 32768
rect 4948 32756 4954 32768
rect 5736 32756 5764 32855
rect 5994 32852 6000 32864
rect 6052 32852 6058 32904
rect 8938 32852 8944 32904
rect 8996 32892 9002 32904
rect 8996 32864 14044 32892
rect 8996 32852 9002 32864
rect 6656 32796 7604 32824
rect 6656 32756 6684 32796
rect 4948 32728 6684 32756
rect 7285 32759 7343 32765
rect 4948 32716 4954 32728
rect 7285 32725 7297 32759
rect 7331 32756 7343 32759
rect 7374 32756 7380 32768
rect 7331 32728 7380 32756
rect 7331 32725 7343 32728
rect 7285 32719 7343 32725
rect 7374 32716 7380 32728
rect 7432 32716 7438 32768
rect 7576 32765 7604 32796
rect 12342 32784 12348 32836
rect 12400 32824 12406 32836
rect 13449 32827 13507 32833
rect 13449 32824 13461 32827
rect 12400 32796 13461 32824
rect 12400 32784 12406 32796
rect 13449 32793 13461 32796
rect 13495 32824 13507 32827
rect 13541 32827 13599 32833
rect 13541 32824 13553 32827
rect 13495 32796 13553 32824
rect 13495 32793 13507 32796
rect 13449 32787 13507 32793
rect 13541 32793 13553 32796
rect 13587 32793 13599 32827
rect 14016 32824 14044 32864
rect 18046 32852 18052 32904
rect 18104 32892 18110 32904
rect 18325 32895 18383 32901
rect 18325 32892 18337 32895
rect 18104 32864 18337 32892
rect 18104 32852 18110 32864
rect 18325 32861 18337 32864
rect 18371 32861 18383 32895
rect 18432 32892 18460 32932
rect 18509 32929 18521 32963
rect 18555 32960 18567 32963
rect 18690 32960 18696 32972
rect 18555 32932 18696 32960
rect 18555 32929 18567 32932
rect 18509 32923 18567 32929
rect 18690 32920 18696 32932
rect 18748 32960 18754 32972
rect 19061 32963 19119 32969
rect 19061 32960 19073 32963
rect 18748 32932 19073 32960
rect 18748 32920 18754 32932
rect 19061 32929 19073 32932
rect 19107 32929 19119 32963
rect 19242 32960 19248 32972
rect 19203 32932 19248 32960
rect 19061 32923 19119 32929
rect 19242 32920 19248 32932
rect 19300 32920 19306 32972
rect 19426 32920 19432 32972
rect 19484 32960 19490 32972
rect 21358 32960 21364 32972
rect 19484 32932 21220 32960
rect 21319 32932 21364 32960
rect 19484 32920 19490 32932
rect 18598 32892 18604 32904
rect 18432 32864 18604 32892
rect 18325 32855 18383 32861
rect 18598 32852 18604 32864
rect 18656 32852 18662 32904
rect 19613 32895 19671 32901
rect 19613 32861 19625 32895
rect 19659 32892 19671 32895
rect 20162 32892 20168 32904
rect 19659 32864 20168 32892
rect 19659 32861 19671 32864
rect 19613 32855 19671 32861
rect 20162 32852 20168 32864
rect 20220 32852 20226 32904
rect 21192 32892 21220 32932
rect 21358 32920 21364 32932
rect 21416 32920 21422 32972
rect 21542 32960 21548 32972
rect 21503 32932 21548 32960
rect 21542 32920 21548 32932
rect 21600 32920 21606 32972
rect 21867 32963 21925 32969
rect 21867 32929 21879 32963
rect 21913 32929 21925 32963
rect 22002 32960 22008 32972
rect 21963 32932 22008 32960
rect 21867 32923 21925 32929
rect 21882 32892 21910 32923
rect 22002 32920 22008 32932
rect 22060 32920 22066 32972
rect 24394 32960 24400 32972
rect 24355 32932 24400 32960
rect 24394 32920 24400 32932
rect 24452 32920 24458 32972
rect 24486 32920 24492 32972
rect 24544 32960 24550 32972
rect 24857 32963 24915 32969
rect 24857 32960 24869 32963
rect 24544 32932 24869 32960
rect 24544 32920 24550 32932
rect 24857 32929 24869 32932
rect 24903 32929 24915 32963
rect 24857 32923 24915 32929
rect 24949 32963 25007 32969
rect 24949 32929 24961 32963
rect 24995 32960 25007 32963
rect 26050 32960 26056 32972
rect 24995 32932 26056 32960
rect 24995 32929 25007 32932
rect 24949 32923 25007 32929
rect 26050 32920 26056 32932
rect 26108 32920 26114 32972
rect 27154 32920 27160 32972
rect 27212 32960 27218 32972
rect 38286 32960 38292 32972
rect 27212 32932 38292 32960
rect 27212 32920 27218 32932
rect 38286 32920 38292 32932
rect 38344 32920 38350 32972
rect 84010 32920 84016 32972
rect 84068 32960 84074 32972
rect 86678 32960 86684 32972
rect 84068 32932 86684 32960
rect 84068 32920 84074 32932
rect 86678 32920 86684 32932
rect 86736 32920 86742 32972
rect 21192 32864 21910 32892
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24210 32892 24216 32904
rect 23900 32864 24216 32892
rect 23900 32852 23906 32864
rect 24210 32852 24216 32864
rect 24268 32852 24274 32904
rect 25501 32895 25559 32901
rect 25501 32861 25513 32895
rect 25547 32892 25559 32895
rect 26326 32892 26332 32904
rect 25547 32864 26332 32892
rect 25547 32861 25559 32864
rect 25501 32855 25559 32861
rect 26326 32852 26332 32864
rect 26384 32852 26390 32904
rect 28810 32852 28816 32904
rect 28868 32892 28874 32904
rect 49326 32892 49332 32904
rect 28868 32864 49332 32892
rect 28868 32852 28874 32864
rect 49326 32852 49332 32864
rect 49384 32852 49390 32904
rect 56594 32824 56600 32836
rect 14016 32796 56600 32824
rect 13541 32787 13599 32793
rect 56594 32784 56600 32796
rect 56652 32784 56658 32836
rect 7561 32759 7619 32765
rect 7561 32725 7573 32759
rect 7607 32756 7619 32759
rect 7742 32756 7748 32768
rect 7607 32728 7748 32756
rect 7607 32725 7619 32728
rect 7561 32719 7619 32725
rect 7742 32716 7748 32728
rect 7800 32716 7806 32768
rect 8297 32759 8355 32765
rect 8297 32725 8309 32759
rect 8343 32756 8355 32759
rect 8662 32756 8668 32768
rect 8343 32728 8668 32756
rect 8343 32725 8355 32728
rect 8297 32719 8355 32725
rect 8662 32716 8668 32728
rect 8720 32716 8726 32768
rect 10042 32716 10048 32768
rect 10100 32756 10106 32768
rect 12526 32756 12532 32768
rect 10100 32728 12532 32756
rect 10100 32716 10106 32728
rect 12526 32716 12532 32728
rect 12584 32756 12590 32768
rect 12713 32759 12771 32765
rect 12713 32756 12725 32759
rect 12584 32728 12725 32756
rect 12584 32716 12590 32728
rect 12713 32725 12725 32728
rect 12759 32725 12771 32759
rect 13906 32756 13912 32768
rect 13867 32728 13912 32756
rect 12713 32719 12771 32725
rect 13906 32716 13912 32728
rect 13964 32716 13970 32768
rect 18046 32716 18052 32768
rect 18104 32756 18110 32768
rect 18141 32759 18199 32765
rect 18141 32756 18153 32759
rect 18104 32728 18153 32756
rect 18104 32716 18110 32728
rect 18141 32725 18153 32728
rect 18187 32725 18199 32759
rect 18141 32719 18199 32725
rect 19242 32716 19248 32768
rect 19300 32756 19306 32768
rect 19889 32759 19947 32765
rect 19889 32756 19901 32759
rect 19300 32728 19901 32756
rect 19300 32716 19306 32728
rect 19889 32725 19901 32728
rect 19935 32756 19947 32759
rect 20346 32756 20352 32768
rect 19935 32728 20352 32756
rect 19935 32725 19947 32728
rect 19889 32719 19947 32725
rect 20346 32716 20352 32728
rect 20404 32716 20410 32768
rect 24210 32716 24216 32768
rect 24268 32756 24274 32768
rect 25869 32759 25927 32765
rect 25869 32756 25881 32759
rect 24268 32728 25881 32756
rect 24268 32716 24274 32728
rect 25869 32725 25881 32728
rect 25915 32756 25927 32759
rect 27798 32756 27804 32768
rect 25915 32728 27804 32756
rect 25915 32725 25927 32728
rect 25869 32719 25927 32725
rect 27798 32716 27804 32728
rect 27856 32716 27862 32768
rect 28258 32716 28264 32768
rect 28316 32756 28322 32768
rect 49234 32756 49240 32768
rect 28316 32728 49240 32756
rect 28316 32716 28322 32728
rect 49234 32716 49240 32728
rect 49292 32716 49298 32768
rect 1104 32666 29256 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 29256 32666
rect 1104 32592 29256 32614
rect 32766 32580 32772 32632
rect 32824 32620 32830 32632
rect 49050 32620 49056 32632
rect 32824 32592 49056 32620
rect 32824 32580 32830 32592
rect 49050 32580 49056 32592
rect 49108 32580 49114 32632
rect 57977 32623 58035 32629
rect 57977 32589 57989 32623
rect 58023 32620 58035 32623
rect 58023 32592 67588 32620
rect 58023 32589 58035 32592
rect 57977 32583 58035 32589
rect 4433 32555 4491 32561
rect 4433 32552 4445 32555
rect 2608 32524 4445 32552
rect 2608 32425 2636 32524
rect 4433 32521 4445 32524
rect 4479 32552 4491 32555
rect 4798 32552 4804 32564
rect 4479 32524 4804 32552
rect 4479 32521 4491 32524
rect 4433 32515 4491 32521
rect 4798 32512 4804 32524
rect 4856 32552 4862 32564
rect 7926 32552 7932 32564
rect 4856 32524 7932 32552
rect 4856 32512 4862 32524
rect 2593 32419 2651 32425
rect 2593 32385 2605 32419
rect 2639 32385 2651 32419
rect 2593 32379 2651 32385
rect 2869 32419 2927 32425
rect 2869 32385 2881 32419
rect 2915 32416 2927 32419
rect 5626 32416 5632 32428
rect 2915 32388 5632 32416
rect 2915 32385 2927 32388
rect 2869 32379 2927 32385
rect 5626 32376 5632 32388
rect 5684 32376 5690 32428
rect 6840 32425 6868 32524
rect 7926 32512 7932 32524
rect 7984 32512 7990 32564
rect 8202 32552 8208 32564
rect 8163 32524 8208 32552
rect 8202 32512 8208 32524
rect 8260 32512 8266 32564
rect 8754 32512 8760 32564
rect 8812 32552 8818 32564
rect 17218 32552 17224 32564
rect 8812 32524 17224 32552
rect 8812 32512 8818 32524
rect 17218 32512 17224 32524
rect 17276 32512 17282 32564
rect 20070 32552 20076 32564
rect 18432 32524 20076 32552
rect 18432 32496 18460 32524
rect 20070 32512 20076 32524
rect 20128 32512 20134 32564
rect 22738 32512 22744 32564
rect 22796 32552 22802 32564
rect 26145 32555 26203 32561
rect 26145 32552 26157 32555
rect 22796 32524 26157 32552
rect 22796 32512 22802 32524
rect 26145 32521 26157 32524
rect 26191 32552 26203 32555
rect 26970 32552 26976 32564
rect 26191 32524 26976 32552
rect 26191 32521 26203 32524
rect 26145 32515 26203 32521
rect 26970 32512 26976 32524
rect 27028 32512 27034 32564
rect 27062 32512 27068 32564
rect 27120 32552 27126 32564
rect 55214 32552 55220 32564
rect 27120 32524 55220 32552
rect 27120 32512 27126 32524
rect 55214 32512 55220 32524
rect 55272 32512 55278 32564
rect 10042 32484 10048 32496
rect 7760 32456 10048 32484
rect 6825 32419 6883 32425
rect 6825 32385 6837 32419
rect 6871 32385 6883 32419
rect 7760 32416 7788 32456
rect 10042 32444 10048 32456
rect 10100 32444 10106 32496
rect 14734 32444 14740 32496
rect 14792 32484 14798 32496
rect 14829 32487 14887 32493
rect 14829 32484 14841 32487
rect 14792 32456 14841 32484
rect 14792 32444 14798 32456
rect 14829 32453 14841 32456
rect 14875 32484 14887 32487
rect 18414 32484 18420 32496
rect 14875 32456 18420 32484
rect 14875 32453 14887 32456
rect 14829 32447 14887 32453
rect 18414 32444 18420 32456
rect 18472 32444 18478 32496
rect 18966 32444 18972 32496
rect 19024 32484 19030 32496
rect 19426 32484 19432 32496
rect 19024 32456 19432 32484
rect 19024 32444 19030 32456
rect 19426 32444 19432 32456
rect 19484 32444 19490 32496
rect 46106 32484 46112 32496
rect 24688 32456 46112 32484
rect 6825 32379 6883 32385
rect 6932 32388 7788 32416
rect 5810 32240 5816 32292
rect 5868 32280 5874 32292
rect 6270 32280 6276 32292
rect 5868 32252 6276 32280
rect 5868 32240 5874 32252
rect 6270 32240 6276 32252
rect 6328 32240 6334 32292
rect 6546 32240 6552 32292
rect 6604 32280 6610 32292
rect 6932 32280 6960 32388
rect 8110 32376 8116 32428
rect 8168 32416 8174 32428
rect 12253 32419 12311 32425
rect 12253 32416 12265 32419
rect 8168 32388 12265 32416
rect 8168 32376 8174 32388
rect 12253 32385 12265 32388
rect 12299 32416 12311 32419
rect 23750 32416 23756 32428
rect 12299 32388 23756 32416
rect 12299 32385 12311 32388
rect 12253 32379 12311 32385
rect 7101 32351 7159 32357
rect 7101 32317 7113 32351
rect 7147 32348 7159 32351
rect 8018 32348 8024 32360
rect 7147 32320 8024 32348
rect 7147 32317 7159 32320
rect 7101 32311 7159 32317
rect 8018 32308 8024 32320
rect 8076 32308 8082 32360
rect 12897 32351 12955 32357
rect 12897 32317 12909 32351
rect 12943 32317 12955 32351
rect 12897 32311 12955 32317
rect 13081 32351 13139 32357
rect 13081 32317 13093 32351
rect 13127 32348 13139 32351
rect 13449 32351 13507 32357
rect 13127 32320 13308 32348
rect 13127 32317 13139 32320
rect 13081 32311 13139 32317
rect 6604 32252 6960 32280
rect 6604 32240 6610 32252
rect 7926 32240 7932 32292
rect 7984 32280 7990 32292
rect 8573 32283 8631 32289
rect 8573 32280 8585 32283
rect 7984 32252 8585 32280
rect 7984 32240 7990 32252
rect 8573 32249 8585 32252
rect 8619 32249 8631 32283
rect 8573 32243 8631 32249
rect 11977 32283 12035 32289
rect 11977 32249 11989 32283
rect 12023 32280 12035 32283
rect 12912 32280 12940 32311
rect 12986 32280 12992 32292
rect 12023 32252 12992 32280
rect 12023 32249 12035 32252
rect 11977 32243 12035 32249
rect 3970 32212 3976 32224
rect 3931 32184 3976 32212
rect 3970 32172 3976 32184
rect 4028 32172 4034 32224
rect 4982 32172 4988 32224
rect 5040 32212 5046 32224
rect 8202 32212 8208 32224
rect 5040 32184 8208 32212
rect 5040 32172 5046 32184
rect 8202 32172 8208 32184
rect 8260 32172 8266 32224
rect 8662 32172 8668 32224
rect 8720 32212 8726 32224
rect 11992 32212 12020 32243
rect 12986 32240 12992 32252
rect 13044 32240 13050 32292
rect 8720 32184 12020 32212
rect 8720 32172 8726 32184
rect 12066 32172 12072 32224
rect 12124 32212 12130 32224
rect 12529 32215 12587 32221
rect 12529 32212 12541 32215
rect 12124 32184 12541 32212
rect 12124 32172 12130 32184
rect 12529 32181 12541 32184
rect 12575 32181 12587 32215
rect 12529 32175 12587 32181
rect 12802 32172 12808 32224
rect 12860 32212 12866 32224
rect 13280 32212 13308 32320
rect 13449 32317 13461 32351
rect 13495 32348 13507 32351
rect 13538 32348 13544 32360
rect 13495 32320 13544 32348
rect 13495 32317 13507 32320
rect 13449 32311 13507 32317
rect 13538 32308 13544 32320
rect 13596 32308 13602 32360
rect 13648 32357 13676 32388
rect 23750 32376 23756 32388
rect 23808 32376 23814 32428
rect 23934 32376 23940 32428
rect 23992 32416 23998 32428
rect 24486 32416 24492 32428
rect 23992 32388 24492 32416
rect 23992 32376 23998 32388
rect 24486 32376 24492 32388
rect 24544 32376 24550 32428
rect 13633 32351 13691 32357
rect 13633 32317 13645 32351
rect 13679 32317 13691 32351
rect 13633 32311 13691 32317
rect 14645 32351 14703 32357
rect 14645 32317 14657 32351
rect 14691 32348 14703 32351
rect 15194 32348 15200 32360
rect 14691 32320 15200 32348
rect 14691 32317 14703 32320
rect 14645 32311 14703 32317
rect 15194 32308 15200 32320
rect 15252 32308 15258 32360
rect 18598 32308 18604 32360
rect 18656 32348 18662 32360
rect 19337 32351 19395 32357
rect 18656 32320 19012 32348
rect 18656 32308 18662 32320
rect 13722 32240 13728 32292
rect 13780 32280 13786 32292
rect 18984 32280 19012 32320
rect 19337 32317 19349 32351
rect 19383 32348 19395 32351
rect 19426 32348 19432 32360
rect 19383 32320 19432 32348
rect 19383 32317 19395 32320
rect 19337 32311 19395 32317
rect 19426 32308 19432 32320
rect 19484 32308 19490 32360
rect 19702 32308 19708 32360
rect 19760 32348 19766 32360
rect 19760 32320 19805 32348
rect 19760 32308 19766 32320
rect 21726 32308 21732 32360
rect 21784 32348 21790 32360
rect 24688 32348 24716 32456
rect 46106 32444 46112 32456
rect 46164 32444 46170 32496
rect 55122 32444 55128 32496
rect 55180 32484 55186 32496
rect 57931 32487 57989 32493
rect 57931 32484 57943 32487
rect 55180 32456 57943 32484
rect 55180 32444 55186 32456
rect 57931 32453 57943 32456
rect 57977 32453 57989 32487
rect 67560 32484 67588 32592
rect 72421 32487 72479 32493
rect 72421 32484 72433 32487
rect 67560 32456 72433 32484
rect 57931 32447 57989 32453
rect 72421 32453 72433 32456
rect 72467 32453 72479 32487
rect 72421 32447 72479 32453
rect 24854 32376 24860 32428
rect 24912 32416 24918 32428
rect 69014 32416 69020 32428
rect 24912 32388 69020 32416
rect 24912 32376 24918 32388
rect 69014 32376 69020 32388
rect 69072 32376 69078 32428
rect 21784 32320 24716 32348
rect 21784 32308 21790 32320
rect 24762 32308 24768 32360
rect 24820 32348 24826 32360
rect 24949 32351 25007 32357
rect 24949 32348 24961 32351
rect 24820 32320 24961 32348
rect 24820 32308 24826 32320
rect 24949 32317 24961 32320
rect 24995 32317 25007 32351
rect 24949 32311 25007 32317
rect 25222 32308 25228 32360
rect 25280 32348 25286 32360
rect 25590 32348 25596 32360
rect 25280 32320 25596 32348
rect 25280 32308 25286 32320
rect 25590 32308 25596 32320
rect 25648 32348 25654 32360
rect 26053 32351 26111 32357
rect 26053 32348 26065 32351
rect 25648 32320 26065 32348
rect 25648 32308 25654 32320
rect 26053 32317 26065 32320
rect 26099 32317 26111 32351
rect 26053 32311 26111 32317
rect 26970 32308 26976 32360
rect 27028 32348 27034 32360
rect 38010 32348 38016 32360
rect 27028 32320 38016 32348
rect 27028 32308 27034 32320
rect 38010 32308 38016 32320
rect 38068 32308 38074 32360
rect 19518 32280 19524 32292
rect 13780 32252 18920 32280
rect 18984 32252 19524 32280
rect 13780 32240 13786 32252
rect 14826 32212 14832 32224
rect 12860 32184 14832 32212
rect 12860 32172 12866 32184
rect 14826 32172 14832 32184
rect 14884 32212 14890 32224
rect 18782 32212 18788 32224
rect 14884 32184 18788 32212
rect 14884 32172 14890 32184
rect 18782 32172 18788 32184
rect 18840 32172 18846 32224
rect 18892 32212 18920 32252
rect 19518 32240 19524 32252
rect 19576 32240 19582 32292
rect 40034 32280 40040 32292
rect 20824 32252 40040 32280
rect 20824 32212 20852 32252
rect 40034 32240 40040 32252
rect 40092 32240 40098 32292
rect 20990 32212 20996 32224
rect 18892 32184 20852 32212
rect 20951 32184 20996 32212
rect 20990 32172 20996 32184
rect 21048 32172 21054 32224
rect 24670 32172 24676 32224
rect 24728 32212 24734 32224
rect 25133 32215 25191 32221
rect 25133 32212 25145 32215
rect 24728 32184 25145 32212
rect 24728 32172 24734 32184
rect 25133 32181 25145 32184
rect 25179 32181 25191 32215
rect 25133 32175 25191 32181
rect 72421 32147 72479 32153
rect 1104 32122 29256 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 29256 32122
rect 72421 32113 72433 32147
rect 72467 32144 72479 32147
rect 84010 32144 84016 32156
rect 72467 32116 84016 32144
rect 72467 32113 72479 32116
rect 72421 32107 72479 32113
rect 84010 32104 84016 32116
rect 84068 32104 84074 32156
rect 1104 32048 29256 32070
rect 4249 32011 4307 32017
rect 4249 31977 4261 32011
rect 4295 32008 4307 32011
rect 4614 32008 4620 32020
rect 4295 31980 4620 32008
rect 4295 31977 4307 31980
rect 4249 31971 4307 31977
rect 4614 31968 4620 31980
rect 4672 31968 4678 32020
rect 5994 31968 6000 32020
rect 6052 32008 6058 32020
rect 7009 32011 7067 32017
rect 7009 32008 7021 32011
rect 6052 31980 7021 32008
rect 6052 31968 6058 31980
rect 7009 31977 7021 31980
rect 7055 31977 7067 32011
rect 7009 31971 7067 31977
rect 7377 32011 7435 32017
rect 7377 31977 7389 32011
rect 7423 32008 7435 32011
rect 8110 32008 8116 32020
rect 7423 31980 8116 32008
rect 7423 31977 7435 31980
rect 7377 31971 7435 31977
rect 7392 31940 7420 31971
rect 8110 31968 8116 31980
rect 8168 31968 8174 32020
rect 8202 31968 8208 32020
rect 8260 32008 8266 32020
rect 16666 32008 16672 32020
rect 8260 31980 16672 32008
rect 8260 31968 8266 31980
rect 16666 31968 16672 31980
rect 16724 31968 16730 32020
rect 18046 32008 18052 32020
rect 18007 31980 18052 32008
rect 18046 31968 18052 31980
rect 18104 31968 18110 32020
rect 19797 32011 19855 32017
rect 19797 31977 19809 32011
rect 19843 32008 19855 32011
rect 21085 32011 21143 32017
rect 21085 32008 21097 32011
rect 19843 31980 21097 32008
rect 19843 31977 19855 31980
rect 19797 31971 19855 31977
rect 21085 31977 21097 31980
rect 21131 32008 21143 32011
rect 23474 32008 23480 32020
rect 21131 31980 23480 32008
rect 21131 31977 21143 31980
rect 21085 31971 21143 31977
rect 12710 31940 12716 31952
rect 7300 31912 7420 31940
rect 8128 31912 12716 31940
rect 4065 31875 4123 31881
rect 4065 31841 4077 31875
rect 4111 31872 4123 31875
rect 4614 31872 4620 31884
rect 4111 31844 4620 31872
rect 4111 31841 4123 31844
rect 4065 31835 4123 31841
rect 4614 31832 4620 31844
rect 4672 31832 4678 31884
rect 5810 31872 5816 31884
rect 5771 31844 5816 31872
rect 5810 31832 5816 31844
rect 5868 31832 5874 31884
rect 5997 31875 6055 31881
rect 5997 31841 6009 31875
rect 6043 31872 6055 31875
rect 6546 31872 6552 31884
rect 6043 31844 6552 31872
rect 6043 31841 6055 31844
rect 5997 31835 6055 31841
rect 6546 31832 6552 31844
rect 6604 31832 6610 31884
rect 6733 31875 6791 31881
rect 6733 31841 6745 31875
rect 6779 31872 6791 31875
rect 7300 31872 7328 31912
rect 6779 31844 7328 31872
rect 6779 31841 6791 31844
rect 6733 31835 6791 31841
rect 7374 31832 7380 31884
rect 7432 31872 7438 31884
rect 8021 31875 8079 31881
rect 8021 31872 8033 31875
rect 7432 31844 8033 31872
rect 7432 31832 7438 31844
rect 8021 31841 8033 31844
rect 8067 31841 8079 31875
rect 8021 31835 8079 31841
rect 3510 31696 3516 31748
rect 3568 31736 3574 31748
rect 8128 31736 8156 31912
rect 12710 31900 12716 31912
rect 12768 31900 12774 31952
rect 12986 31900 12992 31952
rect 13044 31940 13050 31952
rect 19702 31940 19708 31952
rect 13044 31912 19708 31940
rect 13044 31900 13050 31912
rect 19702 31900 19708 31912
rect 19760 31900 19766 31952
rect 11238 31832 11244 31884
rect 11296 31872 11302 31884
rect 12066 31872 12072 31884
rect 11296 31844 12072 31872
rect 11296 31832 11302 31844
rect 12066 31832 12072 31844
rect 12124 31832 12130 31884
rect 12802 31872 12808 31884
rect 12763 31844 12808 31872
rect 12802 31832 12808 31844
rect 12860 31832 12866 31884
rect 13173 31875 13231 31881
rect 13173 31841 13185 31875
rect 13219 31872 13231 31875
rect 18417 31875 18475 31881
rect 13219 31844 13308 31872
rect 13219 31841 13231 31844
rect 13173 31835 13231 31841
rect 8846 31764 8852 31816
rect 8904 31804 8910 31816
rect 12161 31807 12219 31813
rect 12161 31804 12173 31807
rect 8904 31776 12173 31804
rect 8904 31764 8910 31776
rect 12161 31773 12173 31776
rect 12207 31773 12219 31807
rect 12710 31804 12716 31816
rect 12671 31776 12716 31804
rect 12161 31767 12219 31773
rect 12710 31764 12716 31776
rect 12768 31764 12774 31816
rect 12986 31764 12992 31816
rect 13044 31804 13050 31816
rect 13081 31807 13139 31813
rect 13081 31804 13093 31807
rect 13044 31776 13093 31804
rect 13044 31764 13050 31776
rect 13081 31773 13093 31776
rect 13127 31773 13139 31807
rect 13081 31767 13139 31773
rect 3568 31708 8156 31736
rect 13280 31736 13308 31844
rect 18417 31841 18429 31875
rect 18463 31872 18475 31875
rect 18506 31872 18512 31884
rect 18463 31844 18512 31872
rect 18463 31841 18475 31844
rect 18417 31835 18475 31841
rect 18506 31832 18512 31844
rect 18564 31872 18570 31884
rect 18969 31875 19027 31881
rect 18969 31872 18981 31875
rect 18564 31844 18981 31872
rect 18564 31832 18570 31844
rect 18969 31841 18981 31844
rect 19015 31841 19027 31875
rect 19150 31872 19156 31884
rect 19063 31844 19156 31872
rect 18969 31835 19027 31841
rect 19150 31832 19156 31844
rect 19208 31872 19214 31884
rect 19812 31872 19840 31971
rect 23474 31968 23480 31980
rect 23532 31968 23538 32020
rect 24946 32008 24952 32020
rect 24907 31980 24952 32008
rect 24946 31968 24952 31980
rect 25004 31968 25010 32020
rect 27522 31968 27528 32020
rect 27580 32008 27586 32020
rect 27617 32011 27675 32017
rect 27617 32008 27629 32011
rect 27580 31980 27629 32008
rect 27580 31968 27586 31980
rect 27617 31977 27629 31980
rect 27663 32008 27675 32011
rect 48498 32008 48504 32020
rect 27663 31980 32812 32008
rect 27663 31977 27675 31980
rect 27617 31971 27675 31977
rect 20346 31900 20352 31952
rect 20404 31940 20410 31952
rect 22097 31943 22155 31949
rect 22097 31940 22109 31943
rect 20404 31912 22109 31940
rect 20404 31900 20410 31912
rect 22097 31909 22109 31912
rect 22143 31940 22155 31943
rect 22278 31940 22284 31952
rect 22143 31912 22284 31940
rect 22143 31909 22155 31912
rect 22097 31903 22155 31909
rect 22278 31900 22284 31912
rect 22336 31900 22342 31952
rect 27798 31940 27804 31952
rect 27759 31912 27804 31940
rect 27798 31900 27804 31912
rect 27856 31900 27862 31952
rect 32784 31940 32812 31980
rect 48424 31980 48504 32008
rect 48424 31940 48452 31980
rect 48498 31968 48504 31980
rect 48556 31968 48562 32020
rect 32784 31912 48452 31940
rect 20990 31872 20996 31884
rect 19208 31844 19840 31872
rect 20951 31844 20996 31872
rect 19208 31832 19214 31844
rect 20990 31832 20996 31844
rect 21048 31832 21054 31884
rect 21542 31832 21548 31884
rect 21600 31872 21606 31884
rect 22005 31875 22063 31881
rect 22005 31872 22017 31875
rect 21600 31844 22017 31872
rect 21600 31832 21606 31844
rect 22005 31841 22017 31844
rect 22051 31841 22063 31875
rect 22005 31835 22063 31841
rect 24946 31832 24952 31884
rect 25004 31872 25010 31884
rect 25041 31875 25099 31881
rect 25041 31872 25053 31875
rect 25004 31844 25053 31872
rect 25004 31832 25010 31844
rect 25041 31841 25053 31844
rect 25087 31841 25099 31875
rect 25041 31835 25099 31841
rect 27525 31875 27583 31881
rect 27525 31841 27537 31875
rect 27571 31841 27583 31875
rect 27525 31835 27583 31841
rect 13725 31807 13783 31813
rect 13725 31773 13737 31807
rect 13771 31804 13783 31807
rect 13814 31804 13820 31816
rect 13771 31776 13820 31804
rect 13771 31773 13783 31776
rect 13725 31767 13783 31773
rect 13814 31764 13820 31776
rect 13872 31764 13878 31816
rect 18046 31764 18052 31816
rect 18104 31804 18110 31816
rect 18233 31807 18291 31813
rect 18233 31804 18245 31807
rect 18104 31776 18245 31804
rect 18104 31764 18110 31776
rect 18233 31773 18245 31776
rect 18279 31773 18291 31807
rect 18233 31767 18291 31773
rect 20530 31764 20536 31816
rect 20588 31804 20594 31816
rect 27338 31804 27344 31816
rect 20588 31776 27344 31804
rect 20588 31764 20594 31776
rect 27338 31764 27344 31776
rect 27396 31764 27402 31816
rect 27540 31804 27568 31835
rect 27614 31832 27620 31884
rect 27672 31872 27678 31884
rect 27672 31844 29776 31872
rect 27672 31832 27678 31844
rect 27706 31804 27712 31816
rect 27540 31776 27712 31804
rect 27706 31764 27712 31776
rect 27764 31764 27770 31816
rect 29748 31804 29776 31844
rect 43070 31804 43076 31816
rect 29748 31776 43076 31804
rect 43070 31764 43076 31776
rect 43128 31764 43134 31816
rect 86865 31807 86923 31813
rect 86865 31804 86877 31807
rect 57992 31776 59124 31804
rect 13630 31736 13636 31748
rect 13280 31708 13636 31736
rect 3568 31696 3574 31708
rect 13630 31696 13636 31708
rect 13688 31696 13694 31748
rect 15194 31696 15200 31748
rect 15252 31736 15258 31748
rect 16482 31736 16488 31748
rect 15252 31708 16488 31736
rect 15252 31696 15258 31708
rect 16482 31696 16488 31708
rect 16540 31696 16546 31748
rect 19429 31739 19487 31745
rect 19429 31705 19441 31739
rect 19475 31736 19487 31739
rect 19886 31736 19892 31748
rect 19475 31708 19892 31736
rect 19475 31705 19487 31708
rect 19429 31699 19487 31705
rect 19886 31696 19892 31708
rect 19944 31696 19950 31748
rect 57992 31736 58020 31776
rect 24136 31708 58020 31736
rect 8570 31628 8576 31680
rect 8628 31668 8634 31680
rect 8846 31668 8852 31680
rect 8628 31640 8852 31668
rect 8628 31628 8634 31640
rect 8846 31628 8852 31640
rect 8904 31628 8910 31680
rect 12986 31628 12992 31680
rect 13044 31668 13050 31680
rect 13541 31671 13599 31677
rect 13541 31668 13553 31671
rect 13044 31640 13553 31668
rect 13044 31628 13050 31640
rect 13541 31637 13553 31640
rect 13587 31668 13599 31671
rect 13722 31668 13728 31680
rect 13587 31640 13728 31668
rect 13587 31637 13599 31640
rect 13541 31631 13599 31637
rect 13722 31628 13728 31640
rect 13780 31628 13786 31680
rect 16206 31628 16212 31680
rect 16264 31668 16270 31680
rect 24136 31668 24164 31708
rect 16264 31640 24164 31668
rect 16264 31628 16270 31640
rect 24578 31628 24584 31680
rect 24636 31668 24642 31680
rect 25225 31671 25283 31677
rect 25225 31668 25237 31671
rect 24636 31640 25237 31668
rect 24636 31628 24642 31640
rect 25225 31637 25237 31640
rect 25271 31668 25283 31671
rect 26786 31668 26792 31680
rect 25271 31640 26792 31668
rect 25271 31637 25283 31640
rect 25225 31631 25283 31637
rect 26786 31628 26792 31640
rect 26844 31628 26850 31680
rect 59096 31668 59124 31776
rect 77312 31776 86877 31804
rect 77312 31736 77340 31776
rect 86865 31773 86877 31776
rect 86911 31773 86923 31807
rect 86865 31767 86923 31773
rect 77220 31708 77340 31736
rect 77220 31668 77248 31708
rect 59096 31640 77248 31668
rect 59265 31603 59323 31609
rect 59265 31600 59277 31603
rect 1104 31578 29256 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 29256 31578
rect 1104 31504 29256 31526
rect 58452 31572 59277 31600
rect 4433 31467 4491 31473
rect 4433 31433 4445 31467
rect 4479 31464 4491 31467
rect 4890 31464 4896 31476
rect 4479 31436 4896 31464
rect 4479 31433 4491 31436
rect 4433 31427 4491 31433
rect 2866 31328 2872 31340
rect 2827 31300 2872 31328
rect 2866 31288 2872 31300
rect 2924 31288 2930 31340
rect 2593 31263 2651 31269
rect 2593 31229 2605 31263
rect 2639 31260 2651 31263
rect 4448 31260 4476 31427
rect 4890 31424 4896 31436
rect 4948 31424 4954 31476
rect 8018 31464 8024 31476
rect 7979 31436 8024 31464
rect 8018 31424 8024 31436
rect 8076 31424 8082 31476
rect 8389 31467 8447 31473
rect 8389 31433 8401 31467
rect 8435 31464 8447 31467
rect 8662 31464 8668 31476
rect 8435 31436 8668 31464
rect 8435 31433 8447 31436
rect 8389 31427 8447 31433
rect 7466 31356 7472 31408
rect 7524 31396 7530 31408
rect 7650 31396 7656 31408
rect 7524 31368 7656 31396
rect 7524 31356 7530 31368
rect 7650 31356 7656 31368
rect 7708 31356 7714 31408
rect 6270 31288 6276 31340
rect 6328 31328 6334 31340
rect 6917 31331 6975 31337
rect 6917 31328 6929 31331
rect 6328 31300 6929 31328
rect 6328 31288 6334 31300
rect 6917 31297 6929 31300
rect 6963 31297 6975 31331
rect 6917 31291 6975 31297
rect 2639 31232 4476 31260
rect 7009 31263 7067 31269
rect 2639 31229 2651 31232
rect 2593 31223 2651 31229
rect 7009 31229 7021 31263
rect 7055 31260 7067 31263
rect 7561 31263 7619 31269
rect 7561 31260 7573 31263
rect 7055 31232 7573 31260
rect 7055 31229 7067 31232
rect 7009 31223 7067 31229
rect 7561 31229 7573 31232
rect 7607 31260 7619 31263
rect 7650 31260 7656 31272
rect 7607 31232 7656 31260
rect 7607 31229 7619 31232
rect 7561 31223 7619 31229
rect 7650 31220 7656 31232
rect 7708 31220 7714 31272
rect 7745 31263 7803 31269
rect 7745 31229 7757 31263
rect 7791 31260 7803 31263
rect 8404 31260 8432 31427
rect 8662 31424 8668 31436
rect 8720 31424 8726 31476
rect 9585 31467 9643 31473
rect 9585 31433 9597 31467
rect 9631 31464 9643 31467
rect 9766 31464 9772 31476
rect 9631 31436 9772 31464
rect 9631 31433 9643 31436
rect 9585 31427 9643 31433
rect 9766 31424 9772 31436
rect 9824 31424 9830 31476
rect 19242 31424 19248 31476
rect 19300 31464 19306 31476
rect 33502 31464 33508 31476
rect 19300 31436 33508 31464
rect 19300 31424 19306 31436
rect 33502 31424 33508 31436
rect 33560 31424 33566 31476
rect 37277 31467 37335 31473
rect 37277 31433 37289 31467
rect 37323 31464 37335 31467
rect 46845 31467 46903 31473
rect 46845 31464 46857 31467
rect 37323 31436 46857 31464
rect 37323 31433 37335 31436
rect 37277 31427 37335 31433
rect 46845 31433 46857 31436
rect 46891 31433 46903 31467
rect 46845 31427 46903 31433
rect 7791 31232 8432 31260
rect 8496 31368 12848 31396
rect 7791 31229 7803 31232
rect 7745 31223 7803 31229
rect 5074 31152 5080 31204
rect 5132 31192 5138 31204
rect 8496 31192 8524 31368
rect 12820 31328 12848 31368
rect 12894 31356 12900 31408
rect 12952 31396 12958 31408
rect 13081 31399 13139 31405
rect 13081 31396 13093 31399
rect 12952 31368 13093 31396
rect 12952 31356 12958 31368
rect 13081 31365 13093 31368
rect 13127 31365 13139 31399
rect 13081 31359 13139 31365
rect 13170 31356 13176 31408
rect 13228 31396 13234 31408
rect 14185 31399 14243 31405
rect 14185 31396 14197 31399
rect 13228 31368 14197 31396
rect 13228 31356 13234 31368
rect 14185 31365 14197 31368
rect 14231 31365 14243 31399
rect 14185 31359 14243 31365
rect 23753 31399 23811 31405
rect 23753 31365 23765 31399
rect 23799 31396 23811 31399
rect 27338 31396 27344 31408
rect 23799 31368 27344 31396
rect 23799 31365 23811 31368
rect 23753 31359 23811 31365
rect 18046 31328 18052 31340
rect 12820 31300 18052 31328
rect 18046 31288 18052 31300
rect 18104 31288 18110 31340
rect 19426 31288 19432 31340
rect 19484 31288 19490 31340
rect 20162 31328 20168 31340
rect 20123 31300 20168 31328
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 21542 31328 21548 31340
rect 21503 31300 21548 31328
rect 21542 31288 21548 31300
rect 21600 31288 21606 31340
rect 9861 31263 9919 31269
rect 9861 31229 9873 31263
rect 9907 31229 9919 31263
rect 10042 31260 10048 31272
rect 10003 31232 10048 31260
rect 9861 31223 9919 31229
rect 9582 31192 9588 31204
rect 5132 31164 8524 31192
rect 9543 31164 9588 31192
rect 5132 31152 5138 31164
rect 9582 31152 9588 31164
rect 9640 31152 9646 31204
rect 4154 31124 4160 31136
rect 4115 31096 4160 31124
rect 4154 31084 4160 31096
rect 4212 31084 4218 31136
rect 9674 31124 9680 31136
rect 9635 31096 9680 31124
rect 9674 31084 9680 31096
rect 9732 31124 9738 31136
rect 9876 31124 9904 31223
rect 10042 31220 10048 31232
rect 10100 31220 10106 31272
rect 10597 31263 10655 31269
rect 10597 31229 10609 31263
rect 10643 31229 10655 31263
rect 10597 31223 10655 31229
rect 10781 31263 10839 31269
rect 10781 31229 10793 31263
rect 10827 31260 10839 31263
rect 12897 31263 12955 31269
rect 10827 31232 11468 31260
rect 10827 31229 10839 31232
rect 10781 31223 10839 31229
rect 10060 31192 10088 31220
rect 10612 31192 10640 31223
rect 11146 31192 11152 31204
rect 10060 31164 10640 31192
rect 11107 31164 11152 31192
rect 11146 31152 11152 31164
rect 11204 31152 11210 31204
rect 11440 31201 11468 31232
rect 12897 31229 12909 31263
rect 12943 31260 12955 31263
rect 13722 31260 13728 31272
rect 12943 31232 13728 31260
rect 12943 31229 12955 31232
rect 12897 31223 12955 31229
rect 13722 31220 13728 31232
rect 13780 31220 13786 31272
rect 14001 31263 14059 31269
rect 14001 31229 14013 31263
rect 14047 31260 14059 31263
rect 14047 31232 14504 31260
rect 14047 31229 14059 31232
rect 14001 31223 14059 31229
rect 11425 31195 11483 31201
rect 11425 31161 11437 31195
rect 11471 31192 11483 31195
rect 12986 31192 12992 31204
rect 11471 31164 12992 31192
rect 11471 31161 11483 31164
rect 11425 31155 11483 31161
rect 12986 31152 12992 31164
rect 13044 31152 13050 31204
rect 14476 31201 14504 31232
rect 16482 31220 16488 31272
rect 16540 31260 16546 31272
rect 18325 31263 18383 31269
rect 18325 31260 18337 31263
rect 16540 31232 18337 31260
rect 16540 31220 16546 31232
rect 18325 31229 18337 31232
rect 18371 31229 18383 31263
rect 19444 31260 19472 31288
rect 19797 31263 19855 31269
rect 19797 31260 19809 31263
rect 19444 31232 19809 31260
rect 18325 31223 18383 31229
rect 19797 31229 19809 31232
rect 19843 31260 19855 31263
rect 19889 31263 19947 31269
rect 19889 31260 19901 31263
rect 19843 31232 19901 31260
rect 19843 31229 19855 31232
rect 19797 31223 19855 31229
rect 19889 31229 19901 31232
rect 19935 31260 19947 31263
rect 20622 31260 20628 31272
rect 19935 31232 20628 31260
rect 19935 31229 19947 31232
rect 19889 31223 19947 31229
rect 20622 31220 20628 31232
rect 20680 31220 20686 31272
rect 23750 31220 23756 31272
rect 23808 31260 23814 31272
rect 23860 31269 23888 31368
rect 27338 31356 27344 31368
rect 27396 31356 27402 31408
rect 27522 31396 27528 31408
rect 27483 31368 27528 31396
rect 27522 31356 27528 31368
rect 27580 31356 27586 31408
rect 32030 31356 32036 31408
rect 32088 31396 32094 31408
rect 58452 31396 58480 31572
rect 59265 31569 59277 31572
rect 59311 31600 59323 31603
rect 59722 31600 59728 31612
rect 59311 31572 59728 31600
rect 59311 31569 59323 31572
rect 59265 31563 59323 31569
rect 59722 31560 59728 31572
rect 59780 31560 59786 31612
rect 86865 31603 86923 31609
rect 86865 31569 86877 31603
rect 86911 31600 86923 31603
rect 87138 31600 87144 31612
rect 86911 31572 87144 31600
rect 86911 31569 86923 31572
rect 86865 31563 86923 31569
rect 87138 31560 87144 31572
rect 87196 31600 87202 31612
rect 87874 31600 87880 31612
rect 87196 31572 87880 31600
rect 87196 31560 87202 31572
rect 87874 31560 87880 31572
rect 87932 31560 87938 31612
rect 59354 31492 59360 31544
rect 59412 31492 59418 31544
rect 32088 31368 58480 31396
rect 32088 31356 32094 31368
rect 24026 31288 24032 31340
rect 24084 31328 24090 31340
rect 25869 31331 25927 31337
rect 25869 31328 25881 31331
rect 24084 31300 25881 31328
rect 24084 31288 24090 31300
rect 25869 31297 25881 31300
rect 25915 31328 25927 31331
rect 25961 31331 26019 31337
rect 25961 31328 25973 31331
rect 25915 31300 25973 31328
rect 25915 31297 25927 31300
rect 25869 31291 25927 31297
rect 25961 31297 25973 31300
rect 26007 31297 26019 31331
rect 25961 31291 26019 31297
rect 23845 31263 23903 31269
rect 23845 31260 23857 31263
rect 23808 31232 23857 31260
rect 23808 31220 23814 31232
rect 23845 31229 23857 31232
rect 23891 31229 23903 31263
rect 23845 31223 23903 31229
rect 24670 31220 24676 31272
rect 24728 31260 24734 31272
rect 24946 31260 24952 31272
rect 24728 31232 24952 31260
rect 24728 31220 24734 31232
rect 24946 31220 24952 31232
rect 25004 31220 25010 31272
rect 26145 31263 26203 31269
rect 26145 31229 26157 31263
rect 26191 31260 26203 31263
rect 26697 31263 26755 31269
rect 26697 31260 26709 31263
rect 26191 31232 26709 31260
rect 26191 31229 26203 31232
rect 26145 31223 26203 31229
rect 26697 31229 26709 31232
rect 26743 31260 26755 31263
rect 26786 31260 26792 31272
rect 26743 31232 26792 31260
rect 26743 31229 26755 31232
rect 26697 31223 26755 31229
rect 26786 31220 26792 31232
rect 26844 31220 26850 31272
rect 26881 31263 26939 31269
rect 26881 31229 26893 31263
rect 26927 31260 26939 31263
rect 27540 31260 27568 31356
rect 32398 31288 32404 31340
rect 32456 31328 32462 31340
rect 59372 31328 59400 31492
rect 59541 31331 59599 31337
rect 59541 31328 59553 31331
rect 32456 31300 59553 31328
rect 32456 31288 32462 31300
rect 59541 31297 59553 31300
rect 59587 31297 59599 31331
rect 59541 31291 59599 31297
rect 41598 31260 41604 31272
rect 26927 31232 27568 31260
rect 32324 31232 41604 31260
rect 26927 31229 26939 31232
rect 26881 31223 26939 31229
rect 14461 31195 14519 31201
rect 14461 31161 14473 31195
rect 14507 31192 14519 31195
rect 16390 31192 16396 31204
rect 14507 31164 16396 31192
rect 14507 31161 14519 31164
rect 14461 31155 14519 31161
rect 16390 31152 16396 31164
rect 16448 31192 16454 31204
rect 19426 31192 19432 31204
rect 16448 31164 19432 31192
rect 16448 31152 16454 31164
rect 19426 31152 19432 31164
rect 19484 31152 19490 31204
rect 19628 31164 20024 31192
rect 9732 31096 9904 31124
rect 18509 31127 18567 31133
rect 9732 31084 9738 31096
rect 18509 31093 18521 31127
rect 18555 31124 18567 31127
rect 19628 31124 19656 31164
rect 18555 31096 19656 31124
rect 19996 31124 20024 31164
rect 20990 31152 20996 31204
rect 21048 31192 21054 31204
rect 28350 31192 28356 31204
rect 21048 31164 28356 31192
rect 21048 31152 21054 31164
rect 28350 31152 28356 31164
rect 28408 31152 28414 31204
rect 21542 31124 21548 31136
rect 19996 31096 21548 31124
rect 18555 31093 18567 31096
rect 18509 31087 18567 31093
rect 21542 31084 21548 31096
rect 21600 31084 21606 31136
rect 23934 31124 23940 31136
rect 23895 31096 23940 31124
rect 23934 31084 23940 31096
rect 23992 31084 23998 31136
rect 26786 31084 26792 31136
rect 26844 31124 26850 31136
rect 27157 31127 27215 31133
rect 27157 31124 27169 31127
rect 26844 31096 27169 31124
rect 26844 31084 26850 31096
rect 27157 31093 27169 31096
rect 27203 31093 27215 31127
rect 27157 31087 27215 31093
rect 27338 31084 27344 31136
rect 27396 31124 27402 31136
rect 32324 31124 32352 31232
rect 41598 31220 41604 31232
rect 41656 31220 41662 31272
rect 48317 31263 48375 31269
rect 48317 31229 48329 31263
rect 48363 31260 48375 31263
rect 56594 31260 56600 31272
rect 48363 31232 56600 31260
rect 48363 31229 48375 31232
rect 48317 31223 48375 31229
rect 56594 31220 56600 31232
rect 56652 31220 56658 31272
rect 32674 31152 32680 31204
rect 32732 31192 32738 31204
rect 48409 31195 48467 31201
rect 32732 31164 48268 31192
rect 32732 31152 32738 31164
rect 48240 31133 48268 31164
rect 48409 31161 48421 31195
rect 48455 31192 48467 31195
rect 87230 31192 87236 31204
rect 48455 31164 87236 31192
rect 48455 31161 48467 31164
rect 48409 31155 48467 31161
rect 87230 31152 87236 31164
rect 87288 31152 87294 31204
rect 87325 31195 87383 31201
rect 87325 31161 87337 31195
rect 87371 31192 87383 31195
rect 96525 31195 96583 31201
rect 96525 31192 96537 31195
rect 87371 31164 96537 31192
rect 87371 31161 87383 31164
rect 87325 31155 87383 31161
rect 96525 31161 96537 31164
rect 96571 31161 96583 31195
rect 96525 31155 96583 31161
rect 37277 31127 37335 31133
rect 37277 31124 37289 31127
rect 27396 31096 32352 31124
rect 32416 31096 37289 31124
rect 27396 31084 27402 31096
rect 1104 31034 29256 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 29256 31034
rect 1104 30960 29256 30982
rect 2869 30923 2927 30929
rect 2869 30889 2881 30923
rect 2915 30920 2927 30923
rect 2958 30920 2964 30932
rect 2915 30892 2964 30920
rect 2915 30889 2927 30892
rect 2869 30883 2927 30889
rect 2958 30880 2964 30892
rect 3016 30880 3022 30932
rect 4985 30923 5043 30929
rect 4985 30889 4997 30923
rect 5031 30920 5043 30923
rect 20346 30920 20352 30932
rect 5031 30892 20352 30920
rect 5031 30889 5043 30892
rect 4985 30883 5043 30889
rect 2774 30744 2780 30796
rect 2832 30784 2838 30796
rect 2976 30793 3004 30880
rect 2961 30787 3019 30793
rect 2961 30784 2973 30787
rect 2832 30756 2973 30784
rect 2832 30744 2838 30756
rect 2961 30753 2973 30756
rect 3007 30753 3019 30787
rect 2961 30747 3019 30753
rect 3970 30744 3976 30796
rect 4028 30784 4034 30796
rect 4157 30787 4215 30793
rect 4157 30784 4169 30787
rect 4028 30756 4169 30784
rect 4028 30744 4034 30756
rect 4157 30753 4169 30756
rect 4203 30753 4215 30787
rect 4157 30747 4215 30753
rect 4617 30787 4675 30793
rect 4617 30753 4629 30787
rect 4663 30784 4675 30787
rect 5000 30784 5028 30883
rect 20346 30880 20352 30892
rect 20404 30880 20410 30932
rect 20438 30880 20444 30932
rect 20496 30920 20502 30932
rect 25958 30920 25964 30932
rect 20496 30892 25964 30920
rect 20496 30880 20502 30892
rect 25958 30880 25964 30892
rect 26016 30880 26022 30932
rect 27706 30880 27712 30932
rect 27764 30920 27770 30932
rect 27893 30923 27951 30929
rect 27893 30920 27905 30923
rect 27764 30892 27905 30920
rect 27764 30880 27770 30892
rect 27893 30889 27905 30892
rect 27939 30889 27951 30923
rect 27893 30883 27951 30889
rect 6549 30855 6607 30861
rect 6549 30821 6561 30855
rect 6595 30852 6607 30855
rect 9582 30852 9588 30864
rect 6595 30824 9588 30852
rect 6595 30821 6607 30824
rect 6549 30815 6607 30821
rect 4663 30756 5028 30784
rect 5629 30787 5687 30793
rect 4663 30753 4675 30756
rect 4617 30747 4675 30753
rect 5629 30753 5641 30787
rect 5675 30753 5687 30787
rect 5629 30747 5687 30753
rect 6181 30787 6239 30793
rect 6181 30753 6193 30787
rect 6227 30784 6239 30787
rect 6564 30784 6592 30815
rect 9582 30812 9588 30824
rect 9640 30812 9646 30864
rect 12158 30812 12164 30864
rect 12216 30852 12222 30864
rect 16117 30855 16175 30861
rect 16117 30852 16129 30855
rect 12216 30824 16129 30852
rect 12216 30812 12222 30824
rect 16117 30821 16129 30824
rect 16163 30821 16175 30855
rect 16117 30815 16175 30821
rect 17221 30855 17279 30861
rect 17221 30821 17233 30855
rect 17267 30852 17279 30855
rect 17770 30852 17776 30864
rect 17267 30824 17776 30852
rect 17267 30821 17279 30824
rect 17221 30815 17279 30821
rect 6227 30756 6592 30784
rect 6227 30753 6239 30756
rect 6181 30747 6239 30753
rect 4172 30648 4200 30747
rect 4706 30716 4712 30728
rect 4667 30688 4712 30716
rect 4706 30676 4712 30688
rect 4764 30676 4770 30728
rect 5644 30648 5672 30747
rect 7742 30744 7748 30796
rect 7800 30784 7806 30796
rect 10505 30787 10563 30793
rect 10505 30784 10517 30787
rect 7800 30756 10517 30784
rect 7800 30744 7806 30756
rect 10505 30753 10517 30756
rect 10551 30753 10563 30787
rect 10505 30747 10563 30753
rect 10781 30787 10839 30793
rect 10781 30753 10793 30787
rect 10827 30784 10839 30787
rect 11054 30784 11060 30796
rect 10827 30756 11060 30784
rect 10827 30753 10839 30756
rect 10781 30747 10839 30753
rect 6089 30719 6147 30725
rect 6089 30685 6101 30719
rect 6135 30685 6147 30719
rect 10520 30716 10548 30747
rect 11054 30744 11060 30756
rect 11112 30744 11118 30796
rect 12253 30787 12311 30793
rect 12253 30784 12265 30787
rect 11164 30756 12265 30784
rect 11164 30716 11192 30756
rect 12253 30753 12265 30756
rect 12299 30784 12311 30787
rect 13354 30784 13360 30796
rect 12299 30756 13360 30784
rect 12299 30753 12311 30756
rect 12253 30747 12311 30753
rect 13354 30744 13360 30756
rect 13412 30744 13418 30796
rect 13449 30787 13507 30793
rect 13449 30753 13461 30787
rect 13495 30753 13507 30787
rect 13722 30784 13728 30796
rect 13683 30756 13728 30784
rect 13449 30747 13507 30753
rect 10520 30688 11192 30716
rect 12161 30719 12219 30725
rect 6089 30679 6147 30685
rect 12161 30685 12173 30719
rect 12207 30716 12219 30719
rect 12894 30716 12900 30728
rect 12207 30688 12900 30716
rect 12207 30685 12219 30688
rect 12161 30679 12219 30685
rect 5718 30648 5724 30660
rect 4172 30620 5724 30648
rect 5718 30608 5724 30620
rect 5776 30608 5782 30660
rect 3053 30583 3111 30589
rect 3053 30549 3065 30583
rect 3099 30580 3111 30583
rect 4614 30580 4620 30592
rect 3099 30552 4620 30580
rect 3099 30549 3111 30552
rect 3053 30543 3111 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 4890 30540 4896 30592
rect 4948 30580 4954 30592
rect 6104 30580 6132 30679
rect 12894 30676 12900 30688
rect 12952 30676 12958 30728
rect 13464 30716 13492 30747
rect 13722 30744 13728 30756
rect 13780 30744 13786 30796
rect 15010 30716 15016 30728
rect 13464 30688 15016 30716
rect 15010 30676 15016 30688
rect 15068 30676 15074 30728
rect 16132 30716 16160 30815
rect 17770 30812 17776 30824
rect 17828 30812 17834 30864
rect 18046 30852 18052 30864
rect 18007 30824 18052 30852
rect 18046 30812 18052 30824
rect 18104 30812 18110 30864
rect 18966 30812 18972 30864
rect 19024 30852 19030 30864
rect 19024 30824 19104 30852
rect 19024 30812 19030 30824
rect 16298 30744 16304 30796
rect 16356 30784 16362 30796
rect 16485 30787 16543 30793
rect 16485 30784 16497 30787
rect 16356 30756 16497 30784
rect 16356 30744 16362 30756
rect 16485 30753 16497 30756
rect 16531 30753 16543 30787
rect 16485 30747 16543 30753
rect 16632 30787 16690 30793
rect 16632 30753 16644 30787
rect 16678 30784 16690 30787
rect 16758 30784 16764 30796
rect 16678 30756 16764 30784
rect 16678 30753 16690 30756
rect 16632 30747 16690 30753
rect 16758 30744 16764 30756
rect 16816 30744 16822 30796
rect 18693 30787 18751 30793
rect 18693 30753 18705 30787
rect 18739 30784 18751 30787
rect 18874 30784 18880 30796
rect 18739 30756 18880 30784
rect 18739 30753 18751 30756
rect 18693 30747 18751 30753
rect 18874 30744 18880 30756
rect 18932 30744 18938 30796
rect 19076 30793 19104 30824
rect 19150 30812 19156 30864
rect 19208 30852 19214 30864
rect 19208 30824 19288 30852
rect 19208 30812 19214 30824
rect 19260 30793 19288 30824
rect 21634 30812 21640 30864
rect 21692 30852 21698 30864
rect 22646 30852 22652 30864
rect 21692 30824 22652 30852
rect 21692 30812 21698 30824
rect 22646 30812 22652 30824
rect 22704 30852 22710 30864
rect 24026 30852 24032 30864
rect 22704 30824 24032 30852
rect 22704 30812 22710 30824
rect 24026 30812 24032 30824
rect 24084 30812 24090 30864
rect 25590 30852 25596 30864
rect 25551 30824 25596 30852
rect 25590 30812 25596 30824
rect 25648 30812 25654 30864
rect 27522 30812 27528 30864
rect 27580 30852 27586 30864
rect 32416 30852 32444 31096
rect 37277 31093 37289 31096
rect 37323 31093 37335 31127
rect 37277 31087 37335 31093
rect 46843 31127 46901 31133
rect 46843 31093 46855 31127
rect 46889 31124 46901 31127
rect 48133 31127 48191 31133
rect 48133 31124 48145 31127
rect 46889 31096 48145 31124
rect 46889 31093 46901 31096
rect 46843 31087 46901 31093
rect 48133 31093 48145 31096
rect 48179 31093 48191 31127
rect 48133 31087 48191 31093
rect 48225 31127 48283 31133
rect 48225 31093 48237 31127
rect 48271 31093 48283 31127
rect 48225 31087 48283 31093
rect 86862 31084 86868 31136
rect 86920 31124 86926 31136
rect 87414 31124 87420 31136
rect 86920 31096 87420 31124
rect 86920 31084 86926 31096
rect 87414 31084 87420 31096
rect 87472 31084 87478 31136
rect 32490 31016 32496 31068
rect 32548 31056 32554 31068
rect 86126 31056 86132 31068
rect 32548 31028 86132 31056
rect 32548 31016 32554 31028
rect 86126 31016 86132 31028
rect 86184 31056 86190 31068
rect 86954 31056 86960 31068
rect 86184 31028 86960 31056
rect 86184 31016 86190 31028
rect 86954 31016 86960 31028
rect 87012 31016 87018 31068
rect 108298 31056 108304 31068
rect 100588 31028 108304 31056
rect 32582 30948 32588 31000
rect 32640 30988 32646 31000
rect 96525 30991 96583 30997
rect 32640 30960 86172 30988
rect 32640 30948 32646 30960
rect 86144 30920 86172 30960
rect 96525 30957 96537 30991
rect 96571 30988 96583 30991
rect 99285 30991 99343 30997
rect 99285 30988 99297 30991
rect 96571 30960 99297 30988
rect 96571 30957 96583 30960
rect 96525 30951 96583 30957
rect 99285 30957 99297 30960
rect 99331 30957 99343 30991
rect 99285 30951 99343 30957
rect 99377 30991 99435 30997
rect 99377 30957 99389 30991
rect 99423 30988 99435 30991
rect 100588 30988 100616 31028
rect 108298 31016 108304 31028
rect 108356 31016 108362 31068
rect 99423 30960 100616 30988
rect 99423 30957 99435 30960
rect 99377 30951 99435 30957
rect 87046 30920 87052 30932
rect 86144 30892 87052 30920
rect 87046 30880 87052 30892
rect 87104 30880 87110 30932
rect 27580 30824 32444 30852
rect 27580 30812 27586 30824
rect 86218 30812 86224 30864
rect 86276 30852 86282 30864
rect 87325 30855 87383 30861
rect 87325 30852 87337 30855
rect 86276 30824 87337 30852
rect 86276 30812 86282 30824
rect 87325 30821 87337 30824
rect 87371 30821 87383 30855
rect 87325 30815 87383 30821
rect 19061 30787 19119 30793
rect 19061 30753 19073 30787
rect 19107 30753 19119 30787
rect 19061 30747 19119 30753
rect 19245 30787 19303 30793
rect 19245 30753 19257 30787
rect 19291 30784 19303 30787
rect 19337 30787 19395 30793
rect 19337 30784 19349 30787
rect 19291 30756 19349 30784
rect 19291 30753 19303 30756
rect 19245 30747 19303 30753
rect 19337 30753 19349 30756
rect 19383 30753 19395 30787
rect 19337 30747 19395 30753
rect 23937 30787 23995 30793
rect 23937 30753 23949 30787
rect 23983 30784 23995 30787
rect 25222 30784 25228 30796
rect 23983 30756 25228 30784
rect 23983 30753 23995 30756
rect 23937 30747 23995 30753
rect 25222 30744 25228 30756
rect 25280 30784 25286 30796
rect 25685 30787 25743 30793
rect 25685 30784 25697 30787
rect 25280 30756 25697 30784
rect 25280 30744 25286 30756
rect 25685 30753 25697 30756
rect 25731 30753 25743 30787
rect 26786 30784 26792 30796
rect 26747 30756 26792 30784
rect 25685 30747 25743 30753
rect 26786 30744 26792 30756
rect 26844 30744 26850 30796
rect 16853 30719 16911 30725
rect 16853 30716 16865 30719
rect 16132 30688 16865 30716
rect 16853 30685 16865 30688
rect 16899 30685 16911 30719
rect 16853 30679 16911 30685
rect 18785 30719 18843 30725
rect 18785 30685 18797 30719
rect 18831 30716 18843 30719
rect 19521 30719 19579 30725
rect 19521 30716 19533 30719
rect 18831 30688 19533 30716
rect 18831 30685 18843 30688
rect 18785 30679 18843 30685
rect 19076 30660 19104 30688
rect 19521 30685 19533 30688
rect 19567 30685 19579 30719
rect 19521 30679 19579 30685
rect 23474 30676 23480 30728
rect 23532 30716 23538 30728
rect 24213 30719 24271 30725
rect 24213 30716 24225 30719
rect 23532 30688 24225 30716
rect 23532 30676 23538 30688
rect 24213 30685 24225 30688
rect 24259 30685 24271 30719
rect 24213 30679 24271 30685
rect 26513 30719 26571 30725
rect 26513 30685 26525 30719
rect 26559 30685 26571 30719
rect 26513 30679 26571 30685
rect 19058 30608 19064 30660
rect 19116 30608 19122 30660
rect 4948 30552 6132 30580
rect 4948 30540 4954 30552
rect 9214 30540 9220 30592
rect 9272 30580 9278 30592
rect 12158 30580 12164 30592
rect 9272 30552 12164 30580
rect 9272 30540 9278 30552
rect 12158 30540 12164 30552
rect 12216 30540 12222 30592
rect 13265 30583 13323 30589
rect 13265 30549 13277 30583
rect 13311 30580 13323 30583
rect 13354 30580 13360 30592
rect 13311 30552 13360 30580
rect 13311 30549 13323 30552
rect 13265 30543 13323 30549
rect 13354 30540 13360 30552
rect 13412 30540 13418 30592
rect 13909 30583 13967 30589
rect 13909 30549 13921 30583
rect 13955 30580 13967 30583
rect 15194 30580 15200 30592
rect 13955 30552 15200 30580
rect 13955 30549 13967 30552
rect 13909 30543 13967 30549
rect 15194 30540 15200 30552
rect 15252 30540 15258 30592
rect 16393 30583 16451 30589
rect 16393 30549 16405 30583
rect 16439 30580 16451 30583
rect 16666 30580 16672 30592
rect 16439 30552 16672 30580
rect 16439 30549 16451 30552
rect 16393 30543 16451 30549
rect 16666 30540 16672 30552
rect 16724 30580 16730 30592
rect 16761 30583 16819 30589
rect 16761 30580 16773 30583
rect 16724 30552 16773 30580
rect 16724 30540 16730 30552
rect 16761 30549 16773 30552
rect 16807 30549 16819 30583
rect 26528 30580 26556 30679
rect 26970 30580 26976 30592
rect 26528 30552 26976 30580
rect 16761 30543 16819 30549
rect 26970 30540 26976 30552
rect 27028 30580 27034 30592
rect 27246 30580 27252 30592
rect 27028 30552 27252 30580
rect 27028 30540 27034 30552
rect 27246 30540 27252 30552
rect 27304 30580 27310 30592
rect 28261 30583 28319 30589
rect 28261 30580 28273 30583
rect 27304 30552 28273 30580
rect 27304 30540 27310 30552
rect 28261 30549 28273 30552
rect 28307 30549 28319 30583
rect 28261 30543 28319 30549
rect 1104 30490 29256 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 29256 30490
rect 1104 30416 29256 30438
rect 4614 30336 4620 30388
rect 4672 30376 4678 30388
rect 5718 30376 5724 30388
rect 4672 30348 4936 30376
rect 5679 30348 5724 30376
rect 4672 30336 4678 30348
rect 3142 30268 3148 30320
rect 3200 30308 3206 30320
rect 3200 30280 4476 30308
rect 3200 30268 3206 30280
rect 3970 30240 3976 30252
rect 2700 30212 3976 30240
rect 2700 30184 2728 30212
rect 3970 30200 3976 30212
rect 4028 30240 4034 30252
rect 4448 30249 4476 30280
rect 4433 30243 4491 30249
rect 4028 30212 4200 30240
rect 4028 30200 4034 30212
rect 2682 30172 2688 30184
rect 2595 30144 2688 30172
rect 2682 30132 2688 30144
rect 2740 30132 2746 30184
rect 4172 30181 4200 30212
rect 4433 30209 4445 30243
rect 4479 30209 4491 30243
rect 4433 30203 4491 30209
rect 2961 30175 3019 30181
rect 2961 30141 2973 30175
rect 3007 30141 3019 30175
rect 2961 30135 3019 30141
rect 4157 30175 4215 30181
rect 4157 30141 4169 30175
rect 4203 30141 4215 30175
rect 4522 30172 4528 30184
rect 4483 30144 4528 30172
rect 4157 30135 4215 30141
rect 2976 30036 3004 30135
rect 4522 30132 4528 30144
rect 4580 30132 4586 30184
rect 4908 30172 4936 30348
rect 5718 30336 5724 30348
rect 5776 30336 5782 30388
rect 7650 30336 7656 30388
rect 7708 30376 7714 30388
rect 10594 30376 10600 30388
rect 7708 30348 10600 30376
rect 7708 30336 7714 30348
rect 10594 30336 10600 30348
rect 10652 30376 10658 30388
rect 13170 30376 13176 30388
rect 10652 30348 13176 30376
rect 10652 30336 10658 30348
rect 13170 30336 13176 30348
rect 13228 30336 13234 30388
rect 13541 30379 13599 30385
rect 13541 30345 13553 30379
rect 13587 30376 13599 30379
rect 13814 30376 13820 30388
rect 13587 30348 13820 30376
rect 13587 30345 13599 30348
rect 13541 30339 13599 30345
rect 11054 30308 11060 30320
rect 11015 30280 11060 30308
rect 11054 30268 11060 30280
rect 11112 30268 11118 30320
rect 11425 30311 11483 30317
rect 11425 30277 11437 30311
rect 11471 30308 11483 30311
rect 13556 30308 13584 30339
rect 13814 30336 13820 30348
rect 13872 30336 13878 30388
rect 16209 30379 16267 30385
rect 16209 30345 16221 30379
rect 16255 30376 16267 30379
rect 16298 30376 16304 30388
rect 16255 30348 16304 30376
rect 16255 30345 16267 30348
rect 16209 30339 16267 30345
rect 16298 30336 16304 30348
rect 16356 30336 16362 30388
rect 16500 30348 18552 30376
rect 11471 30280 13584 30308
rect 11471 30277 11483 30280
rect 11425 30271 11483 30277
rect 5166 30172 5172 30184
rect 4908 30144 5172 30172
rect 5166 30132 5172 30144
rect 5224 30172 5230 30184
rect 5537 30175 5595 30181
rect 5537 30172 5549 30175
rect 5224 30144 5549 30172
rect 5224 30132 5230 30144
rect 5537 30141 5549 30144
rect 5583 30141 5595 30175
rect 5537 30135 5595 30141
rect 9674 30132 9680 30184
rect 9732 30172 9738 30184
rect 9861 30175 9919 30181
rect 9861 30172 9873 30175
rect 9732 30144 9873 30172
rect 9732 30132 9738 30144
rect 9861 30141 9873 30144
rect 9907 30141 9919 30175
rect 9861 30135 9919 30141
rect 10045 30175 10103 30181
rect 10045 30141 10057 30175
rect 10091 30172 10103 30175
rect 10594 30172 10600 30184
rect 10091 30144 10600 30172
rect 10091 30141 10103 30144
rect 10045 30135 10103 30141
rect 10594 30132 10600 30144
rect 10652 30132 10658 30184
rect 10781 30175 10839 30181
rect 10781 30141 10793 30175
rect 10827 30172 10839 30175
rect 11440 30172 11468 30271
rect 11514 30200 11520 30252
rect 11572 30240 11578 30252
rect 16500 30240 16528 30348
rect 17218 30308 17224 30320
rect 11572 30212 16528 30240
rect 16592 30280 17224 30308
rect 11572 30200 11578 30212
rect 10827 30144 11468 30172
rect 10827 30141 10839 30144
rect 10781 30135 10839 30141
rect 12066 30132 12072 30184
rect 12124 30172 12130 30184
rect 12437 30175 12495 30181
rect 12437 30172 12449 30175
rect 12124 30144 12449 30172
rect 12124 30132 12130 30144
rect 12437 30141 12449 30144
rect 12483 30141 12495 30175
rect 12437 30135 12495 30141
rect 12894 30132 12900 30184
rect 12952 30172 12958 30184
rect 13449 30175 13507 30181
rect 13449 30172 13461 30175
rect 12952 30144 13461 30172
rect 12952 30132 12958 30144
rect 13449 30141 13461 30144
rect 13495 30141 13507 30175
rect 13449 30135 13507 30141
rect 15197 30175 15255 30181
rect 15197 30141 15209 30175
rect 15243 30141 15255 30175
rect 15197 30135 15255 30141
rect 3145 30107 3203 30113
rect 3145 30073 3157 30107
rect 3191 30104 3203 30107
rect 3786 30104 3792 30116
rect 3191 30076 3792 30104
rect 3191 30073 3203 30076
rect 3145 30067 3203 30073
rect 3786 30064 3792 30076
rect 3844 30064 3850 30116
rect 14458 30104 14464 30116
rect 3988 30076 14464 30104
rect 3329 30039 3387 30045
rect 3329 30036 3341 30039
rect 2976 30008 3341 30036
rect 3329 30005 3341 30008
rect 3375 30036 3387 30039
rect 3988 30036 4016 30076
rect 14458 30064 14464 30076
rect 14516 30064 14522 30116
rect 15212 30104 15240 30135
rect 15286 30132 15292 30184
rect 15344 30172 15350 30184
rect 16592 30181 16620 30280
rect 17218 30268 17224 30280
rect 17276 30268 17282 30320
rect 17681 30311 17739 30317
rect 17681 30277 17693 30311
rect 17727 30308 17739 30311
rect 18325 30311 18383 30317
rect 18325 30308 18337 30311
rect 17727 30280 18337 30308
rect 17727 30277 17739 30280
rect 17681 30271 17739 30277
rect 18325 30277 18337 30280
rect 18371 30277 18383 30311
rect 18524 30308 18552 30348
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 25038 30376 25044 30388
rect 19484 30348 25044 30376
rect 19484 30336 19490 30348
rect 19334 30308 19340 30320
rect 18524 30280 19340 30308
rect 18325 30271 18383 30277
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 19812 30317 19840 30348
rect 25038 30336 25044 30348
rect 25096 30336 25102 30388
rect 19797 30311 19855 30317
rect 19797 30277 19809 30311
rect 19843 30277 19855 30311
rect 19797 30271 19855 30277
rect 21082 30268 21088 30320
rect 21140 30308 21146 30320
rect 23661 30311 23719 30317
rect 23661 30308 23673 30311
rect 21140 30280 23673 30308
rect 21140 30268 21146 30280
rect 23661 30277 23673 30280
rect 23707 30308 23719 30311
rect 23707 30280 23888 30308
rect 23707 30277 23719 30280
rect 23661 30271 23719 30277
rect 16758 30200 16764 30252
rect 16816 30240 16822 30252
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 16816 30212 16865 30240
rect 16816 30200 16822 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 17494 30240 17500 30252
rect 16853 30203 16911 30209
rect 16960 30212 17500 30240
rect 16960 30181 16988 30212
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 18230 30249 18236 30252
rect 18196 30243 18236 30249
rect 18196 30209 18208 30243
rect 18196 30203 18236 30209
rect 18230 30200 18236 30203
rect 18288 30200 18294 30252
rect 18414 30200 18420 30252
rect 18472 30240 18478 30252
rect 21269 30243 21327 30249
rect 18472 30212 18517 30240
rect 18472 30200 18478 30212
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 21453 30243 21511 30249
rect 21453 30240 21465 30243
rect 21315 30212 21465 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 21453 30209 21465 30212
rect 21499 30240 21511 30243
rect 21634 30240 21640 30252
rect 21499 30212 21640 30240
rect 21499 30209 21511 30212
rect 21453 30203 21511 30209
rect 21634 30200 21640 30212
rect 21692 30200 21698 30252
rect 22649 30243 22707 30249
rect 22649 30209 22661 30243
rect 22695 30240 22707 30243
rect 23474 30240 23480 30252
rect 22695 30212 23480 30240
rect 22695 30209 22707 30212
rect 22649 30203 22707 30209
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 23860 30249 23888 30280
rect 24486 30268 24492 30320
rect 24544 30308 24550 30320
rect 25409 30311 25467 30317
rect 25409 30308 25421 30311
rect 24544 30280 25421 30308
rect 24544 30268 24550 30280
rect 25409 30277 25421 30280
rect 25455 30308 25467 30311
rect 28810 30308 28816 30320
rect 25455 30280 28816 30308
rect 25455 30277 25467 30280
rect 25409 30271 25467 30277
rect 28810 30268 28816 30280
rect 28868 30268 28874 30320
rect 23845 30243 23903 30249
rect 23845 30209 23857 30243
rect 23891 30209 23903 30243
rect 23845 30203 23903 30209
rect 16393 30175 16451 30181
rect 16393 30172 16405 30175
rect 15344 30144 16405 30172
rect 15344 30132 15350 30144
rect 16393 30141 16405 30144
rect 16439 30141 16451 30175
rect 16393 30135 16451 30141
rect 16577 30175 16635 30181
rect 16577 30141 16589 30175
rect 16623 30141 16635 30175
rect 16577 30135 16635 30141
rect 16945 30175 17003 30181
rect 16945 30141 16957 30175
rect 16991 30141 17003 30175
rect 16945 30135 17003 30141
rect 19334 30132 19340 30184
rect 19392 30172 19398 30184
rect 19613 30175 19671 30181
rect 19613 30172 19625 30175
rect 19392 30144 19625 30172
rect 19392 30132 19398 30144
rect 19613 30141 19625 30144
rect 19659 30141 19671 30175
rect 21542 30172 21548 30184
rect 21503 30144 21548 30172
rect 19613 30135 19671 30141
rect 21542 30132 21548 30144
rect 21600 30172 21606 30184
rect 22097 30175 22155 30181
rect 22097 30172 22109 30175
rect 21600 30144 22109 30172
rect 21600 30132 21606 30144
rect 22097 30141 22109 30144
rect 22143 30141 22155 30175
rect 22097 30135 22155 30141
rect 22281 30175 22339 30181
rect 22281 30141 22293 30175
rect 22327 30172 22339 30175
rect 22738 30172 22744 30184
rect 22327 30144 22744 30172
rect 22327 30141 22339 30144
rect 22281 30135 22339 30141
rect 22738 30132 22744 30144
rect 22796 30132 22802 30184
rect 24029 30175 24087 30181
rect 24029 30141 24041 30175
rect 24075 30141 24087 30175
rect 24486 30172 24492 30184
rect 24447 30144 24492 30172
rect 24029 30135 24087 30141
rect 17218 30104 17224 30116
rect 15212 30076 15424 30104
rect 17179 30076 17224 30104
rect 15396 30048 15424 30076
rect 17218 30064 17224 30076
rect 17276 30064 17282 30116
rect 17681 30107 17739 30113
rect 17681 30104 17693 30107
rect 17328 30076 17693 30104
rect 3375 30008 4016 30036
rect 3375 30005 3387 30008
rect 3329 29999 3387 30005
rect 4522 29996 4528 30048
rect 4580 30036 4586 30048
rect 4893 30039 4951 30045
rect 4893 30036 4905 30039
rect 4580 30008 4905 30036
rect 4580 29996 4586 30008
rect 4893 30005 4905 30008
rect 4939 30036 4951 30039
rect 5534 30036 5540 30048
rect 4939 30008 5540 30036
rect 4939 30005 4951 30008
rect 4893 29999 4951 30005
rect 5534 29996 5540 30008
rect 5592 29996 5598 30048
rect 9766 30036 9772 30048
rect 9727 30008 9772 30036
rect 9766 29996 9772 30008
rect 9824 29996 9830 30048
rect 12529 30039 12587 30045
rect 12529 30005 12541 30039
rect 12575 30036 12587 30039
rect 12986 30036 12992 30048
rect 12575 30008 12992 30036
rect 12575 30005 12587 30008
rect 12529 29999 12587 30005
rect 12986 29996 12992 30008
rect 13044 29996 13050 30048
rect 15010 30036 15016 30048
rect 14971 30008 15016 30036
rect 15010 29996 15016 30008
rect 15068 29996 15074 30048
rect 15378 30036 15384 30048
rect 15339 30008 15384 30036
rect 15378 29996 15384 30008
rect 15436 29996 15442 30048
rect 16666 29996 16672 30048
rect 16724 30036 16730 30048
rect 17328 30036 17356 30076
rect 17681 30073 17693 30076
rect 17727 30104 17739 30107
rect 17773 30107 17831 30113
rect 17773 30104 17785 30107
rect 17727 30076 17785 30104
rect 17727 30073 17739 30076
rect 17681 30067 17739 30073
rect 17773 30073 17785 30076
rect 17819 30073 17831 30107
rect 18046 30104 18052 30116
rect 18007 30076 18052 30104
rect 17773 30067 17831 30073
rect 18046 30064 18052 30076
rect 18104 30064 18110 30116
rect 18322 30064 18328 30116
rect 18380 30104 18386 30116
rect 24044 30104 24072 30135
rect 24486 30132 24492 30144
rect 24544 30132 24550 30184
rect 24578 30132 24584 30184
rect 24636 30172 24642 30184
rect 24636 30144 24681 30172
rect 24636 30132 24642 30144
rect 58434 30132 58440 30184
rect 58492 30172 58498 30184
rect 58894 30172 58900 30184
rect 58492 30144 58900 30172
rect 58492 30132 58498 30144
rect 58894 30132 58900 30144
rect 58952 30132 58958 30184
rect 24596 30104 24624 30132
rect 27062 30104 27068 30116
rect 18380 30076 23980 30104
rect 24044 30076 24624 30104
rect 24688 30076 27068 30104
rect 18380 30064 18386 30076
rect 17494 30036 17500 30048
rect 16724 30008 17356 30036
rect 17455 30008 17500 30036
rect 16724 29996 16730 30008
rect 17494 29996 17500 30008
rect 17552 29996 17558 30048
rect 18690 30036 18696 30048
rect 18651 30008 18696 30036
rect 18690 29996 18696 30008
rect 18748 29996 18754 30048
rect 22738 29996 22744 30048
rect 22796 30036 22802 30048
rect 22833 30039 22891 30045
rect 22833 30036 22845 30039
rect 22796 30008 22845 30036
rect 22796 29996 22802 30008
rect 22833 30005 22845 30008
rect 22879 30005 22891 30039
rect 23952 30036 23980 30076
rect 24688 30036 24716 30076
rect 27062 30064 27068 30076
rect 27120 30064 27126 30116
rect 25038 30036 25044 30048
rect 23952 30008 24716 30036
rect 24999 30008 25044 30036
rect 22833 29999 22891 30005
rect 25038 29996 25044 30008
rect 25096 29996 25102 30048
rect 1104 29946 29256 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 29256 29946
rect 1104 29872 29256 29894
rect 3326 29832 3332 29844
rect 3287 29804 3332 29832
rect 3326 29792 3332 29804
rect 3384 29792 3390 29844
rect 4982 29832 4988 29844
rect 4943 29804 4988 29832
rect 4982 29792 4988 29804
rect 5040 29792 5046 29844
rect 12066 29832 12072 29844
rect 12027 29804 12072 29832
rect 12066 29792 12072 29804
rect 12124 29792 12130 29844
rect 14090 29832 14096 29844
rect 14051 29804 14096 29832
rect 14090 29792 14096 29804
rect 14148 29792 14154 29844
rect 17494 29792 17500 29844
rect 17552 29832 17558 29844
rect 20165 29835 20223 29841
rect 20165 29832 20177 29835
rect 17552 29804 19840 29832
rect 17552 29792 17558 29804
rect 2682 29696 2688 29708
rect 2643 29668 2688 29696
rect 2682 29656 2688 29668
rect 2740 29656 2746 29708
rect 2869 29699 2927 29705
rect 2869 29665 2881 29699
rect 2915 29696 2927 29699
rect 3344 29696 3372 29792
rect 2915 29668 3372 29696
rect 2915 29665 2927 29668
rect 2869 29659 2927 29665
rect 3694 29656 3700 29708
rect 3752 29696 3758 29708
rect 3878 29696 3884 29708
rect 3752 29668 3884 29696
rect 3752 29656 3758 29668
rect 3878 29656 3884 29668
rect 3936 29656 3942 29708
rect 4157 29699 4215 29705
rect 4157 29696 4169 29699
rect 4080 29668 4169 29696
rect 4080 29640 4108 29668
rect 4157 29665 4169 29668
rect 4203 29665 4215 29699
rect 4157 29659 4215 29665
rect 4617 29699 4675 29705
rect 4617 29665 4629 29699
rect 4663 29696 4675 29699
rect 5000 29696 5028 29792
rect 16574 29724 16580 29776
rect 16632 29764 16638 29776
rect 16632 29736 16804 29764
rect 16632 29724 16638 29736
rect 6086 29696 6092 29708
rect 4663 29668 5028 29696
rect 6047 29668 6092 29696
rect 4663 29665 4675 29668
rect 4617 29659 4675 29665
rect 6086 29656 6092 29668
rect 6144 29656 6150 29708
rect 10781 29699 10839 29705
rect 10781 29665 10793 29699
rect 10827 29696 10839 29699
rect 11146 29696 11152 29708
rect 10827 29668 11152 29696
rect 10827 29665 10839 29668
rect 10781 29659 10839 29665
rect 11146 29656 11152 29668
rect 11204 29656 11210 29708
rect 13906 29696 13912 29708
rect 13867 29668 13912 29696
rect 13906 29656 13912 29668
rect 13964 29656 13970 29708
rect 16776 29705 16804 29736
rect 18046 29724 18052 29776
rect 18104 29764 18110 29776
rect 18785 29767 18843 29773
rect 18785 29764 18797 29767
rect 18104 29736 18797 29764
rect 18104 29724 18110 29736
rect 18785 29733 18797 29736
rect 18831 29733 18843 29767
rect 18785 29727 18843 29733
rect 18874 29724 18880 29776
rect 18932 29764 18938 29776
rect 19702 29764 19708 29776
rect 18932 29736 19708 29764
rect 18932 29724 18938 29736
rect 16761 29699 16819 29705
rect 16761 29665 16773 29699
rect 16807 29696 16819 29699
rect 17310 29696 17316 29708
rect 16807 29668 17316 29696
rect 16807 29665 16819 29668
rect 16761 29659 16819 29665
rect 17310 29656 17316 29668
rect 17368 29656 17374 29708
rect 17497 29699 17555 29705
rect 17497 29665 17509 29699
rect 17543 29696 17555 29699
rect 18138 29696 18144 29708
rect 17543 29668 18144 29696
rect 17543 29665 17555 29668
rect 17497 29659 17555 29665
rect 18138 29656 18144 29668
rect 18196 29696 18202 29708
rect 19444 29705 19472 29736
rect 19702 29724 19708 29736
rect 19760 29724 19766 29776
rect 19812 29705 19840 29804
rect 19904 29804 20177 29832
rect 19904 29776 19932 29804
rect 20165 29801 20177 29804
rect 20211 29832 20223 29835
rect 24854 29832 24860 29844
rect 20211 29804 24860 29832
rect 20211 29801 20223 29804
rect 20165 29795 20223 29801
rect 24854 29792 24860 29804
rect 24912 29792 24918 29844
rect 58434 29792 58440 29844
rect 58492 29832 58498 29844
rect 59078 29832 59084 29844
rect 58492 29804 59084 29832
rect 58492 29792 58498 29804
rect 59078 29792 59084 29804
rect 59136 29792 59142 29844
rect 19886 29724 19892 29776
rect 19944 29724 19950 29776
rect 19245 29699 19303 29705
rect 19245 29696 19257 29699
rect 18196 29668 19257 29696
rect 18196 29656 18202 29668
rect 19245 29665 19257 29668
rect 19291 29665 19303 29699
rect 19245 29659 19303 29665
rect 19429 29699 19487 29705
rect 19429 29665 19441 29699
rect 19475 29665 19487 29699
rect 19429 29659 19487 29665
rect 19797 29699 19855 29705
rect 19797 29665 19809 29699
rect 19843 29696 19855 29699
rect 20349 29699 20407 29705
rect 20349 29696 20361 29699
rect 19843 29668 20361 29696
rect 19843 29665 19855 29668
rect 19797 29659 19855 29665
rect 20349 29665 20361 29668
rect 20395 29696 20407 29699
rect 23569 29699 23627 29705
rect 20395 29668 23428 29696
rect 20395 29665 20407 29668
rect 20349 29659 20407 29665
rect 2958 29628 2964 29640
rect 2919 29600 2964 29628
rect 2958 29588 2964 29600
rect 3016 29588 3022 29640
rect 4062 29588 4068 29640
rect 4120 29588 4126 29640
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29597 4583 29631
rect 4525 29591 4583 29597
rect 3050 29520 3056 29572
rect 3108 29560 3114 29572
rect 4540 29560 4568 29591
rect 4798 29588 4804 29640
rect 4856 29628 4862 29640
rect 5813 29631 5871 29637
rect 5813 29628 5825 29631
rect 4856 29600 5825 29628
rect 4856 29588 4862 29600
rect 5813 29597 5825 29600
rect 5859 29628 5871 29631
rect 7561 29631 7619 29637
rect 7561 29628 7573 29631
rect 5859 29600 7573 29628
rect 5859 29597 5871 29600
rect 5813 29591 5871 29597
rect 7561 29597 7573 29600
rect 7607 29628 7619 29631
rect 7926 29628 7932 29640
rect 7607 29600 7932 29628
rect 7607 29597 7619 29600
rect 7561 29591 7619 29597
rect 7926 29588 7932 29600
rect 7984 29628 7990 29640
rect 10321 29631 10379 29637
rect 10321 29628 10333 29631
rect 7984 29600 10333 29628
rect 7984 29588 7990 29600
rect 10321 29597 10333 29600
rect 10367 29628 10379 29631
rect 10505 29631 10563 29637
rect 10505 29628 10517 29631
rect 10367 29600 10517 29628
rect 10367 29597 10379 29600
rect 10321 29591 10379 29597
rect 10505 29597 10517 29600
rect 10551 29597 10563 29631
rect 10505 29591 10563 29597
rect 16577 29631 16635 29637
rect 16577 29597 16589 29631
rect 16623 29597 16635 29631
rect 19705 29631 19763 29637
rect 19705 29628 19717 29631
rect 16577 29591 16635 29597
rect 18616 29600 19717 29628
rect 3108 29532 4568 29560
rect 3108 29520 3114 29532
rect 16592 29504 16620 29591
rect 17494 29520 17500 29572
rect 17552 29560 17558 29572
rect 17681 29563 17739 29569
rect 17681 29560 17693 29563
rect 17552 29532 17693 29560
rect 17552 29520 17558 29532
rect 17681 29529 17693 29532
rect 17727 29529 17739 29563
rect 17681 29523 17739 29529
rect 4982 29452 4988 29504
rect 5040 29492 5046 29504
rect 7193 29495 7251 29501
rect 7193 29492 7205 29495
rect 5040 29464 7205 29492
rect 5040 29452 5046 29464
rect 7193 29461 7205 29464
rect 7239 29461 7251 29495
rect 7193 29455 7251 29461
rect 16485 29495 16543 29501
rect 16485 29461 16497 29495
rect 16531 29492 16543 29495
rect 16574 29492 16580 29504
rect 16531 29464 16580 29492
rect 16531 29461 16543 29464
rect 16485 29455 16543 29461
rect 16574 29452 16580 29464
rect 16632 29452 16638 29504
rect 17310 29452 17316 29504
rect 17368 29492 17374 29504
rect 18049 29495 18107 29501
rect 18049 29492 18061 29495
rect 17368 29464 18061 29492
rect 17368 29452 17374 29464
rect 18049 29461 18061 29464
rect 18095 29492 18107 29495
rect 18233 29495 18291 29501
rect 18233 29492 18245 29495
rect 18095 29464 18245 29492
rect 18095 29461 18107 29464
rect 18049 29455 18107 29461
rect 18233 29461 18245 29464
rect 18279 29461 18291 29495
rect 18233 29455 18291 29461
rect 18414 29452 18420 29504
rect 18472 29492 18478 29504
rect 18616 29501 18644 29600
rect 19705 29597 19717 29600
rect 19751 29597 19763 29631
rect 23293 29631 23351 29637
rect 23293 29628 23305 29631
rect 19705 29591 19763 29597
rect 23124 29600 23305 29628
rect 18601 29495 18659 29501
rect 18601 29492 18613 29495
rect 18472 29464 18613 29492
rect 18472 29452 18478 29464
rect 18601 29461 18613 29464
rect 18647 29461 18659 29495
rect 18601 29455 18659 29461
rect 20622 29452 20628 29504
rect 20680 29492 20686 29504
rect 23124 29501 23152 29600
rect 23293 29597 23305 29600
rect 23339 29597 23351 29631
rect 23400 29628 23428 29668
rect 23569 29665 23581 29699
rect 23615 29696 23627 29699
rect 25038 29696 25044 29708
rect 23615 29668 25044 29696
rect 23615 29665 23627 29668
rect 23569 29659 23627 29665
rect 25038 29656 25044 29668
rect 25096 29656 25102 29708
rect 25866 29628 25872 29640
rect 23400 29600 25872 29628
rect 23293 29591 23351 29597
rect 25866 29588 25872 29600
rect 25924 29588 25930 29640
rect 86218 29520 86224 29572
rect 86276 29560 86282 29572
rect 87230 29560 87236 29572
rect 86276 29532 87236 29560
rect 86276 29520 86282 29532
rect 87230 29520 87236 29532
rect 87288 29520 87294 29572
rect 23109 29495 23167 29501
rect 23109 29492 23121 29495
rect 20680 29464 23121 29492
rect 20680 29452 20686 29464
rect 23109 29461 23121 29464
rect 23155 29461 23167 29495
rect 24670 29492 24676 29504
rect 24631 29464 24676 29492
rect 23109 29455 23167 29461
rect 24670 29452 24676 29464
rect 24728 29452 24734 29504
rect 1104 29402 29256 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 29256 29402
rect 1104 29328 29256 29350
rect 3970 29248 3976 29300
rect 4028 29288 4034 29300
rect 11514 29288 11520 29300
rect 4028 29260 11520 29288
rect 4028 29248 4034 29260
rect 11514 29248 11520 29260
rect 11572 29248 11578 29300
rect 18138 29288 18144 29300
rect 18099 29260 18144 29288
rect 18138 29248 18144 29260
rect 18196 29248 18202 29300
rect 19613 29291 19671 29297
rect 19613 29257 19625 29291
rect 19659 29288 19671 29291
rect 20254 29288 20260 29300
rect 19659 29260 20260 29288
rect 19659 29257 19671 29260
rect 19613 29251 19671 29257
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 24213 29291 24271 29297
rect 24213 29257 24225 29291
rect 24259 29288 24271 29291
rect 24486 29288 24492 29300
rect 24259 29260 24492 29288
rect 24259 29257 24271 29260
rect 24213 29251 24271 29257
rect 24486 29248 24492 29260
rect 24544 29248 24550 29300
rect 26694 29288 26700 29300
rect 25148 29260 26096 29288
rect 26607 29260 26700 29288
rect 5258 29180 5264 29232
rect 5316 29220 5322 29232
rect 5537 29223 5595 29229
rect 5537 29220 5549 29223
rect 5316 29192 5549 29220
rect 5316 29180 5322 29192
rect 5537 29189 5549 29192
rect 5583 29189 5595 29223
rect 5537 29183 5595 29189
rect 18690 29180 18696 29232
rect 18748 29220 18754 29232
rect 25148 29220 25176 29260
rect 18748 29192 25176 29220
rect 26068 29220 26096 29260
rect 26694 29248 26700 29260
rect 26752 29288 26758 29300
rect 28994 29288 29000 29300
rect 26752 29260 29000 29288
rect 26752 29248 26758 29260
rect 28994 29248 29000 29260
rect 29052 29248 29058 29300
rect 31478 29220 31484 29232
rect 26068 29192 31484 29220
rect 18748 29180 18754 29192
rect 31478 29180 31484 29192
rect 31536 29180 31542 29232
rect 8570 29152 8576 29164
rect 4356 29124 8576 29152
rect 4065 29087 4123 29093
rect 4065 29053 4077 29087
rect 4111 29084 4123 29087
rect 4154 29084 4160 29096
rect 4111 29056 4160 29084
rect 4111 29053 4123 29056
rect 4065 29047 4123 29053
rect 4154 29044 4160 29056
rect 4212 29044 4218 29096
rect 4356 29093 4384 29124
rect 8570 29112 8576 29124
rect 8628 29112 8634 29164
rect 12437 29155 12495 29161
rect 12437 29121 12449 29155
rect 12483 29152 12495 29155
rect 13354 29152 13360 29164
rect 12483 29124 13360 29152
rect 12483 29121 12495 29124
rect 12437 29115 12495 29121
rect 13354 29112 13360 29124
rect 13412 29152 13418 29164
rect 14093 29155 14151 29161
rect 13412 29124 13676 29152
rect 13412 29112 13418 29124
rect 4341 29087 4399 29093
rect 4341 29053 4353 29087
rect 4387 29053 4399 29087
rect 4341 29047 4399 29053
rect 5166 29044 5172 29096
rect 5224 29084 5230 29096
rect 5353 29087 5411 29093
rect 5353 29084 5365 29087
rect 5224 29056 5365 29084
rect 5224 29044 5230 29056
rect 5353 29053 5365 29056
rect 5399 29053 5411 29087
rect 5353 29047 5411 29053
rect 12713 29087 12771 29093
rect 12713 29053 12725 29087
rect 12759 29084 12771 29087
rect 13538 29084 13544 29096
rect 12759 29056 13544 29084
rect 12759 29053 12771 29056
rect 12713 29047 12771 29053
rect 13538 29044 13544 29056
rect 13596 29044 13602 29096
rect 13648 29016 13676 29124
rect 14093 29121 14105 29155
rect 14139 29152 14151 29155
rect 16758 29152 16764 29164
rect 14139 29124 16764 29152
rect 14139 29121 14151 29124
rect 14093 29115 14151 29121
rect 14936 29093 14964 29124
rect 16758 29112 16764 29124
rect 16816 29112 16822 29164
rect 25133 29155 25191 29161
rect 25133 29121 25145 29155
rect 25179 29152 25191 29155
rect 26970 29152 26976 29164
rect 25179 29124 26976 29152
rect 25179 29121 25191 29124
rect 25133 29115 25191 29121
rect 26970 29112 26976 29124
rect 27028 29112 27034 29164
rect 14921 29087 14979 29093
rect 14921 29053 14933 29087
rect 14967 29053 14979 29087
rect 14921 29047 14979 29053
rect 15010 29044 15016 29096
rect 15068 29084 15074 29096
rect 16853 29087 16911 29093
rect 16853 29084 16865 29087
rect 15068 29056 16865 29084
rect 15068 29044 15074 29056
rect 16853 29053 16865 29056
rect 16899 29053 16911 29087
rect 16853 29047 16911 29053
rect 18049 29087 18107 29093
rect 18049 29053 18061 29087
rect 18095 29084 18107 29087
rect 18095 29056 18460 29084
rect 18095 29053 18107 29056
rect 18049 29047 18107 29053
rect 14182 29016 14188 29028
rect 13648 28988 14188 29016
rect 14182 28976 14188 28988
rect 14240 28976 14246 29028
rect 18432 28960 18460 29056
rect 19334 29044 19340 29096
rect 19392 29084 19398 29096
rect 19429 29087 19487 29093
rect 19429 29084 19441 29087
rect 19392 29056 19441 29084
rect 19392 29044 19398 29056
rect 19429 29053 19441 29056
rect 19475 29053 19487 29087
rect 19429 29047 19487 29053
rect 24121 29087 24179 29093
rect 24121 29053 24133 29087
rect 24167 29053 24179 29087
rect 25406 29084 25412 29096
rect 25367 29056 25412 29084
rect 24121 29047 24179 29053
rect 24136 29016 24164 29047
rect 25406 29044 25412 29056
rect 25464 29044 25470 29096
rect 24489 29019 24547 29025
rect 24489 29016 24501 29019
rect 24136 28988 24501 29016
rect 24489 28985 24501 28988
rect 24535 29016 24547 29019
rect 24670 29016 24676 29028
rect 24535 28988 24676 29016
rect 24535 28985 24547 28988
rect 24489 28979 24547 28985
rect 24670 28976 24676 28988
rect 24728 28976 24734 29028
rect 3878 28948 3884 28960
rect 3839 28920 3884 28948
rect 3878 28908 3884 28920
rect 3936 28908 3942 28960
rect 5166 28908 5172 28960
rect 5224 28948 5230 28960
rect 9030 28948 9036 28960
rect 5224 28920 9036 28948
rect 5224 28908 5230 28920
rect 9030 28908 9036 28920
rect 9088 28908 9094 28960
rect 15010 28948 15016 28960
rect 14971 28920 15016 28948
rect 15010 28908 15016 28920
rect 15068 28908 15074 28960
rect 16669 28951 16727 28957
rect 16669 28917 16681 28951
rect 16715 28948 16727 28951
rect 17126 28948 17132 28960
rect 16715 28920 17132 28948
rect 16715 28917 16727 28920
rect 16669 28911 16727 28917
rect 17126 28908 17132 28920
rect 17184 28908 17190 28960
rect 18414 28948 18420 28960
rect 18375 28920 18420 28948
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 26970 28948 26976 28960
rect 26931 28920 26976 28948
rect 26970 28908 26976 28920
rect 27028 28908 27034 28960
rect 1104 28858 29256 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 29256 28858
rect 1104 28784 29256 28806
rect 4062 28704 4068 28756
rect 4120 28744 4126 28756
rect 4982 28744 4988 28756
rect 4120 28716 4988 28744
rect 4120 28704 4126 28716
rect 4982 28704 4988 28716
rect 5040 28704 5046 28756
rect 13906 28744 13912 28756
rect 12268 28716 13912 28744
rect 4154 28636 4160 28688
rect 4212 28676 4218 28688
rect 5258 28676 5264 28688
rect 4212 28648 5264 28676
rect 4212 28636 4218 28648
rect 4356 28617 4384 28648
rect 5258 28636 5264 28648
rect 5316 28636 5322 28688
rect 4341 28611 4399 28617
rect 4341 28577 4353 28611
rect 4387 28577 4399 28611
rect 4341 28571 4399 28577
rect 4525 28611 4583 28617
rect 4525 28577 4537 28611
rect 4571 28608 4583 28611
rect 4985 28611 5043 28617
rect 4985 28608 4997 28611
rect 4571 28580 4997 28608
rect 4571 28577 4583 28580
rect 4525 28571 4583 28577
rect 4985 28577 4997 28580
rect 5031 28608 5043 28611
rect 5442 28608 5448 28620
rect 5031 28580 5448 28608
rect 5031 28577 5043 28580
rect 4985 28571 5043 28577
rect 5442 28568 5448 28580
rect 5500 28568 5506 28620
rect 12268 28617 12296 28716
rect 13906 28704 13912 28716
rect 13964 28704 13970 28756
rect 19613 28747 19671 28753
rect 19613 28713 19625 28747
rect 19659 28744 19671 28747
rect 20254 28744 20260 28756
rect 19659 28716 20260 28744
rect 19659 28713 19671 28716
rect 19613 28707 19671 28713
rect 13081 28679 13139 28685
rect 13081 28676 13093 28679
rect 12452 28648 13093 28676
rect 12452 28617 12480 28648
rect 13081 28645 13093 28648
rect 13127 28676 13139 28679
rect 13170 28676 13176 28688
rect 13127 28648 13176 28676
rect 13127 28645 13139 28648
rect 13081 28639 13139 28645
rect 13170 28636 13176 28648
rect 13228 28676 13234 28688
rect 13228 28648 17356 28676
rect 13228 28636 13234 28648
rect 8389 28611 8447 28617
rect 8389 28608 8401 28611
rect 8312 28580 8401 28608
rect 4614 28540 4620 28552
rect 4575 28512 4620 28540
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 5902 28364 5908 28416
rect 5960 28404 5966 28416
rect 6822 28404 6828 28416
rect 5960 28376 6828 28404
rect 5960 28364 5966 28376
rect 6822 28364 6828 28376
rect 6880 28404 6886 28416
rect 8312 28413 8340 28580
rect 8389 28577 8401 28580
rect 8435 28577 8447 28611
rect 8389 28571 8447 28577
rect 11701 28611 11759 28617
rect 11701 28577 11713 28611
rect 11747 28608 11759 28611
rect 12253 28611 12311 28617
rect 12253 28608 12265 28611
rect 11747 28580 12265 28608
rect 11747 28577 11759 28580
rect 11701 28571 11759 28577
rect 12253 28577 12265 28580
rect 12299 28577 12311 28611
rect 12253 28571 12311 28577
rect 12437 28611 12495 28617
rect 12437 28577 12449 28611
rect 12483 28577 12495 28611
rect 13722 28608 13728 28620
rect 13683 28580 13728 28608
rect 12437 28571 12495 28577
rect 13722 28568 13728 28580
rect 13780 28568 13786 28620
rect 11425 28543 11483 28549
rect 11425 28509 11437 28543
rect 11471 28540 11483 28543
rect 11609 28543 11667 28549
rect 11609 28540 11621 28543
rect 11471 28512 11621 28540
rect 11471 28509 11483 28512
rect 11425 28503 11483 28509
rect 11609 28509 11621 28512
rect 11655 28540 11667 28543
rect 11655 28512 11744 28540
rect 11655 28509 11667 28512
rect 11609 28503 11667 28509
rect 11716 28484 11744 28512
rect 12986 28500 12992 28552
rect 13044 28540 13050 28552
rect 16574 28540 16580 28552
rect 13044 28512 16580 28540
rect 13044 28500 13050 28512
rect 16574 28500 16580 28512
rect 16632 28500 16638 28552
rect 17221 28543 17279 28549
rect 17221 28540 17233 28543
rect 17144 28512 17233 28540
rect 11698 28432 11704 28484
rect 11756 28432 11762 28484
rect 12618 28472 12624 28484
rect 12579 28444 12624 28472
rect 12618 28432 12624 28444
rect 12676 28432 12682 28484
rect 13906 28472 13912 28484
rect 13867 28444 13912 28472
rect 13906 28432 13912 28444
rect 13964 28432 13970 28484
rect 17144 28416 17172 28512
rect 17221 28509 17233 28512
rect 17267 28509 17279 28543
rect 17328 28540 17356 28648
rect 17494 28608 17500 28620
rect 17455 28580 17500 28608
rect 17494 28568 17500 28580
rect 17552 28568 17558 28620
rect 19720 28617 19748 28716
rect 20254 28704 20260 28716
rect 20312 28704 20318 28756
rect 19705 28611 19763 28617
rect 19705 28577 19717 28611
rect 19751 28577 19763 28611
rect 19705 28571 19763 28577
rect 25409 28611 25467 28617
rect 25409 28577 25421 28611
rect 25455 28608 25467 28611
rect 26694 28608 26700 28620
rect 25455 28580 26700 28608
rect 25455 28577 25467 28580
rect 25409 28571 25467 28577
rect 26694 28568 26700 28580
rect 26752 28568 26758 28620
rect 27341 28611 27399 28617
rect 27341 28577 27353 28611
rect 27387 28608 27399 28611
rect 28074 28608 28080 28620
rect 27387 28580 28080 28608
rect 27387 28577 27399 28580
rect 27341 28571 27399 28577
rect 28074 28568 28080 28580
rect 28132 28568 28138 28620
rect 28626 28540 28632 28552
rect 17328 28512 28632 28540
rect 17221 28503 17279 28509
rect 28626 28500 28632 28512
rect 28684 28500 28690 28552
rect 8297 28407 8355 28413
rect 8297 28404 8309 28407
rect 6880 28376 8309 28404
rect 6880 28364 6886 28376
rect 8297 28373 8309 28376
rect 8343 28373 8355 28407
rect 8478 28404 8484 28416
rect 8439 28376 8484 28404
rect 8297 28367 8355 28373
rect 8478 28364 8484 28376
rect 8536 28364 8542 28416
rect 17126 28404 17132 28416
rect 17087 28376 17132 28404
rect 17126 28364 17132 28376
rect 17184 28364 17190 28416
rect 18414 28364 18420 28416
rect 18472 28404 18478 28416
rect 18601 28407 18659 28413
rect 18601 28404 18613 28407
rect 18472 28376 18613 28404
rect 18472 28364 18478 28376
rect 18601 28373 18613 28376
rect 18647 28373 18659 28407
rect 19886 28404 19892 28416
rect 19847 28376 19892 28404
rect 18601 28367 18659 28373
rect 19886 28364 19892 28376
rect 19944 28364 19950 28416
rect 25222 28364 25228 28416
rect 25280 28404 25286 28416
rect 25501 28407 25559 28413
rect 25501 28404 25513 28407
rect 25280 28376 25513 28404
rect 25280 28364 25286 28376
rect 25501 28373 25513 28376
rect 25547 28373 25559 28407
rect 27430 28404 27436 28416
rect 27391 28376 27436 28404
rect 25501 28367 25559 28373
rect 27430 28364 27436 28376
rect 27488 28364 27494 28416
rect 1104 28314 29256 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 29256 28314
rect 1104 28240 29256 28262
rect 8478 28160 8484 28212
rect 8536 28200 8542 28212
rect 18322 28200 18328 28212
rect 8536 28172 18328 28200
rect 8536 28160 8542 28172
rect 2869 28067 2927 28073
rect 2869 28033 2881 28067
rect 2915 28064 2927 28067
rect 3602 28064 3608 28076
rect 2915 28036 3608 28064
rect 2915 28033 2927 28036
rect 2869 28027 2927 28033
rect 3602 28024 3608 28036
rect 3660 28024 3666 28076
rect 9324 28073 9352 28172
rect 18322 28160 18328 28172
rect 18380 28160 18386 28212
rect 20714 28160 20720 28212
rect 20772 28200 20778 28212
rect 20990 28200 20996 28212
rect 20772 28172 20996 28200
rect 20772 28160 20778 28172
rect 20990 28160 20996 28172
rect 21048 28160 21054 28212
rect 28074 28200 28080 28212
rect 27987 28172 28080 28200
rect 28074 28160 28080 28172
rect 28132 28200 28138 28212
rect 28902 28200 28908 28212
rect 28132 28172 28908 28200
rect 28132 28160 28138 28172
rect 28902 28160 28908 28172
rect 28960 28160 28966 28212
rect 86218 28160 86224 28212
rect 86276 28200 86282 28212
rect 87046 28200 87052 28212
rect 86276 28172 87052 28200
rect 86276 28160 86282 28172
rect 87046 28160 87052 28172
rect 87104 28160 87110 28212
rect 9858 28132 9864 28144
rect 9819 28104 9864 28132
rect 9858 28092 9864 28104
rect 9916 28092 9922 28144
rect 11330 28132 11336 28144
rect 11291 28104 11336 28132
rect 11330 28092 11336 28104
rect 11388 28092 11394 28144
rect 16666 28132 16672 28144
rect 11440 28104 16672 28132
rect 9309 28067 9367 28073
rect 5644 28036 9260 28064
rect 2590 27996 2596 28008
rect 2551 27968 2596 27996
rect 2590 27956 2596 27968
rect 2648 27956 2654 28008
rect 5258 27996 5264 28008
rect 5219 27968 5264 27996
rect 5258 27956 5264 27968
rect 5316 27956 5322 28008
rect 5644 28005 5672 28036
rect 5629 27999 5687 28005
rect 5629 27965 5641 27999
rect 5675 27965 5687 27999
rect 5629 27959 5687 27965
rect 7561 27999 7619 28005
rect 7561 27965 7573 27999
rect 7607 27996 7619 27999
rect 8478 27996 8484 28008
rect 7607 27968 8484 27996
rect 7607 27965 7619 27968
rect 7561 27959 7619 27965
rect 8478 27956 8484 27968
rect 8536 27956 8542 28008
rect 3602 27888 3608 27940
rect 3660 27928 3666 27940
rect 8754 27928 8760 27940
rect 3660 27900 5212 27928
rect 8715 27900 8760 27928
rect 3660 27888 3666 27900
rect 4154 27860 4160 27872
rect 4115 27832 4160 27860
rect 4154 27820 4160 27832
rect 4212 27820 4218 27872
rect 4433 27863 4491 27869
rect 4433 27829 4445 27863
rect 4479 27860 4491 27863
rect 4798 27860 4804 27872
rect 4479 27832 4804 27860
rect 4479 27829 4491 27832
rect 4433 27823 4491 27829
rect 4798 27820 4804 27832
rect 4856 27820 4862 27872
rect 5184 27869 5212 27900
rect 8754 27888 8760 27900
rect 8812 27888 8818 27940
rect 9232 27928 9260 28036
rect 9309 28033 9321 28067
rect 9355 28033 9367 28067
rect 9309 28027 9367 28033
rect 9398 27956 9404 28008
rect 9456 28005 9462 28008
rect 9456 27999 9505 28005
rect 9456 27965 9459 27999
rect 9493 27965 9505 27999
rect 9456 27959 9505 27965
rect 9585 27999 9643 28005
rect 9585 27965 9597 27999
rect 9631 27996 9643 27999
rect 9674 27996 9680 28008
rect 9631 27968 9680 27996
rect 9631 27965 9643 27968
rect 9585 27959 9643 27965
rect 9456 27956 9462 27959
rect 9674 27956 9680 27968
rect 9732 27996 9738 28008
rect 9876 27996 9904 28092
rect 9732 27968 9904 27996
rect 10965 27999 11023 28005
rect 9732 27956 9738 27968
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11348 27996 11376 28092
rect 11011 27968 11376 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11238 27928 11244 27940
rect 9232 27900 11244 27928
rect 11238 27888 11244 27900
rect 11296 27888 11302 27940
rect 5169 27863 5227 27869
rect 5169 27829 5181 27863
rect 5215 27829 5227 27863
rect 7650 27860 7656 27872
rect 7611 27832 7656 27860
rect 5169 27823 5227 27829
rect 7650 27820 7656 27832
rect 7708 27820 7714 27872
rect 11146 27860 11152 27872
rect 11059 27832 11152 27860
rect 11146 27820 11152 27832
rect 11204 27860 11210 27872
rect 11440 27860 11468 28104
rect 16666 28092 16672 28104
rect 16724 28092 16730 28144
rect 25406 28132 25412 28144
rect 25367 28104 25412 28132
rect 25406 28092 25412 28104
rect 25464 28092 25470 28144
rect 13630 28064 13636 28076
rect 13591 28036 13636 28064
rect 13630 28024 13636 28036
rect 13688 28024 13694 28076
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 19705 28067 19763 28073
rect 19705 28064 19717 28067
rect 19484 28036 19717 28064
rect 19484 28024 19490 28036
rect 19705 28033 19717 28036
rect 19751 28033 19763 28067
rect 19705 28027 19763 28033
rect 26513 28067 26571 28073
rect 26513 28033 26525 28067
rect 26559 28064 26571 28067
rect 26970 28064 26976 28076
rect 26559 28036 26976 28064
rect 26559 28033 26571 28036
rect 26513 28027 26571 28033
rect 26970 28024 26976 28036
rect 27028 28064 27034 28076
rect 28261 28067 28319 28073
rect 28261 28064 28273 28067
rect 27028 28036 28273 28064
rect 27028 28024 27034 28036
rect 28261 28033 28273 28036
rect 28307 28033 28319 28067
rect 28261 28027 28319 28033
rect 58434 28024 58440 28076
rect 58492 28064 58498 28076
rect 59538 28064 59544 28076
rect 58492 28036 59544 28064
rect 58492 28024 58498 28036
rect 59538 28024 59544 28036
rect 59596 28024 59602 28076
rect 12253 27999 12311 28005
rect 12253 27965 12265 27999
rect 12299 27996 12311 27999
rect 12437 27999 12495 28005
rect 12437 27996 12449 27999
rect 12299 27968 12449 27996
rect 12299 27965 12311 27968
rect 12253 27959 12311 27965
rect 12437 27965 12449 27968
rect 12483 27965 12495 27999
rect 12437 27959 12495 27965
rect 12621 27999 12679 28005
rect 12621 27965 12633 27999
rect 12667 27965 12679 27999
rect 13078 27996 13084 28008
rect 13039 27968 13084 27996
rect 12621 27959 12679 27965
rect 11204 27832 11468 27860
rect 12452 27860 12480 27959
rect 12636 27928 12664 27959
rect 13078 27956 13084 27968
rect 13136 27956 13142 28008
rect 13173 27999 13231 28005
rect 13173 27965 13185 27999
rect 13219 27996 13231 27999
rect 13906 27996 13912 28008
rect 13219 27968 13912 27996
rect 13219 27965 13231 27968
rect 13173 27959 13231 27965
rect 13188 27928 13216 27959
rect 13906 27956 13912 27968
rect 13964 27956 13970 28008
rect 16390 27956 16396 28008
rect 16448 27996 16454 28008
rect 19886 27996 19892 28008
rect 16448 27968 19892 27996
rect 16448 27956 16454 27968
rect 19886 27956 19892 27968
rect 19944 27996 19950 28008
rect 20441 27999 20499 28005
rect 20441 27996 20453 27999
rect 19944 27968 20453 27996
rect 19944 27956 19950 27968
rect 20441 27965 20453 27968
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 20625 27999 20683 28005
rect 20625 27965 20637 27999
rect 20671 27996 20683 27999
rect 23934 27996 23940 28008
rect 20671 27968 23940 27996
rect 20671 27965 20683 27968
rect 20625 27959 20683 27965
rect 23934 27956 23940 27968
rect 23992 27956 23998 28008
rect 24305 27999 24363 28005
rect 24305 27996 24317 27999
rect 24136 27968 24317 27996
rect 12636 27900 13216 27928
rect 16574 27888 16580 27940
rect 16632 27928 16638 27940
rect 20990 27928 20996 27940
rect 16632 27900 19656 27928
rect 20951 27900 20996 27928
rect 16632 27888 16638 27900
rect 12986 27860 12992 27872
rect 12452 27832 12992 27860
rect 11204 27820 11210 27832
rect 12986 27820 12992 27832
rect 13044 27820 13050 27872
rect 13078 27820 13084 27872
rect 13136 27860 13142 27872
rect 15010 27860 15016 27872
rect 13136 27832 15016 27860
rect 13136 27820 13142 27832
rect 15010 27820 15016 27832
rect 15068 27820 15074 27872
rect 19426 27820 19432 27872
rect 19484 27860 19490 27872
rect 19521 27863 19579 27869
rect 19521 27860 19533 27863
rect 19484 27832 19533 27860
rect 19484 27820 19490 27832
rect 19521 27829 19533 27832
rect 19567 27829 19579 27863
rect 19628 27860 19656 27900
rect 20990 27888 20996 27900
rect 21048 27888 21054 27940
rect 24136 27869 24164 27968
rect 24305 27965 24317 27968
rect 24351 27965 24363 27999
rect 24305 27959 24363 27965
rect 24489 27999 24547 28005
rect 24489 27965 24501 27999
rect 24535 27965 24547 27999
rect 24489 27959 24547 27965
rect 25041 27999 25099 28005
rect 25041 27965 25053 27999
rect 25087 27996 25099 27999
rect 25222 27996 25228 28008
rect 25087 27968 25121 27996
rect 25183 27968 25228 27996
rect 25087 27965 25099 27968
rect 25041 27959 25099 27965
rect 24504 27928 24532 27959
rect 25056 27928 25084 27959
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 26789 27999 26847 28005
rect 26789 27965 26801 27999
rect 26835 27996 26847 27999
rect 27798 27996 27804 28008
rect 26835 27968 27804 27996
rect 26835 27965 26847 27968
rect 26789 27959 26847 27965
rect 27798 27956 27804 27968
rect 27856 27956 27862 28008
rect 26602 27928 26608 27940
rect 24504 27900 26608 27928
rect 26602 27888 26608 27900
rect 26660 27888 26666 27940
rect 59538 27928 59544 27940
rect 59499 27900 59544 27928
rect 59538 27888 59544 27900
rect 59596 27888 59602 27940
rect 24121 27863 24179 27869
rect 24121 27860 24133 27863
rect 19628 27832 24133 27860
rect 19521 27823 19579 27829
rect 24121 27829 24133 27832
rect 24167 27829 24179 27863
rect 24121 27823 24179 27829
rect 1104 27770 29256 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 29256 27770
rect 1104 27696 29256 27718
rect 8478 27656 8484 27668
rect 8439 27628 8484 27656
rect 8478 27616 8484 27628
rect 8536 27616 8542 27668
rect 9306 27656 9312 27668
rect 8956 27628 9312 27656
rect 5258 27588 5264 27600
rect 4356 27560 5264 27588
rect 4356 27529 4384 27560
rect 5258 27548 5264 27560
rect 5316 27548 5322 27600
rect 8754 27588 8760 27600
rect 8036 27560 8760 27588
rect 4341 27523 4399 27529
rect 4341 27489 4353 27523
rect 4387 27489 4399 27523
rect 4341 27483 4399 27489
rect 4525 27523 4583 27529
rect 4525 27489 4537 27523
rect 4571 27520 4583 27523
rect 4985 27523 5043 27529
rect 4985 27520 4997 27523
rect 4571 27492 4997 27520
rect 4571 27489 4583 27492
rect 4525 27483 4583 27489
rect 4985 27489 4997 27492
rect 5031 27520 5043 27523
rect 5074 27520 5080 27532
rect 5031 27492 5080 27520
rect 5031 27489 5043 27492
rect 4985 27483 5043 27489
rect 5074 27480 5080 27492
rect 5132 27480 5138 27532
rect 8036 27529 8064 27560
rect 8754 27548 8760 27560
rect 8812 27548 8818 27600
rect 8956 27597 8984 27628
rect 9306 27616 9312 27628
rect 9364 27656 9370 27668
rect 11146 27656 11152 27668
rect 9364 27628 11152 27656
rect 9364 27616 9370 27628
rect 11146 27616 11152 27628
rect 11204 27616 11210 27668
rect 12066 27616 12072 27668
rect 12124 27656 12130 27668
rect 13722 27656 13728 27668
rect 12124 27628 13728 27656
rect 12124 27616 12130 27628
rect 13722 27616 13728 27628
rect 13780 27616 13786 27668
rect 26602 27616 26608 27668
rect 26660 27656 26666 27668
rect 28994 27656 29000 27668
rect 26660 27628 29000 27656
rect 26660 27616 26666 27628
rect 28994 27616 29000 27628
rect 29052 27616 29058 27668
rect 59265 27659 59323 27665
rect 59265 27625 59277 27659
rect 59311 27656 59323 27659
rect 59354 27656 59360 27668
rect 59311 27628 59360 27656
rect 59311 27625 59323 27628
rect 59265 27619 59323 27625
rect 59354 27616 59360 27628
rect 59412 27616 59418 27668
rect 8941 27591 8999 27597
rect 8941 27557 8953 27591
rect 8987 27557 8999 27591
rect 17310 27588 17316 27600
rect 8941 27551 8999 27557
rect 15856 27560 17316 27588
rect 8021 27523 8079 27529
rect 8021 27489 8033 27523
rect 8067 27489 8079 27523
rect 8021 27483 8079 27489
rect 8297 27523 8355 27529
rect 8297 27489 8309 27523
rect 8343 27520 8355 27523
rect 8956 27520 8984 27551
rect 9122 27520 9128 27532
rect 8343 27492 8984 27520
rect 9083 27492 9128 27520
rect 8343 27489 8355 27492
rect 8297 27483 8355 27489
rect 9122 27480 9128 27492
rect 9180 27480 9186 27532
rect 10594 27520 10600 27532
rect 10555 27492 10600 27520
rect 10594 27480 10600 27492
rect 10652 27480 10658 27532
rect 11793 27523 11851 27529
rect 11793 27489 11805 27523
rect 11839 27520 11851 27523
rect 12618 27520 12624 27532
rect 11839 27492 12624 27520
rect 11839 27489 11851 27492
rect 11793 27483 11851 27489
rect 12618 27480 12624 27492
rect 12676 27480 12682 27532
rect 15856 27529 15884 27560
rect 17310 27548 17316 27560
rect 17368 27548 17374 27600
rect 24854 27548 24860 27600
rect 24912 27588 24918 27600
rect 25130 27588 25136 27600
rect 24912 27560 25136 27588
rect 24912 27548 24918 27560
rect 25130 27548 25136 27560
rect 25188 27548 25194 27600
rect 27798 27588 27804 27600
rect 27759 27560 27804 27588
rect 27798 27548 27804 27560
rect 27856 27548 27862 27600
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27489 15899 27523
rect 15841 27483 15899 27489
rect 15930 27480 15936 27532
rect 15988 27520 15994 27532
rect 16390 27520 16396 27532
rect 15988 27492 16033 27520
rect 16351 27492 16396 27520
rect 15988 27480 15994 27492
rect 16390 27480 16396 27492
rect 16448 27480 16454 27532
rect 16577 27523 16635 27529
rect 16577 27489 16589 27523
rect 16623 27520 16635 27523
rect 16623 27492 16988 27520
rect 16623 27489 16635 27492
rect 16577 27483 16635 27489
rect 2866 27412 2872 27464
rect 2924 27452 2930 27464
rect 4617 27455 4675 27461
rect 4617 27452 4629 27455
rect 2924 27424 4629 27452
rect 2924 27412 2930 27424
rect 4617 27421 4629 27424
rect 4663 27421 4675 27455
rect 4617 27415 4675 27421
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27452 8171 27455
rect 9140 27452 9168 27480
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 8159 27424 9168 27452
rect 11348 27424 11529 27452
rect 8159 27421 8171 27424
rect 8113 27415 8171 27421
rect 3510 27344 3516 27396
rect 3568 27384 3574 27396
rect 10962 27384 10968 27396
rect 3568 27356 10968 27384
rect 3568 27344 3574 27356
rect 10962 27344 10968 27356
rect 11020 27344 11026 27396
rect 9582 27276 9588 27328
rect 9640 27316 9646 27328
rect 11348 27325 11376 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 11698 27412 11704 27464
rect 11756 27452 11762 27464
rect 15565 27455 15623 27461
rect 15565 27452 15577 27455
rect 11756 27424 15577 27452
rect 11756 27412 11762 27424
rect 15565 27421 15577 27424
rect 15611 27452 15623 27455
rect 15948 27452 15976 27480
rect 15611 27424 15976 27452
rect 15611 27421 15623 27424
rect 15565 27415 15623 27421
rect 16960 27328 16988 27492
rect 20990 27480 20996 27532
rect 21048 27520 21054 27532
rect 21177 27523 21235 27529
rect 21177 27520 21189 27523
rect 21048 27492 21189 27520
rect 21048 27480 21054 27492
rect 21177 27489 21189 27492
rect 21223 27489 21235 27523
rect 21177 27483 21235 27489
rect 23201 27523 23259 27529
rect 23201 27489 23213 27523
rect 23247 27520 23259 27523
rect 23501 27523 23559 27529
rect 23501 27520 23513 27523
rect 23247 27492 23513 27520
rect 23247 27489 23259 27492
rect 23201 27483 23259 27489
rect 23501 27489 23513 27492
rect 23547 27520 23559 27523
rect 24118 27520 24124 27532
rect 23547 27492 24124 27520
rect 23547 27489 23559 27492
rect 23501 27483 23559 27489
rect 24118 27480 24124 27492
rect 24176 27480 24182 27532
rect 26694 27520 26700 27532
rect 26655 27492 26700 27520
rect 26694 27480 26700 27492
rect 26752 27520 26758 27532
rect 27249 27523 27307 27529
rect 27249 27520 27261 27523
rect 26752 27492 27261 27520
rect 26752 27480 26758 27492
rect 27249 27489 27261 27492
rect 27295 27489 27307 27523
rect 27430 27520 27436 27532
rect 27391 27492 27436 27520
rect 27249 27483 27307 27489
rect 27430 27480 27436 27492
rect 27488 27480 27494 27532
rect 17126 27412 17132 27464
rect 17184 27452 17190 27464
rect 20622 27452 20628 27464
rect 17184 27424 20628 27452
rect 17184 27412 17190 27424
rect 20622 27412 20628 27424
rect 20680 27452 20686 27464
rect 20717 27455 20775 27461
rect 20717 27452 20729 27455
rect 20680 27424 20729 27452
rect 20680 27412 20686 27424
rect 20717 27421 20729 27424
rect 20763 27452 20775 27455
rect 20901 27455 20959 27461
rect 20901 27452 20913 27455
rect 20763 27424 20913 27452
rect 20763 27421 20775 27424
rect 20717 27415 20775 27421
rect 20901 27421 20913 27424
rect 20947 27421 20959 27455
rect 20901 27415 20959 27421
rect 22278 27412 22284 27464
rect 22336 27452 22342 27464
rect 22557 27455 22615 27461
rect 22557 27452 22569 27455
rect 22336 27424 22569 27452
rect 22336 27412 22342 27424
rect 22557 27421 22569 27424
rect 22603 27452 22615 27455
rect 23750 27452 23756 27464
rect 22603 27424 23756 27452
rect 22603 27421 22615 27424
rect 22557 27415 22615 27421
rect 23750 27412 23756 27424
rect 23808 27412 23814 27464
rect 26513 27455 26571 27461
rect 26513 27452 26525 27455
rect 26252 27424 26525 27452
rect 26252 27328 26280 27424
rect 26513 27421 26525 27424
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 10413 27319 10471 27325
rect 10413 27316 10425 27319
rect 9640 27288 10425 27316
rect 9640 27276 9646 27288
rect 10413 27285 10425 27288
rect 10459 27316 10471 27319
rect 11333 27319 11391 27325
rect 11333 27316 11345 27319
rect 10459 27288 11345 27316
rect 10459 27285 10471 27288
rect 10413 27279 10471 27285
rect 11333 27285 11345 27288
rect 11379 27285 11391 27319
rect 13078 27316 13084 27328
rect 13039 27288 13084 27316
rect 11333 27279 11391 27285
rect 13078 27276 13084 27288
rect 13136 27276 13142 27328
rect 16850 27316 16856 27328
rect 16811 27288 16856 27316
rect 16850 27276 16856 27288
rect 16908 27276 16914 27328
rect 16942 27276 16948 27328
rect 17000 27316 17006 27328
rect 17129 27319 17187 27325
rect 17129 27316 17141 27319
rect 17000 27288 17141 27316
rect 17000 27276 17006 27288
rect 17129 27285 17141 27288
rect 17175 27285 17187 27319
rect 17129 27279 17187 27285
rect 17862 27276 17868 27328
rect 17920 27316 17926 27328
rect 23201 27319 23259 27325
rect 23201 27316 23213 27319
rect 17920 27288 23213 27316
rect 17920 27276 17926 27288
rect 23201 27285 23213 27288
rect 23247 27316 23259 27319
rect 23293 27319 23351 27325
rect 23293 27316 23305 27319
rect 23247 27288 23305 27316
rect 23247 27285 23259 27288
rect 23201 27279 23259 27285
rect 23293 27285 23305 27288
rect 23339 27285 23351 27319
rect 23566 27316 23572 27328
rect 23527 27288 23572 27316
rect 23293 27279 23351 27285
rect 23566 27276 23572 27288
rect 23624 27276 23630 27328
rect 26234 27316 26240 27328
rect 26195 27288 26240 27316
rect 26234 27276 26240 27288
rect 26292 27276 26298 27328
rect 1104 27226 29256 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 29256 27226
rect 1104 27152 29256 27174
rect 11241 27115 11299 27121
rect 11241 27081 11253 27115
rect 11287 27112 11299 27115
rect 11330 27112 11336 27124
rect 11287 27084 11336 27112
rect 11287 27081 11299 27084
rect 11241 27075 11299 27081
rect 2590 26976 2596 26988
rect 2551 26948 2596 26976
rect 2590 26936 2596 26948
rect 2648 26936 2654 26988
rect 2866 26976 2872 26988
rect 2827 26948 2872 26976
rect 2866 26936 2872 26948
rect 2924 26936 2930 26988
rect 7745 26979 7803 26985
rect 7745 26945 7757 26979
rect 7791 26976 7803 26979
rect 9398 26976 9404 26988
rect 7791 26948 9404 26976
rect 7791 26945 7803 26948
rect 7745 26939 7803 26945
rect 9398 26936 9404 26948
rect 9456 26976 9462 26988
rect 9677 26979 9735 26985
rect 9677 26976 9689 26979
rect 9456 26948 9689 26976
rect 9456 26936 9462 26948
rect 9677 26945 9689 26948
rect 9723 26976 9735 26979
rect 9723 26948 10548 26976
rect 9723 26945 9735 26948
rect 9677 26939 9735 26945
rect 2608 26908 2636 26936
rect 4246 26908 4252 26920
rect 2608 26880 4252 26908
rect 4246 26868 4252 26880
rect 4304 26908 4310 26920
rect 4341 26911 4399 26917
rect 4341 26908 4353 26911
rect 4304 26880 4353 26908
rect 4304 26868 4310 26880
rect 4341 26877 4353 26880
rect 4387 26908 4399 26911
rect 4798 26908 4804 26920
rect 4387 26880 4804 26908
rect 4387 26877 4399 26880
rect 4341 26871 4399 26877
rect 4798 26868 4804 26880
rect 4856 26868 4862 26920
rect 7653 26911 7711 26917
rect 7653 26908 7665 26911
rect 7576 26880 7665 26908
rect 7576 26784 7604 26880
rect 7653 26877 7665 26880
rect 7699 26877 7711 26911
rect 8570 26908 8576 26920
rect 8483 26880 8576 26908
rect 7653 26871 7711 26877
rect 8570 26868 8576 26880
rect 8628 26908 8634 26920
rect 9214 26908 9220 26920
rect 8628 26880 9220 26908
rect 8628 26868 8634 26880
rect 9214 26868 9220 26880
rect 9272 26868 9278 26920
rect 10520 26917 10548 26948
rect 9493 26911 9551 26917
rect 9493 26877 9505 26911
rect 9539 26877 9551 26911
rect 9493 26871 9551 26877
rect 10505 26911 10563 26917
rect 10505 26877 10517 26911
rect 10551 26877 10563 26911
rect 10505 26871 10563 26877
rect 10689 26911 10747 26917
rect 10689 26877 10701 26911
rect 10735 26908 10747 26911
rect 11256 26908 11284 27075
rect 11330 27072 11336 27084
rect 11388 27072 11394 27124
rect 13170 27112 13176 27124
rect 13131 27084 13176 27112
rect 13170 27072 13176 27084
rect 13228 27072 13234 27124
rect 15930 27072 15936 27124
rect 15988 27112 15994 27124
rect 26234 27112 26240 27124
rect 15988 27084 26240 27112
rect 15988 27072 15994 27084
rect 26234 27072 26240 27084
rect 26292 27072 26298 27124
rect 26602 27112 26608 27124
rect 26563 27084 26608 27112
rect 26602 27072 26608 27084
rect 26660 27072 26666 27124
rect 14182 26976 14188 26988
rect 14095 26948 14188 26976
rect 14182 26936 14188 26948
rect 14240 26976 14246 26988
rect 14277 26979 14335 26985
rect 14277 26976 14289 26979
rect 14240 26948 14289 26976
rect 14240 26936 14246 26948
rect 14277 26945 14289 26948
rect 14323 26945 14335 26979
rect 14277 26939 14335 26945
rect 14553 26979 14611 26985
rect 14553 26945 14565 26979
rect 14599 26976 14611 26979
rect 16850 26976 16856 26988
rect 14599 26948 16856 26976
rect 14599 26945 14611 26948
rect 14553 26939 14611 26945
rect 16850 26936 16856 26948
rect 16908 26936 16914 26988
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26976 20683 26979
rect 20671 26948 21036 26976
rect 20671 26945 20683 26948
rect 20625 26939 20683 26945
rect 13078 26908 13084 26920
rect 10735 26880 11284 26908
rect 13039 26880 13084 26908
rect 10735 26877 10747 26880
rect 10689 26871 10747 26877
rect 8386 26800 8392 26852
rect 8444 26840 8450 26852
rect 8665 26843 8723 26849
rect 8665 26840 8677 26843
rect 8444 26812 8677 26840
rect 8444 26800 8450 26812
rect 8665 26809 8677 26812
rect 8711 26809 8723 26843
rect 9508 26840 9536 26871
rect 13078 26868 13084 26880
rect 13136 26868 13142 26920
rect 16761 26911 16819 26917
rect 16761 26908 16773 26911
rect 15672 26880 16773 26908
rect 9861 26843 9919 26849
rect 9861 26840 9873 26843
rect 9508 26812 9873 26840
rect 8665 26803 8723 26809
rect 9861 26809 9873 26812
rect 9907 26840 9919 26843
rect 12342 26840 12348 26852
rect 9907 26812 12348 26840
rect 9907 26809 9919 26812
rect 9861 26803 9919 26809
rect 12342 26800 12348 26812
rect 12400 26800 12406 26852
rect 15672 26784 15700 26880
rect 16761 26877 16773 26880
rect 16807 26877 16819 26911
rect 16761 26871 16819 26877
rect 20806 26868 20812 26920
rect 20864 26908 20870 26920
rect 21008 26917 21036 26948
rect 22186 26936 22192 26988
rect 22244 26976 22250 26988
rect 31018 26976 31024 26988
rect 22244 26948 31024 26976
rect 22244 26936 22250 26948
rect 31018 26936 31024 26948
rect 31076 26936 31082 26988
rect 87046 26936 87052 26988
rect 87104 26976 87110 26988
rect 87322 26976 87328 26988
rect 87104 26948 87328 26976
rect 87104 26936 87110 26948
rect 87322 26936 87328 26948
rect 87380 26936 87386 26988
rect 20901 26911 20959 26917
rect 20901 26908 20913 26911
rect 20864 26880 20913 26908
rect 20864 26868 20870 26880
rect 20901 26877 20913 26880
rect 20947 26877 20959 26911
rect 20901 26871 20959 26877
rect 20993 26911 21051 26917
rect 20993 26877 21005 26911
rect 21039 26908 21051 26911
rect 21082 26908 21088 26920
rect 21039 26880 21088 26908
rect 21039 26877 21051 26880
rect 20993 26871 21051 26877
rect 20916 26840 20944 26871
rect 21082 26868 21088 26880
rect 21140 26868 21146 26920
rect 21453 26911 21511 26917
rect 21453 26877 21465 26911
rect 21499 26908 21511 26911
rect 21542 26908 21548 26920
rect 21499 26880 21548 26908
rect 21499 26877 21511 26880
rect 21453 26871 21511 26877
rect 21468 26840 21496 26871
rect 21542 26868 21548 26880
rect 21600 26868 21606 26920
rect 21637 26911 21695 26917
rect 21637 26877 21649 26911
rect 21683 26908 21695 26911
rect 25041 26911 25099 26917
rect 21683 26880 22048 26908
rect 21683 26877 21695 26880
rect 21637 26871 21695 26877
rect 20916 26812 21496 26840
rect 4154 26772 4160 26784
rect 4115 26744 4160 26772
rect 4154 26732 4160 26744
rect 4212 26732 4218 26784
rect 7558 26772 7564 26784
rect 7519 26744 7564 26772
rect 7558 26732 7564 26744
rect 7616 26732 7622 26784
rect 10781 26775 10839 26781
rect 10781 26741 10793 26775
rect 10827 26772 10839 26775
rect 11790 26772 11796 26784
rect 10827 26744 11796 26772
rect 10827 26741 10839 26744
rect 10781 26735 10839 26741
rect 11790 26732 11796 26744
rect 11848 26732 11854 26784
rect 15654 26772 15660 26784
rect 15615 26744 15660 26772
rect 15654 26732 15660 26744
rect 15712 26732 15718 26784
rect 16850 26772 16856 26784
rect 16811 26744 16856 26772
rect 16850 26732 16856 26744
rect 16908 26732 16914 26784
rect 21542 26732 21548 26784
rect 21600 26772 21606 26784
rect 21913 26775 21971 26781
rect 21913 26772 21925 26775
rect 21600 26744 21925 26772
rect 21600 26732 21606 26744
rect 21913 26741 21925 26744
rect 21959 26741 21971 26775
rect 22020 26772 22048 26880
rect 25041 26877 25053 26911
rect 25087 26877 25099 26911
rect 25314 26908 25320 26920
rect 25275 26880 25320 26908
rect 25041 26871 25099 26877
rect 22281 26775 22339 26781
rect 22281 26772 22293 26775
rect 22020 26744 22293 26772
rect 21913 26735 21971 26741
rect 22281 26741 22293 26744
rect 22327 26772 22339 26775
rect 22370 26772 22376 26784
rect 22327 26744 22376 26772
rect 22327 26741 22339 26744
rect 22281 26735 22339 26741
rect 22370 26732 22376 26744
rect 22428 26732 22434 26784
rect 24949 26775 25007 26781
rect 24949 26741 24961 26775
rect 24995 26772 25007 26775
rect 25056 26772 25084 26871
rect 25314 26868 25320 26880
rect 25372 26868 25378 26920
rect 58434 26800 58440 26852
rect 58492 26840 58498 26852
rect 59354 26840 59360 26852
rect 58492 26812 59360 26840
rect 58492 26800 58498 26812
rect 59354 26800 59360 26812
rect 59412 26800 59418 26852
rect 25130 26772 25136 26784
rect 24995 26744 25136 26772
rect 24995 26741 25007 26744
rect 24949 26735 25007 26741
rect 25130 26732 25136 26744
rect 25188 26732 25194 26784
rect 86218 26732 86224 26784
rect 86276 26772 86282 26784
rect 87230 26772 87236 26784
rect 86276 26744 87236 26772
rect 86276 26732 86282 26744
rect 87230 26732 87236 26744
rect 87288 26732 87294 26784
rect 1104 26682 29256 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 29256 26682
rect 1104 26608 29256 26630
rect 58434 26596 58440 26648
rect 58492 26636 58498 26648
rect 59446 26636 59452 26648
rect 58492 26608 59452 26636
rect 58492 26596 58498 26608
rect 59446 26596 59452 26608
rect 59504 26596 59510 26648
rect 5902 26528 5908 26580
rect 5960 26568 5966 26580
rect 6822 26568 6828 26580
rect 5960 26540 6828 26568
rect 5960 26528 5966 26540
rect 6822 26528 6828 26540
rect 6880 26568 6886 26580
rect 7929 26571 7987 26577
rect 7929 26568 7941 26571
rect 6880 26540 7941 26568
rect 6880 26528 6886 26540
rect 7929 26537 7941 26540
rect 7975 26537 7987 26571
rect 7929 26531 7987 26537
rect 16850 26528 16856 26580
rect 16908 26568 16914 26580
rect 22186 26568 22192 26580
rect 16908 26540 22192 26568
rect 16908 26528 16914 26540
rect 22186 26528 22192 26540
rect 22244 26528 22250 26580
rect 22370 26528 22376 26580
rect 22428 26568 22434 26580
rect 23845 26571 23903 26577
rect 23845 26568 23857 26571
rect 22428 26540 23857 26568
rect 22428 26528 22434 26540
rect 23845 26537 23857 26540
rect 23891 26568 23903 26571
rect 27154 26568 27160 26580
rect 23891 26540 27160 26568
rect 23891 26537 23903 26540
rect 23845 26531 23903 26537
rect 27154 26528 27160 26540
rect 27212 26528 27218 26580
rect 17586 26460 17592 26512
rect 17644 26500 17650 26512
rect 17862 26500 17868 26512
rect 17644 26472 17868 26500
rect 17644 26460 17650 26472
rect 17862 26460 17868 26472
rect 17920 26460 17926 26512
rect 4341 26435 4399 26441
rect 4341 26401 4353 26435
rect 4387 26432 4399 26435
rect 4614 26432 4620 26444
rect 4387 26404 4620 26432
rect 4387 26401 4399 26404
rect 4341 26395 4399 26401
rect 4614 26392 4620 26404
rect 4672 26392 4678 26444
rect 6825 26435 6883 26441
rect 6825 26401 6837 26435
rect 6871 26432 6883 26435
rect 7650 26432 7656 26444
rect 6871 26404 7656 26432
rect 6871 26401 6883 26404
rect 6825 26395 6883 26401
rect 7650 26392 7656 26404
rect 7708 26392 7714 26444
rect 16209 26435 16267 26441
rect 16209 26401 16221 26435
rect 16255 26432 16267 26435
rect 17126 26432 17132 26444
rect 16255 26404 17132 26432
rect 16255 26401 16267 26404
rect 16209 26395 16267 26401
rect 17126 26392 17132 26404
rect 17184 26432 17190 26444
rect 21542 26432 21548 26444
rect 17184 26404 17816 26432
rect 21503 26404 21548 26432
rect 17184 26392 17190 26404
rect 4065 26367 4123 26373
rect 4065 26333 4077 26367
rect 4111 26364 4123 26367
rect 4246 26364 4252 26376
rect 4111 26336 4252 26364
rect 4111 26333 4123 26336
rect 4065 26327 4123 26333
rect 4246 26324 4252 26336
rect 4304 26364 4310 26376
rect 5813 26367 5871 26373
rect 5813 26364 5825 26367
rect 4304 26336 5825 26364
rect 4304 26324 4310 26336
rect 5813 26333 5825 26336
rect 5859 26364 5871 26367
rect 6549 26367 6607 26373
rect 6549 26364 6561 26367
rect 5859 26336 6561 26364
rect 5859 26333 5871 26336
rect 5813 26327 5871 26333
rect 6549 26333 6561 26336
rect 6595 26364 6607 26367
rect 8297 26367 8355 26373
rect 8297 26364 8309 26367
rect 6595 26336 8309 26364
rect 6595 26333 6607 26336
rect 6549 26327 6607 26333
rect 8297 26333 8309 26336
rect 8343 26364 8355 26367
rect 9582 26364 9588 26376
rect 8343 26336 9588 26364
rect 8343 26333 8355 26336
rect 8297 26327 8355 26333
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 16485 26367 16543 26373
rect 16485 26333 16497 26367
rect 16531 26364 16543 26367
rect 16666 26364 16672 26376
rect 16531 26336 16672 26364
rect 16531 26333 16543 26336
rect 16485 26327 16543 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17788 26308 17816 26404
rect 21542 26392 21548 26404
rect 21600 26392 21606 26444
rect 22925 26435 22983 26441
rect 22925 26401 22937 26435
rect 22971 26432 22983 26435
rect 23753 26435 23811 26441
rect 23753 26432 23765 26435
rect 22971 26404 23765 26432
rect 22971 26401 22983 26404
rect 22925 26395 22983 26401
rect 23753 26401 23765 26404
rect 23799 26401 23811 26435
rect 23753 26395 23811 26401
rect 25409 26435 25467 26441
rect 25409 26401 25421 26435
rect 25455 26432 25467 26435
rect 26602 26432 26608 26444
rect 25455 26404 26608 26432
rect 25455 26401 25467 26404
rect 25409 26395 25467 26401
rect 26602 26392 26608 26404
rect 26660 26392 26666 26444
rect 26697 26435 26755 26441
rect 26697 26401 26709 26435
rect 26743 26432 26755 26435
rect 27798 26432 27804 26444
rect 26743 26404 27804 26432
rect 26743 26401 26755 26404
rect 26697 26395 26755 26401
rect 27798 26392 27804 26404
rect 27856 26392 27862 26444
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26333 21327 26367
rect 21269 26327 21327 26333
rect 17770 26256 17776 26308
rect 17828 26296 17834 26308
rect 17957 26299 18015 26305
rect 17957 26296 17969 26299
rect 17828 26268 17969 26296
rect 17828 26256 17834 26268
rect 17957 26265 17969 26268
rect 18003 26296 18015 26299
rect 21085 26299 21143 26305
rect 21085 26296 21097 26299
rect 18003 26268 21097 26296
rect 18003 26265 18015 26268
rect 17957 26259 18015 26265
rect 21085 26265 21097 26268
rect 21131 26296 21143 26299
rect 21284 26296 21312 26327
rect 21131 26268 21312 26296
rect 21131 26265 21143 26268
rect 21085 26259 21143 26265
rect 3510 26188 3516 26240
rect 3568 26228 3574 26240
rect 5445 26231 5503 26237
rect 5445 26228 5457 26231
rect 3568 26200 5457 26228
rect 3568 26188 3574 26200
rect 5445 26197 5457 26200
rect 5491 26197 5503 26231
rect 25498 26228 25504 26240
rect 25459 26200 25504 26228
rect 5445 26191 5503 26197
rect 25498 26188 25504 26200
rect 25556 26188 25562 26240
rect 26786 26228 26792 26240
rect 26747 26200 26792 26228
rect 26786 26188 26792 26200
rect 26844 26188 26850 26240
rect 1104 26138 29256 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 29256 26138
rect 1104 26064 29256 26086
rect 3970 25984 3976 26036
rect 4028 26024 4034 26036
rect 6270 26024 6276 26036
rect 4028 25996 6276 26024
rect 4028 25984 4034 25996
rect 6270 25984 6276 25996
rect 6328 25984 6334 26036
rect 7469 26027 7527 26033
rect 7469 25993 7481 26027
rect 7515 26024 7527 26027
rect 8570 26024 8576 26036
rect 7515 25996 8576 26024
rect 7515 25993 7527 25996
rect 7469 25987 7527 25993
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 9306 26024 9312 26036
rect 9267 25996 9312 26024
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 17129 26027 17187 26033
rect 17129 25993 17141 26027
rect 17175 26024 17187 26027
rect 23566 26024 23572 26036
rect 17175 25996 23572 26024
rect 17175 25993 17187 25996
rect 17129 25987 17187 25993
rect 8110 25956 8116 25968
rect 7208 25928 8116 25956
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25888 2927 25891
rect 7208 25888 7236 25928
rect 8110 25916 8116 25928
rect 8168 25916 8174 25968
rect 8481 25959 8539 25965
rect 8481 25925 8493 25959
rect 8527 25956 8539 25959
rect 8662 25956 8668 25968
rect 8527 25928 8668 25956
rect 8527 25925 8539 25928
rect 8481 25919 8539 25925
rect 8662 25916 8668 25928
rect 8720 25956 8726 25968
rect 9401 25959 9459 25965
rect 9401 25956 9413 25959
rect 8720 25928 9413 25956
rect 8720 25916 8726 25928
rect 9401 25925 9413 25928
rect 9447 25925 9459 25959
rect 9401 25919 9459 25925
rect 11974 25916 11980 25968
rect 12032 25956 12038 25968
rect 16666 25956 16672 25968
rect 12032 25928 15792 25956
rect 16627 25928 16672 25956
rect 12032 25916 12038 25928
rect 2915 25860 7236 25888
rect 2915 25857 2927 25860
rect 2869 25851 2927 25857
rect 7282 25848 7288 25900
rect 7340 25888 7346 25900
rect 15381 25891 15439 25897
rect 15381 25888 15393 25891
rect 7340 25860 15393 25888
rect 7340 25848 7346 25860
rect 15381 25857 15393 25860
rect 15427 25888 15439 25891
rect 15565 25891 15623 25897
rect 15565 25888 15577 25891
rect 15427 25860 15577 25888
rect 15427 25857 15439 25860
rect 15381 25851 15439 25857
rect 15565 25857 15577 25860
rect 15611 25857 15623 25891
rect 15565 25851 15623 25857
rect 15764 25888 15792 25928
rect 16666 25916 16672 25928
rect 16724 25916 16730 25968
rect 15764 25860 15976 25888
rect 2590 25820 2596 25832
rect 2551 25792 2596 25820
rect 2590 25780 2596 25792
rect 2648 25780 2654 25832
rect 7006 25780 7012 25832
rect 7064 25820 7070 25832
rect 7377 25823 7435 25829
rect 7377 25820 7389 25823
rect 7064 25792 7389 25820
rect 7064 25780 7070 25792
rect 7377 25789 7389 25792
rect 7423 25789 7435 25823
rect 8386 25820 8392 25832
rect 8347 25792 8392 25820
rect 7377 25783 7435 25789
rect 8386 25780 8392 25792
rect 8444 25780 8450 25832
rect 8662 25820 8668 25832
rect 8575 25792 8668 25820
rect 8662 25780 8668 25792
rect 8720 25820 8726 25832
rect 9306 25820 9312 25832
rect 8720 25792 9312 25820
rect 8720 25780 8726 25792
rect 9306 25780 9312 25792
rect 9364 25780 9370 25832
rect 10965 25823 11023 25829
rect 10965 25789 10977 25823
rect 11011 25820 11023 25823
rect 11011 25792 11192 25820
rect 11011 25789 11023 25792
rect 10965 25783 11023 25789
rect 4154 25684 4160 25696
rect 4115 25656 4160 25684
rect 4154 25644 4160 25656
rect 4212 25644 4218 25696
rect 4433 25687 4491 25693
rect 4433 25653 4445 25687
rect 4479 25684 4491 25687
rect 5442 25684 5448 25696
rect 4479 25656 5448 25684
rect 4479 25653 4491 25656
rect 4433 25647 4491 25653
rect 5442 25644 5448 25656
rect 5500 25644 5506 25696
rect 7742 25644 7748 25696
rect 7800 25684 7806 25696
rect 8849 25687 8907 25693
rect 8849 25684 8861 25687
rect 7800 25656 8861 25684
rect 7800 25644 7806 25656
rect 8849 25653 8861 25656
rect 8895 25653 8907 25687
rect 8849 25647 8907 25653
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 10594 25684 10600 25696
rect 10008 25656 10600 25684
rect 10008 25644 10014 25656
rect 10594 25644 10600 25656
rect 10652 25684 10658 25696
rect 11164 25693 11192 25792
rect 15580 25752 15608 25851
rect 15764 25829 15792 25860
rect 15749 25823 15807 25829
rect 15749 25789 15761 25823
rect 15795 25789 15807 25823
rect 15948 25820 15976 25860
rect 16298 25820 16304 25832
rect 15948 25792 16304 25820
rect 15749 25783 15807 25789
rect 16298 25780 16304 25792
rect 16356 25780 16362 25832
rect 16485 25823 16543 25829
rect 16485 25789 16497 25823
rect 16531 25820 16543 25823
rect 17144 25820 17172 25987
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 25133 26027 25191 26033
rect 25133 25993 25145 26027
rect 25179 26024 25191 26027
rect 25314 26024 25320 26036
rect 25179 25996 25320 26024
rect 25179 25993 25191 25996
rect 25133 25987 25191 25993
rect 25314 25984 25320 25996
rect 25372 25984 25378 26036
rect 27798 26024 27804 26036
rect 27711 25996 27804 26024
rect 27798 25984 27804 25996
rect 27856 26024 27862 26036
rect 28902 26024 28908 26036
rect 27856 25996 28908 26024
rect 27856 25984 27862 25996
rect 28902 25984 28908 25996
rect 28960 25984 28966 26036
rect 16531 25792 17172 25820
rect 16531 25789 16543 25792
rect 16485 25783 16543 25789
rect 17954 25780 17960 25832
rect 18012 25820 18018 25832
rect 18049 25823 18107 25829
rect 18049 25820 18061 25823
rect 18012 25792 18061 25820
rect 18012 25780 18018 25792
rect 18049 25789 18061 25792
rect 18095 25789 18107 25823
rect 18049 25783 18107 25789
rect 23937 25823 23995 25829
rect 23937 25789 23949 25823
rect 23983 25789 23995 25823
rect 24118 25820 24124 25832
rect 24079 25792 24124 25820
rect 23937 25783 23995 25789
rect 19426 25752 19432 25764
rect 15580 25724 19432 25752
rect 19426 25712 19432 25724
rect 19484 25752 19490 25764
rect 23753 25755 23811 25761
rect 23753 25752 23765 25755
rect 19484 25724 23765 25752
rect 19484 25712 19490 25724
rect 23753 25721 23765 25724
rect 23799 25752 23811 25755
rect 23952 25752 23980 25783
rect 24118 25780 24124 25792
rect 24176 25820 24182 25832
rect 24673 25823 24731 25829
rect 24673 25820 24685 25823
rect 24176 25792 24685 25820
rect 24176 25780 24182 25792
rect 24673 25789 24685 25792
rect 24719 25789 24731 25823
rect 24673 25783 24731 25789
rect 24857 25823 24915 25829
rect 24857 25789 24869 25823
rect 24903 25820 24915 25823
rect 25498 25820 25504 25832
rect 24903 25792 25504 25820
rect 24903 25789 24915 25792
rect 24857 25783 24915 25789
rect 25498 25780 25504 25792
rect 25556 25780 25562 25832
rect 26237 25823 26295 25829
rect 26237 25820 26249 25823
rect 26068 25792 26249 25820
rect 23799 25724 23980 25752
rect 23799 25721 23811 25724
rect 23753 25715 23811 25721
rect 10781 25687 10839 25693
rect 10781 25684 10793 25687
rect 10652 25656 10793 25684
rect 10652 25644 10658 25656
rect 10781 25653 10793 25656
rect 10827 25653 10839 25687
rect 10781 25647 10839 25653
rect 11149 25687 11207 25693
rect 11149 25653 11161 25687
rect 11195 25684 11207 25687
rect 15378 25684 15384 25696
rect 11195 25656 15384 25684
rect 11195 25653 11207 25656
rect 11149 25647 11207 25653
rect 15378 25644 15384 25656
rect 15436 25684 15442 25696
rect 15930 25684 15936 25696
rect 15436 25656 15936 25684
rect 15436 25644 15442 25656
rect 15930 25644 15936 25656
rect 15988 25644 15994 25696
rect 18138 25684 18144 25696
rect 18099 25656 18144 25684
rect 18138 25644 18144 25656
rect 18196 25644 18202 25696
rect 25222 25644 25228 25696
rect 25280 25684 25286 25696
rect 26068 25693 26096 25792
rect 26237 25789 26249 25792
rect 26283 25789 26295 25823
rect 26510 25820 26516 25832
rect 26471 25792 26516 25820
rect 26237 25783 26295 25789
rect 26510 25780 26516 25792
rect 26568 25780 26574 25832
rect 26053 25687 26111 25693
rect 26053 25684 26065 25687
rect 25280 25656 26065 25684
rect 25280 25644 25286 25656
rect 26053 25653 26065 25656
rect 26099 25653 26111 25687
rect 26053 25647 26111 25653
rect 1104 25594 29256 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 29256 25594
rect 86218 25576 86224 25628
rect 86276 25616 86282 25628
rect 87138 25616 87144 25628
rect 86276 25588 87144 25616
rect 86276 25576 86282 25588
rect 87138 25576 87144 25588
rect 87196 25576 87202 25628
rect 1104 25520 29256 25542
rect 11054 25440 11060 25492
rect 11112 25480 11118 25492
rect 11974 25480 11980 25492
rect 11112 25452 11980 25480
rect 11112 25440 11118 25452
rect 11974 25440 11980 25452
rect 12032 25440 12038 25492
rect 20806 25480 20812 25492
rect 17328 25452 20812 25480
rect 6917 25347 6975 25353
rect 6917 25313 6929 25347
rect 6963 25344 6975 25347
rect 7006 25344 7012 25356
rect 6963 25316 7012 25344
rect 6963 25313 6975 25316
rect 6917 25307 6975 25313
rect 7006 25304 7012 25316
rect 7064 25304 7070 25356
rect 7742 25344 7748 25356
rect 7703 25316 7748 25344
rect 7742 25304 7748 25316
rect 7800 25304 7806 25356
rect 11793 25347 11851 25353
rect 11793 25313 11805 25347
rect 11839 25344 11851 25347
rect 11974 25344 11980 25356
rect 11839 25316 11980 25344
rect 11839 25313 11851 25316
rect 11793 25307 11851 25313
rect 11974 25304 11980 25316
rect 12032 25304 12038 25356
rect 16298 25304 16304 25356
rect 16356 25344 16362 25356
rect 17328 25353 17356 25452
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 25409 25483 25467 25489
rect 25409 25449 25421 25483
rect 25455 25480 25467 25483
rect 26510 25480 26516 25492
rect 25455 25452 26516 25480
rect 25455 25449 25467 25452
rect 25409 25443 25467 25449
rect 26510 25440 26516 25452
rect 26568 25440 26574 25492
rect 18138 25372 18144 25424
rect 18196 25412 18202 25424
rect 28258 25412 28264 25424
rect 18196 25384 28264 25412
rect 18196 25372 18202 25384
rect 28258 25372 28264 25384
rect 28316 25372 28322 25424
rect 16761 25347 16819 25353
rect 16761 25344 16773 25347
rect 16356 25316 16773 25344
rect 16356 25304 16362 25316
rect 16761 25313 16773 25316
rect 16807 25313 16819 25347
rect 16761 25307 16819 25313
rect 17313 25347 17371 25353
rect 17313 25313 17325 25347
rect 17359 25313 17371 25347
rect 17313 25307 17371 25313
rect 17497 25347 17555 25353
rect 17497 25313 17509 25347
rect 17543 25344 17555 25347
rect 17862 25344 17868 25356
rect 17543 25316 17868 25344
rect 17543 25313 17555 25316
rect 17497 25307 17555 25313
rect 17862 25304 17868 25316
rect 17920 25304 17926 25356
rect 23566 25304 23572 25356
rect 23624 25344 23630 25356
rect 24118 25344 24124 25356
rect 23624 25316 24124 25344
rect 23624 25304 23630 25316
rect 24118 25304 24124 25316
rect 24176 25344 24182 25356
rect 24397 25347 24455 25353
rect 24397 25344 24409 25347
rect 24176 25316 24409 25344
rect 24176 25304 24182 25316
rect 24397 25313 24409 25316
rect 24443 25344 24455 25347
rect 24949 25347 25007 25353
rect 24949 25344 24961 25347
rect 24443 25316 24961 25344
rect 24443 25313 24455 25316
rect 24397 25307 24455 25313
rect 24949 25313 24961 25316
rect 24995 25313 25007 25347
rect 24949 25307 25007 25313
rect 25133 25347 25191 25353
rect 25133 25313 25145 25347
rect 25179 25344 25191 25347
rect 26786 25344 26792 25356
rect 25179 25316 26792 25344
rect 25179 25313 25191 25316
rect 25133 25307 25191 25313
rect 26786 25304 26792 25316
rect 26844 25304 26850 25356
rect 5261 25279 5319 25285
rect 5261 25245 5273 25279
rect 5307 25245 5319 25279
rect 5261 25239 5319 25245
rect 5537 25279 5595 25285
rect 5537 25245 5549 25279
rect 5583 25276 5595 25279
rect 7837 25279 7895 25285
rect 7837 25276 7849 25279
rect 5583 25248 7849 25276
rect 5583 25245 5595 25248
rect 5537 25239 5595 25245
rect 7837 25245 7849 25248
rect 7883 25245 7895 25279
rect 16482 25276 16488 25288
rect 16443 25248 16488 25276
rect 7837 25239 7895 25245
rect 5276 25140 5304 25239
rect 16482 25236 16488 25248
rect 16540 25276 16546 25288
rect 16577 25279 16635 25285
rect 16577 25276 16589 25279
rect 16540 25248 16589 25276
rect 16540 25236 16546 25248
rect 16577 25245 16589 25248
rect 16623 25245 16635 25279
rect 24213 25279 24271 25285
rect 24213 25276 24225 25279
rect 16577 25239 16635 25245
rect 24044 25248 24225 25276
rect 24044 25152 24072 25248
rect 24213 25245 24225 25248
rect 24259 25245 24271 25279
rect 24213 25239 24271 25245
rect 5442 25140 5448 25152
rect 5276 25112 5448 25140
rect 5442 25100 5448 25112
rect 5500 25140 5506 25152
rect 7101 25143 7159 25149
rect 7101 25140 7113 25143
rect 5500 25112 7113 25140
rect 5500 25100 5506 25112
rect 7101 25109 7113 25112
rect 7147 25140 7159 25143
rect 8294 25140 8300 25152
rect 7147 25112 8300 25140
rect 7147 25109 7159 25112
rect 7101 25103 7159 25109
rect 8294 25100 8300 25112
rect 8352 25100 8358 25152
rect 17773 25143 17831 25149
rect 17773 25109 17785 25143
rect 17819 25140 17831 25143
rect 18322 25140 18328 25152
rect 17819 25112 18328 25140
rect 17819 25109 17831 25112
rect 17773 25103 17831 25109
rect 18322 25100 18328 25112
rect 18380 25100 18386 25152
rect 24026 25140 24032 25152
rect 23987 25112 24032 25140
rect 24026 25100 24032 25112
rect 24084 25100 24090 25152
rect 1104 25050 29256 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 29256 25050
rect 1104 24976 29256 24998
rect 13170 24936 13176 24948
rect 13131 24908 13176 24936
rect 13170 24896 13176 24908
rect 13228 24936 13234 24948
rect 14182 24936 14188 24948
rect 13228 24908 14188 24936
rect 13228 24896 13234 24908
rect 14182 24896 14188 24908
rect 14240 24896 14246 24948
rect 10428 24840 11192 24868
rect 2869 24803 2927 24809
rect 2869 24769 2881 24803
rect 2915 24800 2927 24803
rect 3602 24800 3608 24812
rect 2915 24772 3608 24800
rect 2915 24769 2927 24772
rect 2869 24763 2927 24769
rect 3602 24760 3608 24772
rect 3660 24760 3666 24812
rect 8297 24803 8355 24809
rect 8297 24800 8309 24803
rect 7852 24772 8309 24800
rect 7852 24744 7880 24772
rect 8297 24769 8309 24772
rect 8343 24769 8355 24803
rect 8297 24763 8355 24769
rect 10045 24803 10103 24809
rect 10045 24769 10057 24803
rect 10091 24800 10103 24803
rect 10428 24800 10456 24840
rect 10091 24772 10456 24800
rect 11164 24800 11192 24840
rect 12342 24828 12348 24880
rect 12400 24868 12406 24880
rect 13354 24868 13360 24880
rect 12400 24840 13360 24868
rect 12400 24828 12406 24840
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 28994 24868 29000 24880
rect 13648 24840 14688 24868
rect 13538 24800 13544 24812
rect 11164 24772 13544 24800
rect 10091 24769 10103 24772
rect 10045 24763 10103 24769
rect 2590 24732 2596 24744
rect 2551 24704 2596 24732
rect 2590 24692 2596 24704
rect 2648 24692 2654 24744
rect 7466 24732 7472 24744
rect 7427 24704 7472 24732
rect 7466 24692 7472 24704
rect 7524 24692 7530 24744
rect 7561 24735 7619 24741
rect 7561 24701 7573 24735
rect 7607 24701 7619 24735
rect 7834 24732 7840 24744
rect 7795 24704 7840 24732
rect 7561 24695 7619 24701
rect 4249 24667 4307 24673
rect 4249 24633 4261 24667
rect 4295 24664 4307 24667
rect 4614 24664 4620 24676
rect 4295 24636 4620 24664
rect 4295 24633 4307 24636
rect 4249 24627 4307 24633
rect 4614 24624 4620 24636
rect 4672 24624 4678 24676
rect 5718 24624 5724 24676
rect 5776 24664 5782 24676
rect 6825 24667 6883 24673
rect 6825 24664 6837 24667
rect 5776 24636 6837 24664
rect 5776 24624 5782 24636
rect 6825 24633 6837 24636
rect 6871 24633 6883 24667
rect 7576 24664 7604 24695
rect 7834 24692 7840 24704
rect 7892 24692 7898 24744
rect 8018 24732 8024 24744
rect 7979 24704 8024 24732
rect 8018 24692 8024 24704
rect 8076 24692 8082 24744
rect 8113 24735 8171 24741
rect 8113 24701 8125 24735
rect 8159 24732 8171 24735
rect 8662 24732 8668 24744
rect 8159 24704 8668 24732
rect 8159 24701 8171 24704
rect 8113 24695 8171 24701
rect 8128 24664 8156 24695
rect 8662 24692 8668 24704
rect 8720 24692 8726 24744
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24732 9459 24735
rect 9950 24732 9956 24744
rect 9447 24704 9956 24732
rect 9447 24701 9459 24704
rect 9401 24695 9459 24701
rect 9950 24692 9956 24704
rect 10008 24692 10014 24744
rect 7576 24636 8156 24664
rect 6825 24627 6883 24633
rect 8202 24624 8208 24676
rect 8260 24664 8266 24676
rect 9861 24667 9919 24673
rect 9861 24664 9873 24667
rect 8260 24636 9873 24664
rect 8260 24624 8266 24636
rect 9861 24633 9873 24636
rect 9907 24664 9919 24667
rect 10060 24664 10088 24763
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 13648 24809 13676 24840
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24769 13691 24803
rect 14660 24800 14688 24840
rect 26344 24840 29000 24868
rect 15654 24800 15660 24812
rect 14660 24772 15660 24800
rect 13633 24763 13691 24769
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 18322 24800 18328 24812
rect 18283 24772 18328 24800
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 19484 24772 19717 24800
rect 19484 24760 19490 24772
rect 19705 24769 19717 24772
rect 19751 24800 19763 24803
rect 20530 24800 20536 24812
rect 19751 24772 20536 24800
rect 19751 24769 19763 24772
rect 19705 24763 19763 24769
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 25501 24803 25559 24809
rect 25501 24769 25513 24803
rect 25547 24800 25559 24803
rect 26344 24800 26372 24840
rect 28994 24828 29000 24840
rect 29052 24828 29058 24880
rect 25547 24772 26372 24800
rect 25547 24769 25559 24772
rect 25501 24763 25559 24769
rect 10229 24735 10287 24741
rect 10229 24701 10241 24735
rect 10275 24701 10287 24735
rect 10229 24695 10287 24701
rect 10781 24735 10839 24741
rect 10781 24701 10793 24735
rect 10827 24701 10839 24735
rect 10781 24695 10839 24701
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 11011 24704 11652 24732
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 9907 24636 10088 24664
rect 10244 24664 10272 24695
rect 10796 24664 10824 24695
rect 11054 24664 11060 24676
rect 10244 24636 11060 24664
rect 9907 24633 9919 24636
rect 9861 24627 9919 24633
rect 11054 24624 11060 24636
rect 11112 24624 11118 24676
rect 4433 24599 4491 24605
rect 4433 24565 4445 24599
rect 4479 24596 4491 24599
rect 5442 24596 5448 24608
rect 4479 24568 5448 24596
rect 4479 24565 4491 24568
rect 4433 24559 4491 24565
rect 5442 24556 5448 24568
rect 5500 24556 5506 24608
rect 9217 24599 9275 24605
rect 9217 24565 9229 24599
rect 9263 24596 9275 24599
rect 9582 24596 9588 24608
rect 9263 24568 9588 24596
rect 9263 24565 9275 24568
rect 9217 24559 9275 24565
rect 9582 24556 9588 24568
rect 9640 24556 9646 24608
rect 9950 24556 9956 24608
rect 10008 24596 10014 24608
rect 11624 24605 11652 24704
rect 11698 24692 11704 24744
rect 11756 24732 11762 24744
rect 12437 24735 12495 24741
rect 12437 24732 12449 24735
rect 11756 24704 12449 24732
rect 11756 24692 11762 24704
rect 12437 24701 12449 24704
rect 12483 24701 12495 24735
rect 12437 24695 12495 24701
rect 13710 24735 13768 24741
rect 13710 24701 13722 24735
rect 13756 24701 13768 24735
rect 14182 24732 14188 24744
rect 14143 24704 14188 24732
rect 13710 24695 13768 24701
rect 13740 24608 13768 24695
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 15887 24735 15945 24741
rect 15887 24732 15899 24735
rect 14332 24704 14377 24732
rect 15764 24704 15899 24732
rect 14332 24692 14338 24704
rect 15764 24664 15792 24704
rect 15887 24701 15899 24704
rect 15933 24701 15945 24735
rect 16022 24732 16028 24744
rect 15983 24704 16028 24732
rect 15887 24695 15945 24701
rect 16022 24692 16028 24704
rect 16080 24692 16086 24744
rect 16485 24735 16543 24741
rect 16485 24701 16497 24735
rect 16531 24701 16543 24735
rect 16485 24695 16543 24701
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24701 16727 24735
rect 16669 24695 16727 24701
rect 16390 24664 16396 24676
rect 15764 24636 16396 24664
rect 16390 24624 16396 24636
rect 16448 24664 16454 24676
rect 16500 24664 16528 24695
rect 16448 24636 16528 24664
rect 16684 24664 16712 24695
rect 16942 24692 16948 24744
rect 17000 24732 17006 24744
rect 17865 24735 17923 24741
rect 17865 24732 17877 24735
rect 17000 24704 17877 24732
rect 17000 24692 17006 24704
rect 17865 24701 17877 24704
rect 17911 24732 17923 24735
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 17911 24704 18061 24732
rect 17911 24701 17923 24704
rect 17865 24695 17923 24701
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24701 23903 24735
rect 23845 24695 23903 24701
rect 24121 24735 24179 24741
rect 24121 24701 24133 24735
rect 24167 24732 24179 24735
rect 24486 24732 24492 24744
rect 24167 24704 24492 24732
rect 24167 24701 24179 24704
rect 24121 24695 24179 24701
rect 17313 24667 17371 24673
rect 17313 24664 17325 24667
rect 16684 24636 17325 24664
rect 16448 24624 16454 24636
rect 17313 24633 17325 24636
rect 17359 24664 17371 24667
rect 18138 24664 18144 24676
rect 17359 24636 18144 24664
rect 17359 24633 17371 24636
rect 17313 24627 17371 24633
rect 18138 24624 18144 24636
rect 18196 24624 18202 24676
rect 11241 24599 11299 24605
rect 11241 24596 11253 24599
rect 10008 24568 11253 24596
rect 10008 24556 10014 24568
rect 11241 24565 11253 24568
rect 11287 24565 11299 24599
rect 11241 24559 11299 24565
rect 11609 24599 11667 24605
rect 11609 24565 11621 24599
rect 11655 24596 11667 24599
rect 12529 24599 12587 24605
rect 12529 24596 12541 24599
rect 11655 24568 12541 24596
rect 11655 24565 11667 24568
rect 11609 24559 11667 24565
rect 12529 24565 12541 24568
rect 12575 24596 12587 24599
rect 13078 24596 13084 24608
rect 12575 24568 13084 24596
rect 12575 24565 12587 24568
rect 12529 24559 12587 24565
rect 13078 24556 13084 24568
rect 13136 24556 13142 24608
rect 13722 24556 13728 24608
rect 13780 24556 13786 24608
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14240 24568 14749 24596
rect 14240 24556 14246 24568
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 14737 24559 14795 24565
rect 15657 24599 15715 24605
rect 15657 24565 15669 24599
rect 15703 24596 15715 24599
rect 16022 24596 16028 24608
rect 15703 24568 16028 24596
rect 15703 24565 15715 24568
rect 15657 24559 15715 24565
rect 16022 24556 16028 24568
rect 16080 24556 16086 24608
rect 16850 24556 16856 24608
rect 16908 24596 16914 24608
rect 16945 24599 17003 24605
rect 16945 24596 16957 24599
rect 16908 24568 16957 24596
rect 16908 24556 16914 24568
rect 16945 24565 16957 24568
rect 16991 24565 17003 24599
rect 16945 24559 17003 24565
rect 20714 24556 20720 24608
rect 20772 24596 20778 24608
rect 23753 24599 23811 24605
rect 23753 24596 23765 24599
rect 20772 24568 23765 24596
rect 20772 24556 20778 24568
rect 23753 24565 23765 24568
rect 23799 24596 23811 24599
rect 23860 24596 23888 24695
rect 24486 24692 24492 24704
rect 24544 24692 24550 24744
rect 26344 24741 26372 24772
rect 26329 24735 26387 24741
rect 26329 24701 26341 24735
rect 26375 24701 26387 24735
rect 26329 24695 26387 24701
rect 25222 24596 25228 24608
rect 23799 24568 25228 24596
rect 23799 24565 23811 24568
rect 23753 24559 23811 24565
rect 25222 24556 25228 24568
rect 25280 24556 25286 24608
rect 25314 24556 25320 24608
rect 25372 24596 25378 24608
rect 26421 24599 26479 24605
rect 26421 24596 26433 24599
rect 25372 24568 26433 24596
rect 25372 24556 25378 24568
rect 26421 24565 26433 24568
rect 26467 24565 26479 24599
rect 26421 24559 26479 24565
rect 1104 24506 29256 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 29256 24506
rect 1104 24432 29256 24454
rect 3970 24352 3976 24404
rect 4028 24392 4034 24404
rect 9766 24392 9772 24404
rect 4028 24364 9772 24392
rect 4028 24352 4034 24364
rect 9766 24352 9772 24364
rect 9824 24352 9830 24404
rect 13538 24352 13544 24404
rect 13596 24392 13602 24404
rect 16022 24392 16028 24404
rect 13596 24364 16028 24392
rect 13596 24352 13602 24364
rect 16022 24352 16028 24364
rect 16080 24352 16086 24404
rect 16482 24352 16488 24404
rect 16540 24392 16546 24404
rect 23109 24395 23167 24401
rect 23109 24392 23121 24395
rect 16540 24364 23121 24392
rect 16540 24352 16546 24364
rect 23109 24361 23121 24364
rect 23155 24361 23167 24395
rect 24486 24392 24492 24404
rect 24447 24364 24492 24392
rect 23109 24355 23167 24361
rect 13998 24284 14004 24336
rect 14056 24324 14062 24336
rect 16500 24324 16528 24352
rect 19889 24327 19947 24333
rect 19889 24324 19901 24327
rect 14056 24296 16528 24324
rect 19720 24296 19901 24324
rect 14056 24284 14062 24296
rect 5353 24259 5411 24265
rect 5353 24225 5365 24259
rect 5399 24256 5411 24259
rect 5442 24256 5448 24268
rect 5399 24228 5448 24256
rect 5399 24225 5411 24228
rect 5353 24219 5411 24225
rect 5442 24216 5448 24228
rect 5500 24216 5506 24268
rect 9950 24256 9956 24268
rect 9911 24228 9956 24256
rect 9950 24216 9956 24228
rect 10008 24216 10014 24268
rect 15473 24259 15531 24265
rect 15473 24225 15485 24259
rect 15519 24256 15531 24259
rect 15838 24256 15844 24268
rect 15519 24228 15844 24256
rect 15519 24225 15531 24228
rect 15473 24219 15531 24225
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 16850 24256 16856 24268
rect 16811 24228 16856 24256
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 19720 24265 19748 24296
rect 19889 24293 19901 24296
rect 19935 24324 19947 24327
rect 20990 24324 20996 24336
rect 19935 24296 20996 24324
rect 19935 24293 19947 24296
rect 19889 24287 19947 24293
rect 20990 24284 20996 24296
rect 21048 24324 21054 24336
rect 21048 24296 23060 24324
rect 21048 24284 21054 24296
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24225 19763 24259
rect 19705 24219 19763 24225
rect 22189 24259 22247 24265
rect 22189 24225 22201 24259
rect 22235 24225 22247 24259
rect 22189 24219 22247 24225
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24188 5687 24191
rect 5810 24188 5816 24200
rect 5675 24160 5816 24188
rect 5675 24157 5687 24160
rect 5629 24151 5687 24157
rect 5810 24148 5816 24160
rect 5868 24148 5874 24200
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24188 7251 24191
rect 8294 24188 8300 24200
rect 7239 24160 8300 24188
rect 7239 24157 7251 24160
rect 7193 24151 7251 24157
rect 8294 24148 8300 24160
rect 8352 24188 8358 24200
rect 9493 24191 9551 24197
rect 9493 24188 9505 24191
rect 8352 24160 9505 24188
rect 8352 24148 8358 24160
rect 9493 24157 9505 24160
rect 9539 24188 9551 24191
rect 9582 24188 9588 24200
rect 9539 24160 9588 24188
rect 9539 24157 9551 24160
rect 9493 24151 9551 24157
rect 9582 24148 9588 24160
rect 9640 24188 9646 24200
rect 9677 24191 9735 24197
rect 9677 24188 9689 24191
rect 9640 24160 9689 24188
rect 9640 24148 9646 24160
rect 9677 24157 9689 24160
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 15565 24191 15623 24197
rect 15565 24157 15577 24191
rect 15611 24188 15623 24191
rect 15746 24188 15752 24200
rect 15611 24160 15752 24188
rect 15611 24157 15623 24160
rect 15565 24151 15623 24157
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 16577 24191 16635 24197
rect 16577 24157 16589 24191
rect 16623 24188 16635 24191
rect 16758 24188 16764 24200
rect 16623 24160 16764 24188
rect 16623 24157 16635 24160
rect 16577 24151 16635 24157
rect 16758 24148 16764 24160
rect 16816 24188 16822 24200
rect 17770 24188 17776 24200
rect 16816 24160 17776 24188
rect 16816 24148 16822 24160
rect 17770 24148 17776 24160
rect 17828 24188 17834 24200
rect 18325 24191 18383 24197
rect 18325 24188 18337 24191
rect 17828 24160 18337 24188
rect 17828 24148 17834 24160
rect 18325 24157 18337 24160
rect 18371 24188 18383 24191
rect 20714 24188 20720 24200
rect 18371 24160 20720 24188
rect 18371 24157 18383 24160
rect 18325 24151 18383 24157
rect 20714 24148 20720 24160
rect 20772 24148 20778 24200
rect 19521 24123 19579 24129
rect 19521 24120 19533 24123
rect 17512 24092 19533 24120
rect 6914 24052 6920 24064
rect 6875 24024 6920 24052
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 11146 24012 11152 24064
rect 11204 24052 11210 24064
rect 11241 24055 11299 24061
rect 11241 24052 11253 24055
rect 11204 24024 11253 24052
rect 11204 24012 11210 24024
rect 11241 24021 11253 24024
rect 11287 24052 11299 24055
rect 11698 24052 11704 24064
rect 11287 24024 11704 24052
rect 11287 24021 11299 24024
rect 11241 24015 11299 24021
rect 11698 24012 11704 24024
rect 11756 24012 11762 24064
rect 15838 24052 15844 24064
rect 15799 24024 15844 24052
rect 15838 24012 15844 24024
rect 15896 24012 15902 24064
rect 15930 24012 15936 24064
rect 15988 24052 15994 24064
rect 17512 24052 17540 24092
rect 19521 24089 19533 24092
rect 19567 24089 19579 24123
rect 19521 24083 19579 24089
rect 22097 24123 22155 24129
rect 22097 24089 22109 24123
rect 22143 24120 22155 24123
rect 22204 24120 22232 24219
rect 23032 24188 23060 24296
rect 23124 24256 23152 24355
rect 24486 24352 24492 24364
rect 24544 24352 24550 24404
rect 28629 24395 28687 24401
rect 28629 24361 28641 24395
rect 28675 24392 28687 24395
rect 28718 24392 28724 24404
rect 28675 24364 28724 24392
rect 28675 24361 28687 24364
rect 28629 24355 28687 24361
rect 28718 24352 28724 24364
rect 28776 24352 28782 24404
rect 28353 24327 28411 24333
rect 28353 24324 28365 24327
rect 23400 24296 28365 24324
rect 23293 24259 23351 24265
rect 23293 24256 23305 24259
rect 23124 24228 23305 24256
rect 23293 24225 23305 24228
rect 23339 24225 23351 24259
rect 23293 24219 23351 24225
rect 23400 24188 23428 24296
rect 28353 24293 28365 24296
rect 28399 24293 28411 24327
rect 28353 24287 28411 24293
rect 23477 24259 23535 24265
rect 23477 24225 23489 24259
rect 23523 24256 23535 24259
rect 23566 24256 23572 24268
rect 23523 24228 23572 24256
rect 23523 24225 23535 24228
rect 23477 24219 23535 24225
rect 23566 24216 23572 24228
rect 23624 24216 23630 24268
rect 24029 24259 24087 24265
rect 24029 24225 24041 24259
rect 24075 24256 24087 24259
rect 24118 24256 24124 24268
rect 24075 24228 24124 24256
rect 24075 24225 24087 24228
rect 24029 24219 24087 24225
rect 24118 24216 24124 24228
rect 24176 24216 24182 24268
rect 24213 24259 24271 24265
rect 24213 24225 24225 24259
rect 24259 24256 24271 24259
rect 25314 24256 25320 24268
rect 24259 24228 25320 24256
rect 24259 24225 24271 24228
rect 24213 24219 24271 24225
rect 25314 24216 25320 24228
rect 25372 24216 25378 24268
rect 26510 24256 26516 24268
rect 26471 24228 26516 24256
rect 26510 24216 26516 24228
rect 26568 24216 26574 24268
rect 27341 24259 27399 24265
rect 27341 24225 27353 24259
rect 27387 24225 27399 24259
rect 28736 24256 28764 24352
rect 28905 24259 28963 24265
rect 28905 24256 28917 24259
rect 28736 24228 28917 24256
rect 27341 24219 27399 24225
rect 28905 24225 28917 24228
rect 28951 24225 28963 24259
rect 28905 24219 28963 24225
rect 23032 24160 23428 24188
rect 22462 24120 22468 24132
rect 22143 24092 22468 24120
rect 22143 24089 22155 24092
rect 22097 24083 22155 24089
rect 22462 24080 22468 24092
rect 22520 24080 22526 24132
rect 17954 24052 17960 24064
rect 15988 24024 17540 24052
rect 17915 24024 17960 24052
rect 15988 24012 15994 24024
rect 17954 24012 17960 24024
rect 18012 24012 18018 24064
rect 22373 24055 22431 24061
rect 22373 24021 22385 24055
rect 22419 24052 22431 24055
rect 23584 24052 23612 24216
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 27356 24188 27384 24219
rect 86218 24216 86224 24268
rect 86276 24256 86282 24268
rect 86954 24256 86960 24268
rect 86276 24228 86960 24256
rect 86276 24216 86282 24228
rect 86954 24216 86960 24228
rect 87012 24216 87018 24268
rect 28994 24188 29000 24200
rect 26292 24160 29000 24188
rect 26292 24148 26298 24160
rect 28994 24148 29000 24160
rect 29052 24148 29058 24200
rect 25038 24080 25044 24132
rect 25096 24120 25102 24132
rect 27433 24123 27491 24129
rect 27433 24120 27445 24123
rect 25096 24092 27445 24120
rect 25096 24080 25102 24092
rect 27433 24089 27445 24092
rect 27479 24089 27491 24123
rect 27433 24083 27491 24089
rect 28353 24123 28411 24129
rect 28353 24089 28365 24123
rect 28399 24120 28411 24123
rect 28721 24123 28779 24129
rect 28721 24120 28733 24123
rect 28399 24092 28733 24120
rect 28399 24089 28411 24092
rect 28353 24083 28411 24089
rect 28721 24089 28733 24092
rect 28767 24089 28779 24123
rect 28721 24083 28779 24089
rect 26694 24052 26700 24064
rect 22419 24024 23612 24052
rect 26655 24024 26700 24052
rect 22419 24021 22431 24024
rect 22373 24015 22431 24021
rect 26694 24012 26700 24024
rect 26752 24012 26758 24064
rect 1104 23962 29256 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 29256 23962
rect 1104 23888 29256 23910
rect 4433 23851 4491 23857
rect 4433 23817 4445 23851
rect 4479 23848 4491 23851
rect 5442 23848 5448 23860
rect 4479 23820 5448 23848
rect 4479 23817 4491 23820
rect 4433 23811 4491 23817
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 5810 23848 5816 23860
rect 5771 23820 5816 23848
rect 5810 23808 5816 23820
rect 5868 23808 5874 23860
rect 11241 23851 11299 23857
rect 11241 23817 11253 23851
rect 11287 23848 11299 23851
rect 12342 23848 12348 23860
rect 11287 23820 12348 23848
rect 11287 23817 11299 23820
rect 11241 23811 11299 23817
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 14090 23848 14096 23860
rect 14003 23820 14096 23848
rect 14090 23808 14096 23820
rect 14148 23848 14154 23860
rect 16942 23848 16948 23860
rect 14148 23820 16948 23848
rect 14148 23808 14154 23820
rect 16942 23808 16948 23820
rect 17000 23808 17006 23860
rect 18046 23808 18052 23860
rect 18104 23848 18110 23860
rect 18417 23851 18475 23857
rect 18417 23848 18429 23851
rect 18104 23820 18429 23848
rect 18104 23808 18110 23820
rect 18417 23817 18429 23820
rect 18463 23848 18475 23851
rect 19426 23848 19432 23860
rect 18463 23820 19432 23848
rect 18463 23817 18475 23820
rect 18417 23811 18475 23817
rect 19426 23808 19432 23820
rect 19484 23808 19490 23860
rect 23937 23851 23995 23857
rect 23937 23817 23949 23851
rect 23983 23848 23995 23851
rect 26234 23848 26240 23860
rect 23983 23820 26096 23848
rect 26195 23820 26240 23848
rect 23983 23817 23995 23820
rect 23937 23811 23995 23817
rect 9582 23740 9588 23792
rect 9640 23780 9646 23792
rect 10413 23783 10471 23789
rect 10413 23780 10425 23783
rect 9640 23752 10425 23780
rect 9640 23740 9646 23752
rect 10413 23749 10425 23752
rect 10459 23780 10471 23783
rect 14108 23780 14136 23808
rect 10459 23752 14136 23780
rect 10459 23749 10471 23752
rect 10413 23743 10471 23749
rect 16022 23740 16028 23792
rect 16080 23780 16086 23792
rect 24026 23780 24032 23792
rect 16080 23752 24032 23780
rect 16080 23740 16086 23752
rect 24026 23740 24032 23752
rect 24084 23740 24090 23792
rect 26068 23780 26096 23820
rect 26234 23808 26240 23820
rect 26292 23808 26298 23860
rect 28629 23851 28687 23857
rect 28629 23817 28641 23851
rect 28675 23848 28687 23851
rect 28718 23848 28724 23860
rect 28675 23820 28724 23848
rect 28675 23817 28687 23820
rect 28629 23811 28687 23817
rect 28718 23808 28724 23820
rect 28776 23808 28782 23860
rect 26510 23780 26516 23792
rect 26068 23752 26516 23780
rect 26510 23740 26516 23752
rect 26568 23740 26574 23792
rect 2869 23715 2927 23721
rect 2869 23681 2881 23715
rect 2915 23712 2927 23715
rect 3878 23712 3884 23724
rect 2915 23684 3884 23712
rect 2915 23681 2927 23684
rect 2869 23675 2927 23681
rect 3878 23672 3884 23684
rect 3936 23672 3942 23724
rect 7466 23712 7472 23724
rect 7427 23684 7472 23712
rect 7466 23672 7472 23684
rect 7524 23672 7530 23724
rect 8573 23715 8631 23721
rect 8573 23681 8585 23715
rect 8619 23712 8631 23715
rect 9600 23712 9628 23740
rect 8619 23684 9628 23712
rect 8619 23681 8631 23684
rect 8573 23675 8631 23681
rect 13078 23672 13084 23724
rect 13136 23712 13142 23724
rect 26878 23712 26884 23724
rect 13136 23684 26884 23712
rect 13136 23672 13142 23684
rect 26878 23672 26884 23684
rect 26936 23672 26942 23724
rect 2590 23644 2596 23656
rect 2551 23616 2596 23644
rect 2590 23604 2596 23616
rect 2648 23604 2654 23656
rect 5718 23644 5724 23656
rect 5679 23616 5724 23644
rect 5718 23604 5724 23616
rect 5776 23604 5782 23656
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 7101 23647 7159 23653
rect 7101 23644 7113 23647
rect 6972 23616 7113 23644
rect 6972 23604 6978 23616
rect 7101 23613 7113 23616
rect 7147 23613 7159 23647
rect 7101 23607 7159 23613
rect 7377 23647 7435 23653
rect 7377 23613 7389 23647
rect 7423 23644 7435 23647
rect 7926 23644 7932 23656
rect 7423 23616 7932 23644
rect 7423 23613 7435 23616
rect 7377 23607 7435 23613
rect 7116 23576 7144 23607
rect 7926 23604 7932 23616
rect 7984 23604 7990 23656
rect 8846 23644 8852 23656
rect 8807 23616 8852 23644
rect 8846 23604 8852 23616
rect 8904 23604 8910 23656
rect 11057 23647 11115 23653
rect 11057 23613 11069 23647
rect 11103 23644 11115 23647
rect 11103 23616 11137 23644
rect 11103 23613 11115 23616
rect 11057 23607 11115 23613
rect 10226 23576 10232 23588
rect 7116 23548 7788 23576
rect 10187 23548 10232 23576
rect 7760 23520 7788 23548
rect 10226 23536 10232 23548
rect 10284 23536 10290 23588
rect 10965 23579 11023 23585
rect 10965 23545 10977 23579
rect 11011 23576 11023 23579
rect 11072 23576 11100 23607
rect 14090 23604 14096 23656
rect 14148 23644 14154 23656
rect 14185 23647 14243 23653
rect 14185 23644 14197 23647
rect 14148 23616 14197 23644
rect 14148 23604 14154 23616
rect 14185 23613 14197 23616
rect 14231 23613 14243 23647
rect 14185 23607 14243 23613
rect 14461 23647 14519 23653
rect 14461 23613 14473 23647
rect 14507 23644 14519 23647
rect 14826 23644 14832 23656
rect 14507 23616 14832 23644
rect 14507 23613 14519 23616
rect 14461 23607 14519 23613
rect 14826 23604 14832 23616
rect 14884 23604 14890 23656
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 21821 23647 21879 23653
rect 21821 23613 21833 23647
rect 21867 23644 21879 23647
rect 21867 23616 22232 23644
rect 21867 23613 21879 23616
rect 21821 23607 21879 23613
rect 11330 23576 11336 23588
rect 11011 23548 11336 23576
rect 11011 23545 11023 23548
rect 10965 23539 11023 23545
rect 11330 23536 11336 23548
rect 11388 23536 11394 23588
rect 15838 23576 15844 23588
rect 15799 23548 15844 23576
rect 15838 23536 15844 23548
rect 15896 23536 15902 23588
rect 3970 23508 3976 23520
rect 3931 23480 3976 23508
rect 3970 23468 3976 23480
rect 4028 23468 4034 23520
rect 7742 23508 7748 23520
rect 7703 23480 7748 23508
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 17862 23468 17868 23520
rect 17920 23508 17926 23520
rect 18141 23511 18199 23517
rect 18141 23508 18153 23511
rect 17920 23480 18153 23508
rect 17920 23468 17926 23480
rect 18141 23477 18153 23480
rect 18187 23477 18199 23511
rect 21910 23508 21916 23520
rect 21871 23480 21916 23508
rect 18141 23471 18199 23477
rect 21910 23468 21916 23480
rect 21968 23468 21974 23520
rect 22204 23517 22232 23616
rect 22462 23604 22468 23656
rect 22520 23644 22526 23656
rect 23753 23647 23811 23653
rect 23753 23644 23765 23647
rect 22520 23616 23765 23644
rect 22520 23604 22526 23616
rect 23753 23613 23765 23616
rect 23799 23644 23811 23647
rect 24673 23647 24731 23653
rect 23799 23616 24256 23644
rect 23799 23613 23811 23616
rect 23753 23607 23811 23613
rect 24228 23520 24256 23616
rect 24673 23613 24685 23647
rect 24719 23613 24731 23647
rect 24673 23607 24731 23613
rect 24949 23647 25007 23653
rect 24949 23613 24961 23647
rect 24995 23644 25007 23647
rect 25406 23644 25412 23656
rect 24995 23616 25412 23644
rect 24995 23613 25007 23616
rect 24949 23607 25007 23613
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 22554 23508 22560 23520
rect 22235 23480 22560 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 24210 23508 24216 23520
rect 24171 23480 24216 23508
rect 24210 23468 24216 23480
rect 24268 23468 24274 23520
rect 24581 23511 24639 23517
rect 24581 23477 24593 23511
rect 24627 23508 24639 23511
rect 24688 23508 24716 23607
rect 25406 23604 25412 23616
rect 25464 23604 25470 23656
rect 58434 23604 58440 23656
rect 58492 23644 58498 23656
rect 58986 23644 58992 23656
rect 58492 23616 58992 23644
rect 58492 23604 58498 23616
rect 58986 23604 58992 23616
rect 59044 23604 59050 23656
rect 27065 23579 27123 23585
rect 27065 23545 27077 23579
rect 27111 23576 27123 23579
rect 27154 23576 27160 23588
rect 27111 23548 27160 23576
rect 27111 23545 27123 23548
rect 27065 23539 27123 23545
rect 27154 23536 27160 23548
rect 27212 23536 27218 23588
rect 25222 23508 25228 23520
rect 24627 23480 25228 23508
rect 24627 23477 24639 23480
rect 24581 23471 24639 23477
rect 25222 23468 25228 23480
rect 25280 23468 25286 23520
rect 1104 23418 29256 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 29256 23418
rect 1104 23344 29256 23366
rect 10226 23264 10232 23316
rect 10284 23304 10290 23316
rect 32030 23304 32036 23316
rect 10284 23276 32036 23304
rect 10284 23264 10290 23276
rect 32030 23264 32036 23276
rect 32088 23264 32094 23316
rect 10686 23196 10692 23248
rect 10744 23236 10750 23248
rect 11974 23236 11980 23248
rect 10744 23208 11744 23236
rect 11935 23208 11980 23236
rect 10744 23196 10750 23208
rect 11716 23180 11744 23208
rect 11974 23196 11980 23208
rect 12032 23196 12038 23248
rect 15105 23239 15163 23245
rect 15105 23205 15117 23239
rect 15151 23236 15163 23239
rect 15194 23236 15200 23248
rect 15151 23208 15200 23236
rect 15151 23205 15163 23208
rect 15105 23199 15163 23205
rect 15194 23196 15200 23208
rect 15252 23236 15258 23248
rect 20714 23236 20720 23248
rect 15252 23208 16344 23236
rect 20675 23208 20720 23236
rect 15252 23196 15258 23208
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23137 11575 23171
rect 11517 23131 11575 23137
rect 3326 23060 3332 23112
rect 3384 23100 3390 23112
rect 4614 23100 4620 23112
rect 3384 23072 4620 23100
rect 3384 23060 3390 23072
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 11532 23100 11560 23131
rect 11698 23128 11704 23180
rect 11756 23168 11762 23180
rect 12158 23168 12164 23180
rect 11756 23140 11801 23168
rect 11900 23140 12164 23168
rect 11756 23128 11762 23140
rect 11900 23100 11928 23140
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 16316 23177 16344 23208
rect 20714 23196 20720 23208
rect 20772 23236 20778 23248
rect 22554 23236 22560 23248
rect 20772 23208 20944 23236
rect 22515 23208 22560 23236
rect 20772 23196 20778 23208
rect 14185 23171 14243 23177
rect 14185 23168 14197 23171
rect 14016 23140 14197 23168
rect 14016 23109 14044 23140
rect 14185 23137 14197 23140
rect 14231 23137 14243 23171
rect 15933 23171 15991 23177
rect 15933 23168 15945 23171
rect 14185 23131 14243 23137
rect 14844 23140 15945 23168
rect 14001 23103 14059 23109
rect 14001 23100 14013 23103
rect 11532 23072 11928 23100
rect 11992 23072 14013 23100
rect 9674 22924 9680 22976
rect 9732 22964 9738 22976
rect 11992 22964 12020 23072
rect 14001 23069 14013 23072
rect 14047 23069 14059 23103
rect 14001 23063 14059 23069
rect 12158 22964 12164 22976
rect 9732 22936 12020 22964
rect 12119 22936 12164 22964
rect 9732 22924 9738 22936
rect 12158 22924 12164 22936
rect 12216 22924 12222 22976
rect 13722 22924 13728 22976
rect 13780 22964 13786 22976
rect 14274 22964 14280 22976
rect 13780 22936 14280 22964
rect 13780 22924 13786 22936
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14734 22924 14740 22976
rect 14792 22964 14798 22976
rect 14844 22973 14872 23140
rect 15933 23137 15945 23140
rect 15979 23137 15991 23171
rect 15933 23131 15991 23137
rect 16301 23171 16359 23177
rect 16301 23137 16313 23171
rect 16347 23137 16359 23171
rect 16301 23131 16359 23137
rect 16485 23171 16543 23177
rect 16485 23137 16497 23171
rect 16531 23168 16543 23171
rect 17862 23168 17868 23180
rect 16531 23140 17868 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 20916 23177 20944 23208
rect 22554 23196 22560 23208
rect 22612 23196 22618 23248
rect 24118 23196 24124 23248
rect 24176 23196 24182 23248
rect 25406 23236 25412 23248
rect 24872 23208 25268 23236
rect 25367 23208 25412 23236
rect 20901 23171 20959 23177
rect 20901 23137 20913 23171
rect 20947 23137 20959 23171
rect 24136 23168 24164 23196
rect 24872 23177 24900 23208
rect 24305 23171 24363 23177
rect 24305 23168 24317 23171
rect 24136 23140 24317 23168
rect 20901 23131 20959 23137
rect 24305 23137 24317 23140
rect 24351 23168 24363 23171
rect 24857 23171 24915 23177
rect 24857 23168 24869 23171
rect 24351 23140 24869 23168
rect 24351 23137 24363 23140
rect 24305 23131 24363 23137
rect 24857 23137 24869 23140
rect 24903 23137 24915 23171
rect 25038 23168 25044 23180
rect 24999 23140 25044 23168
rect 24857 23131 24915 23137
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 25240 23168 25268 23208
rect 25406 23196 25412 23208
rect 25464 23196 25470 23248
rect 26694 23168 26700 23180
rect 25240 23140 26700 23168
rect 26694 23128 26700 23140
rect 26752 23168 26758 23180
rect 27249 23171 27307 23177
rect 27249 23168 27261 23171
rect 26752 23140 27261 23168
rect 26752 23128 26758 23140
rect 27249 23137 27261 23140
rect 27295 23137 27307 23171
rect 27249 23131 27307 23137
rect 27433 23171 27491 23177
rect 27433 23137 27445 23171
rect 27479 23168 27491 23171
rect 27706 23168 27712 23180
rect 27479 23140 27712 23168
rect 27479 23137 27491 23140
rect 27433 23131 27491 23137
rect 27706 23128 27712 23140
rect 27764 23128 27770 23180
rect 15746 23100 15752 23112
rect 15707 23072 15752 23100
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 21174 23100 21180 23112
rect 21135 23072 21180 23100
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 23937 23103 23995 23109
rect 23937 23100 23949 23103
rect 22572 23072 23949 23100
rect 14829 22967 14887 22973
rect 14829 22964 14841 22967
rect 14792 22936 14841 22964
rect 14792 22924 14798 22936
rect 14829 22933 14841 22936
rect 14875 22933 14887 22967
rect 14829 22927 14887 22933
rect 15470 22924 15476 22976
rect 15528 22964 15534 22976
rect 15565 22967 15623 22973
rect 15565 22964 15577 22967
rect 15528 22936 15577 22964
rect 15528 22924 15534 22936
rect 15565 22933 15577 22936
rect 15611 22933 15623 22967
rect 15565 22927 15623 22933
rect 21082 22924 21088 22976
rect 21140 22964 21146 22976
rect 22572 22964 22600 23072
rect 23937 23069 23949 23072
rect 23983 23100 23995 23103
rect 24121 23103 24179 23109
rect 24121 23100 24133 23103
rect 23983 23072 24133 23100
rect 23983 23069 23995 23072
rect 23937 23063 23995 23069
rect 24121 23069 24133 23072
rect 24167 23069 24179 23103
rect 26513 23103 26571 23109
rect 26513 23100 26525 23103
rect 24121 23063 24179 23069
rect 26252 23072 26525 23100
rect 21140 22936 22600 22964
rect 21140 22924 21146 22936
rect 22646 22924 22652 22976
rect 22704 22964 22710 22976
rect 26252 22973 26280 23072
rect 26513 23069 26525 23072
rect 26559 23069 26571 23103
rect 26513 23063 26571 23069
rect 26237 22967 26295 22973
rect 26237 22964 26249 22967
rect 22704 22936 26249 22964
rect 22704 22924 22710 22936
rect 26237 22933 26249 22936
rect 26283 22933 26295 22967
rect 26237 22927 26295 22933
rect 26786 22924 26792 22976
rect 26844 22964 26850 22976
rect 27709 22967 27767 22973
rect 27709 22964 27721 22967
rect 26844 22936 27721 22964
rect 26844 22924 26850 22936
rect 27709 22933 27721 22936
rect 27755 22933 27767 22967
rect 27709 22927 27767 22933
rect 1104 22874 29256 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 29256 22874
rect 1104 22800 29256 22822
rect 4062 22720 4068 22772
rect 4120 22760 4126 22772
rect 25314 22760 25320 22772
rect 4120 22732 25320 22760
rect 4120 22720 4126 22732
rect 25314 22720 25320 22732
rect 25372 22720 25378 22772
rect 27614 22720 27620 22772
rect 27672 22760 27678 22772
rect 28077 22763 28135 22769
rect 28077 22760 28089 22763
rect 27672 22732 28089 22760
rect 27672 22720 27678 22732
rect 28077 22729 28089 22732
rect 28123 22760 28135 22763
rect 29086 22760 29092 22772
rect 28123 22732 29092 22760
rect 28123 22729 28135 22732
rect 28077 22723 28135 22729
rect 29086 22720 29092 22732
rect 29144 22720 29150 22772
rect 4617 22695 4675 22701
rect 4617 22661 4629 22695
rect 4663 22692 4675 22695
rect 4798 22692 4804 22704
rect 4663 22664 4804 22692
rect 4663 22661 4675 22664
rect 4617 22655 4675 22661
rect 4798 22652 4804 22664
rect 4856 22692 4862 22704
rect 5442 22692 5448 22704
rect 4856 22664 5448 22692
rect 4856 22652 4862 22664
rect 5442 22652 5448 22664
rect 5500 22652 5506 22704
rect 9582 22652 9588 22704
rect 9640 22692 9646 22704
rect 10045 22695 10103 22701
rect 10045 22692 10057 22695
rect 9640 22664 10057 22692
rect 9640 22652 9646 22664
rect 10045 22661 10057 22664
rect 10091 22661 10103 22695
rect 14826 22692 14832 22704
rect 14787 22664 14832 22692
rect 10045 22655 10103 22661
rect 14826 22652 14832 22664
rect 14884 22652 14890 22704
rect 21174 22692 21180 22704
rect 21135 22664 21180 22692
rect 21174 22652 21180 22664
rect 21232 22652 21238 22704
rect 2869 22627 2927 22633
rect 2869 22593 2881 22627
rect 2915 22624 2927 22627
rect 4433 22627 4491 22633
rect 4433 22624 4445 22627
rect 2915 22596 4445 22624
rect 2915 22593 2927 22596
rect 2869 22587 2927 22593
rect 4433 22593 4445 22596
rect 4479 22624 4491 22627
rect 5166 22624 5172 22636
rect 4479 22596 5172 22624
rect 4479 22593 4491 22596
rect 4433 22587 4491 22593
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 5350 22584 5356 22636
rect 5408 22624 5414 22636
rect 5718 22624 5724 22636
rect 5408 22596 5724 22624
rect 5408 22584 5414 22596
rect 5718 22584 5724 22596
rect 5776 22584 5782 22636
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22624 8355 22627
rect 9600 22624 9628 22652
rect 8343 22596 9628 22624
rect 13633 22627 13691 22633
rect 8343 22593 8355 22596
rect 8297 22587 8355 22593
rect 13633 22593 13645 22627
rect 13679 22624 13691 22627
rect 13679 22596 14044 22624
rect 13679 22593 13691 22596
rect 13633 22587 13691 22593
rect 14016 22568 14044 22596
rect 17972 22596 20484 22624
rect 2590 22556 2596 22568
rect 2551 22528 2596 22556
rect 2590 22516 2596 22528
rect 2648 22516 2654 22568
rect 8570 22556 8576 22568
rect 8531 22528 8576 22556
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 13722 22516 13728 22568
rect 13780 22556 13786 22568
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 13780 22528 13921 22556
rect 13780 22516 13786 22528
rect 13909 22525 13921 22528
rect 13955 22525 13967 22559
rect 13909 22519 13967 22525
rect 9950 22488 9956 22500
rect 9911 22460 9956 22488
rect 9950 22448 9956 22460
rect 10008 22448 10014 22500
rect 13924 22488 13952 22519
rect 13998 22516 14004 22568
rect 14056 22556 14062 22568
rect 14366 22556 14372 22568
rect 14056 22528 14372 22556
rect 14056 22516 14062 22528
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 14461 22559 14519 22565
rect 14461 22525 14473 22559
rect 14507 22525 14519 22559
rect 14461 22519 14519 22525
rect 14645 22559 14703 22565
rect 14645 22525 14657 22559
rect 14691 22556 14703 22559
rect 15746 22556 15752 22568
rect 14691 22528 15752 22556
rect 14691 22525 14703 22528
rect 14645 22519 14703 22525
rect 14476 22488 14504 22519
rect 15746 22516 15752 22528
rect 15804 22516 15810 22568
rect 17972 22488 18000 22596
rect 20272 22565 20300 22596
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22556 18107 22559
rect 20257 22559 20315 22565
rect 18095 22528 18460 22556
rect 18095 22525 18107 22528
rect 18049 22519 18107 22525
rect 13924 22460 18000 22488
rect 2866 22380 2872 22432
rect 2924 22420 2930 22432
rect 3973 22423 4031 22429
rect 3973 22420 3985 22423
rect 2924 22392 3985 22420
rect 2924 22380 2930 22392
rect 3973 22389 3985 22392
rect 4019 22389 4031 22423
rect 3973 22383 4031 22389
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 18432 22429 18460 22528
rect 20257 22525 20269 22559
rect 20303 22525 20315 22559
rect 20257 22519 20315 22525
rect 20349 22559 20407 22565
rect 20349 22525 20361 22559
rect 20395 22525 20407 22559
rect 20456 22556 20484 22596
rect 25222 22584 25228 22636
rect 25280 22624 25286 22636
rect 26421 22627 26479 22633
rect 26421 22624 26433 22627
rect 25280 22596 26433 22624
rect 25280 22584 25286 22596
rect 26421 22593 26433 22596
rect 26467 22624 26479 22627
rect 26513 22627 26571 22633
rect 26513 22624 26525 22627
rect 26467 22596 26525 22624
rect 26467 22593 26479 22596
rect 26421 22587 26479 22593
rect 26513 22593 26525 22596
rect 26559 22593 26571 22627
rect 26786 22624 26792 22636
rect 26747 22596 26792 22624
rect 26513 22587 26571 22593
rect 26786 22584 26792 22596
rect 26844 22584 26850 22636
rect 20806 22556 20812 22568
rect 20456 22528 20812 22556
rect 20349 22519 20407 22525
rect 18690 22448 18696 22500
rect 18748 22488 18754 22500
rect 19981 22491 20039 22497
rect 19981 22488 19993 22491
rect 18748 22460 19993 22488
rect 18748 22448 18754 22460
rect 19981 22457 19993 22460
rect 20027 22488 20039 22491
rect 20364 22488 20392 22519
rect 20806 22516 20812 22528
rect 20864 22516 20870 22568
rect 20993 22559 21051 22565
rect 20993 22525 21005 22559
rect 21039 22556 21051 22559
rect 21634 22556 21640 22568
rect 21039 22528 21640 22556
rect 21039 22525 21051 22528
rect 20993 22519 21051 22525
rect 21634 22516 21640 22528
rect 21692 22556 21698 22568
rect 21910 22556 21916 22568
rect 21692 22528 21916 22556
rect 21692 22516 21698 22528
rect 21910 22516 21916 22528
rect 21968 22516 21974 22568
rect 21082 22488 21088 22500
rect 20027 22460 21088 22488
rect 20027 22457 20039 22460
rect 19981 22451 20039 22457
rect 21082 22448 21088 22460
rect 21140 22448 21146 22500
rect 18141 22423 18199 22429
rect 18141 22420 18153 22423
rect 16724 22392 18153 22420
rect 16724 22380 16730 22392
rect 18141 22389 18153 22392
rect 18187 22389 18199 22423
rect 18141 22383 18199 22389
rect 18417 22423 18475 22429
rect 18417 22389 18429 22423
rect 18463 22420 18475 22423
rect 18598 22420 18604 22432
rect 18463 22392 18604 22420
rect 18463 22389 18475 22392
rect 18417 22383 18475 22389
rect 18598 22380 18604 22392
rect 18656 22380 18662 22432
rect 1104 22330 29256 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 29256 22330
rect 1104 22256 29256 22278
rect 8570 22216 8576 22228
rect 8531 22188 8576 22216
rect 8570 22176 8576 22188
rect 8628 22176 8634 22228
rect 18598 22148 18604 22160
rect 18559 22120 18604 22148
rect 18598 22108 18604 22120
rect 18656 22108 18662 22160
rect 22281 22151 22339 22157
rect 22281 22148 22293 22151
rect 22112 22120 22293 22148
rect 7561 22083 7619 22089
rect 7561 22049 7573 22083
rect 7607 22080 7619 22083
rect 8110 22080 8116 22092
rect 7607 22052 8116 22080
rect 7607 22049 7619 22052
rect 7561 22043 7619 22049
rect 8110 22040 8116 22052
rect 8168 22040 8174 22092
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22080 8355 22083
rect 9677 22083 9735 22089
rect 8343 22052 9628 22080
rect 8343 22049 8355 22052
rect 8297 22043 8355 22049
rect 7282 21972 7288 22024
rect 7340 22012 7346 22024
rect 7377 22015 7435 22021
rect 7377 22012 7389 22015
rect 7340 21984 7389 22012
rect 7340 21972 7346 21984
rect 7377 21981 7389 21984
rect 7423 21981 7435 22015
rect 9600 22012 9628 22052
rect 9677 22049 9689 22083
rect 9723 22080 9735 22083
rect 10045 22083 10103 22089
rect 10045 22080 10057 22083
rect 9723 22052 10057 22080
rect 9723 22049 9735 22052
rect 9677 22043 9735 22049
rect 10045 22049 10057 22052
rect 10091 22080 10103 22083
rect 10226 22080 10232 22092
rect 10091 22052 10232 22080
rect 10091 22049 10103 22052
rect 10045 22043 10103 22049
rect 10226 22040 10232 22052
rect 10284 22040 10290 22092
rect 11330 22040 11336 22092
rect 11388 22080 11394 22092
rect 11974 22080 11980 22092
rect 11388 22052 11980 22080
rect 11388 22040 11394 22052
rect 11974 22040 11980 22052
rect 12032 22080 12038 22092
rect 12161 22083 12219 22089
rect 12161 22080 12173 22083
rect 12032 22052 12173 22080
rect 12032 22040 12038 22052
rect 12161 22049 12173 22052
rect 12207 22049 12219 22083
rect 16758 22080 16764 22092
rect 16719 22052 16764 22080
rect 12161 22043 12219 22049
rect 16758 22040 16764 22052
rect 16816 22080 16822 22092
rect 22112 22089 22140 22120
rect 22281 22117 22293 22120
rect 22327 22148 22339 22151
rect 22370 22148 22376 22160
rect 22327 22120 22376 22148
rect 22327 22117 22339 22120
rect 22281 22111 22339 22117
rect 22370 22108 22376 22120
rect 22428 22108 22434 22160
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 16816 22052 16957 22080
rect 16816 22040 16822 22052
rect 16945 22049 16957 22052
rect 16991 22049 17003 22083
rect 20441 22083 20499 22089
rect 20441 22080 20453 22083
rect 16945 22043 17003 22049
rect 17052 22052 20453 22080
rect 9766 22012 9772 22024
rect 9600 21984 9772 22012
rect 7377 21975 7435 21981
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 17052 22012 17080 22052
rect 20441 22049 20453 22052
rect 20487 22049 20499 22083
rect 21545 22083 21603 22089
rect 21545 22080 21557 22083
rect 20441 22043 20499 22049
rect 21100 22052 21557 22080
rect 17218 22012 17224 22024
rect 15151 21984 17080 22012
rect 17179 21984 17224 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 17218 21972 17224 21984
rect 17276 21972 17282 22024
rect 4062 21904 4068 21956
rect 4120 21944 4126 21956
rect 20456 21944 20484 22043
rect 21100 22024 21128 22052
rect 21545 22049 21557 22052
rect 21591 22049 21603 22083
rect 21545 22043 21603 22049
rect 21913 22083 21971 22089
rect 21913 22049 21925 22083
rect 21959 22049 21971 22083
rect 21913 22043 21971 22049
rect 22097 22083 22155 22089
rect 22097 22049 22109 22083
rect 22143 22049 22155 22083
rect 27614 22080 27620 22092
rect 27575 22052 27620 22080
rect 22097 22043 22155 22049
rect 20714 21972 20720 22024
rect 20772 22012 20778 22024
rect 20901 22015 20959 22021
rect 20901 22012 20913 22015
rect 20772 21984 20913 22012
rect 20772 21972 20778 21984
rect 20901 21981 20913 21984
rect 20947 21981 20959 22015
rect 20901 21975 20959 21981
rect 21082 21972 21088 22024
rect 21140 21972 21146 22024
rect 21634 22012 21640 22024
rect 21595 21984 21640 22012
rect 21634 21972 21640 21984
rect 21692 21972 21698 22024
rect 21928 22012 21956 22043
rect 27614 22040 27620 22052
rect 27672 22040 27678 22092
rect 27706 22040 27712 22092
rect 27764 22080 27770 22092
rect 27764 22052 27809 22080
rect 27764 22040 27770 22052
rect 59354 22040 59360 22092
rect 59412 22080 59418 22092
rect 59538 22080 59544 22092
rect 59412 22052 59544 22080
rect 59412 22040 59418 22052
rect 59538 22040 59544 22052
rect 59596 22040 59602 22092
rect 21836 21984 21956 22012
rect 21174 21944 21180 21956
rect 4120 21916 16160 21944
rect 20456 21916 21180 21944
rect 4120 21904 4126 21916
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 7193 21879 7251 21885
rect 7193 21876 7205 21879
rect 6972 21848 7205 21876
rect 6972 21836 6978 21848
rect 7193 21845 7205 21848
rect 7239 21876 7251 21879
rect 7282 21876 7288 21888
rect 7239 21848 7288 21876
rect 7239 21845 7251 21848
rect 7193 21839 7251 21845
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 9030 21836 9036 21888
rect 9088 21876 9094 21888
rect 9769 21879 9827 21885
rect 9769 21876 9781 21879
rect 9088 21848 9781 21876
rect 9088 21836 9094 21848
rect 9769 21845 9781 21848
rect 9815 21845 9827 21879
rect 11974 21876 11980 21888
rect 11935 21848 11980 21876
rect 9769 21839 9827 21845
rect 11974 21836 11980 21848
rect 12032 21836 12038 21888
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 12345 21879 12403 21885
rect 12345 21876 12357 21879
rect 12216 21848 12357 21876
rect 12216 21836 12222 21848
rect 12345 21845 12357 21848
rect 12391 21876 12403 21879
rect 15105 21879 15163 21885
rect 15105 21876 15117 21879
rect 12391 21848 15117 21876
rect 12391 21845 12403 21848
rect 12345 21839 12403 21845
rect 15105 21845 15117 21848
rect 15151 21845 15163 21879
rect 16132 21876 16160 21916
rect 21174 21904 21180 21916
rect 21232 21944 21238 21956
rect 21836 21944 21864 21984
rect 21232 21916 21864 21944
rect 21232 21904 21238 21916
rect 19794 21876 19800 21888
rect 16132 21848 19800 21876
rect 15105 21839 15163 21845
rect 19794 21836 19800 21848
rect 19852 21836 19858 21888
rect 20717 21879 20775 21885
rect 20717 21845 20729 21879
rect 20763 21876 20775 21879
rect 21082 21876 21088 21888
rect 20763 21848 21088 21876
rect 20763 21845 20775 21848
rect 20717 21839 20775 21845
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 1104 21786 29256 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 29256 21786
rect 1104 21712 29256 21734
rect 3602 21632 3608 21684
rect 3660 21672 3666 21684
rect 3973 21675 4031 21681
rect 3973 21672 3985 21675
rect 3660 21644 3985 21672
rect 3660 21632 3666 21644
rect 3973 21641 3985 21644
rect 4019 21641 4031 21675
rect 3973 21635 4031 21641
rect 4617 21675 4675 21681
rect 4617 21641 4629 21675
rect 4663 21672 4675 21675
rect 4798 21672 4804 21684
rect 4663 21644 4804 21672
rect 4663 21641 4675 21644
rect 4617 21635 4675 21641
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 8772 21644 9628 21672
rect 8772 21604 8800 21644
rect 4356 21576 8800 21604
rect 2590 21468 2596 21480
rect 2551 21440 2596 21468
rect 2590 21428 2596 21440
rect 2648 21428 2654 21480
rect 4356 21477 4384 21576
rect 8846 21564 8852 21616
rect 8904 21604 8910 21616
rect 9033 21607 9091 21613
rect 9033 21604 9045 21607
rect 8904 21576 9045 21604
rect 8904 21564 8910 21576
rect 9033 21573 9045 21576
rect 9079 21573 9091 21607
rect 9600 21604 9628 21644
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 10321 21675 10379 21681
rect 10321 21672 10333 21675
rect 9732 21644 10333 21672
rect 9732 21632 9738 21644
rect 10321 21641 10333 21644
rect 10367 21641 10379 21675
rect 10321 21635 10379 21641
rect 12713 21675 12771 21681
rect 12713 21641 12725 21675
rect 12759 21672 12771 21675
rect 14090 21672 14096 21684
rect 12759 21644 14096 21672
rect 12759 21641 12771 21644
rect 12713 21635 12771 21641
rect 11238 21604 11244 21616
rect 9600 21576 11244 21604
rect 9033 21567 9091 21573
rect 11238 21564 11244 21576
rect 11296 21564 11302 21616
rect 8202 21536 8208 21548
rect 7944 21508 8208 21536
rect 7944 21477 7972 21508
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 11882 21536 11888 21548
rect 11164 21508 11888 21536
rect 2869 21471 2927 21477
rect 2869 21437 2881 21471
rect 2915 21468 2927 21471
rect 4341 21471 4399 21477
rect 4341 21468 4353 21471
rect 2915 21440 4353 21468
rect 2915 21437 2927 21440
rect 2869 21431 2927 21437
rect 4341 21437 4353 21440
rect 4387 21437 4399 21471
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 4341 21431 4399 21437
rect 7760 21440 7941 21468
rect 7098 21292 7104 21344
rect 7156 21332 7162 21344
rect 7760 21341 7788 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 8110 21468 8116 21480
rect 8023 21440 8116 21468
rect 7929 21431 7987 21437
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21468 8907 21471
rect 9030 21468 9036 21480
rect 8895 21440 9036 21468
rect 8895 21437 8907 21440
rect 8849 21431 8907 21437
rect 8128 21400 8156 21428
rect 8680 21400 8708 21431
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 10137 21471 10195 21477
rect 10137 21437 10149 21471
rect 10183 21468 10195 21471
rect 10870 21468 10876 21480
rect 10183 21440 10876 21468
rect 10183 21437 10195 21440
rect 10137 21431 10195 21437
rect 10870 21428 10876 21440
rect 10928 21428 10934 21480
rect 11164 21468 11192 21508
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 12820 21545 12848 21644
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 16945 21675 17003 21681
rect 16945 21641 16957 21675
rect 16991 21672 17003 21675
rect 17218 21672 17224 21684
rect 16991 21644 17224 21672
rect 16991 21641 17003 21644
rect 16945 21635 17003 21641
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 19334 21672 19340 21684
rect 19295 21644 19340 21672
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 22646 21604 22652 21616
rect 21284 21576 22652 21604
rect 21284 21548 21312 21576
rect 22646 21564 22652 21576
rect 22704 21564 22710 21616
rect 12805 21539 12863 21545
rect 12805 21505 12817 21539
rect 12851 21505 12863 21539
rect 21266 21536 21272 21548
rect 21227 21508 21272 21536
rect 12805 21499 12863 21505
rect 21266 21496 21272 21508
rect 21324 21496 21330 21548
rect 11229 21471 11287 21477
rect 11229 21468 11241 21471
rect 11164 21440 11241 21468
rect 11229 21437 11241 21440
rect 11275 21437 11287 21471
rect 13078 21468 13084 21480
rect 13039 21440 13084 21468
rect 11229 21431 11287 21437
rect 13078 21428 13084 21440
rect 13136 21428 13142 21480
rect 13170 21428 13176 21480
rect 13228 21468 13234 21480
rect 15565 21471 15623 21477
rect 15565 21468 15577 21471
rect 13228 21440 15577 21468
rect 13228 21428 13234 21440
rect 15565 21437 15577 21440
rect 15611 21468 15623 21471
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 15611 21440 15761 21468
rect 15611 21437 15623 21440
rect 15565 21431 15623 21437
rect 15749 21437 15761 21440
rect 15795 21437 15807 21471
rect 15749 21431 15807 21437
rect 15933 21471 15991 21477
rect 15933 21437 15945 21471
rect 15979 21468 15991 21471
rect 16485 21471 16543 21477
rect 16485 21468 16497 21471
rect 15979 21440 16497 21468
rect 15979 21437 15991 21440
rect 15933 21431 15991 21437
rect 16485 21437 16497 21440
rect 16531 21437 16543 21471
rect 16666 21468 16672 21480
rect 16627 21440 16672 21468
rect 16485 21431 16543 21437
rect 14458 21400 14464 21412
rect 8128 21372 11468 21400
rect 14419 21372 14464 21400
rect 11440 21341 11468 21372
rect 14458 21360 14464 21372
rect 14516 21360 14522 21412
rect 16500 21400 16528 21431
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 19245 21471 19303 21477
rect 19245 21468 19257 21471
rect 18840 21440 19257 21468
rect 18840 21428 18846 21440
rect 19245 21437 19257 21440
rect 19291 21437 19303 21471
rect 19245 21431 19303 21437
rect 20806 21428 20812 21480
rect 20864 21468 20870 21480
rect 21453 21471 21511 21477
rect 21453 21468 21465 21471
rect 20864 21440 21465 21468
rect 20864 21428 20870 21440
rect 21453 21437 21465 21440
rect 21499 21437 21511 21471
rect 22002 21468 22008 21480
rect 21963 21440 22008 21468
rect 21453 21431 21511 21437
rect 22002 21428 22008 21440
rect 22060 21428 22066 21480
rect 22094 21428 22100 21480
rect 22152 21468 22158 21480
rect 22189 21471 22247 21477
rect 22189 21468 22201 21471
rect 22152 21440 22201 21468
rect 22152 21428 22158 21440
rect 22189 21437 22201 21440
rect 22235 21468 22247 21471
rect 23661 21471 23719 21477
rect 22235 21440 22784 21468
rect 22235 21437 22247 21440
rect 22189 21431 22247 21437
rect 16758 21400 16764 21412
rect 16500 21372 16764 21400
rect 16758 21360 16764 21372
rect 16816 21360 16822 21412
rect 22557 21403 22615 21409
rect 22557 21369 22569 21403
rect 22603 21400 22615 21403
rect 22646 21400 22652 21412
rect 22603 21372 22652 21400
rect 22603 21369 22615 21372
rect 22557 21363 22615 21369
rect 22646 21360 22652 21372
rect 22704 21360 22710 21412
rect 22756 21400 22784 21440
rect 23661 21437 23673 21471
rect 23707 21468 23719 21471
rect 23707 21440 23980 21468
rect 23707 21437 23719 21440
rect 23661 21431 23719 21437
rect 23753 21403 23811 21409
rect 23753 21400 23765 21403
rect 22756 21372 23765 21400
rect 23753 21369 23765 21372
rect 23799 21369 23811 21403
rect 23753 21363 23811 21369
rect 23952 21344 23980 21440
rect 7745 21335 7803 21341
rect 7745 21332 7757 21335
rect 7156 21304 7757 21332
rect 7156 21292 7162 21304
rect 7745 21301 7757 21304
rect 7791 21301 7803 21335
rect 7745 21295 7803 21301
rect 11425 21335 11483 21341
rect 11425 21301 11437 21335
rect 11471 21332 11483 21335
rect 12434 21332 12440 21344
rect 11471 21304 12440 21332
rect 11471 21301 11483 21304
rect 11425 21295 11483 21301
rect 12434 21292 12440 21304
rect 12492 21292 12498 21344
rect 21177 21335 21235 21341
rect 21177 21301 21189 21335
rect 21223 21332 21235 21335
rect 21266 21332 21272 21344
rect 21223 21304 21272 21332
rect 21223 21301 21235 21304
rect 21177 21295 21235 21301
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 23934 21332 23940 21344
rect 23895 21304 23940 21332
rect 23934 21292 23940 21304
rect 23992 21292 23998 21344
rect 1104 21242 29256 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 29256 21242
rect 1104 21168 29256 21190
rect 9766 21128 9772 21140
rect 9727 21100 9772 21128
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 9950 21128 9956 21140
rect 9911 21100 9956 21128
rect 9950 21088 9956 21100
rect 10008 21088 10014 21140
rect 11606 21128 11612 21140
rect 11567 21100 11612 21128
rect 11606 21088 11612 21100
rect 11664 21088 11670 21140
rect 14277 21131 14335 21137
rect 14277 21097 14289 21131
rect 14323 21128 14335 21131
rect 14458 21128 14464 21140
rect 14323 21100 14464 21128
rect 14323 21097 14335 21100
rect 14277 21091 14335 21097
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 26142 21128 26148 21140
rect 22480 21100 26148 21128
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9968 20992 9996 21088
rect 12989 21063 13047 21069
rect 12989 21029 13001 21063
rect 13035 21060 13047 21063
rect 13078 21060 13084 21072
rect 13035 21032 13084 21060
rect 13035 21029 13047 21032
rect 12989 21023 13047 21029
rect 13078 21020 13084 21032
rect 13136 21020 13142 21072
rect 22480 21060 22508 21100
rect 26142 21088 26148 21100
rect 26200 21088 26206 21140
rect 27893 21131 27951 21137
rect 27893 21097 27905 21131
rect 27939 21128 27951 21131
rect 27982 21128 27988 21140
rect 27939 21100 27988 21128
rect 27939 21097 27951 21100
rect 27893 21091 27951 21097
rect 27982 21088 27988 21100
rect 28040 21088 28046 21140
rect 14568 21032 22508 21060
rect 10686 20992 10692 21004
rect 9723 20964 9996 20992
rect 10647 20964 10692 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 10686 20952 10692 20964
rect 10744 20952 10750 21004
rect 11606 20952 11612 21004
rect 11664 20992 11670 21004
rect 11701 20995 11759 21001
rect 11701 20992 11713 20995
rect 11664 20964 11713 20992
rect 11664 20952 11670 20964
rect 11701 20961 11713 20964
rect 11747 20961 11759 20995
rect 11882 20992 11888 21004
rect 11843 20964 11888 20992
rect 11701 20955 11759 20961
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 12621 20995 12679 21001
rect 12492 20964 12537 20992
rect 12492 20952 12498 20964
rect 12621 20961 12633 20995
rect 12667 20992 12679 20995
rect 12894 20992 12900 21004
rect 12667 20964 12900 20992
rect 12667 20961 12679 20964
rect 12621 20955 12679 20961
rect 12894 20952 12900 20964
rect 12952 20952 12958 21004
rect 13909 20995 13967 21001
rect 13909 20961 13921 20995
rect 13955 20992 13967 20995
rect 14458 20992 14464 21004
rect 13955 20964 14464 20992
rect 13955 20961 13967 20964
rect 13909 20955 13967 20961
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 4062 20884 4068 20936
rect 4120 20924 4126 20936
rect 12912 20924 12940 20952
rect 14001 20927 14059 20933
rect 14001 20924 14013 20927
rect 4120 20896 12112 20924
rect 12912 20896 14013 20924
rect 4120 20884 4126 20896
rect 11054 20816 11060 20868
rect 11112 20856 11118 20868
rect 12084 20856 12112 20896
rect 14001 20893 14013 20896
rect 14047 20893 14059 20927
rect 14001 20887 14059 20893
rect 14568 20856 14596 21032
rect 15010 20952 15016 21004
rect 15068 20992 15074 21004
rect 15749 20995 15807 21001
rect 15749 20992 15761 20995
rect 15068 20964 15761 20992
rect 15068 20952 15074 20964
rect 15749 20961 15761 20964
rect 15795 20961 15807 20995
rect 15749 20955 15807 20961
rect 15933 20995 15991 21001
rect 15933 20961 15945 20995
rect 15979 20961 15991 20995
rect 16301 20995 16359 21001
rect 16301 20992 16313 20995
rect 15933 20955 15991 20961
rect 16224 20964 16313 20992
rect 15286 20924 15292 20936
rect 15247 20896 15292 20924
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 15013 20859 15071 20865
rect 15013 20856 15025 20859
rect 11112 20828 11652 20856
rect 12084 20828 14596 20856
rect 14660 20828 15025 20856
rect 11112 20816 11118 20828
rect 10781 20791 10839 20797
rect 10781 20757 10793 20791
rect 10827 20788 10839 20791
rect 10962 20788 10968 20800
rect 10827 20760 10968 20788
rect 10827 20757 10839 20760
rect 10781 20751 10839 20757
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 11624 20788 11652 20828
rect 11974 20788 11980 20800
rect 11624 20760 11980 20788
rect 11974 20748 11980 20760
rect 12032 20788 12038 20800
rect 14660 20788 14688 20828
rect 15013 20825 15025 20828
rect 15059 20856 15071 20859
rect 15194 20856 15200 20868
rect 15059 20828 15200 20856
rect 15059 20825 15071 20828
rect 15013 20819 15071 20825
rect 15194 20816 15200 20828
rect 15252 20856 15258 20868
rect 15948 20856 15976 20955
rect 15252 20828 15976 20856
rect 16224 20924 16252 20964
rect 16301 20961 16313 20964
rect 16347 20961 16359 20995
rect 16301 20955 16359 20961
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20992 16543 20995
rect 16666 20992 16672 21004
rect 16531 20964 16672 20992
rect 16531 20961 16543 20964
rect 16485 20955 16543 20961
rect 16666 20952 16672 20964
rect 16724 20952 16730 21004
rect 16758 20952 16764 21004
rect 16816 20992 16822 21004
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 16816 20964 19257 20992
rect 16816 20952 16822 20964
rect 19245 20961 19257 20964
rect 19291 20961 19303 20995
rect 22646 20992 22652 21004
rect 22607 20964 22652 20992
rect 19245 20955 19303 20961
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 21082 20924 21088 20936
rect 16224 20896 21088 20924
rect 15252 20816 15258 20828
rect 12032 20760 14688 20788
rect 12032 20748 12038 20760
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 14829 20791 14887 20797
rect 14829 20788 14841 20791
rect 14792 20760 14841 20788
rect 14792 20748 14798 20760
rect 14829 20757 14841 20760
rect 14875 20788 14887 20791
rect 16224 20788 16252 20896
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 22373 20927 22431 20933
rect 22373 20893 22385 20927
rect 22419 20893 22431 20927
rect 26513 20927 26571 20933
rect 26513 20924 26525 20927
rect 22373 20887 22431 20893
rect 26252 20896 26525 20924
rect 14875 20760 16252 20788
rect 19429 20791 19487 20797
rect 14875 20757 14887 20760
rect 14829 20751 14887 20757
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 22002 20788 22008 20800
rect 19475 20760 22008 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 22002 20748 22008 20760
rect 22060 20748 22066 20800
rect 22388 20788 22416 20887
rect 26252 20868 26280 20896
rect 26513 20893 26525 20896
rect 26559 20893 26571 20927
rect 26786 20924 26792 20936
rect 26747 20896 26792 20924
rect 26513 20887 26571 20893
rect 26786 20884 26792 20896
rect 26844 20884 26850 20936
rect 24121 20859 24179 20865
rect 24121 20856 24133 20859
rect 23768 20828 24133 20856
rect 23768 20788 23796 20828
rect 24121 20825 24133 20828
rect 24167 20856 24179 20859
rect 26234 20856 26240 20868
rect 24167 20828 26240 20856
rect 24167 20825 24179 20828
rect 24121 20819 24179 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 23934 20788 23940 20800
rect 22388 20760 23796 20788
rect 23895 20760 23940 20788
rect 23934 20748 23940 20760
rect 23992 20748 23998 20800
rect 1104 20698 29256 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 29256 20698
rect 1104 20624 29256 20646
rect 2590 20584 2596 20596
rect 2503 20556 2596 20584
rect 2590 20544 2596 20556
rect 2648 20584 2654 20596
rect 4433 20587 4491 20593
rect 4433 20584 4445 20587
rect 2648 20556 4445 20584
rect 2648 20544 2654 20556
rect 4433 20553 4445 20556
rect 4479 20584 4491 20587
rect 4798 20584 4804 20596
rect 4479 20556 4804 20584
rect 4479 20553 4491 20556
rect 4433 20547 4491 20553
rect 4798 20544 4804 20556
rect 4856 20544 4862 20596
rect 11882 20544 11888 20596
rect 11940 20584 11946 20596
rect 12621 20587 12679 20593
rect 12621 20584 12633 20587
rect 11940 20556 12633 20584
rect 11940 20544 11946 20556
rect 12621 20553 12633 20556
rect 12667 20584 12679 20587
rect 16758 20584 16764 20596
rect 12667 20556 16764 20584
rect 12667 20553 12679 20556
rect 12621 20547 12679 20553
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 20809 20587 20867 20593
rect 20809 20584 20821 20587
rect 20680 20556 20821 20584
rect 20680 20544 20686 20556
rect 20809 20553 20821 20556
rect 20855 20553 20867 20587
rect 21174 20584 21180 20596
rect 21135 20556 21180 20584
rect 20809 20547 20867 20553
rect 21174 20544 21180 20556
rect 21232 20544 21238 20596
rect 22738 20544 22744 20596
rect 22796 20584 22802 20596
rect 22833 20587 22891 20593
rect 22833 20584 22845 20587
rect 22796 20556 22845 20584
rect 22796 20544 22802 20556
rect 22833 20553 22845 20556
rect 22879 20553 22891 20587
rect 22833 20547 22891 20553
rect 25777 20587 25835 20593
rect 25777 20553 25789 20587
rect 25823 20584 25835 20587
rect 26234 20584 26240 20596
rect 25823 20556 26240 20584
rect 25823 20553 25835 20556
rect 25777 20547 25835 20553
rect 26234 20544 26240 20556
rect 26292 20544 26298 20596
rect 27433 20587 27491 20593
rect 27433 20553 27445 20587
rect 27479 20584 27491 20587
rect 27522 20584 27528 20596
rect 27479 20556 27528 20584
rect 27479 20553 27491 20556
rect 27433 20547 27491 20553
rect 27522 20544 27528 20556
rect 27580 20584 27586 20596
rect 27890 20584 27896 20596
rect 27580 20556 27896 20584
rect 27580 20544 27586 20556
rect 27890 20544 27896 20556
rect 27948 20544 27954 20596
rect 2608 20457 2636 20544
rect 18782 20476 18788 20528
rect 18840 20516 18846 20528
rect 18840 20488 20484 20516
rect 18840 20476 18846 20488
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20417 2651 20451
rect 2593 20411 2651 20417
rect 18892 20420 19932 20448
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20380 2927 20383
rect 3142 20380 3148 20392
rect 2915 20352 3148 20380
rect 2915 20349 2927 20352
rect 2869 20343 2927 20349
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 10686 20380 10692 20392
rect 10647 20352 10692 20380
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 10870 20340 10876 20392
rect 10928 20380 10934 20392
rect 12437 20383 12495 20389
rect 10928 20352 10973 20380
rect 10928 20340 10934 20352
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12710 20380 12716 20392
rect 12483 20352 12716 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12710 20340 12716 20352
rect 12768 20340 12774 20392
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20380 14795 20383
rect 15286 20380 15292 20392
rect 14783 20352 15292 20380
rect 14783 20349 14795 20352
rect 14737 20343 14795 20349
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 11241 20315 11299 20321
rect 11241 20281 11253 20315
rect 11287 20312 11299 20315
rect 16942 20312 16948 20324
rect 11287 20284 16948 20312
rect 11287 20281 11299 20284
rect 11241 20275 11299 20281
rect 16942 20272 16948 20284
rect 17000 20312 17006 20324
rect 18782 20312 18788 20324
rect 17000 20284 18788 20312
rect 17000 20272 17006 20284
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 3326 20204 3332 20256
rect 3384 20244 3390 20256
rect 3973 20247 4031 20253
rect 3973 20244 3985 20247
rect 3384 20216 3985 20244
rect 3384 20204 3390 20216
rect 3973 20213 3985 20216
rect 4019 20213 4031 20247
rect 14826 20244 14832 20256
rect 14787 20216 14832 20244
rect 3973 20207 4031 20213
rect 14826 20204 14832 20216
rect 14884 20204 14890 20256
rect 18138 20204 18144 20256
rect 18196 20244 18202 20256
rect 18892 20253 18920 20420
rect 19904 20389 19932 20420
rect 19705 20383 19763 20389
rect 19705 20349 19717 20383
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 19889 20383 19947 20389
rect 19889 20349 19901 20383
rect 19935 20349 19947 20383
rect 20162 20380 20168 20392
rect 20123 20352 20168 20380
rect 19889 20343 19947 20349
rect 19245 20315 19303 20321
rect 19245 20281 19257 20315
rect 19291 20312 19303 20315
rect 19426 20312 19432 20324
rect 19291 20284 19432 20312
rect 19291 20281 19303 20284
rect 19245 20275 19303 20281
rect 19426 20272 19432 20284
rect 19484 20272 19490 20324
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18196 20216 18889 20244
rect 18196 20204 18202 20216
rect 18877 20213 18889 20216
rect 18923 20213 18935 20247
rect 19150 20244 19156 20256
rect 19111 20216 19156 20244
rect 18877 20207 18935 20213
rect 19150 20204 19156 20216
rect 19208 20244 19214 20256
rect 19720 20244 19748 20343
rect 20162 20340 20168 20352
rect 20220 20340 20226 20392
rect 20456 20380 20484 20488
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20640 20448 20668 20544
rect 21082 20476 21088 20528
rect 21140 20516 21146 20528
rect 21361 20519 21419 20525
rect 21361 20516 21373 20519
rect 21140 20488 21373 20516
rect 21140 20476 21146 20488
rect 21361 20485 21373 20488
rect 21407 20485 21419 20519
rect 21361 20479 21419 20485
rect 20579 20420 20668 20448
rect 21376 20448 21404 20479
rect 22002 20476 22008 20528
rect 22060 20516 22066 20528
rect 25314 20516 25320 20528
rect 22060 20488 25320 20516
rect 22060 20476 22066 20488
rect 25314 20476 25320 20488
rect 25372 20476 25378 20528
rect 21376 20420 21772 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20717 20383 20775 20389
rect 20717 20380 20729 20383
rect 20456 20352 20729 20380
rect 20717 20349 20729 20352
rect 20763 20349 20775 20383
rect 20717 20343 20775 20349
rect 21174 20340 21180 20392
rect 21232 20380 21238 20392
rect 21744 20380 21772 20420
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22152 20420 22197 20448
rect 22152 20408 22158 20420
rect 25406 20408 25412 20460
rect 25464 20448 25470 20460
rect 26145 20451 26203 20457
rect 26145 20448 26157 20451
rect 25464 20420 26157 20448
rect 25464 20408 25470 20420
rect 26145 20417 26157 20420
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 22189 20383 22247 20389
rect 22189 20380 22201 20383
rect 21232 20352 21680 20380
rect 21744 20352 22201 20380
rect 21232 20340 21238 20352
rect 19978 20272 19984 20324
rect 20036 20312 20042 20324
rect 21545 20315 21603 20321
rect 21545 20312 21557 20315
rect 20036 20284 21557 20312
rect 20036 20272 20042 20284
rect 21545 20281 21557 20284
rect 21591 20281 21603 20315
rect 21545 20275 21603 20281
rect 19208 20216 19748 20244
rect 21652 20244 21680 20352
rect 22189 20349 22201 20352
rect 22235 20349 22247 20383
rect 22189 20343 22247 20349
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22738 20380 22744 20392
rect 22699 20352 22744 20380
rect 22557 20343 22615 20349
rect 22572 20244 22600 20343
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 25869 20383 25927 20389
rect 25869 20349 25881 20383
rect 25915 20380 25927 20383
rect 26234 20380 26240 20392
rect 25915 20352 26240 20380
rect 25915 20349 25927 20352
rect 25869 20343 25927 20349
rect 26234 20340 26240 20352
rect 26292 20340 26298 20392
rect 58434 20272 58440 20324
rect 58492 20312 58498 20324
rect 59170 20312 59176 20324
rect 58492 20284 59176 20312
rect 58492 20272 58498 20284
rect 59170 20272 59176 20284
rect 59228 20272 59234 20324
rect 23750 20244 23756 20256
rect 21652 20216 23756 20244
rect 19208 20204 19214 20216
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 1104 20154 29256 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 29256 20154
rect 1104 20080 29256 20102
rect 2774 20000 2780 20052
rect 2832 20040 2838 20052
rect 4801 20043 4859 20049
rect 2832 20012 2877 20040
rect 2832 20000 2838 20012
rect 4801 20009 4813 20043
rect 4847 20009 4859 20043
rect 4801 20003 4859 20009
rect 5997 20043 6055 20049
rect 5997 20009 6009 20043
rect 6043 20040 6055 20043
rect 11425 20043 11483 20049
rect 11425 20040 11437 20043
rect 6043 20012 11437 20040
rect 6043 20009 6055 20012
rect 5997 20003 6055 20009
rect 11425 20009 11437 20012
rect 11471 20009 11483 20043
rect 11425 20003 11483 20009
rect 12897 20043 12955 20049
rect 12897 20009 12909 20043
rect 12943 20040 12955 20043
rect 13722 20040 13728 20052
rect 12943 20012 13728 20040
rect 12943 20009 12955 20012
rect 12897 20003 12955 20009
rect 2792 19904 2820 20000
rect 4816 19972 4844 20003
rect 11054 19972 11060 19984
rect 4816 19944 11060 19972
rect 11054 19932 11060 19944
rect 11112 19932 11118 19984
rect 11440 19972 11468 20003
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 16758 20000 16764 20052
rect 16816 20040 16822 20052
rect 17221 20043 17279 20049
rect 17221 20040 17233 20043
rect 16816 20012 17233 20040
rect 16816 20000 16822 20012
rect 17221 20009 17233 20012
rect 17267 20040 17279 20043
rect 21358 20040 21364 20052
rect 17267 20012 21364 20040
rect 17267 20009 17279 20012
rect 17221 20003 17279 20009
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 25406 20040 25412 20052
rect 25367 20012 25412 20040
rect 25406 20000 25412 20012
rect 25464 20000 25470 20052
rect 27522 20040 27528 20052
rect 27483 20012 27528 20040
rect 27522 20000 27528 20012
rect 27580 20000 27586 20052
rect 14734 19972 14740 19984
rect 11440 19944 14740 19972
rect 2869 19907 2927 19913
rect 2869 19904 2881 19907
rect 2792 19876 2881 19904
rect 2869 19873 2881 19876
rect 2915 19873 2927 19907
rect 4614 19904 4620 19916
rect 4575 19876 4620 19904
rect 2869 19867 2927 19873
rect 4614 19864 4620 19876
rect 4672 19864 4678 19916
rect 5810 19904 5816 19916
rect 5771 19876 5816 19904
rect 5810 19864 5816 19876
rect 5868 19864 5874 19916
rect 9490 19904 9496 19916
rect 9451 19876 9496 19904
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 9766 19904 9772 19916
rect 9727 19876 9772 19904
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 10042 19904 10048 19916
rect 10003 19876 10048 19904
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10502 19904 10508 19916
rect 10463 19876 10508 19904
rect 10502 19864 10508 19876
rect 10560 19864 10566 19916
rect 11440 19904 11468 19944
rect 14734 19932 14740 19944
rect 14792 19932 14798 19984
rect 25685 19975 25743 19981
rect 25685 19972 25697 19975
rect 24964 19944 25697 19972
rect 11609 19907 11667 19913
rect 11609 19904 11621 19907
rect 11440 19876 11621 19904
rect 11609 19873 11621 19876
rect 11655 19873 11667 19907
rect 12710 19904 12716 19916
rect 12671 19876 12716 19904
rect 11609 19867 11667 19873
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 16025 19907 16083 19913
rect 16025 19904 16037 19907
rect 15335 19876 16037 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 16025 19873 16037 19876
rect 16071 19873 16083 19907
rect 16025 19867 16083 19873
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19873 16267 19907
rect 16209 19867 16267 19873
rect 16485 19907 16543 19913
rect 16485 19873 16497 19907
rect 16531 19904 16543 19907
rect 17034 19904 17040 19916
rect 16531 19876 17040 19904
rect 16531 19873 16543 19876
rect 16485 19867 16543 19873
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 15013 19839 15071 19845
rect 15013 19836 15025 19839
rect 11296 19808 15025 19836
rect 11296 19796 11302 19808
rect 15013 19805 15025 19808
rect 15059 19805 15071 19839
rect 15562 19836 15568 19848
rect 15523 19808 15568 19836
rect 15013 19799 15071 19805
rect 9766 19728 9772 19780
rect 9824 19768 9830 19780
rect 10505 19771 10563 19777
rect 10505 19768 10517 19771
rect 9824 19740 10517 19768
rect 9824 19728 9830 19740
rect 10505 19737 10517 19740
rect 10551 19737 10563 19771
rect 15028 19768 15056 19799
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 16224 19768 16252 19867
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 24397 19907 24455 19913
rect 24397 19873 24409 19907
rect 24443 19904 24455 19907
rect 24854 19904 24860 19916
rect 24443 19876 24860 19904
rect 24443 19873 24455 19876
rect 24397 19867 24455 19873
rect 24854 19864 24860 19876
rect 24912 19904 24918 19916
rect 24964 19913 24992 19944
rect 25685 19941 25697 19944
rect 25731 19972 25743 19975
rect 25774 19972 25780 19984
rect 25731 19944 25780 19972
rect 25731 19941 25743 19944
rect 25685 19935 25743 19941
rect 25774 19932 25780 19944
rect 25832 19972 25838 19984
rect 25869 19975 25927 19981
rect 25869 19972 25881 19975
rect 25832 19944 25881 19972
rect 25832 19932 25838 19944
rect 25869 19941 25881 19944
rect 25915 19941 25927 19975
rect 25869 19935 25927 19941
rect 24949 19907 25007 19913
rect 24949 19904 24961 19907
rect 24912 19876 24961 19904
rect 24912 19864 24918 19876
rect 24949 19873 24961 19876
rect 24995 19873 25007 19907
rect 24949 19867 25007 19873
rect 25133 19907 25191 19913
rect 25133 19873 25145 19907
rect 25179 19904 25191 19907
rect 25406 19904 25412 19916
rect 25179 19876 25412 19904
rect 25179 19873 25191 19876
rect 25133 19867 25191 19873
rect 25406 19864 25412 19876
rect 25464 19904 25470 19916
rect 26605 19907 26663 19913
rect 25464 19876 26004 19904
rect 25464 19864 25470 19876
rect 16758 19836 16764 19848
rect 16719 19808 16764 19836
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 16942 19836 16948 19848
rect 16903 19808 16948 19836
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 24305 19839 24363 19845
rect 24305 19805 24317 19839
rect 24351 19805 24363 19839
rect 24305 19799 24363 19805
rect 18138 19768 18144 19780
rect 15028 19740 18144 19768
rect 10505 19731 10563 19737
rect 18138 19728 18144 19740
rect 18196 19728 18202 19780
rect 24121 19771 24179 19777
rect 24121 19737 24133 19771
rect 24167 19768 24179 19771
rect 24320 19768 24348 19799
rect 24762 19768 24768 19780
rect 24167 19740 24768 19768
rect 24167 19737 24179 19740
rect 24121 19731 24179 19737
rect 24762 19728 24768 19740
rect 24820 19728 24826 19780
rect 25976 19768 26004 19876
rect 26605 19873 26617 19907
rect 26651 19873 26663 19907
rect 27540 19904 27568 20000
rect 27617 19907 27675 19913
rect 27617 19904 27629 19907
rect 27540 19876 27629 19904
rect 26605 19867 26663 19873
rect 27617 19873 27629 19876
rect 27663 19873 27675 19907
rect 27617 19867 27675 19873
rect 26620 19836 26648 19867
rect 26973 19839 27031 19845
rect 26973 19836 26985 19839
rect 26620 19808 26985 19836
rect 26973 19805 26985 19808
rect 27019 19836 27031 19839
rect 27982 19836 27988 19848
rect 27019 19808 27988 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 27709 19771 27767 19777
rect 27709 19768 27721 19771
rect 25976 19740 27721 19768
rect 27709 19737 27721 19740
rect 27755 19737 27767 19771
rect 27709 19731 27767 19737
rect 3053 19703 3111 19709
rect 3053 19669 3065 19703
rect 3099 19700 3111 19703
rect 4062 19700 4068 19712
rect 3099 19672 4068 19700
rect 3099 19669 3111 19672
rect 3053 19663 3111 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 10042 19660 10048 19712
rect 10100 19700 10106 19712
rect 10318 19700 10324 19712
rect 10100 19672 10324 19700
rect 10100 19660 10106 19672
rect 10318 19660 10324 19672
rect 10376 19700 10382 19712
rect 10965 19703 11023 19709
rect 10965 19700 10977 19703
rect 10376 19672 10977 19700
rect 10376 19660 10382 19672
rect 10965 19669 10977 19672
rect 11011 19700 11023 19703
rect 11790 19700 11796 19712
rect 11011 19672 11796 19700
rect 11011 19669 11023 19672
rect 10965 19663 11023 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 14918 19700 14924 19712
rect 14424 19672 14924 19700
rect 14424 19660 14430 19672
rect 14918 19660 14924 19672
rect 14976 19700 14982 19712
rect 15289 19703 15347 19709
rect 15289 19700 15301 19703
rect 14976 19672 15301 19700
rect 14976 19660 14982 19672
rect 15289 19669 15301 19672
rect 15335 19700 15347 19703
rect 15381 19703 15439 19709
rect 15381 19700 15393 19703
rect 15335 19672 15393 19700
rect 15335 19669 15347 19672
rect 15289 19663 15347 19669
rect 15381 19669 15393 19672
rect 15427 19669 15439 19703
rect 26694 19700 26700 19712
rect 26655 19672 26700 19700
rect 15381 19663 15439 19669
rect 26694 19660 26700 19672
rect 26752 19660 26758 19712
rect 1104 19610 29256 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 29256 19610
rect 1104 19536 29256 19558
rect 10318 19496 10324 19508
rect 10279 19468 10324 19496
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 11149 19499 11207 19505
rect 11149 19465 11161 19499
rect 11195 19496 11207 19499
rect 11238 19496 11244 19508
rect 11195 19468 11244 19496
rect 11195 19465 11207 19468
rect 11149 19459 11207 19465
rect 11238 19456 11244 19468
rect 11296 19456 11302 19508
rect 16758 19496 16764 19508
rect 16719 19468 16764 19496
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 20680 19468 20729 19496
rect 20680 19456 20686 19468
rect 20717 19465 20729 19468
rect 20763 19496 20775 19499
rect 20898 19496 20904 19508
rect 20763 19468 20904 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 10336 19428 10364 19456
rect 9692 19400 10364 19428
rect 7926 19360 7932 19372
rect 7887 19332 7932 19360
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 9088 19332 9137 19360
rect 9088 19320 9094 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 9692 19360 9720 19400
rect 10134 19360 10140 19372
rect 9125 19323 9183 19329
rect 9600 19332 9720 19360
rect 10095 19332 10140 19360
rect 2590 19292 2596 19304
rect 2551 19264 2596 19292
rect 2590 19252 2596 19264
rect 2648 19252 2654 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 2958 19292 2964 19304
rect 2915 19264 2964 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 5261 19295 5319 19301
rect 5261 19261 5273 19295
rect 5307 19292 5319 19295
rect 5813 19295 5871 19301
rect 5813 19292 5825 19295
rect 5307 19264 5825 19292
rect 5307 19261 5319 19264
rect 5261 19255 5319 19261
rect 5813 19261 5825 19264
rect 5859 19292 5871 19295
rect 5902 19292 5908 19304
rect 5859 19264 5908 19292
rect 5859 19261 5871 19264
rect 5813 19255 5871 19261
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 9600 19301 9628 19332
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 15473 19363 15531 19369
rect 15120 19332 15332 19360
rect 7101 19295 7159 19301
rect 7101 19261 7113 19295
rect 7147 19292 7159 19295
rect 9585 19295 9643 19301
rect 7147 19264 7604 19292
rect 7147 19261 7159 19264
rect 7101 19255 7159 19261
rect 7576 19236 7604 19264
rect 9585 19261 9597 19295
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 9861 19295 9919 19301
rect 9861 19292 9873 19295
rect 9732 19264 9873 19292
rect 9732 19252 9738 19264
rect 9861 19261 9873 19264
rect 9907 19292 9919 19295
rect 10502 19292 10508 19304
rect 9907 19264 10508 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 10962 19292 10968 19304
rect 10923 19264 10968 19292
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 15120 19292 15148 19332
rect 11112 19264 15148 19292
rect 15197 19295 15255 19301
rect 11112 19252 11118 19264
rect 15197 19261 15209 19295
rect 15243 19261 15255 19295
rect 15304 19292 15332 19332
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 15562 19360 15568 19372
rect 15519 19332 15568 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 17586 19292 17592 19304
rect 15304 19264 17592 19292
rect 15197 19255 15255 19261
rect 4341 19227 4399 19233
rect 4341 19224 4353 19227
rect 3528 19196 4353 19224
rect 2590 19116 2596 19168
rect 2648 19156 2654 19168
rect 3528 19156 3556 19196
rect 4341 19193 4353 19196
rect 4387 19193 4399 19227
rect 4341 19187 4399 19193
rect 4890 19184 4896 19236
rect 4948 19224 4954 19236
rect 5077 19227 5135 19233
rect 5077 19224 5089 19227
rect 4948 19196 5089 19224
rect 4948 19184 4954 19196
rect 5077 19193 5089 19196
rect 5123 19193 5135 19227
rect 5626 19224 5632 19236
rect 5587 19196 5632 19224
rect 5077 19187 5135 19193
rect 5626 19184 5632 19196
rect 5684 19184 5690 19236
rect 7190 19224 7196 19236
rect 7151 19196 7196 19224
rect 7190 19184 7196 19196
rect 7248 19184 7254 19236
rect 7558 19224 7564 19236
rect 7519 19196 7564 19224
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 8941 19227 8999 19233
rect 8941 19193 8953 19227
rect 8987 19224 8999 19227
rect 9692 19224 9720 19252
rect 8987 19196 9720 19224
rect 8987 19193 8999 19196
rect 8941 19187 8999 19193
rect 3970 19156 3976 19168
rect 2648 19128 3556 19156
rect 3931 19128 3976 19156
rect 2648 19116 2654 19128
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 7374 19156 7380 19168
rect 7335 19128 7380 19156
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 7469 19159 7527 19165
rect 7469 19125 7481 19159
rect 7515 19156 7527 19159
rect 8570 19156 8576 19168
rect 7515 19128 8576 19156
rect 7515 19125 7527 19128
rect 7469 19119 7527 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 15105 19159 15163 19165
rect 15105 19125 15117 19159
rect 15151 19156 15163 19159
rect 15212 19156 15240 19255
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19168 19264 19349 19292
rect 17862 19156 17868 19168
rect 15151 19128 17868 19156
rect 15151 19125 15163 19128
rect 15105 19119 15163 19125
rect 17862 19116 17868 19128
rect 17920 19156 17926 19168
rect 19168 19165 19196 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19337 19255 19395 19261
rect 19426 19252 19432 19304
rect 19484 19292 19490 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19484 19264 19625 19292
rect 19484 19252 19490 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19261 25283 19295
rect 25225 19255 25283 19261
rect 25317 19295 25375 19301
rect 25317 19261 25329 19295
rect 25363 19261 25375 19295
rect 25682 19292 25688 19304
rect 25643 19264 25688 19292
rect 25317 19255 25375 19261
rect 24854 19184 24860 19236
rect 24912 19224 24918 19236
rect 25240 19224 25268 19255
rect 24912 19196 25268 19224
rect 24912 19184 24918 19196
rect 19153 19159 19211 19165
rect 19153 19156 19165 19159
rect 17920 19128 19165 19156
rect 17920 19116 17926 19128
rect 19153 19125 19165 19128
rect 19199 19125 19211 19159
rect 24946 19156 24952 19168
rect 24907 19128 24952 19156
rect 19153 19119 19211 19125
rect 24946 19116 24952 19128
rect 25004 19156 25010 19168
rect 25332 19156 25360 19255
rect 25682 19252 25688 19264
rect 25740 19252 25746 19304
rect 25774 19252 25780 19304
rect 25832 19292 25838 19304
rect 26513 19295 26571 19301
rect 26513 19292 26525 19295
rect 25832 19264 26525 19292
rect 25832 19252 25838 19264
rect 26513 19261 26525 19264
rect 26559 19292 26571 19295
rect 26697 19295 26755 19301
rect 26697 19292 26709 19295
rect 26559 19264 26709 19292
rect 26559 19261 26571 19264
rect 26513 19255 26571 19261
rect 26697 19261 26709 19264
rect 26743 19261 26755 19295
rect 26697 19255 26755 19261
rect 26329 19227 26387 19233
rect 26329 19193 26341 19227
rect 26375 19224 26387 19227
rect 26786 19224 26792 19236
rect 26375 19196 26792 19224
rect 26375 19193 26387 19196
rect 26329 19187 26387 19193
rect 26786 19184 26792 19196
rect 26844 19184 26850 19236
rect 25004 19128 25360 19156
rect 25004 19116 25010 19128
rect 25682 19116 25688 19168
rect 25740 19156 25746 19168
rect 26694 19156 26700 19168
rect 25740 19128 26700 19156
rect 25740 19116 25746 19128
rect 26694 19116 26700 19128
rect 26752 19116 26758 19168
rect 1104 19066 29256 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 29256 19066
rect 1104 18992 29256 19014
rect 4154 18952 4160 18964
rect 4115 18924 4160 18952
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 10244 18924 10609 18952
rect 4172 18816 4200 18912
rect 4525 18887 4583 18893
rect 4525 18853 4537 18887
rect 4571 18884 4583 18887
rect 5626 18884 5632 18896
rect 4571 18856 5632 18884
rect 4571 18853 4583 18856
rect 4525 18847 4583 18853
rect 5626 18844 5632 18856
rect 5684 18844 5690 18896
rect 9674 18844 9680 18896
rect 9732 18884 9738 18896
rect 9861 18887 9919 18893
rect 9861 18884 9873 18887
rect 9732 18856 9873 18884
rect 9732 18844 9738 18856
rect 9861 18853 9873 18856
rect 9907 18853 9919 18887
rect 9861 18847 9919 18853
rect 10045 18887 10103 18893
rect 10045 18853 10057 18887
rect 10091 18884 10103 18887
rect 10244 18884 10272 18924
rect 10597 18921 10609 18924
rect 10643 18952 10655 18955
rect 11054 18952 11060 18964
rect 10643 18924 11060 18952
rect 10643 18921 10655 18924
rect 10597 18915 10655 18921
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 11330 18912 11336 18964
rect 11388 18952 11394 18964
rect 11517 18955 11575 18961
rect 11517 18952 11529 18955
rect 11388 18924 11529 18952
rect 11388 18912 11394 18924
rect 11517 18921 11529 18924
rect 11563 18921 11575 18955
rect 11517 18915 11575 18921
rect 16209 18955 16267 18961
rect 16209 18921 16221 18955
rect 16255 18952 16267 18955
rect 18414 18952 18420 18964
rect 16255 18924 18420 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 10410 18884 10416 18896
rect 10091 18856 10272 18884
rect 10371 18856 10416 18884
rect 10091 18853 10103 18856
rect 10045 18847 10103 18853
rect 10410 18844 10416 18856
rect 10468 18844 10474 18896
rect 10962 18844 10968 18896
rect 11020 18884 11026 18896
rect 11609 18887 11667 18893
rect 11609 18884 11621 18887
rect 11020 18856 11621 18884
rect 11020 18844 11026 18856
rect 11609 18853 11621 18856
rect 11655 18884 11667 18887
rect 12158 18884 12164 18896
rect 11655 18856 12164 18884
rect 11655 18853 11667 18856
rect 11609 18847 11667 18853
rect 12158 18844 12164 18856
rect 12216 18844 12222 18896
rect 16224 18884 16252 18915
rect 18414 18912 18420 18924
rect 18472 18912 18478 18964
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 23845 18955 23903 18961
rect 23845 18952 23857 18955
rect 23808 18924 23857 18952
rect 23808 18912 23814 18924
rect 23845 18921 23857 18924
rect 23891 18952 23903 18955
rect 23891 18924 25268 18952
rect 23891 18921 23903 18924
rect 23845 18915 23903 18921
rect 18138 18884 18144 18896
rect 12360 18856 14228 18884
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 4172 18788 4353 18816
rect 4341 18785 4353 18788
rect 4387 18785 4399 18819
rect 4341 18779 4399 18785
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 5074 18816 5080 18828
rect 4663 18788 5080 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 4356 18748 4384 18779
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 9953 18819 10011 18825
rect 9953 18816 9965 18819
rect 8628 18788 9965 18816
rect 8628 18776 8634 18788
rect 9953 18785 9965 18788
rect 9999 18816 10011 18819
rect 11330 18816 11336 18828
rect 9999 18788 11336 18816
rect 9999 18785 10011 18788
rect 9953 18779 10011 18785
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12360 18816 12388 18856
rect 12023 18788 12388 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 6362 18748 6368 18760
rect 4356 18720 6368 18748
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 7190 18708 7196 18760
rect 7248 18748 7254 18760
rect 8846 18748 8852 18760
rect 7248 18720 8852 18748
rect 7248 18708 7254 18720
rect 8846 18708 8852 18720
rect 8904 18748 8910 18760
rect 9677 18751 9735 18757
rect 9677 18748 9689 18751
rect 8904 18720 9689 18748
rect 8904 18708 8910 18720
rect 9677 18717 9689 18720
rect 9723 18748 9735 18751
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 9723 18720 11253 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 11241 18711 11299 18717
rect 3418 18640 3424 18692
rect 3476 18680 3482 18692
rect 3476 18652 5120 18680
rect 3476 18640 3482 18652
rect 4801 18615 4859 18621
rect 4801 18581 4813 18615
rect 4847 18612 4859 18615
rect 4982 18612 4988 18624
rect 4847 18584 4988 18612
rect 4847 18581 4859 18584
rect 4801 18575 4859 18581
rect 4982 18572 4988 18584
rect 5040 18572 5046 18624
rect 5092 18612 5120 18652
rect 9214 18640 9220 18692
rect 9272 18680 9278 18692
rect 10410 18680 10416 18692
rect 9272 18652 10416 18680
rect 9272 18640 9278 18652
rect 10410 18640 10416 18652
rect 10468 18640 10474 18692
rect 10778 18640 10784 18692
rect 10836 18680 10842 18692
rect 11440 18680 11468 18779
rect 10836 18652 11468 18680
rect 14200 18680 14228 18856
rect 15488 18856 16252 18884
rect 18099 18856 18144 18884
rect 15488 18825 15516 18856
rect 18138 18844 18144 18856
rect 18196 18884 18202 18896
rect 20162 18884 20168 18896
rect 18196 18856 19196 18884
rect 18196 18844 18202 18856
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18785 15531 18819
rect 15473 18779 15531 18785
rect 15565 18819 15623 18825
rect 15565 18785 15577 18819
rect 15611 18816 15623 18819
rect 16390 18816 16396 18828
rect 15611 18788 16396 18816
rect 15611 18785 15623 18788
rect 15565 18779 15623 18785
rect 14274 18708 14280 18760
rect 14332 18748 14338 18760
rect 15580 18748 15608 18779
rect 16390 18776 16396 18788
rect 16448 18816 16454 18828
rect 16853 18819 16911 18825
rect 16853 18816 16865 18819
rect 16448 18788 16865 18816
rect 16448 18776 16454 18788
rect 16853 18785 16865 18788
rect 16899 18785 16911 18819
rect 16853 18779 16911 18785
rect 18417 18819 18475 18825
rect 18417 18785 18429 18819
rect 18463 18816 18475 18819
rect 18966 18816 18972 18828
rect 18463 18788 18972 18816
rect 18463 18785 18475 18788
rect 18417 18779 18475 18785
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 19168 18825 19196 18856
rect 19444 18856 20168 18884
rect 19444 18828 19472 18856
rect 20162 18844 20168 18856
rect 20220 18844 20226 18896
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18785 19211 18819
rect 19426 18816 19432 18828
rect 19387 18788 19432 18816
rect 19153 18779 19211 18785
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18816 19855 18819
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 19843 18788 20085 18816
rect 19843 18785 19855 18788
rect 19797 18779 19855 18785
rect 20073 18785 20085 18788
rect 20119 18816 20131 18819
rect 21174 18816 21180 18828
rect 20119 18788 21180 18816
rect 20119 18785 20131 18788
rect 20073 18779 20131 18785
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 24026 18776 24032 18828
rect 24084 18816 24090 18828
rect 25240 18825 25268 18924
rect 24857 18819 24915 18825
rect 24857 18816 24869 18819
rect 24084 18788 24869 18816
rect 24084 18776 24090 18788
rect 24857 18785 24869 18788
rect 24903 18785 24915 18819
rect 24857 18779 24915 18785
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 18506 18748 18512 18760
rect 14332 18720 15608 18748
rect 18467 18720 18512 18748
rect 14332 18708 14338 18720
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 19889 18751 19947 18757
rect 19889 18748 19901 18751
rect 18840 18720 19901 18748
rect 18840 18708 18846 18720
rect 19889 18717 19901 18720
rect 19935 18717 19947 18751
rect 24210 18748 24216 18760
rect 24171 18720 24216 18748
rect 19889 18711 19947 18717
rect 24210 18708 24216 18720
rect 24268 18708 24274 18760
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 24118 18680 24124 18692
rect 14200 18652 24124 18680
rect 10836 18640 10842 18652
rect 24118 18640 24124 18652
rect 24176 18640 24182 18692
rect 24964 18680 24992 18711
rect 25038 18708 25044 18760
rect 25096 18748 25102 18760
rect 25133 18751 25191 18757
rect 25133 18748 25145 18751
rect 25096 18720 25145 18748
rect 25096 18708 25102 18720
rect 25133 18717 25145 18720
rect 25179 18717 25191 18751
rect 25133 18711 25191 18717
rect 25774 18680 25780 18692
rect 24964 18652 25780 18680
rect 25774 18640 25780 18652
rect 25832 18640 25838 18692
rect 14458 18612 14464 18624
rect 5092 18584 14464 18612
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 15746 18612 15752 18624
rect 15707 18584 15752 18612
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 17034 18612 17040 18624
rect 16995 18584 17040 18612
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 21726 18612 21732 18624
rect 17184 18584 21732 18612
rect 17184 18572 17190 18584
rect 21726 18572 21732 18584
rect 21784 18572 21790 18624
rect 24026 18612 24032 18624
rect 23987 18584 24032 18612
rect 24026 18572 24032 18584
rect 24084 18572 24090 18624
rect 1104 18522 29256 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 29256 18522
rect 1104 18448 29256 18470
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 5132 18380 13952 18408
rect 5132 18368 5138 18380
rect 7009 18343 7067 18349
rect 7009 18309 7021 18343
rect 7055 18340 7067 18343
rect 7190 18340 7196 18352
rect 7055 18312 7196 18340
rect 7055 18309 7067 18312
rect 7009 18303 7067 18309
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 7282 18300 7288 18352
rect 7340 18340 7346 18352
rect 12434 18340 12440 18352
rect 7340 18312 12440 18340
rect 7340 18300 7346 18312
rect 12434 18300 12440 18312
rect 12492 18340 12498 18352
rect 13538 18340 13544 18352
rect 12492 18312 13544 18340
rect 12492 18300 12498 18312
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 13630 18300 13636 18352
rect 13688 18340 13694 18352
rect 13725 18343 13783 18349
rect 13725 18340 13737 18343
rect 13688 18312 13737 18340
rect 13688 18300 13694 18312
rect 13725 18309 13737 18312
rect 13771 18309 13783 18343
rect 13924 18340 13952 18380
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 15105 18411 15163 18417
rect 15105 18408 15117 18411
rect 14884 18380 15117 18408
rect 14884 18368 14890 18380
rect 15105 18377 15117 18380
rect 15151 18377 15163 18411
rect 15105 18371 15163 18377
rect 15194 18368 15200 18420
rect 15252 18408 15258 18420
rect 24026 18408 24032 18420
rect 15252 18380 24032 18408
rect 15252 18368 15258 18380
rect 24026 18368 24032 18380
rect 24084 18368 24090 18420
rect 25314 18368 25320 18420
rect 25372 18408 25378 18420
rect 25866 18408 25872 18420
rect 25372 18380 25872 18408
rect 25372 18368 25378 18380
rect 25866 18368 25872 18380
rect 25924 18368 25930 18420
rect 27706 18408 27712 18420
rect 27667 18380 27712 18408
rect 27706 18368 27712 18380
rect 27764 18368 27770 18420
rect 15289 18343 15347 18349
rect 15289 18340 15301 18343
rect 13924 18312 15301 18340
rect 13725 18303 13783 18309
rect 15289 18309 15301 18312
rect 15335 18309 15347 18343
rect 21174 18340 21180 18352
rect 21135 18312 21180 18340
rect 15289 18303 15347 18309
rect 21174 18300 21180 18312
rect 21232 18300 21238 18352
rect 25774 18300 25780 18352
rect 25832 18340 25838 18352
rect 27433 18343 27491 18349
rect 27433 18340 27445 18343
rect 25832 18312 27445 18340
rect 25832 18300 25838 18312
rect 27433 18309 27445 18312
rect 27479 18309 27491 18343
rect 27433 18303 27491 18309
rect 2685 18275 2743 18281
rect 2685 18241 2697 18275
rect 2731 18272 2743 18275
rect 3697 18275 3755 18281
rect 3697 18272 3709 18275
rect 2731 18244 3709 18272
rect 2731 18241 2743 18244
rect 2685 18235 2743 18241
rect 3697 18241 3709 18244
rect 3743 18272 3755 18275
rect 5810 18272 5816 18284
rect 3743 18244 5304 18272
rect 5771 18244 5816 18272
rect 3743 18241 3755 18244
rect 3697 18235 3755 18241
rect 5276 18216 5304 18244
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 8846 18232 8852 18284
rect 8904 18272 8910 18284
rect 9493 18275 9551 18281
rect 9493 18272 9505 18275
rect 8904 18244 9505 18272
rect 8904 18232 8910 18244
rect 9493 18241 9505 18244
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 18506 18232 18512 18284
rect 18564 18272 18570 18284
rect 20073 18275 20131 18281
rect 20073 18272 20085 18275
rect 18564 18244 20085 18272
rect 18564 18232 18570 18244
rect 20073 18241 20085 18244
rect 20119 18241 20131 18275
rect 32766 18272 32772 18284
rect 20073 18235 20131 18241
rect 26252 18244 32772 18272
rect 2501 18207 2559 18213
rect 2501 18173 2513 18207
rect 2547 18204 2559 18207
rect 2593 18207 2651 18213
rect 2593 18204 2605 18207
rect 2547 18176 2605 18204
rect 2547 18173 2559 18176
rect 2501 18167 2559 18173
rect 2593 18173 2605 18176
rect 2639 18173 2651 18207
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 2593 18167 2651 18173
rect 3252 18176 3617 18204
rect 2608 18136 2636 18167
rect 3142 18136 3148 18148
rect 2608 18108 3148 18136
rect 3142 18096 3148 18108
rect 3200 18096 3206 18148
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3252 18077 3280 18176
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 3605 18167 3663 18173
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18173 3939 18207
rect 5166 18204 5172 18216
rect 5127 18176 5172 18204
rect 3881 18167 3939 18173
rect 3237 18071 3295 18077
rect 3237 18068 3249 18071
rect 3016 18040 3249 18068
rect 3016 18028 3022 18040
rect 3237 18037 3249 18040
rect 3283 18037 3295 18071
rect 3418 18068 3424 18080
rect 3379 18040 3424 18068
rect 3237 18031 3295 18037
rect 3418 18028 3424 18040
rect 3476 18068 3482 18080
rect 3896 18068 3924 18167
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5445 18207 5503 18213
rect 5316 18176 5361 18204
rect 5316 18164 5322 18176
rect 5445 18173 5457 18207
rect 5491 18204 5503 18207
rect 6270 18204 6276 18216
rect 5491 18176 6276 18204
rect 5491 18173 5503 18176
rect 5445 18167 5503 18173
rect 6270 18164 6276 18176
rect 6328 18204 6334 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6328 18176 6837 18204
rect 6328 18164 6334 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 7926 18204 7932 18216
rect 7887 18176 7932 18204
rect 6825 18167 6883 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 9769 18207 9827 18213
rect 9769 18204 9781 18207
rect 8628 18176 9781 18204
rect 8628 18164 8634 18176
rect 9769 18173 9781 18176
rect 9815 18173 9827 18207
rect 11146 18204 11152 18216
rect 9769 18167 9827 18173
rect 9876 18176 11152 18204
rect 9876 18145 9904 18176
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13446 18204 13452 18216
rect 13407 18176 13452 18204
rect 13446 18164 13452 18176
rect 13504 18164 13510 18216
rect 13538 18164 13544 18216
rect 13596 18204 13602 18216
rect 15010 18213 15016 18216
rect 13725 18207 13783 18213
rect 13725 18204 13737 18207
rect 13596 18176 13737 18204
rect 13596 18164 13602 18176
rect 13725 18173 13737 18176
rect 13771 18173 13783 18207
rect 13725 18167 13783 18173
rect 14976 18207 15016 18213
rect 14976 18173 14988 18207
rect 14976 18167 15016 18173
rect 15010 18164 15016 18167
rect 15068 18164 15074 18216
rect 15168 18207 15226 18213
rect 15168 18173 15180 18207
rect 15214 18204 15226 18207
rect 16390 18204 16396 18216
rect 15214 18173 15240 18204
rect 16351 18176 16396 18204
rect 15168 18167 15240 18173
rect 4341 18139 4399 18145
rect 4341 18105 4353 18139
rect 4387 18136 4399 18139
rect 9861 18139 9919 18145
rect 4387 18108 9352 18136
rect 4387 18105 4399 18108
rect 4341 18099 4399 18105
rect 8110 18068 8116 18080
rect 3476 18040 3924 18068
rect 8071 18040 8116 18068
rect 3476 18028 3482 18040
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 9324 18068 9352 18108
rect 9508 18108 9812 18136
rect 9508 18068 9536 18108
rect 9674 18068 9680 18080
rect 9324 18040 9536 18068
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 9784 18068 9812 18108
rect 9861 18105 9873 18139
rect 9907 18105 9919 18139
rect 9861 18099 9919 18105
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 10229 18139 10287 18145
rect 10229 18136 10241 18139
rect 10100 18108 10241 18136
rect 10100 18096 10106 18108
rect 10229 18105 10241 18108
rect 10275 18105 10287 18139
rect 10229 18099 10287 18105
rect 13170 18096 13176 18148
rect 13228 18136 13234 18148
rect 14829 18139 14887 18145
rect 14829 18136 14841 18139
rect 13228 18108 14841 18136
rect 13228 18096 13234 18108
rect 14829 18105 14841 18108
rect 14875 18105 14887 18139
rect 15212 18136 15240 18167
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18204 19579 18207
rect 19797 18207 19855 18213
rect 19797 18204 19809 18207
rect 19567 18176 19809 18204
rect 19567 18173 19579 18176
rect 19521 18167 19579 18173
rect 19797 18173 19809 18176
rect 19843 18173 19855 18207
rect 19797 18167 19855 18173
rect 24762 18164 24768 18216
rect 24820 18204 24826 18216
rect 24949 18207 25007 18213
rect 24949 18204 24961 18207
rect 24820 18176 24961 18204
rect 24820 18164 24826 18176
rect 24949 18173 24961 18176
rect 24995 18204 25007 18207
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 24995 18176 25145 18204
rect 24995 18173 25007 18176
rect 24949 18167 25007 18173
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25314 18204 25320 18216
rect 25275 18176 25320 18204
rect 25133 18167 25191 18173
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 25774 18204 25780 18216
rect 25735 18176 25780 18204
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 25866 18164 25872 18216
rect 25924 18204 25930 18216
rect 25924 18176 25969 18204
rect 25924 18164 25930 18176
rect 15746 18136 15752 18148
rect 15212 18108 15752 18136
rect 14829 18099 14887 18105
rect 15746 18096 15752 18108
rect 15804 18096 15810 18148
rect 18966 18096 18972 18148
rect 19024 18136 19030 18148
rect 19024 18108 19932 18136
rect 19024 18096 19030 18108
rect 10870 18068 10876 18080
rect 9784 18040 10876 18068
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11790 18028 11796 18080
rect 11848 18068 11854 18080
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 11848 18040 12817 18068
rect 11848 18028 11854 18040
rect 12805 18037 12817 18040
rect 12851 18068 12863 18071
rect 13446 18068 13452 18080
rect 12851 18040 13452 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 13446 18028 13452 18040
rect 13504 18068 13510 18080
rect 15194 18068 15200 18080
rect 13504 18040 15200 18068
rect 13504 18028 13510 18040
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 16577 18071 16635 18077
rect 16577 18037 16589 18071
rect 16623 18068 16635 18071
rect 16666 18068 16672 18080
rect 16623 18040 16672 18068
rect 16623 18037 16635 18040
rect 16577 18031 16635 18037
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 19521 18071 19579 18077
rect 19521 18068 19533 18071
rect 17920 18040 19533 18068
rect 17920 18028 17926 18040
rect 19521 18037 19533 18040
rect 19567 18068 19579 18071
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19567 18040 19625 18068
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 19904 18068 19932 18108
rect 21174 18096 21180 18148
rect 21232 18136 21238 18148
rect 26252 18136 26280 18244
rect 32766 18232 32772 18244
rect 32824 18232 32830 18284
rect 27341 18207 27399 18213
rect 27341 18173 27353 18207
rect 27387 18204 27399 18207
rect 27706 18204 27712 18216
rect 27387 18176 27712 18204
rect 27387 18173 27399 18176
rect 27341 18167 27399 18173
rect 27706 18164 27712 18176
rect 27764 18164 27770 18216
rect 26418 18136 26424 18148
rect 21232 18108 26280 18136
rect 26379 18108 26424 18136
rect 21232 18096 21238 18108
rect 26418 18096 26424 18108
rect 26476 18096 26482 18148
rect 21542 18068 21548 18080
rect 19904 18040 21548 18068
rect 19613 18031 19671 18037
rect 21542 18028 21548 18040
rect 21600 18068 21606 18080
rect 24762 18068 24768 18080
rect 21600 18040 24768 18068
rect 21600 18028 21606 18040
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 1104 17978 29256 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 29256 17978
rect 1104 17904 29256 17926
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 4614 17864 4620 17876
rect 4571 17836 4620 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 8570 17864 8576 17876
rect 8531 17836 8576 17864
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 9214 17824 9220 17876
rect 9272 17864 9278 17876
rect 10413 17867 10471 17873
rect 10413 17864 10425 17867
rect 9272 17836 10425 17864
rect 9272 17824 9278 17836
rect 10413 17833 10425 17836
rect 10459 17864 10471 17867
rect 10778 17864 10784 17876
rect 10459 17836 10784 17864
rect 10459 17833 10471 17836
rect 10413 17827 10471 17833
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 12710 17864 12716 17876
rect 10980 17836 12716 17864
rect 5166 17756 5172 17808
rect 5224 17796 5230 17808
rect 6733 17799 6791 17805
rect 5224 17768 6592 17796
rect 5224 17756 5230 17768
rect 2958 17728 2964 17740
rect 2919 17700 2964 17728
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4614 17728 4620 17740
rect 4387 17700 4620 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17660 3111 17663
rect 4080 17660 4108 17691
rect 4614 17688 4620 17700
rect 4672 17728 4678 17740
rect 5994 17728 6000 17740
rect 4672 17700 5212 17728
rect 5955 17700 6000 17728
rect 4672 17688 4678 17700
rect 5074 17660 5080 17672
rect 3099 17632 5080 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 4157 17595 4215 17601
rect 4157 17561 4169 17595
rect 4203 17561 4215 17595
rect 4157 17555 4215 17561
rect 2869 17527 2927 17533
rect 2869 17493 2881 17527
rect 2915 17524 2927 17527
rect 2958 17524 2964 17536
rect 2915 17496 2964 17524
rect 2915 17493 2927 17496
rect 2869 17487 2927 17493
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 3694 17524 3700 17536
rect 3200 17496 3700 17524
rect 3200 17484 3206 17496
rect 3694 17484 3700 17496
rect 3752 17524 3758 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3752 17496 3801 17524
rect 3752 17484 3758 17496
rect 3789 17493 3801 17496
rect 3835 17524 3847 17527
rect 4172 17524 4200 17555
rect 3835 17496 4200 17524
rect 5184 17524 5212 17700
rect 5994 17688 6000 17700
rect 6052 17688 6058 17740
rect 6270 17728 6276 17740
rect 6231 17700 6276 17728
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 6564 17728 6592 17768
rect 6733 17765 6745 17799
rect 6779 17796 6791 17799
rect 7926 17796 7932 17808
rect 6779 17768 7932 17796
rect 6779 17765 6791 17768
rect 6733 17759 6791 17765
rect 7926 17756 7932 17768
rect 7984 17756 7990 17808
rect 10502 17796 10508 17808
rect 9140 17768 10508 17796
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 6564 17700 8401 17728
rect 8389 17697 8401 17700
rect 8435 17728 8447 17731
rect 9030 17728 9036 17740
rect 8435 17700 9036 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 6012 17660 6040 17688
rect 9140 17660 9168 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 10597 17799 10655 17805
rect 10597 17765 10609 17799
rect 10643 17796 10655 17799
rect 10870 17796 10876 17808
rect 10643 17768 10876 17796
rect 10643 17765 10655 17768
rect 10597 17759 10655 17765
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 10980 17805 11008 17836
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 23017 17867 23075 17873
rect 23017 17833 23029 17867
rect 23063 17864 23075 17867
rect 23842 17864 23848 17876
rect 23063 17836 23848 17864
rect 23063 17833 23075 17836
rect 23017 17827 23075 17833
rect 10965 17799 11023 17805
rect 10965 17765 10977 17799
rect 11011 17765 11023 17799
rect 10965 17759 11023 17765
rect 11054 17756 11060 17808
rect 11112 17796 11118 17808
rect 11977 17799 12035 17805
rect 11977 17796 11989 17799
rect 11112 17768 11989 17796
rect 11112 17756 11118 17768
rect 11977 17765 11989 17768
rect 12023 17765 12035 17799
rect 12158 17796 12164 17808
rect 12119 17768 12164 17796
rect 11977 17759 12035 17765
rect 12158 17756 12164 17768
rect 12216 17756 12222 17808
rect 18690 17796 18696 17808
rect 16592 17768 18696 17796
rect 9674 17728 9680 17740
rect 6012 17632 9168 17660
rect 9232 17700 9680 17728
rect 5350 17552 5356 17604
rect 5408 17592 5414 17604
rect 6089 17595 6147 17601
rect 6089 17592 6101 17595
rect 5408 17564 6101 17592
rect 5408 17552 5414 17564
rect 6089 17561 6101 17564
rect 6135 17592 6147 17595
rect 9232 17592 9260 17700
rect 9674 17688 9680 17700
rect 9732 17728 9738 17740
rect 10410 17728 10416 17740
rect 9732 17700 10416 17728
rect 9732 17688 9738 17700
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17728 11207 17731
rect 11238 17728 11244 17740
rect 11195 17700 11244 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 16592 17737 16620 17768
rect 18690 17756 18696 17768
rect 18748 17756 18754 17808
rect 21545 17799 21603 17805
rect 21545 17796 21557 17799
rect 20916 17768 21557 17796
rect 20916 17740 20944 17768
rect 21545 17765 21557 17768
rect 21591 17765 21603 17799
rect 21545 17759 21603 17765
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11388 17700 12081 17728
rect 11388 17688 11394 17700
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17697 16635 17731
rect 16577 17691 16635 17697
rect 16669 17731 16727 17737
rect 16669 17697 16681 17731
rect 16715 17697 16727 17731
rect 16853 17731 16911 17737
rect 16853 17728 16865 17731
rect 16669 17691 16727 17697
rect 16776 17700 16865 17728
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 6135 17564 9260 17592
rect 9600 17632 10241 17660
rect 6135 17561 6147 17564
rect 6089 17555 6147 17561
rect 9600 17524 9628 17632
rect 10229 17629 10241 17632
rect 10275 17660 10287 17663
rect 10870 17660 10876 17672
rect 10275 17632 10876 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10870 17620 10876 17632
rect 10928 17660 10934 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 10928 17632 11805 17660
rect 10928 17620 10934 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12618 17660 12624 17672
rect 12575 17632 12624 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 12618 17620 12624 17632
rect 12676 17620 12682 17672
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 16040 17592 16068 17623
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 16684 17660 16712 17691
rect 16540 17632 16712 17660
rect 16540 17620 16546 17632
rect 9732 17564 16068 17592
rect 9732 17552 9738 17564
rect 5184 17496 9628 17524
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 15102 17524 15108 17536
rect 10560 17496 15108 17524
rect 10560 17484 10566 17496
rect 15102 17484 15108 17496
rect 15160 17524 15166 17536
rect 16776 17524 16804 17700
rect 16853 17697 16865 17700
rect 16899 17697 16911 17731
rect 16853 17691 16911 17697
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 17954 17728 17960 17740
rect 17359 17700 17960 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 20714 17728 20720 17740
rect 19843 17700 20720 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 20714 17688 20720 17700
rect 20772 17688 20778 17740
rect 20898 17728 20904 17740
rect 20859 17700 20904 17728
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 20993 17731 21051 17737
rect 20993 17697 21005 17731
rect 21039 17697 21051 17731
rect 22370 17728 22376 17740
rect 22331 17700 22376 17728
rect 20993 17691 21051 17697
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17092 17632 17417 17660
rect 17092 17620 17098 17632
rect 17405 17629 17417 17632
rect 17451 17660 17463 17663
rect 19426 17660 19432 17672
rect 17451 17632 19432 17660
rect 17451 17629 17463 17632
rect 17405 17623 17463 17629
rect 19426 17620 19432 17632
rect 19484 17660 19490 17672
rect 21008 17660 21036 17691
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 21450 17660 21456 17672
rect 19484 17632 21036 17660
rect 21411 17632 21456 17660
rect 19484 17620 19490 17632
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22281 17663 22339 17669
rect 22281 17629 22293 17663
rect 22327 17660 22339 17663
rect 23032 17660 23060 17827
rect 23842 17824 23848 17836
rect 23900 17824 23906 17876
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24121 17867 24179 17873
rect 24121 17864 24133 17867
rect 24084 17836 24133 17864
rect 24084 17824 24090 17836
rect 24121 17833 24133 17836
rect 24167 17864 24179 17867
rect 26234 17864 26240 17876
rect 24167 17836 25360 17864
rect 26195 17836 26240 17864
rect 24167 17833 24179 17836
rect 24121 17827 24179 17833
rect 23750 17756 23756 17808
rect 23808 17796 23814 17808
rect 23937 17799 23995 17805
rect 23937 17796 23949 17799
rect 23808 17768 23949 17796
rect 23808 17756 23814 17768
rect 23937 17765 23949 17768
rect 23983 17765 23995 17799
rect 23937 17759 23995 17765
rect 23952 17728 23980 17759
rect 25332 17737 25360 17836
rect 26234 17824 26240 17836
rect 26292 17824 26298 17876
rect 27706 17824 27712 17876
rect 27764 17864 27770 17876
rect 27893 17867 27951 17873
rect 27893 17864 27905 17867
rect 27764 17836 27905 17864
rect 27764 17824 27770 17836
rect 27893 17833 27905 17836
rect 27939 17833 27951 17867
rect 27893 17827 27951 17833
rect 24949 17731 25007 17737
rect 24949 17728 24961 17731
rect 23952 17700 24961 17728
rect 24949 17697 24961 17700
rect 24995 17697 25007 17731
rect 24949 17691 25007 17697
rect 25317 17731 25375 17737
rect 25317 17697 25329 17731
rect 25363 17697 25375 17731
rect 25317 17691 25375 17697
rect 25501 17731 25559 17737
rect 25501 17697 25513 17731
rect 25547 17728 25559 17731
rect 26326 17728 26332 17740
rect 25547 17700 26332 17728
rect 25547 17697 25559 17700
rect 25501 17691 25559 17697
rect 26326 17688 26332 17700
rect 26384 17688 26390 17740
rect 26418 17688 26424 17740
rect 26476 17728 26482 17740
rect 26789 17731 26847 17737
rect 26789 17728 26801 17731
rect 26476 17700 26801 17728
rect 26476 17688 26482 17700
rect 26789 17697 26801 17700
rect 26835 17697 26847 17731
rect 26789 17691 26847 17697
rect 22327 17632 23060 17660
rect 22327 17629 22339 17632
rect 22281 17623 22339 17629
rect 23658 17620 23664 17672
rect 23716 17660 23722 17672
rect 24305 17663 24363 17669
rect 24305 17660 24317 17663
rect 23716 17632 24317 17660
rect 23716 17620 23722 17632
rect 24305 17629 24317 17632
rect 24351 17629 24363 17663
rect 24305 17623 24363 17629
rect 25041 17663 25099 17669
rect 25041 17629 25053 17663
rect 25087 17660 25099 17663
rect 25682 17660 25688 17672
rect 25087 17632 25688 17660
rect 25087 17629 25099 17632
rect 25041 17623 25099 17629
rect 25682 17620 25688 17632
rect 25740 17620 25746 17672
rect 26234 17620 26240 17672
rect 26292 17660 26298 17672
rect 26513 17663 26571 17669
rect 26513 17660 26525 17663
rect 26292 17632 26525 17660
rect 26292 17620 26298 17632
rect 26513 17629 26525 17632
rect 26559 17629 26571 17663
rect 26513 17623 26571 17629
rect 17494 17552 17500 17604
rect 17552 17592 17558 17604
rect 22186 17592 22192 17604
rect 17552 17564 22192 17592
rect 17552 17552 17558 17564
rect 22186 17552 22192 17564
rect 22244 17552 22250 17604
rect 15160 17496 16804 17524
rect 19889 17527 19947 17533
rect 15160 17484 15166 17496
rect 19889 17493 19901 17527
rect 19935 17524 19947 17527
rect 20898 17524 20904 17536
rect 19935 17496 20904 17524
rect 19935 17493 19947 17496
rect 19889 17487 19947 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 22557 17527 22615 17533
rect 22557 17524 22569 17527
rect 22152 17496 22569 17524
rect 22152 17484 22158 17496
rect 22557 17493 22569 17496
rect 22603 17493 22615 17527
rect 22557 17487 22615 17493
rect 1104 17434 29256 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 29256 17434
rect 1104 17360 29256 17382
rect 3418 17280 3424 17332
rect 3476 17320 3482 17332
rect 5537 17323 5595 17329
rect 5537 17320 5549 17323
rect 3476 17292 5549 17320
rect 3476 17280 3482 17292
rect 5537 17289 5549 17292
rect 5583 17289 5595 17323
rect 5537 17283 5595 17289
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6270 17320 6276 17332
rect 5859 17292 6276 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 3237 17255 3295 17261
rect 3237 17221 3249 17255
rect 3283 17252 3295 17255
rect 3283 17224 4476 17252
rect 3283 17221 3295 17224
rect 3237 17215 3295 17221
rect 3053 17119 3111 17125
rect 3053 17085 3065 17119
rect 3099 17116 3111 17119
rect 3418 17116 3424 17128
rect 3099 17088 3424 17116
rect 3099 17085 3111 17088
rect 3053 17079 3111 17085
rect 3068 16992 3096 17079
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 4154 17116 4160 17128
rect 4115 17088 4160 17116
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 4448 17125 4476 17224
rect 4433 17119 4491 17125
rect 4304 17088 4349 17116
rect 4304 17076 4310 17088
rect 4433 17085 4445 17119
rect 4479 17116 4491 17119
rect 4614 17116 4620 17128
rect 4479 17088 4620 17116
rect 4479 17085 4491 17088
rect 4433 17079 4491 17085
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 4890 17116 4896 17128
rect 4803 17088 4896 17116
rect 4890 17076 4896 17088
rect 4948 17116 4954 17128
rect 5552 17116 5580 17283
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 12713 17323 12771 17329
rect 12713 17320 12725 17323
rect 9640 17292 12725 17320
rect 9640 17280 9646 17292
rect 8846 17212 8852 17264
rect 8904 17252 8910 17264
rect 9398 17252 9404 17264
rect 8904 17224 9404 17252
rect 8904 17212 8910 17224
rect 9398 17212 9404 17224
rect 9456 17212 9462 17264
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 9048 17156 9689 17184
rect 9048 17128 9076 17156
rect 9677 17153 9689 17156
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17184 10011 17187
rect 11425 17187 11483 17193
rect 11425 17184 11437 17187
rect 9999 17156 11437 17184
rect 9999 17153 10011 17156
rect 9953 17147 10011 17153
rect 11425 17153 11437 17156
rect 11471 17153 11483 17187
rect 11425 17147 11483 17153
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 4948 17088 5488 17116
rect 5552 17088 5733 17116
rect 4948 17076 4954 17088
rect 4172 17048 4200 17076
rect 5166 17048 5172 17060
rect 4172 17020 5172 17048
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 5460 17048 5488 17088
rect 5721 17085 5733 17088
rect 5767 17085 5779 17119
rect 9030 17116 9036 17128
rect 8991 17088 9036 17116
rect 5721 17079 5779 17085
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 9214 17116 9220 17128
rect 9175 17088 9220 17116
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 9398 17116 9404 17128
rect 9359 17088 9404 17116
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 10870 17116 10876 17128
rect 10831 17088 10876 17116
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 10962 17076 10968 17128
rect 11020 17116 11026 17128
rect 11020 17088 11113 17116
rect 11020 17076 11026 17088
rect 7282 17048 7288 17060
rect 5460 17020 7288 17048
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 8573 17051 8631 17057
rect 8573 17017 8585 17051
rect 8619 17048 8631 17051
rect 9858 17048 9864 17060
rect 8619 17020 9864 17048
rect 8619 17017 8631 17020
rect 8573 17011 8631 17017
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 10410 17008 10416 17060
rect 10468 17048 10474 17060
rect 10980 17048 11008 17076
rect 10468 17020 11008 17048
rect 11440 17048 11468 17147
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17116 12495 17119
rect 12544 17116 12572 17292
rect 12713 17289 12725 17292
rect 12759 17289 12771 17323
rect 16850 17320 16856 17332
rect 16811 17292 16856 17320
rect 12713 17283 12771 17289
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 21174 17280 21180 17332
rect 21232 17320 21238 17332
rect 21361 17323 21419 17329
rect 21361 17320 21373 17323
rect 21232 17292 21373 17320
rect 21232 17280 21238 17292
rect 21361 17289 21373 17292
rect 21407 17289 21419 17323
rect 21818 17320 21824 17332
rect 21779 17292 21824 17320
rect 21361 17283 21419 17289
rect 16758 17252 16764 17264
rect 16592 17224 16764 17252
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17184 14059 17187
rect 14645 17187 14703 17193
rect 14047 17156 14228 17184
rect 14047 17153 14059 17156
rect 14001 17147 14059 17153
rect 12483 17088 12572 17116
rect 13817 17119 13875 17125
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 14090 17116 14096 17128
rect 13863 17088 14096 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 14200 17125 14228 17156
rect 14645 17153 14657 17187
rect 14691 17184 14703 17187
rect 15010 17184 15016 17196
rect 14691 17156 15016 17184
rect 14691 17153 14703 17156
rect 14645 17147 14703 17153
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 16592 17193 16620 17224
rect 16758 17212 16764 17224
rect 16816 17252 16822 17264
rect 17221 17255 17279 17261
rect 17221 17252 17233 17255
rect 16816 17224 17233 17252
rect 16816 17212 16822 17224
rect 17221 17221 17233 17224
rect 17267 17221 17279 17255
rect 17221 17215 17279 17221
rect 16577 17187 16635 17193
rect 16577 17153 16589 17187
rect 16623 17153 16635 17187
rect 21376 17184 21404 17283
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 16577 17147 16635 17153
rect 16684 17156 20300 17184
rect 21376 17156 21557 17184
rect 16684 17128 16712 17156
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17116 14243 17119
rect 14366 17116 14372 17128
rect 14231 17088 14372 17116
rect 14231 17085 14243 17088
rect 14185 17079 14243 17085
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 15470 17116 15476 17128
rect 15431 17088 15476 17116
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 20272 17125 20300 17156
rect 21545 17153 21557 17156
rect 21591 17153 21603 17187
rect 21545 17147 21603 17153
rect 24946 17144 24952 17196
rect 25004 17184 25010 17196
rect 25222 17184 25228 17196
rect 25004 17156 25228 17184
rect 25004 17144 25010 17156
rect 25222 17144 25228 17156
rect 25280 17184 25286 17196
rect 25409 17187 25467 17193
rect 25409 17184 25421 17187
rect 25280 17156 25421 17184
rect 25280 17144 25286 17156
rect 25409 17153 25421 17156
rect 25455 17153 25467 17187
rect 25409 17147 25467 17153
rect 20165 17119 20223 17125
rect 16724 17088 16769 17116
rect 16724 17076 16730 17088
rect 20165 17085 20177 17119
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 20257 17119 20315 17125
rect 20257 17085 20269 17119
rect 20303 17116 20315 17119
rect 21637 17119 21695 17125
rect 21637 17116 21649 17119
rect 20303 17088 21649 17116
rect 20303 17085 20315 17088
rect 20257 17079 20315 17085
rect 21637 17085 21649 17088
rect 21683 17116 21695 17119
rect 22370 17116 22376 17128
rect 21683 17088 22376 17116
rect 21683 17085 21695 17088
rect 21637 17079 21695 17085
rect 15194 17048 15200 17060
rect 11440 17020 15200 17048
rect 10468 17008 10474 17020
rect 15194 17008 15200 17020
rect 15252 17008 15258 17060
rect 2961 16983 3019 16989
rect 2961 16949 2973 16983
rect 3007 16980 3019 16983
rect 3050 16980 3056 16992
rect 3007 16952 3056 16980
rect 3007 16949 3019 16952
rect 2961 16943 3019 16949
rect 3050 16940 3056 16952
rect 3108 16940 3114 16992
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 8938 16980 8944 16992
rect 4120 16952 8944 16980
rect 4120 16940 4126 16952
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 12526 16980 12532 16992
rect 12487 16952 12532 16980
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 15562 16980 15568 16992
rect 15523 16952 15568 16980
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 20180 16980 20208 17079
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 25314 17076 25320 17128
rect 25372 17116 25378 17128
rect 25593 17119 25651 17125
rect 25593 17116 25605 17119
rect 25372 17088 25605 17116
rect 25372 17076 25378 17088
rect 25593 17085 25605 17088
rect 25639 17116 25651 17119
rect 26145 17119 26203 17125
rect 26145 17116 26157 17119
rect 25639 17088 26157 17116
rect 25639 17085 25651 17088
rect 25593 17079 25651 17085
rect 26145 17085 26157 17088
rect 26191 17085 26203 17119
rect 26326 17116 26332 17128
rect 26239 17088 26332 17116
rect 26145 17079 26203 17085
rect 26326 17076 26332 17088
rect 26384 17116 26390 17128
rect 27246 17116 27252 17128
rect 26384 17088 27252 17116
rect 26384 17076 26390 17088
rect 27246 17076 27252 17088
rect 27304 17076 27310 17128
rect 20717 17051 20775 17057
rect 20717 17017 20729 17051
rect 20763 17048 20775 17051
rect 21082 17048 21088 17060
rect 20763 17020 21088 17048
rect 20763 17017 20775 17020
rect 20717 17011 20775 17017
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 24670 17048 24676 17060
rect 21192 17020 24676 17048
rect 20901 16983 20959 16989
rect 20901 16980 20913 16983
rect 20180 16952 20913 16980
rect 20901 16949 20913 16952
rect 20947 16980 20959 16983
rect 21192 16980 21220 17020
rect 24670 17008 24676 17020
rect 24728 17008 24734 17060
rect 26697 17051 26755 17057
rect 26697 17017 26709 17051
rect 26743 17048 26755 17051
rect 26786 17048 26792 17060
rect 26743 17020 26792 17048
rect 26743 17017 26755 17020
rect 26697 17011 26755 17017
rect 26786 17008 26792 17020
rect 26844 17008 26850 17060
rect 20947 16952 21220 16980
rect 20947 16949 20959 16952
rect 20901 16943 20959 16949
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 22554 16980 22560 16992
rect 21784 16952 22560 16980
rect 21784 16940 21790 16952
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 25222 16980 25228 16992
rect 25183 16952 25228 16980
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 1104 16890 29256 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 29256 16890
rect 1104 16816 29256 16838
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 4154 16776 4160 16788
rect 3099 16748 4160 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 5350 16776 5356 16788
rect 4304 16748 4349 16776
rect 5311 16748 5356 16776
rect 4304 16736 4310 16748
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 13173 16779 13231 16785
rect 13173 16776 13185 16779
rect 12452 16748 13185 16776
rect 4264 16708 4292 16736
rect 7374 16708 7380 16720
rect 4264 16680 7380 16708
rect 7374 16668 7380 16680
rect 7432 16708 7438 16720
rect 9214 16708 9220 16720
rect 7432 16680 9220 16708
rect 7432 16668 7438 16680
rect 9214 16668 9220 16680
rect 9272 16668 9278 16720
rect 9490 16708 9496 16720
rect 9403 16680 9496 16708
rect 9490 16668 9496 16680
rect 9548 16708 9554 16720
rect 9548 16680 10548 16708
rect 9548 16668 9554 16680
rect 10520 16652 10548 16680
rect 10612 16680 11376 16708
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16609 2927 16643
rect 2869 16603 2927 16609
rect 2777 16439 2835 16445
rect 2777 16405 2789 16439
rect 2823 16436 2835 16439
rect 2884 16436 2912 16603
rect 3694 16600 3700 16652
rect 3752 16640 3758 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3752 16612 4077 16640
rect 3752 16600 3758 16612
rect 4065 16609 4077 16612
rect 4111 16640 4123 16643
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 4111 16612 4445 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16640 5227 16643
rect 5258 16640 5264 16652
rect 5215 16612 5264 16640
rect 5215 16609 5227 16612
rect 5169 16603 5227 16609
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10042 16640 10048 16652
rect 10003 16612 10048 16640
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 10134 16600 10140 16652
rect 10192 16640 10198 16652
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 10192 16612 10241 16640
rect 10192 16600 10198 16612
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10502 16640 10508 16652
rect 10463 16612 10508 16640
rect 10229 16603 10287 16609
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 10612 16649 10640 16680
rect 11348 16652 11376 16680
rect 10597 16643 10655 16649
rect 10597 16609 10609 16643
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 11330 16640 11336 16652
rect 10744 16612 11008 16640
rect 11291 16612 11336 16640
rect 10744 16600 10750 16612
rect 10980 16581 11008 16612
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11422 16600 11428 16652
rect 11480 16640 11486 16652
rect 12452 16640 12480 16748
rect 13173 16745 13185 16748
rect 13219 16776 13231 16779
rect 13219 16748 13400 16776
rect 13219 16745 13231 16748
rect 13173 16739 13231 16745
rect 13372 16708 13400 16748
rect 15102 16736 15108 16788
rect 15160 16776 15166 16788
rect 17494 16776 17500 16788
rect 15160 16748 16712 16776
rect 17455 16748 17500 16776
rect 15160 16736 15166 16748
rect 14366 16708 14372 16720
rect 13372 16680 14372 16708
rect 13262 16640 13268 16652
rect 11480 16612 12480 16640
rect 13223 16612 13268 16640
rect 11480 16600 11486 16612
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13372 16649 13400 16680
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 15194 16668 15200 16720
rect 15252 16708 15258 16720
rect 16482 16708 16488 16720
rect 15252 16680 16488 16708
rect 15252 16668 15258 16680
rect 16482 16668 16488 16680
rect 16540 16708 16546 16720
rect 16540 16680 16620 16708
rect 16540 16668 16546 16680
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16609 13415 16643
rect 15841 16643 15899 16649
rect 15841 16640 15853 16643
rect 13357 16603 13415 16609
rect 13464 16612 15853 16640
rect 10965 16575 11023 16581
rect 10965 16541 10977 16575
rect 11011 16541 11023 16575
rect 10965 16535 11023 16541
rect 12342 16532 12348 16584
rect 12400 16572 12406 16584
rect 13464 16572 13492 16612
rect 15841 16609 15853 16612
rect 15887 16609 15899 16643
rect 16390 16640 16396 16652
rect 16351 16612 16396 16640
rect 15841 16603 15899 16609
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 16592 16649 16620 16680
rect 16684 16649 16712 16748
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 20625 16779 20683 16785
rect 20625 16776 20637 16779
rect 18012 16748 20637 16776
rect 18012 16736 18018 16748
rect 20625 16745 20637 16748
rect 20671 16776 20683 16779
rect 21910 16776 21916 16788
rect 20671 16748 21916 16776
rect 20671 16745 20683 16748
rect 20625 16739 20683 16745
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 22554 16776 22560 16788
rect 22515 16748 22560 16776
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 16669 16643 16727 16649
rect 16669 16609 16681 16643
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 17129 16643 17187 16649
rect 16816 16612 17080 16640
rect 16816 16600 16822 16612
rect 13814 16572 13820 16584
rect 12400 16544 13492 16572
rect 13775 16544 13820 16572
rect 12400 16532 12406 16544
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 14090 16532 14096 16584
rect 14148 16572 14154 16584
rect 14274 16572 14280 16584
rect 14148 16544 14280 16572
rect 14148 16532 14154 16544
rect 14274 16532 14280 16544
rect 14332 16572 14338 16584
rect 16942 16572 16948 16584
rect 14332 16544 16948 16572
rect 14332 16532 14338 16544
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17052 16572 17080 16612
rect 17129 16609 17141 16643
rect 17175 16640 17187 16643
rect 17512 16640 17540 16736
rect 19978 16708 19984 16720
rect 19812 16680 19984 16708
rect 19812 16649 19840 16680
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 17175 16612 17540 16640
rect 19797 16643 19855 16649
rect 17175 16609 17187 16612
rect 17129 16603 17187 16609
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 19889 16643 19947 16649
rect 19889 16609 19901 16643
rect 19935 16640 19947 16643
rect 20806 16640 20812 16652
rect 19935 16612 20812 16640
rect 19935 16609 19947 16612
rect 19889 16603 19947 16609
rect 20806 16600 20812 16612
rect 20864 16600 20870 16652
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21082 16640 21088 16652
rect 20956 16612 21001 16640
rect 21043 16612 21088 16640
rect 20956 16600 20962 16612
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21174 16600 21180 16652
rect 21232 16640 21238 16652
rect 21453 16643 21511 16649
rect 21453 16640 21465 16643
rect 21232 16612 21465 16640
rect 21232 16600 21238 16612
rect 21453 16609 21465 16612
rect 21499 16609 21511 16643
rect 21726 16640 21732 16652
rect 21687 16612 21732 16640
rect 21453 16603 21511 16609
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 21910 16640 21916 16652
rect 21871 16612 21916 16640
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16640 23259 16643
rect 24210 16640 24216 16652
rect 23247 16612 24216 16640
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 24210 16600 24216 16612
rect 24268 16600 24274 16652
rect 17221 16575 17279 16581
rect 17221 16572 17233 16575
rect 17052 16544 17233 16572
rect 17221 16541 17233 16544
rect 17267 16541 17279 16575
rect 32674 16572 32680 16584
rect 17221 16535 17279 16541
rect 17328 16544 32680 16572
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 16298 16504 16304 16516
rect 3936 16476 16304 16504
rect 3936 16464 3942 16476
rect 16298 16464 16304 16476
rect 16356 16464 16362 16516
rect 2958 16436 2964 16448
rect 2823 16408 2964 16436
rect 2823 16405 2835 16408
rect 2777 16399 2835 16405
rect 2958 16396 2964 16408
rect 3016 16396 3022 16448
rect 12250 16396 12256 16448
rect 12308 16436 12314 16448
rect 12897 16439 12955 16445
rect 12897 16436 12909 16439
rect 12308 16408 12909 16436
rect 12308 16396 12314 16408
rect 12897 16405 12909 16408
rect 12943 16436 12955 16439
rect 13262 16436 13268 16448
rect 12943 16408 13268 16436
rect 12943 16405 12955 16408
rect 12897 16399 12955 16405
rect 13262 16396 13268 16408
rect 13320 16436 13326 16448
rect 17328 16436 17356 16544
rect 32674 16532 32680 16544
rect 32732 16532 32738 16584
rect 17770 16464 17776 16516
rect 17828 16504 17834 16516
rect 32490 16504 32496 16516
rect 17828 16476 32496 16504
rect 17828 16464 17834 16476
rect 32490 16464 32496 16476
rect 32548 16464 32554 16516
rect 13320 16408 17356 16436
rect 13320 16396 13326 16408
rect 20622 16396 20628 16448
rect 20680 16436 20686 16448
rect 22281 16439 22339 16445
rect 22281 16436 22293 16439
rect 20680 16408 22293 16436
rect 20680 16396 20686 16408
rect 22281 16405 22293 16408
rect 22327 16405 22339 16439
rect 23290 16436 23296 16448
rect 23251 16408 23296 16436
rect 22281 16399 22339 16405
rect 23290 16396 23296 16408
rect 23348 16396 23354 16448
rect 1104 16346 29256 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 29256 16346
rect 1104 16272 29256 16294
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5994 16232 6000 16244
rect 5307 16204 6000 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 13170 16232 13176 16244
rect 13131 16204 13176 16232
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 21174 16232 21180 16244
rect 16080 16204 21180 16232
rect 16080 16192 16086 16204
rect 21174 16192 21180 16204
rect 21232 16232 21238 16244
rect 21634 16232 21640 16244
rect 21232 16204 21640 16232
rect 21232 16192 21238 16204
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 27246 16232 27252 16244
rect 27207 16204 27252 16232
rect 27246 16192 27252 16204
rect 27304 16192 27310 16244
rect 16298 16124 16304 16176
rect 16356 16164 16362 16176
rect 20070 16164 20076 16176
rect 16356 16136 20076 16164
rect 16356 16124 16362 16136
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 32582 16164 32588 16176
rect 20180 16136 32588 16164
rect 2590 16096 2596 16108
rect 2551 16068 2596 16096
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 2866 16096 2872 16108
rect 2827 16068 2872 16096
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16096 9275 16099
rect 12342 16096 12348 16108
rect 9263 16068 12348 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 12342 16056 12348 16068
rect 12400 16056 12406 16108
rect 12526 16056 12532 16108
rect 12584 16096 12590 16108
rect 13633 16099 13691 16105
rect 13633 16096 13645 16099
rect 12584 16068 13645 16096
rect 12584 16056 12590 16068
rect 13633 16065 13645 16068
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 13964 16068 14197 16096
rect 13964 16056 13970 16068
rect 14185 16065 14197 16068
rect 14231 16096 14243 16099
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 14231 16068 15669 16096
rect 14231 16065 14243 16068
rect 14185 16059 14243 16065
rect 15657 16065 15669 16068
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 5074 16028 5080 16040
rect 5035 16000 5080 16028
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 7006 16028 7012 16040
rect 6967 16000 7012 16028
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 9306 15988 9312 16040
rect 9364 16028 9370 16040
rect 9401 16031 9459 16037
rect 9401 16028 9413 16031
rect 9364 16000 9413 16028
rect 9364 15988 9370 16000
rect 9401 15997 9413 16000
rect 9447 15997 9459 16031
rect 9766 16028 9772 16040
rect 9727 16000 9772 16028
rect 9401 15991 9459 15997
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 6825 15963 6883 15969
rect 6825 15929 6837 15963
rect 6871 15960 6883 15963
rect 7282 15960 7288 15972
rect 6871 15932 7288 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 7282 15920 7288 15932
rect 7340 15920 7346 15972
rect 3970 15892 3976 15904
rect 3931 15864 3976 15892
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 4246 15852 4252 15904
rect 4304 15892 4310 15904
rect 4341 15895 4399 15901
rect 4341 15892 4353 15895
rect 4304 15864 4353 15892
rect 4304 15852 4310 15864
rect 4341 15861 4353 15864
rect 4387 15861 4399 15895
rect 4341 15855 4399 15861
rect 6730 15852 6736 15904
rect 6788 15892 6794 15904
rect 7101 15895 7159 15901
rect 7101 15892 7113 15895
rect 6788 15864 7113 15892
rect 6788 15852 6794 15864
rect 7101 15861 7113 15864
rect 7147 15861 7159 15895
rect 7101 15855 7159 15861
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8812 15864 9137 15892
rect 8812 15852 8818 15864
rect 9125 15861 9137 15864
rect 9171 15892 9183 15895
rect 9968 15892 9996 15991
rect 10152 15960 10180 15991
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 10689 16031 10747 16037
rect 10689 16028 10701 16031
rect 10652 16000 10701 16028
rect 10652 15988 10658 16000
rect 10689 15997 10701 16000
rect 10735 15997 10747 16031
rect 10689 15991 10747 15997
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 12768 16000 13737 16028
rect 12768 15988 12774 16000
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 14090 16028 14096 16040
rect 14051 16000 14096 16028
rect 13725 15991 13783 15997
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 15102 16028 15108 16040
rect 15063 16000 15108 16028
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 15252 16000 15297 16028
rect 15252 15988 15258 16000
rect 10873 15963 10931 15969
rect 10873 15960 10885 15963
rect 10152 15932 10885 15960
rect 10873 15929 10885 15932
rect 10919 15960 10931 15963
rect 11330 15960 11336 15972
rect 10919 15932 11336 15960
rect 10919 15929 10931 15932
rect 10873 15923 10931 15929
rect 11330 15920 11336 15932
rect 11388 15960 11394 15972
rect 17126 15960 17132 15972
rect 11388 15932 17132 15960
rect 11388 15920 11394 15932
rect 17126 15920 17132 15932
rect 17184 15920 17190 15972
rect 20180 15892 20208 16136
rect 32582 16124 32588 16136
rect 32640 16124 32646 16176
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 21177 16099 21235 16105
rect 21177 16096 21189 16099
rect 20864 16068 21189 16096
rect 20864 16056 20870 16068
rect 21177 16065 21189 16068
rect 21223 16065 21235 16099
rect 22002 16096 22008 16108
rect 21177 16059 21235 16065
rect 21560 16068 22008 16096
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 16028 20775 16031
rect 20990 16028 20996 16040
rect 20763 16000 20996 16028
rect 20763 15997 20775 16000
rect 20717 15991 20775 15997
rect 20990 15988 20996 16000
rect 21048 15988 21054 16040
rect 21560 16037 21588 16068
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 21545 16031 21603 16037
rect 21545 15997 21557 16031
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 21729 16031 21787 16037
rect 21729 16028 21741 16031
rect 21692 16000 21741 16028
rect 21692 15988 21698 16000
rect 21729 15997 21741 16000
rect 21775 15997 21787 16031
rect 21910 16028 21916 16040
rect 21871 16000 21916 16028
rect 21729 15991 21787 15997
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 22189 16031 22247 16037
rect 22189 15997 22201 16031
rect 22235 16028 22247 16031
rect 22554 16028 22560 16040
rect 22235 16000 22560 16028
rect 22235 15997 22247 16000
rect 22189 15991 22247 15997
rect 20530 15960 20536 15972
rect 20443 15932 20536 15960
rect 20530 15920 20536 15932
rect 20588 15960 20594 15972
rect 21928 15960 21956 15988
rect 20588 15932 21956 15960
rect 20588 15920 20594 15932
rect 22002 15920 22008 15972
rect 22060 15960 22066 15972
rect 22204 15960 22232 15991
rect 22554 15988 22560 16000
rect 22612 15988 22618 16040
rect 23658 16028 23664 16040
rect 23619 16000 23664 16028
rect 23658 15988 23664 16000
rect 23716 15988 23722 16040
rect 27157 16031 27215 16037
rect 27157 15997 27169 16031
rect 27203 16028 27215 16031
rect 27203 16000 27568 16028
rect 27203 15997 27215 16000
rect 27157 15991 27215 15997
rect 22060 15932 22232 15960
rect 22060 15920 22066 15932
rect 27540 15904 27568 16000
rect 20806 15892 20812 15904
rect 9171 15864 20208 15892
rect 20767 15864 20812 15892
rect 9171 15861 9183 15864
rect 9125 15855 9183 15861
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22557 15895 22615 15901
rect 22557 15892 22569 15895
rect 22152 15864 22569 15892
rect 22152 15852 22158 15864
rect 22557 15861 22569 15864
rect 22603 15861 22615 15895
rect 22557 15855 22615 15861
rect 22922 15852 22928 15904
rect 22980 15892 22986 15904
rect 23753 15895 23811 15901
rect 23753 15892 23765 15895
rect 22980 15864 23765 15892
rect 22980 15852 22986 15864
rect 23753 15861 23765 15864
rect 23799 15861 23811 15895
rect 27522 15892 27528 15904
rect 27483 15864 27528 15892
rect 23753 15855 23811 15861
rect 27522 15852 27528 15864
rect 27580 15852 27586 15904
rect 1104 15802 29256 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 29256 15802
rect 1104 15728 29256 15750
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 4120 15660 5457 15688
rect 4120 15648 4126 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6362 15688 6368 15700
rect 5592 15660 6368 15688
rect 5592 15648 5598 15660
rect 6362 15648 6368 15660
rect 6420 15688 6426 15700
rect 8754 15688 8760 15700
rect 6420 15660 6592 15688
rect 8715 15660 8760 15688
rect 6420 15648 6426 15660
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4706 15552 4712 15564
rect 4387 15524 4712 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4706 15512 4712 15524
rect 4764 15552 4770 15564
rect 6564 15561 6592 15660
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 11422 15688 11428 15700
rect 10183 15660 11428 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 6730 15620 6736 15632
rect 6691 15592 6736 15620
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 4764 15524 5825 15552
rect 4764 15512 4770 15524
rect 5813 15521 5825 15524
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15552 8447 15555
rect 8772 15552 8800 15648
rect 8435 15524 8800 15552
rect 9677 15555 9735 15561
rect 8435 15521 8447 15524
rect 8389 15515 8447 15521
rect 9677 15521 9689 15555
rect 9723 15552 9735 15555
rect 9858 15552 9864 15564
rect 9723 15524 9864 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 2648 15456 4077 15484
rect 2648 15444 2654 15456
rect 4065 15453 4077 15456
rect 4111 15484 4123 15487
rect 4246 15484 4252 15496
rect 4111 15456 4252 15484
rect 4111 15453 4123 15456
rect 4065 15447 4123 15453
rect 4246 15444 4252 15456
rect 4304 15484 4310 15496
rect 4522 15484 4528 15496
rect 4304 15456 4528 15484
rect 4304 15444 4310 15456
rect 4522 15444 4528 15456
rect 4580 15484 4586 15496
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 4580 15456 6009 15484
rect 4580 15444 4586 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 6840 15484 6868 15515
rect 9858 15512 9864 15524
rect 9916 15552 9922 15564
rect 10152 15552 10180 15651
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 12710 15688 12716 15700
rect 12671 15660 12716 15688
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 15381 15691 15439 15697
rect 15381 15688 15393 15691
rect 14424 15660 15393 15688
rect 14424 15648 14430 15660
rect 15381 15657 15393 15660
rect 15427 15688 15439 15691
rect 15427 15660 16988 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 13630 15620 13636 15632
rect 13591 15592 13636 15620
rect 13630 15580 13636 15592
rect 13688 15580 13694 15632
rect 16850 15620 16856 15632
rect 15856 15592 16856 15620
rect 9916 15524 10180 15552
rect 9916 15512 9922 15524
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 13814 15561 13820 15564
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12492 15524 12633 15552
rect 12492 15512 12498 15524
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 13780 15555 13820 15561
rect 13780 15521 13792 15555
rect 13780 15515 13820 15521
rect 13814 15512 13820 15515
rect 13872 15512 13878 15564
rect 15473 15555 15531 15561
rect 13924 15524 15424 15552
rect 6840 15456 11928 15484
rect 5997 15447 6055 15453
rect 6178 15376 6184 15428
rect 6236 15416 6242 15428
rect 9861 15419 9919 15425
rect 6236 15388 7052 15416
rect 6236 15376 6242 15388
rect 7024 15357 7052 15388
rect 9861 15385 9873 15419
rect 9907 15416 9919 15419
rect 11330 15416 11336 15428
rect 9907 15388 11336 15416
rect 9907 15385 9919 15388
rect 9861 15379 9919 15385
rect 11330 15376 11336 15388
rect 11388 15376 11394 15428
rect 11900 15416 11928 15456
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 13924 15484 13952 15524
rect 13596 15456 13952 15484
rect 14001 15487 14059 15493
rect 13596 15444 13602 15456
rect 14001 15453 14013 15487
rect 14047 15484 14059 15487
rect 14458 15484 14464 15496
rect 14047 15456 14464 15484
rect 14047 15453 14059 15456
rect 14001 15447 14059 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 15396 15484 15424 15524
rect 15473 15521 15485 15555
rect 15519 15552 15531 15555
rect 15562 15552 15568 15564
rect 15519 15524 15568 15552
rect 15519 15521 15531 15524
rect 15473 15515 15531 15521
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 15856 15561 15884 15592
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 15841 15555 15899 15561
rect 15841 15521 15853 15555
rect 15887 15521 15899 15555
rect 16022 15552 16028 15564
rect 15935 15524 16028 15552
rect 15841 15515 15899 15521
rect 16022 15512 16028 15524
rect 16080 15512 16086 15564
rect 16206 15552 16212 15564
rect 16167 15524 16212 15552
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15552 16543 15555
rect 16960 15552 16988 15660
rect 17126 15648 17132 15700
rect 17184 15688 17190 15700
rect 20993 15691 21051 15697
rect 20993 15688 21005 15691
rect 17184 15660 21005 15688
rect 17184 15648 17190 15660
rect 20993 15657 21005 15660
rect 21039 15688 21051 15691
rect 21082 15688 21088 15700
rect 21039 15660 21088 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 21082 15648 21088 15660
rect 21140 15688 21146 15700
rect 21453 15691 21511 15697
rect 21453 15688 21465 15691
rect 21140 15660 21465 15688
rect 21140 15648 21146 15660
rect 21453 15657 21465 15660
rect 21499 15688 21511 15691
rect 22002 15688 22008 15700
rect 21499 15660 22008 15688
rect 21499 15657 21511 15660
rect 21453 15651 21511 15657
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 24118 15648 24124 15700
rect 24176 15688 24182 15700
rect 24673 15691 24731 15697
rect 24673 15688 24685 15691
rect 24176 15660 24685 15688
rect 24176 15648 24182 15660
rect 24673 15657 24685 15660
rect 24719 15657 24731 15691
rect 26234 15688 26240 15700
rect 26195 15660 26240 15688
rect 24673 15651 24731 15657
rect 21634 15580 21640 15632
rect 21692 15620 21698 15632
rect 21692 15592 22232 15620
rect 21692 15580 21698 15592
rect 17954 15552 17960 15564
rect 16531 15524 17960 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 21818 15552 21824 15564
rect 21779 15524 21824 15552
rect 21818 15512 21824 15524
rect 21876 15512 21882 15564
rect 22204 15561 22232 15592
rect 22388 15592 23428 15620
rect 22388 15561 22416 15592
rect 22189 15555 22247 15561
rect 22189 15521 22201 15555
rect 22235 15521 22247 15555
rect 22189 15515 22247 15521
rect 22373 15555 22431 15561
rect 22373 15521 22385 15555
rect 22419 15521 22431 15555
rect 22554 15552 22560 15564
rect 22515 15524 22560 15552
rect 22373 15515 22431 15521
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 16040 15484 16068 15512
rect 15396 15456 16068 15484
rect 16224 15484 16252 15512
rect 17037 15487 17095 15493
rect 17037 15484 17049 15487
rect 16224 15456 17049 15484
rect 17037 15453 17049 15456
rect 17083 15453 17095 15487
rect 17037 15447 17095 15453
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 23290 15484 23296 15496
rect 21683 15456 23296 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 14093 15419 14151 15425
rect 14093 15416 14105 15419
rect 11900 15388 14105 15416
rect 14093 15385 14105 15388
rect 14139 15385 14151 15419
rect 14093 15379 14151 15385
rect 15194 15376 15200 15428
rect 15252 15416 15258 15428
rect 23017 15419 23075 15425
rect 23017 15416 23029 15419
rect 15252 15388 23029 15416
rect 15252 15376 15258 15388
rect 23017 15385 23029 15388
rect 23063 15385 23075 15419
rect 23017 15379 23075 15385
rect 23201 15419 23259 15425
rect 23201 15385 23213 15419
rect 23247 15416 23259 15419
rect 23400 15416 23428 15592
rect 24688 15552 24716 15651
rect 26234 15648 26240 15660
rect 26292 15648 26298 15700
rect 24857 15555 24915 15561
rect 24857 15552 24869 15555
rect 24688 15524 24869 15552
rect 24857 15521 24869 15524
rect 24903 15521 24915 15555
rect 26252 15552 26280 15648
rect 27522 15580 27528 15632
rect 27580 15620 27586 15632
rect 28169 15623 28227 15629
rect 28169 15620 28181 15623
rect 27580 15592 28181 15620
rect 27580 15580 27586 15592
rect 28169 15589 28181 15592
rect 28215 15620 28227 15623
rect 32398 15620 32404 15632
rect 28215 15592 32404 15620
rect 28215 15589 28227 15592
rect 28169 15583 28227 15589
rect 32398 15580 32404 15592
rect 32456 15580 32462 15632
rect 26513 15555 26571 15561
rect 26513 15552 26525 15555
rect 26252 15524 26525 15552
rect 24857 15515 24915 15521
rect 26513 15521 26525 15524
rect 26559 15521 26571 15555
rect 26786 15552 26792 15564
rect 26747 15524 26792 15552
rect 26513 15515 26571 15521
rect 26786 15512 26792 15524
rect 26844 15512 26850 15564
rect 24854 15416 24860 15428
rect 23247 15388 24860 15416
rect 23247 15385 23259 15388
rect 23201 15379 23259 15385
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 7009 15351 7067 15357
rect 7009 15317 7021 15351
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 7984 15320 8493 15348
rect 7984 15308 7990 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 8481 15311 8539 15317
rect 13909 15351 13967 15357
rect 13909 15317 13921 15351
rect 13955 15348 13967 15351
rect 14182 15348 14188 15360
rect 13955 15320 14188 15348
rect 13955 15317 13967 15320
rect 13909 15311 13967 15317
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 16850 15348 16856 15360
rect 16811 15320 16856 15348
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 25041 15351 25099 15357
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 25682 15348 25688 15360
rect 25087 15320 25688 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 25682 15308 25688 15320
rect 25740 15308 25746 15360
rect 1104 15258 29256 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 29256 15258
rect 1104 15184 29256 15206
rect 58434 15172 58440 15224
rect 58492 15212 58498 15224
rect 59354 15212 59360 15224
rect 58492 15184 59360 15212
rect 58492 15172 58498 15184
rect 59354 15172 59360 15184
rect 59412 15172 59418 15224
rect 4890 15104 4896 15156
rect 4948 15144 4954 15156
rect 25498 15144 25504 15156
rect 4948 15116 25504 15144
rect 4948 15104 4954 15116
rect 25498 15104 25504 15116
rect 25556 15104 25562 15156
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 4341 15079 4399 15085
rect 4341 15076 4353 15079
rect 3844 15048 4353 15076
rect 3844 15036 3850 15048
rect 4341 15045 4353 15048
rect 4387 15045 4399 15079
rect 4614 15076 4620 15088
rect 4575 15048 4620 15076
rect 4341 15039 4399 15045
rect 4614 15036 4620 15048
rect 4672 15076 4678 15088
rect 4672 15048 7604 15076
rect 4672 15036 4678 15048
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3804 15008 3832 15036
rect 7576 15017 7604 15048
rect 8754 15036 8760 15088
rect 8812 15076 8818 15088
rect 8941 15079 8999 15085
rect 8941 15076 8953 15079
rect 8812 15048 8953 15076
rect 8812 15036 8818 15048
rect 8941 15045 8953 15048
rect 8987 15045 8999 15079
rect 8941 15039 8999 15045
rect 2915 14980 3832 15008
rect 7561 15011 7619 15017
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 7561 14977 7573 15011
rect 7607 15008 7619 15011
rect 9309 15011 9367 15017
rect 9309 15008 9321 15011
rect 7607 14980 9321 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 9309 14977 9321 14980
rect 9355 14977 9367 15011
rect 9309 14971 9367 14977
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19705 15011 19763 15017
rect 19705 15008 19717 15011
rect 19392 14980 19717 15008
rect 19392 14968 19398 14980
rect 19705 14977 19717 14980
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20772 14980 21097 15008
rect 20772 14968 20778 14980
rect 21085 14977 21097 14980
rect 21131 15008 21143 15011
rect 21726 15008 21732 15020
rect 21131 14980 21732 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21726 14968 21732 14980
rect 21784 14968 21790 15020
rect 24762 14968 24768 15020
rect 24820 15008 24826 15020
rect 25409 15011 25467 15017
rect 25409 15008 25421 15011
rect 24820 14980 25421 15008
rect 24820 14968 24826 14980
rect 25409 14977 25421 14980
rect 25455 15008 25467 15011
rect 25501 15011 25559 15017
rect 25501 15008 25513 15011
rect 25455 14980 25513 15008
rect 25455 14977 25467 14980
rect 25409 14971 25467 14977
rect 25501 14977 25513 14980
rect 25547 14977 25559 15011
rect 27801 15011 27859 15017
rect 27801 15008 27813 15011
rect 25501 14971 25559 14977
rect 26620 14980 27813 15008
rect 7834 14940 7840 14952
rect 7795 14912 7840 14940
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12986 14940 12992 14952
rect 12207 14912 12992 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14940 13139 14943
rect 13906 14940 13912 14952
rect 13127 14912 13912 14940
rect 13127 14909 13139 14912
rect 13081 14903 13139 14909
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14909 14243 14943
rect 14366 14940 14372 14952
rect 14327 14912 14372 14940
rect 14185 14903 14243 14909
rect 14200 14816 14228 14903
rect 14366 14900 14372 14912
rect 14424 14940 14430 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 14424 14912 14933 14940
rect 14424 14900 14430 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 14921 14903 14979 14909
rect 15105 14943 15163 14949
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15654 14940 15660 14952
rect 15151 14912 15660 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 19352 14912 19441 14940
rect 3970 14804 3976 14816
rect 3931 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11977 14807 12035 14813
rect 11977 14804 11989 14807
rect 11020 14776 11989 14804
rect 11020 14764 11026 14776
rect 11977 14773 11989 14776
rect 12023 14804 12035 14807
rect 12710 14804 12716 14816
rect 12023 14776 12716 14804
rect 12023 14773 12035 14776
rect 11977 14767 12035 14773
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 13538 14804 13544 14816
rect 13311 14776 13544 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14093 14807 14151 14813
rect 14093 14773 14105 14807
rect 14139 14804 14151 14807
rect 14182 14804 14188 14816
rect 14139 14776 14188 14804
rect 14139 14773 14151 14776
rect 14093 14767 14151 14773
rect 14182 14764 14188 14776
rect 14240 14804 14246 14816
rect 14918 14804 14924 14816
rect 14240 14776 14924 14804
rect 14240 14764 14246 14776
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 15010 14764 15016 14816
rect 15068 14804 15074 14816
rect 15381 14807 15439 14813
rect 15381 14804 15393 14807
rect 15068 14776 15393 14804
rect 15068 14764 15074 14776
rect 15381 14773 15393 14776
rect 15427 14773 15439 14807
rect 15381 14767 15439 14773
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 17862 14804 17868 14816
rect 16724 14776 17868 14804
rect 16724 14764 16730 14776
rect 17862 14764 17868 14776
rect 17920 14804 17926 14816
rect 19352 14813 19380 14912
rect 19429 14909 19441 14912
rect 19475 14909 19487 14943
rect 25682 14940 25688 14952
rect 25643 14912 25688 14940
rect 19429 14903 19487 14909
rect 25682 14900 25688 14912
rect 25740 14900 25746 14952
rect 26237 14943 26295 14949
rect 26237 14909 26249 14943
rect 26283 14909 26295 14943
rect 26237 14903 26295 14909
rect 26421 14943 26479 14949
rect 26421 14909 26433 14943
rect 26467 14940 26479 14943
rect 26620 14940 26648 14980
rect 27801 14977 27813 14980
rect 27847 14977 27859 15011
rect 27801 14971 27859 14977
rect 26467 14912 26648 14940
rect 27709 14943 27767 14949
rect 26467 14909 26479 14912
rect 26421 14903 26479 14909
rect 27709 14909 27721 14943
rect 27755 14940 27767 14943
rect 29086 14940 29092 14952
rect 27755 14912 29092 14940
rect 27755 14909 27767 14912
rect 27709 14903 27767 14909
rect 25700 14872 25728 14900
rect 26252 14872 26280 14903
rect 29086 14900 29092 14912
rect 29144 14900 29150 14952
rect 26786 14872 26792 14884
rect 25700 14844 26280 14872
rect 26747 14844 26792 14872
rect 26786 14832 26792 14844
rect 26844 14832 26850 14884
rect 86218 14832 86224 14884
rect 86276 14872 86282 14884
rect 87138 14872 87144 14884
rect 86276 14844 87144 14872
rect 86276 14832 86282 14844
rect 87138 14832 87144 14844
rect 87196 14832 87202 14884
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 17920 14776 19349 14804
rect 17920 14764 17926 14776
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 19337 14767 19395 14773
rect 1104 14714 29256 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 29256 14714
rect 1104 14640 29256 14662
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9548 14572 9965 14600
rect 9548 14560 9554 14572
rect 9769 14535 9827 14541
rect 9769 14532 9781 14535
rect 7944 14504 9781 14532
rect 7190 14464 7196 14476
rect 7151 14436 7196 14464
rect 7190 14424 7196 14436
rect 7248 14464 7254 14476
rect 7944 14473 7972 14504
rect 9769 14501 9781 14504
rect 9815 14501 9827 14535
rect 9769 14495 9827 14501
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7248 14436 7757 14464
rect 7248 14424 7254 14436
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14433 7987 14467
rect 7929 14427 7987 14433
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 9876 14464 9904 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 12897 14603 12955 14609
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 14366 14600 14372 14612
rect 12943 14572 14372 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 15933 14603 15991 14609
rect 15933 14569 15945 14603
rect 15979 14600 15991 14603
rect 16206 14600 16212 14612
rect 15979 14572 16212 14600
rect 15979 14569 15991 14572
rect 15933 14563 15991 14569
rect 9723 14436 9904 14464
rect 11517 14467 11575 14473
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 11517 14433 11529 14467
rect 11563 14464 11575 14467
rect 12618 14464 12624 14476
rect 11563 14436 12624 14464
rect 11563 14433 11575 14436
rect 11517 14427 11575 14433
rect 12618 14424 12624 14436
rect 12676 14464 12682 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12676 14436 12725 14464
rect 12676 14424 12682 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 13906 14464 13912 14476
rect 13867 14436 13912 14464
rect 12713 14427 12771 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 14369 14467 14427 14473
rect 14369 14433 14381 14467
rect 14415 14464 14427 14467
rect 14458 14464 14464 14476
rect 14415 14436 14464 14464
rect 14415 14433 14427 14436
rect 14369 14427 14427 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14464 15623 14467
rect 15948 14464 15976 14563
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 20165 14603 20223 14609
rect 20165 14569 20177 14603
rect 20211 14600 20223 14603
rect 20714 14600 20720 14612
rect 20211 14572 20720 14600
rect 20211 14569 20223 14572
rect 20165 14563 20223 14569
rect 15611 14436 15976 14464
rect 19797 14467 19855 14473
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 19797 14433 19809 14467
rect 19843 14464 19855 14467
rect 20180 14464 20208 14563
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 26234 14600 26240 14612
rect 26195 14572 26240 14600
rect 26234 14560 26240 14572
rect 26292 14560 26298 14612
rect 22922 14532 22928 14544
rect 22204 14504 22928 14532
rect 19843 14436 20208 14464
rect 21913 14467 21971 14473
rect 19843 14433 19855 14436
rect 19797 14427 19855 14433
rect 21913 14433 21925 14467
rect 21959 14464 21971 14467
rect 22204 14464 22232 14504
rect 22922 14492 22928 14504
rect 22980 14492 22986 14544
rect 21959 14436 22232 14464
rect 22281 14467 22339 14473
rect 21959 14433 21971 14436
rect 21913 14427 21971 14433
rect 22281 14433 22293 14467
rect 22327 14464 22339 14467
rect 26252 14464 26280 14560
rect 28169 14535 28227 14541
rect 28169 14501 28181 14535
rect 28215 14532 28227 14535
rect 29086 14532 29092 14544
rect 28215 14504 29092 14532
rect 28215 14501 28227 14504
rect 28169 14495 28227 14501
rect 29086 14492 29092 14504
rect 29144 14492 29150 14544
rect 26513 14467 26571 14473
rect 26513 14464 26525 14467
rect 22327 14436 22692 14464
rect 26252 14436 26525 14464
rect 22327 14433 22339 14436
rect 22281 14427 22339 14433
rect 7009 14399 7067 14405
rect 7009 14365 7021 14399
rect 7055 14365 7067 14399
rect 13814 14396 13820 14408
rect 13775 14368 13820 14396
rect 7009 14359 7067 14365
rect 7024 14272 7052 14359
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 21821 14399 21879 14405
rect 21821 14396 21833 14399
rect 21508 14368 21833 14396
rect 21508 14356 21514 14368
rect 21821 14365 21833 14368
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 22002 14356 22008 14408
rect 22060 14396 22066 14408
rect 22373 14399 22431 14405
rect 22373 14396 22385 14399
rect 22060 14368 22385 14396
rect 22060 14356 22066 14368
rect 22373 14365 22385 14368
rect 22419 14365 22431 14399
rect 22373 14359 22431 14365
rect 8110 14328 8116 14340
rect 8071 14300 8116 14328
rect 8110 14288 8116 14300
rect 8168 14288 8174 14340
rect 16942 14288 16948 14340
rect 17000 14328 17006 14340
rect 21361 14331 21419 14337
rect 21361 14328 21373 14331
rect 17000 14300 21373 14328
rect 17000 14288 17006 14300
rect 21361 14297 21373 14300
rect 21407 14297 21419 14331
rect 21361 14291 21419 14297
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14260 6975 14263
rect 7006 14260 7012 14272
rect 6963 14232 7012 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12526 14260 12532 14272
rect 11747 14232 12532 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 19058 14220 19064 14272
rect 19116 14260 19122 14272
rect 22664 14269 22692 14436
rect 26513 14433 26525 14436
rect 26559 14433 26571 14467
rect 26786 14464 26792 14476
rect 26747 14436 26792 14464
rect 26513 14427 26571 14433
rect 26786 14424 26792 14436
rect 26844 14424 26850 14476
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19116 14232 19901 14260
rect 19116 14220 19122 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 19889 14223 19947 14229
rect 22649 14263 22707 14269
rect 22649 14229 22661 14263
rect 22695 14260 22707 14263
rect 24026 14260 24032 14272
rect 22695 14232 24032 14260
rect 22695 14229 22707 14232
rect 22649 14223 22707 14229
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 1104 14170 29256 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 29256 14170
rect 1104 14096 29256 14118
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 4798 14056 4804 14068
rect 4479 14028 4804 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13920 2927 13923
rect 4448 13920 4476 14019
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 16942 14056 16948 14068
rect 8260 14028 16948 14056
rect 8260 14016 8266 14028
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 19334 14056 19340 14068
rect 19295 14028 19340 14056
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 4614 13988 4620 14000
rect 4575 13960 4620 13988
rect 4614 13948 4620 13960
rect 4672 13988 4678 14000
rect 4672 13960 7880 13988
rect 4672 13948 4678 13960
rect 7852 13929 7880 13960
rect 12710 13948 12716 14000
rect 12768 13988 12774 14000
rect 14553 13991 14611 13997
rect 14553 13988 14565 13991
rect 12768 13960 14565 13988
rect 12768 13948 12774 13960
rect 14553 13957 14565 13960
rect 14599 13988 14611 13991
rect 18782 13988 18788 14000
rect 14599 13960 14780 13988
rect 14599 13957 14611 13960
rect 14553 13951 14611 13957
rect 2915 13892 4476 13920
rect 7837 13923 7895 13929
rect 2915 13889 2927 13892
rect 2869 13883 2927 13889
rect 7837 13889 7849 13923
rect 7883 13889 7895 13923
rect 8110 13920 8116 13932
rect 8071 13892 8116 13920
rect 7837 13883 7895 13889
rect 7852 13852 7880 13883
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 9490 13920 9496 13932
rect 9451 13892 9496 13920
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 14752 13929 14780 13960
rect 18156 13960 18788 13988
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 15010 13920 15016 13932
rect 14971 13892 15016 13920
rect 14737 13883 14795 13889
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 7852 13824 9597 13852
rect 9585 13821 9597 13824
rect 9631 13852 9643 13855
rect 10962 13852 10968 13864
rect 9631 13824 10968 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 14752 13852 14780 13883
rect 15010 13880 15016 13892
rect 15068 13880 15074 13932
rect 16206 13920 16212 13932
rect 16167 13892 16212 13920
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 17770 13852 17776 13864
rect 14752 13824 16436 13852
rect 17731 13824 17776 13852
rect 16408 13784 16436 13824
rect 17770 13812 17776 13824
rect 17828 13852 17834 13864
rect 18156 13861 18184 13960
rect 18782 13948 18788 13960
rect 18840 13948 18846 14000
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 23032 13892 23765 13920
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 17828 13824 18153 13852
rect 17828 13812 17834 13824
rect 18141 13821 18153 13824
rect 18187 13821 18199 13855
rect 18141 13815 18199 13821
rect 18325 13855 18383 13861
rect 18325 13821 18337 13855
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 18877 13855 18935 13861
rect 18877 13821 18889 13855
rect 18923 13821 18935 13855
rect 19058 13852 19064 13864
rect 19019 13824 19064 13852
rect 18877 13815 18935 13821
rect 16666 13784 16672 13796
rect 16408 13756 16672 13784
rect 16666 13744 16672 13756
rect 16724 13744 16730 13796
rect 16758 13744 16764 13796
rect 16816 13784 16822 13796
rect 18340 13784 18368 13815
rect 18892 13784 18920 13815
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 19260 13824 21189 13852
rect 16816 13756 18920 13784
rect 16816 13744 16822 13756
rect 3970 13716 3976 13728
rect 3931 13688 3976 13716
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 19150 13716 19156 13728
rect 4120 13688 19156 13716
rect 4120 13676 4126 13688
rect 19150 13676 19156 13688
rect 19208 13716 19214 13728
rect 19260 13716 19288 13824
rect 21177 13821 21189 13824
rect 21223 13852 21235 13855
rect 21358 13852 21364 13864
rect 21223 13824 21364 13852
rect 21223 13821 21235 13824
rect 21177 13815 21235 13821
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 21545 13855 21603 13861
rect 21545 13821 21557 13855
rect 21591 13821 21603 13855
rect 21545 13815 21603 13821
rect 22097 13855 22155 13861
rect 22097 13821 22109 13855
rect 22143 13821 22155 13855
rect 22097 13815 22155 13821
rect 22281 13855 22339 13861
rect 22281 13821 22293 13855
rect 22327 13852 22339 13855
rect 23032 13852 23060 13892
rect 23753 13889 23765 13892
rect 23799 13889 23811 13923
rect 24026 13920 24032 13932
rect 23987 13892 24032 13920
rect 23753 13883 23811 13889
rect 24026 13880 24032 13892
rect 24084 13880 24090 13932
rect 22327 13824 23060 13852
rect 23661 13855 23719 13861
rect 22327 13821 22339 13824
rect 22281 13815 22339 13821
rect 23661 13821 23673 13855
rect 23707 13852 23719 13855
rect 24044 13852 24072 13880
rect 23707 13824 24072 13852
rect 27617 13855 27675 13861
rect 23707 13821 23719 13824
rect 23661 13815 23719 13821
rect 27617 13821 27629 13855
rect 27663 13852 27675 13855
rect 28074 13852 28080 13864
rect 27663 13824 28080 13852
rect 27663 13821 27675 13824
rect 27617 13815 27675 13821
rect 21560 13784 21588 13815
rect 22002 13784 22008 13796
rect 21560 13756 22008 13784
rect 22002 13744 22008 13756
rect 22060 13784 22066 13796
rect 22112 13784 22140 13815
rect 28074 13812 28080 13824
rect 28132 13852 28138 13864
rect 28994 13852 29000 13864
rect 28132 13824 29000 13852
rect 28132 13812 28138 13824
rect 28994 13812 29000 13824
rect 29052 13812 29058 13864
rect 22646 13784 22652 13796
rect 22060 13756 22140 13784
rect 22607 13756 22652 13784
rect 22060 13744 22066 13756
rect 22646 13744 22652 13756
rect 22704 13744 22710 13796
rect 27706 13716 27712 13728
rect 19208 13688 19288 13716
rect 27667 13688 27712 13716
rect 19208 13676 19214 13688
rect 27706 13676 27712 13688
rect 27764 13676 27770 13728
rect 1104 13626 29256 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 29256 13626
rect 1104 13552 29256 13574
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 7892 13484 8033 13512
rect 7892 13472 7898 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 11606 13512 11612 13524
rect 8021 13475 8079 13481
rect 8128 13484 11612 13512
rect 6822 13404 6828 13456
rect 6880 13444 6886 13456
rect 8128 13444 8156 13484
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13044 13484 13553 13512
rect 13044 13472 13050 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 13541 13475 13599 13481
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 20806 13512 20812 13524
rect 13955 13484 20812 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 6880 13416 8156 13444
rect 6880 13404 6886 13416
rect 5718 13376 5724 13388
rect 5679 13348 5724 13376
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 7009 13379 7067 13385
rect 7009 13376 7021 13379
rect 5920 13348 7021 13376
rect 5920 13249 5948 13348
rect 7009 13345 7021 13348
rect 7055 13376 7067 13379
rect 7190 13376 7196 13388
rect 7055 13348 7196 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7190 13336 7196 13348
rect 7248 13376 7254 13388
rect 7558 13376 7564 13388
rect 7248 13348 7564 13376
rect 7248 13336 7254 13348
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7745 13379 7803 13385
rect 7745 13345 7757 13379
rect 7791 13376 7803 13379
rect 7926 13376 7932 13388
rect 7791 13348 7932 13376
rect 7791 13345 7803 13348
rect 7745 13339 7803 13345
rect 7926 13336 7932 13348
rect 7984 13336 7990 13388
rect 10962 13376 10968 13388
rect 10923 13348 10968 13376
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 13725 13379 13783 13385
rect 13725 13345 13737 13379
rect 13771 13376 13783 13379
rect 13924 13376 13952 13475
rect 20806 13472 20812 13484
rect 20864 13472 20870 13524
rect 21358 13472 21364 13524
rect 21416 13512 21422 13524
rect 25222 13512 25228 13524
rect 21416 13484 25228 13512
rect 21416 13472 21422 13484
rect 25222 13472 25228 13484
rect 25280 13512 25286 13524
rect 26145 13515 26203 13521
rect 26145 13512 26157 13515
rect 25280 13484 26157 13512
rect 25280 13472 25286 13484
rect 26145 13481 26157 13484
rect 26191 13512 26203 13515
rect 26237 13515 26295 13521
rect 26237 13512 26249 13515
rect 26191 13484 26249 13512
rect 26191 13481 26203 13484
rect 26145 13475 26203 13481
rect 26237 13481 26249 13484
rect 26283 13481 26295 13515
rect 26237 13475 26295 13481
rect 16666 13444 16672 13456
rect 16627 13416 16672 13444
rect 16666 13404 16672 13416
rect 16724 13444 16730 13456
rect 18509 13447 18567 13453
rect 16724 13416 16896 13444
rect 16724 13404 16730 13416
rect 16868 13385 16896 13416
rect 18509 13413 18521 13447
rect 18555 13444 18567 13447
rect 19334 13444 19340 13456
rect 18555 13416 19340 13444
rect 18555 13413 18567 13416
rect 18509 13407 18567 13413
rect 19334 13404 19340 13416
rect 19392 13444 19398 13456
rect 20530 13444 20536 13456
rect 19392 13416 20536 13444
rect 19392 13404 19398 13416
rect 20530 13404 20536 13416
rect 20588 13404 20594 13456
rect 24026 13444 24032 13456
rect 23987 13416 24032 13444
rect 24026 13404 24032 13416
rect 24084 13404 24090 13456
rect 13771 13348 13952 13376
rect 16853 13379 16911 13385
rect 13771 13345 13783 13348
rect 13725 13339 13783 13345
rect 16853 13345 16865 13379
rect 16899 13345 16911 13379
rect 22646 13376 22652 13388
rect 22607 13348 22652 13376
rect 16853 13339 16911 13345
rect 22646 13336 22652 13348
rect 22704 13336 22710 13388
rect 25130 13336 25136 13388
rect 25188 13376 25194 13388
rect 25682 13376 25688 13388
rect 25188 13348 25688 13376
rect 25188 13336 25194 13348
rect 25682 13336 25688 13348
rect 25740 13376 25746 13388
rect 26697 13379 26755 13385
rect 26697 13376 26709 13379
rect 25740 13348 26709 13376
rect 25740 13336 25746 13348
rect 26697 13345 26709 13348
rect 26743 13376 26755 13379
rect 27249 13379 27307 13385
rect 27249 13376 27261 13379
rect 26743 13348 27261 13376
rect 26743 13345 26755 13348
rect 26697 13339 26755 13345
rect 27249 13345 27261 13348
rect 27295 13345 27307 13379
rect 27249 13339 27307 13345
rect 27433 13379 27491 13385
rect 27433 13345 27445 13379
rect 27479 13376 27491 13379
rect 27706 13376 27712 13388
rect 27479 13348 27712 13376
rect 27479 13345 27491 13348
rect 27433 13339 27491 13345
rect 27706 13336 27712 13348
rect 27764 13336 27770 13388
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6656 13280 6837 13308
rect 5905 13243 5963 13249
rect 5905 13209 5917 13243
rect 5951 13209 5963 13243
rect 5905 13203 5963 13209
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 6656 13181 6684 13280
rect 6825 13277 6837 13280
rect 6871 13308 6883 13311
rect 6914 13308 6920 13320
rect 6871 13280 6920 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 11238 13308 11244 13320
rect 11199 13280 11244 13308
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 12618 13308 12624 13320
rect 12531 13280 12624 13308
rect 12618 13268 12624 13280
rect 12676 13308 12682 13320
rect 14274 13308 14280 13320
rect 12676 13280 14280 13308
rect 12676 13268 12682 13280
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 22370 13308 22376 13320
rect 22283 13280 22376 13308
rect 22370 13268 22376 13280
rect 22428 13308 22434 13320
rect 23382 13308 23388 13320
rect 22428 13280 23388 13308
rect 22428 13268 22434 13280
rect 23382 13268 23388 13280
rect 23440 13308 23446 13320
rect 26145 13311 26203 13317
rect 23440 13280 24256 13308
rect 23440 13268 23446 13280
rect 24228 13249 24256 13280
rect 26145 13277 26157 13311
rect 26191 13308 26203 13311
rect 26513 13311 26571 13317
rect 26513 13308 26525 13311
rect 26191 13280 26525 13308
rect 26191 13277 26203 13280
rect 26145 13271 26203 13277
rect 26513 13277 26525 13280
rect 26559 13277 26571 13311
rect 26513 13271 26571 13277
rect 24213 13243 24271 13249
rect 24213 13209 24225 13243
rect 24259 13240 24271 13243
rect 26234 13240 26240 13252
rect 24259 13212 26240 13240
rect 24259 13209 24271 13212
rect 24213 13203 24271 13209
rect 26234 13200 26240 13212
rect 26292 13200 26298 13252
rect 6641 13175 6699 13181
rect 6641 13172 6653 13175
rect 3752 13144 6653 13172
rect 3752 13132 3758 13144
rect 6641 13141 6653 13144
rect 6687 13141 6699 13175
rect 6641 13135 6699 13141
rect 8846 13132 8852 13184
rect 8904 13172 8910 13184
rect 12250 13172 12256 13184
rect 8904 13144 12256 13172
rect 8904 13132 8910 13144
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12710 13172 12716 13184
rect 12671 13144 12716 13172
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 26786 13132 26792 13184
rect 26844 13172 26850 13184
rect 27709 13175 27767 13181
rect 27709 13172 27721 13175
rect 26844 13144 27721 13172
rect 26844 13132 26850 13144
rect 27709 13141 27721 13144
rect 27755 13141 27767 13175
rect 27709 13135 27767 13141
rect 1104 13082 29256 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 29256 13082
rect 1104 13008 29256 13030
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 5442 12968 5448 12980
rect 4479 12940 5448 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 4448 12832 4476 12931
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 18417 12971 18475 12977
rect 7208 12940 10364 12968
rect 2915 12804 4476 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 6604 12804 6653 12832
rect 6604 12792 6610 12804
rect 6641 12801 6653 12804
rect 6687 12832 6699 12835
rect 6822 12832 6828 12844
rect 6687 12804 6828 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 5718 12724 5724 12776
rect 5776 12764 5782 12776
rect 7009 12767 7067 12773
rect 7009 12764 7021 12767
rect 5776 12736 7021 12764
rect 5776 12724 5782 12736
rect 7009 12733 7021 12736
rect 7055 12764 7067 12767
rect 7208 12764 7236 12940
rect 7466 12860 7472 12912
rect 7524 12900 7530 12912
rect 9953 12903 10011 12909
rect 9953 12900 9965 12903
rect 7524 12872 9965 12900
rect 7524 12860 7530 12872
rect 9953 12869 9965 12872
rect 9999 12900 10011 12903
rect 9999 12872 10180 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 10152 12841 10180 12872
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 7558 12764 7564 12776
rect 7055 12736 7236 12764
rect 7519 12736 7564 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 7760 12696 7788 12727
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8904 12736 9045 12764
rect 8904 12724 8910 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 9125 12699 9183 12705
rect 9125 12696 9137 12699
rect 7760 12668 9137 12696
rect 9125 12665 9137 12668
rect 9171 12665 9183 12699
rect 10152 12696 10180 12795
rect 10336 12773 10364 12940
rect 18417 12937 18429 12971
rect 18463 12968 18475 12971
rect 19334 12968 19340 12980
rect 18463 12940 19340 12968
rect 18463 12937 18475 12940
rect 18417 12931 18475 12937
rect 11238 12900 11244 12912
rect 11199 12872 11244 12900
rect 11238 12860 11244 12872
rect 11296 12860 11302 12912
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12764 10379 12767
rect 10870 12764 10876 12776
rect 10367 12736 10876 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 11057 12767 11115 12773
rect 11057 12733 11069 12767
rect 11103 12764 11115 12767
rect 11974 12764 11980 12776
rect 11103 12736 11980 12764
rect 11103 12733 11115 12736
rect 11057 12727 11115 12733
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12425 12767 12483 12773
rect 12425 12733 12437 12767
rect 12471 12764 12483 12767
rect 12526 12764 12532 12776
rect 12471 12736 12532 12764
rect 12471 12733 12483 12736
rect 12425 12727 12483 12733
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18432 12764 18460 12931
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 21542 12968 21548 12980
rect 21315 12940 21548 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 21376 12841 21404 12940
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 24854 12928 24860 12980
rect 24912 12968 24918 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 24912 12940 25053 12968
rect 24912 12928 24918 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 25041 12931 25099 12937
rect 25501 12971 25559 12977
rect 25501 12937 25513 12971
rect 25547 12968 25559 12971
rect 26234 12968 26240 12980
rect 25547 12940 26240 12968
rect 25547 12937 25559 12940
rect 25501 12931 25559 12937
rect 26234 12928 26240 12940
rect 26292 12968 26298 12980
rect 26329 12971 26387 12977
rect 26329 12968 26341 12971
rect 26292 12940 26341 12968
rect 26292 12928 26298 12940
rect 26329 12937 26341 12940
rect 26375 12937 26387 12971
rect 28074 12968 28080 12980
rect 28035 12940 28080 12968
rect 26329 12931 26387 12937
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 21232 12804 21373 12832
rect 21232 12792 21238 12804
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12832 22707 12835
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 22695 12804 23949 12832
rect 22695 12801 22707 12804
rect 22649 12795 22707 12801
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 26344 12832 26372 12931
rect 28074 12928 28080 12940
rect 28132 12928 28138 12980
rect 26510 12832 26516 12844
rect 26344 12804 26516 12832
rect 23937 12795 23995 12801
rect 26510 12792 26516 12804
rect 26568 12792 26574 12844
rect 26786 12832 26792 12844
rect 26747 12804 26792 12832
rect 26786 12792 26792 12804
rect 26844 12792 26850 12844
rect 18095 12736 18460 12764
rect 21545 12767 21603 12773
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 21545 12733 21557 12767
rect 21591 12733 21603 12767
rect 21545 12727 21603 12733
rect 22097 12767 22155 12773
rect 22097 12733 22109 12767
rect 22143 12733 22155 12767
rect 22278 12764 22284 12776
rect 22239 12736 22284 12764
rect 22097 12727 22155 12733
rect 12894 12696 12900 12708
rect 10152 12668 12900 12696
rect 9125 12659 9183 12665
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 21560 12696 21588 12727
rect 22002 12696 22008 12708
rect 17052 12668 22008 12696
rect 17052 12640 17080 12668
rect 22002 12656 22008 12668
rect 22060 12696 22066 12708
rect 22112 12696 22140 12727
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 23661 12767 23719 12773
rect 23661 12764 23673 12767
rect 23440 12736 23673 12764
rect 23440 12724 23446 12736
rect 23661 12733 23673 12736
rect 23707 12733 23719 12767
rect 23661 12727 23719 12733
rect 22060 12668 22140 12696
rect 22060 12656 22066 12668
rect 4154 12628 4160 12640
rect 4115 12600 4160 12628
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4614 12628 4620 12640
rect 4575 12600 4620 12628
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 8018 12628 8024 12640
rect 7979 12600 8024 12628
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 10870 12588 10876 12640
rect 10928 12628 10934 12640
rect 12526 12628 12532 12640
rect 10928 12600 12532 12628
rect 10928 12588 10934 12600
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12621 12631 12679 12637
rect 12621 12597 12633 12631
rect 12667 12628 12679 12631
rect 17034 12628 17040 12640
rect 12667 12600 17040 12628
rect 12667 12597 12679 12600
rect 12621 12591 12679 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 18138 12628 18144 12640
rect 18099 12600 18144 12628
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 1104 12538 29256 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 29256 12538
rect 1104 12464 29256 12486
rect 7929 12427 7987 12433
rect 7929 12393 7941 12427
rect 7975 12424 7987 12427
rect 8846 12424 8852 12436
rect 7975 12396 8852 12424
rect 7975 12393 7987 12396
rect 7929 12387 7987 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 11974 12424 11980 12436
rect 11935 12396 11980 12424
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12084 12396 13308 12424
rect 12084 12356 12112 12396
rect 7300 12328 12112 12356
rect 12253 12359 12311 12365
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 7300 12288 7328 12328
rect 12253 12325 12265 12359
rect 12299 12356 12311 12359
rect 12618 12356 12624 12368
rect 12299 12328 12624 12356
rect 12299 12325 12311 12328
rect 12253 12319 12311 12325
rect 4120 12260 7328 12288
rect 11885 12291 11943 12297
rect 4120 12248 4126 12260
rect 11885 12257 11897 12291
rect 11931 12288 11943 12291
rect 12268 12288 12296 12319
rect 12618 12316 12624 12328
rect 12676 12316 12682 12368
rect 13280 12356 13308 12396
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17184 12396 17509 12424
rect 17184 12384 17190 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 17497 12387 17555 12393
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 22925 12427 22983 12433
rect 22925 12424 22937 12427
rect 22336 12396 22937 12424
rect 22336 12384 22342 12396
rect 22925 12393 22937 12396
rect 22971 12393 22983 12427
rect 22925 12387 22983 12393
rect 23201 12427 23259 12433
rect 23201 12393 23213 12427
rect 23247 12424 23259 12427
rect 24854 12424 24860 12436
rect 23247 12396 24860 12424
rect 23247 12393 23259 12396
rect 23201 12387 23259 12393
rect 21174 12356 21180 12368
rect 13280 12328 21180 12356
rect 21174 12316 21180 12328
rect 21232 12316 21238 12368
rect 11931 12260 12296 12288
rect 11931 12257 11943 12260
rect 11885 12251 11943 12257
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 13044 12260 13093 12288
rect 13044 12248 13050 12260
rect 13081 12257 13093 12260
rect 13127 12257 13139 12291
rect 13538 12288 13544 12300
rect 13499 12260 13544 12288
rect 13081 12251 13139 12257
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 14424 12260 16497 12288
rect 14424 12248 14430 12260
rect 16485 12257 16497 12260
rect 16531 12288 16543 12291
rect 16666 12288 16672 12300
rect 16531 12260 16672 12288
rect 16531 12257 16543 12260
rect 16485 12251 16543 12257
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 17034 12288 17040 12300
rect 16995 12260 17040 12288
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17221 12291 17279 12297
rect 17221 12257 17233 12291
rect 17267 12288 17279 12291
rect 18138 12288 18144 12300
rect 17267 12260 18144 12288
rect 17267 12257 17279 12260
rect 17221 12251 17279 12257
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 22833 12291 22891 12297
rect 22833 12257 22845 12291
rect 22879 12288 22891 12291
rect 23216 12288 23244 12387
rect 24854 12384 24860 12396
rect 24912 12384 24918 12436
rect 22879 12260 23244 12288
rect 22879 12257 22891 12260
rect 22833 12251 22891 12257
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 8018 12220 8024 12232
rect 6687 12192 8024 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 6380 12084 6408 12183
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 12584 12192 16037 12220
rect 12584 12180 12590 12192
rect 16025 12189 16037 12192
rect 16071 12220 16083 12223
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 16071 12192 16313 12220
rect 16071 12189 16083 12192
rect 16025 12183 16083 12189
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 22094 12152 22100 12164
rect 12676 12124 22100 12152
rect 12676 12112 12682 12124
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 4672 12056 8125 12084
rect 4672 12044 4678 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 12894 12084 12900 12096
rect 12855 12056 12900 12084
rect 8113 12047 8171 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 13633 12087 13691 12093
rect 13633 12084 13645 12087
rect 13504 12056 13645 12084
rect 13504 12044 13510 12056
rect 13633 12053 13645 12056
rect 13679 12053 13691 12087
rect 13633 12047 13691 12053
rect 16025 12087 16083 12093
rect 16025 12053 16037 12087
rect 16071 12084 16083 12087
rect 16209 12087 16267 12093
rect 16209 12084 16221 12087
rect 16071 12056 16221 12084
rect 16071 12053 16083 12056
rect 16025 12047 16083 12053
rect 16209 12053 16221 12056
rect 16255 12084 16267 12087
rect 21266 12084 21272 12096
rect 16255 12056 21272 12084
rect 16255 12053 16267 12056
rect 16209 12047 16267 12053
rect 21266 12044 21272 12056
rect 21324 12044 21330 12096
rect 1104 11994 29256 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 29256 11994
rect 1104 11920 29256 11942
rect 6914 11840 6920 11892
rect 6972 11880 6978 11892
rect 7561 11883 7619 11889
rect 7561 11880 7573 11883
rect 6972 11852 7573 11880
rect 6972 11840 6978 11852
rect 7561 11849 7573 11852
rect 7607 11880 7619 11883
rect 8202 11880 8208 11892
rect 7607 11852 8208 11880
rect 7607 11849 7619 11852
rect 7561 11843 7619 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 12526 11880 12532 11892
rect 8312 11852 12532 11880
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 8312 11812 8340 11852
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 12710 11880 12716 11892
rect 12671 11852 12716 11880
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 12894 11840 12900 11892
rect 12952 11880 12958 11892
rect 15010 11880 15016 11892
rect 12952 11852 15016 11880
rect 12952 11840 12958 11852
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21726 11880 21732 11892
rect 20772 11852 21732 11880
rect 20772 11840 20778 11852
rect 21726 11840 21732 11852
rect 21784 11880 21790 11892
rect 29638 11880 29644 11892
rect 21784 11852 29644 11880
rect 21784 11840 21790 11852
rect 29638 11840 29644 11852
rect 29696 11840 29702 11892
rect 4028 11784 8340 11812
rect 4028 11772 4034 11784
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 2915 11716 7389 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 12728 11744 12756 11840
rect 24489 11815 24547 11821
rect 24489 11812 24501 11815
rect 24320 11784 24501 11812
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12728 11716 12909 11744
rect 7377 11707 7435 11713
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11744 18659 11747
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 18647 11716 20545 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 20533 11713 20545 11716
rect 20579 11744 20591 11747
rect 24320 11744 24348 11784
rect 24489 11781 24501 11784
rect 24535 11781 24547 11815
rect 24489 11775 24547 11781
rect 24857 11747 24915 11753
rect 24857 11744 24869 11747
rect 20579 11716 20852 11744
rect 20579 11713 20591 11716
rect 20533 11707 20591 11713
rect 2590 11676 2596 11688
rect 2551 11648 2596 11676
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 6840 11608 6868 11639
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 6972 11648 7017 11676
rect 6972 11636 6978 11648
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7984 11648 8217 11676
rect 7984 11636 7990 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 10594 11676 10600 11688
rect 8343 11648 10600 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 10594 11636 10600 11648
rect 10652 11636 10658 11688
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11676 13231 11679
rect 15378 11676 15384 11688
rect 13219 11648 15384 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 20349 11679 20407 11685
rect 20349 11676 20361 11679
rect 18923 11648 20361 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 20349 11645 20361 11648
rect 20395 11676 20407 11679
rect 20714 11676 20720 11688
rect 20395 11648 20720 11676
rect 20395 11645 20407 11648
rect 20349 11639 20407 11645
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 20824 11676 20852 11716
rect 24320 11716 24869 11744
rect 22370 11676 22376 11688
rect 20824 11648 22376 11676
rect 22370 11636 22376 11648
rect 22428 11676 22434 11688
rect 24320 11685 24348 11716
rect 24857 11713 24869 11716
rect 24903 11713 24915 11747
rect 25130 11744 25136 11756
rect 25091 11716 25136 11744
rect 24857 11707 24915 11713
rect 25130 11704 25136 11716
rect 25188 11704 25194 11756
rect 24305 11679 24363 11685
rect 24305 11676 24317 11679
rect 22428 11648 24317 11676
rect 22428 11636 22434 11648
rect 24305 11645 24317 11648
rect 24351 11645 24363 11679
rect 24305 11639 24363 11645
rect 24394 11636 24400 11688
rect 24452 11676 24458 11688
rect 24673 11679 24731 11685
rect 24673 11676 24685 11679
rect 24452 11648 24685 11676
rect 24452 11636 24458 11648
rect 24673 11645 24685 11648
rect 24719 11645 24731 11679
rect 24673 11639 24731 11645
rect 7944 11608 7972 11636
rect 6840 11580 7972 11608
rect 8110 11568 8116 11620
rect 8168 11608 8174 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 8168 11580 8769 11608
rect 8168 11568 8174 11580
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 14090 11568 14096 11620
rect 14148 11608 14154 11620
rect 14550 11608 14556 11620
rect 14148 11580 14556 11608
rect 14148 11568 14154 11580
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 4154 11540 4160 11552
rect 4115 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4433 11543 4491 11549
rect 4433 11509 4445 11543
rect 4479 11540 4491 11543
rect 4614 11540 4620 11552
rect 4479 11512 4620 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 11330 11540 11336 11552
rect 5592 11512 11336 11540
rect 5592 11500 5598 11512
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 18598 11500 18604 11552
rect 18656 11540 18662 11552
rect 19981 11543 20039 11549
rect 19981 11540 19993 11543
rect 18656 11512 19993 11540
rect 18656 11500 18662 11512
rect 19981 11509 19993 11512
rect 20027 11509 20039 11543
rect 26234 11540 26240 11552
rect 26195 11512 26240 11540
rect 19981 11503 20039 11509
rect 26234 11500 26240 11512
rect 26292 11500 26298 11552
rect 1104 11450 29256 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 29256 11450
rect 1104 11376 29256 11398
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5534 11336 5540 11348
rect 5307 11308 5540 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5368 11209 5396 11308
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 10686 11336 10692 11348
rect 6564 11308 10692 11336
rect 6564 11209 6592 11308
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 12621 11339 12679 11345
rect 12621 11305 12633 11339
rect 12667 11336 12679 11339
rect 12710 11336 12716 11348
rect 12667 11308 12716 11336
rect 12667 11305 12679 11308
rect 12621 11299 12679 11305
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13872 11308 14105 11336
rect 13872 11296 13878 11308
rect 14093 11305 14105 11308
rect 14139 11336 14151 11339
rect 14458 11336 14464 11348
rect 14139 11308 14464 11336
rect 14139 11305 14151 11308
rect 14093 11299 14151 11305
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 15378 11336 15384 11348
rect 15339 11308 15384 11336
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 18233 11339 18291 11345
rect 18233 11305 18245 11339
rect 18279 11336 18291 11339
rect 20073 11339 20131 11345
rect 20073 11336 20085 11339
rect 18279 11308 20085 11336
rect 18279 11305 18291 11308
rect 18233 11299 18291 11305
rect 20073 11305 20085 11308
rect 20119 11336 20131 11339
rect 21082 11336 21088 11348
rect 20119 11308 21088 11336
rect 20119 11305 20131 11308
rect 20073 11299 20131 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 8021 11271 8079 11277
rect 8021 11237 8033 11271
rect 8067 11268 8079 11271
rect 9122 11268 9128 11280
rect 8067 11240 9128 11268
rect 8067 11237 8079 11240
rect 8021 11231 8079 11237
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11169 6607 11203
rect 7926 11200 7932 11212
rect 7887 11172 7932 11200
rect 6549 11163 6607 11169
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 8159 11172 8769 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 8757 11169 8769 11172
rect 8803 11200 8815 11203
rect 12618 11200 12624 11212
rect 8803 11172 12624 11200
rect 8803 11169 8815 11172
rect 8757 11163 8815 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 12728 11209 12756 11296
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11169 12771 11203
rect 12713 11163 12771 11169
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 14608 11172 15945 11200
rect 14608 11160 14614 11172
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11200 16359 11203
rect 18598 11200 18604 11212
rect 16347 11172 18460 11200
rect 18559 11172 18604 11200
rect 16347 11169 16359 11172
rect 16301 11163 16359 11169
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 5552 11104 6469 11132
rect 2958 11024 2964 11076
rect 3016 11064 3022 11076
rect 5552 11073 5580 11104
rect 6457 11101 6469 11104
rect 6503 11132 6515 11135
rect 7944 11132 7972 11160
rect 6503 11104 7972 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8076 11104 8585 11132
rect 8076 11092 8082 11104
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13814 11132 13820 11144
rect 13035 11104 13820 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 16206 11132 16212 11144
rect 15887 11104 15921 11132
rect 16167 11104 16212 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 5537 11067 5595 11073
rect 3016 11036 5488 11064
rect 3016 11024 3022 11036
rect 5460 10996 5488 11036
rect 5537 11033 5549 11067
rect 5583 11033 5595 11067
rect 5537 11027 5595 11033
rect 5644 11036 6776 11064
rect 5644 10996 5672 11036
rect 6748 11005 6776 11036
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 15856 11064 15884 11095
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 18012 11104 18245 11132
rect 18012 11092 18018 11104
rect 18233 11101 18245 11104
rect 18279 11132 18291 11135
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 18279 11104 18337 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18432 11132 18460 11172
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 23753 11203 23811 11209
rect 23753 11200 23765 11203
rect 22020 11172 23765 11200
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 18432 11104 19717 11132
rect 18325 11095 18383 11101
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 21082 11092 21088 11144
rect 21140 11132 21146 11144
rect 22020 11141 22048 11172
rect 23753 11169 23765 11172
rect 23799 11169 23811 11203
rect 23753 11163 23811 11169
rect 22005 11135 22063 11141
rect 22005 11132 22017 11135
rect 21140 11104 22017 11132
rect 21140 11092 21146 11104
rect 22005 11101 22017 11104
rect 22051 11101 22063 11135
rect 22278 11132 22284 11144
rect 22239 11104 22284 11132
rect 22005 11095 22063 11101
rect 22278 11092 22284 11104
rect 22336 11092 22342 11144
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 15344 11036 16589 11064
rect 15344 11024 15350 11036
rect 16577 11033 16589 11036
rect 16623 11033 16635 11067
rect 16577 11027 16635 11033
rect 5460 10968 5672 10996
rect 6733 10999 6791 11005
rect 6733 10965 6745 10999
rect 6779 10965 6791 10999
rect 6733 10959 6791 10965
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 17770 10996 17776 11008
rect 6880 10968 17776 10996
rect 6880 10956 6886 10968
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 23566 10996 23572 11008
rect 23527 10968 23572 10996
rect 23566 10956 23572 10968
rect 23624 10956 23630 11008
rect 1104 10906 29256 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 29256 10906
rect 1104 10832 29256 10854
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 6822 10792 6828 10804
rect 4028 10764 6828 10792
rect 4028 10752 4034 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7377 10795 7435 10801
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 7926 10792 7932 10804
rect 7423 10764 7932 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8297 10795 8355 10801
rect 8297 10761 8309 10795
rect 8343 10792 8355 10795
rect 15194 10792 15200 10804
rect 8343 10764 15200 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 8113 10659 8171 10665
rect 8113 10656 8125 10659
rect 2915 10628 8125 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 8113 10625 8125 10628
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 2590 10588 2596 10600
rect 2551 10560 2596 10588
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 8312 10588 8340 10755
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 22278 10752 22284 10804
rect 22336 10792 22342 10804
rect 22465 10795 22523 10801
rect 22465 10792 22477 10795
rect 22336 10764 22477 10792
rect 22336 10752 22342 10764
rect 22465 10761 22477 10764
rect 22511 10761 22523 10795
rect 22465 10755 22523 10761
rect 13814 10656 13820 10668
rect 13775 10628 13820 10656
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10625 14611 10659
rect 23566 10656 23572 10668
rect 14553 10619 14611 10625
rect 14844 10628 23572 10656
rect 14458 10588 14464 10600
rect 7699 10560 8340 10588
rect 14419 10560 14464 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 7558 10520 7564 10532
rect 7519 10492 7564 10520
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 4154 10452 4160 10464
rect 4115 10424 4160 10452
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4614 10452 4620 10464
rect 4479 10424 4620 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 14568 10452 14596 10619
rect 14844 10597 14872 10628
rect 23566 10616 23572 10628
rect 23624 10616 23630 10668
rect 25869 10659 25927 10665
rect 25869 10625 25881 10659
rect 25915 10656 25927 10659
rect 26234 10656 26240 10668
rect 25915 10628 26240 10656
rect 25915 10625 25927 10628
rect 25869 10619 25927 10625
rect 26234 10616 26240 10628
rect 26292 10616 26298 10668
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10557 14887 10591
rect 14829 10551 14887 10557
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15841 10591 15899 10597
rect 15841 10588 15853 10591
rect 15059 10560 15853 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15841 10557 15853 10560
rect 15887 10588 15899 10591
rect 16206 10588 16212 10600
rect 15887 10560 16212 10588
rect 15887 10557 15899 10560
rect 15841 10551 15899 10557
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 21082 10588 21088 10600
rect 21043 10560 21088 10588
rect 21082 10548 21088 10560
rect 21140 10548 21146 10600
rect 21358 10588 21364 10600
rect 21319 10560 21364 10588
rect 21358 10548 21364 10560
rect 21416 10548 21422 10600
rect 25501 10591 25559 10597
rect 25501 10557 25513 10591
rect 25547 10588 25559 10591
rect 25593 10591 25651 10597
rect 25593 10588 25605 10591
rect 25547 10560 25605 10588
rect 25547 10557 25559 10560
rect 25501 10551 25559 10557
rect 25593 10557 25605 10560
rect 25639 10588 25651 10591
rect 26510 10588 26516 10600
rect 25639 10560 26516 10588
rect 25639 10557 25651 10560
rect 25593 10551 25651 10557
rect 26510 10548 26516 10560
rect 26568 10548 26574 10600
rect 15194 10452 15200 10464
rect 14568 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 16025 10455 16083 10461
rect 16025 10421 16037 10455
rect 16071 10452 16083 10455
rect 16482 10452 16488 10464
rect 16071 10424 16488 10452
rect 16071 10421 16083 10424
rect 16025 10415 16083 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 21100 10452 21128 10548
rect 22833 10455 22891 10461
rect 22833 10452 22845 10455
rect 21100 10424 22845 10452
rect 22833 10421 22845 10424
rect 22879 10421 22891 10455
rect 22833 10415 22891 10421
rect 26786 10412 26792 10464
rect 26844 10452 26850 10464
rect 26973 10455 27031 10461
rect 26973 10452 26985 10455
rect 26844 10424 26985 10452
rect 26844 10412 26850 10424
rect 26973 10421 26985 10424
rect 27019 10421 27031 10455
rect 26973 10415 27031 10421
rect 1104 10362 29256 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 29256 10362
rect 1104 10288 29256 10310
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 7616 10220 8493 10248
rect 7616 10208 7622 10220
rect 8481 10217 8493 10220
rect 8527 10217 8539 10251
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 8481 10211 8539 10217
rect 11330 10208 11336 10220
rect 11388 10248 11394 10260
rect 12437 10251 12495 10257
rect 12437 10248 12449 10251
rect 11388 10220 11560 10248
rect 11388 10208 11394 10220
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 6822 10112 6828 10124
rect 5767 10084 6828 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6822 10072 6828 10084
rect 6880 10112 6886 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 6880 10084 7481 10112
rect 6880 10072 6886 10084
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10112 8263 10115
rect 8294 10112 8300 10124
rect 8251 10084 8300 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 11532 10121 11560 10220
rect 11808 10220 12449 10248
rect 11808 10121 11836 10220
rect 12437 10217 12449 10220
rect 12483 10248 12495 10251
rect 15010 10248 15016 10260
rect 12483 10220 14872 10248
rect 14971 10220 15016 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10081 8447 10115
rect 8389 10075 8447 10081
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10044 6055 10047
rect 6914 10044 6920 10056
rect 6043 10016 6920 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 8404 10044 8432 10075
rect 7392 10016 8432 10044
rect 11716 10044 11744 10075
rect 12526 10044 12532 10056
rect 11716 10016 12532 10044
rect 7392 9920 7420 10016
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 14844 10044 14872 10220
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 16448 10220 16681 10248
rect 16448 10208 16454 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 21358 10208 21364 10260
rect 21416 10248 21422 10260
rect 21545 10251 21603 10257
rect 21545 10248 21557 10251
rect 21416 10220 21557 10248
rect 21416 10208 21422 10220
rect 21545 10217 21557 10220
rect 21591 10217 21603 10251
rect 21726 10248 21732 10260
rect 21687 10220 21732 10248
rect 21545 10211 21603 10217
rect 21726 10208 21732 10220
rect 21784 10208 21790 10260
rect 15028 10112 15056 10208
rect 20622 10180 20628 10192
rect 16224 10152 20628 10180
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 15028 10084 15301 10112
rect 15289 10081 15301 10084
rect 15335 10081 15347 10115
rect 16224 10112 16252 10152
rect 20622 10140 20628 10152
rect 20680 10140 20686 10192
rect 15289 10075 15347 10081
rect 15396 10084 16252 10112
rect 20901 10115 20959 10121
rect 15396 10044 15424 10084
rect 20901 10081 20913 10115
rect 20947 10112 20959 10115
rect 21744 10112 21772 10208
rect 20947 10084 21772 10112
rect 26329 10115 26387 10121
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 26329 10081 26341 10115
rect 26375 10112 26387 10115
rect 26510 10112 26516 10124
rect 26375 10084 26516 10112
rect 26375 10081 26387 10084
rect 26329 10075 26387 10081
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 26786 10112 26792 10124
rect 26747 10084 26792 10112
rect 26786 10072 26792 10084
rect 26844 10072 26850 10124
rect 15562 10044 15568 10056
rect 14844 10016 15424 10044
rect 15523 10016 15568 10044
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7374 9908 7380 9920
rect 7331 9880 7380 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11112 9880 11989 9908
rect 11112 9868 11118 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 27890 9908 27896 9920
rect 27851 9880 27896 9908
rect 11977 9871 12035 9877
rect 27890 9868 27896 9880
rect 27948 9868 27954 9920
rect 1104 9818 29256 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 29256 9818
rect 1104 9744 29256 9766
rect 9122 9704 9128 9716
rect 9083 9676 9128 9704
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 11388 9676 12173 9704
rect 11388 9664 11394 9676
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 12161 9667 12219 9673
rect 26237 9707 26295 9713
rect 26237 9673 26249 9707
rect 26283 9704 26295 9707
rect 26510 9704 26516 9716
rect 26283 9676 26516 9704
rect 26283 9673 26295 9676
rect 26237 9667 26295 9673
rect 8018 9636 8024 9648
rect 4632 9608 8024 9636
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 4632 9568 4660 9608
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 12176 9636 12204 9667
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12176 9608 12449 9636
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 12437 9599 12495 9605
rect 13354 9596 13360 9648
rect 13412 9636 13418 9648
rect 13412 9608 16160 9636
rect 13412 9596 13418 9608
rect 16132 9580 16160 9608
rect 20806 9596 20812 9648
rect 20864 9636 20870 9648
rect 24213 9639 24271 9645
rect 24213 9636 24225 9639
rect 20864 9608 24225 9636
rect 20864 9596 20870 9608
rect 24213 9605 24225 9608
rect 24259 9605 24271 9639
rect 24394 9636 24400 9648
rect 24355 9608 24400 9636
rect 24213 9599 24271 9605
rect 6914 9568 6920 9580
rect 2915 9540 4660 9568
rect 6875 9540 6920 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 7432 9540 7757 9568
rect 7432 9528 7438 9540
rect 7745 9537 7757 9540
rect 7791 9537 7803 9571
rect 8205 9571 8263 9577
rect 8205 9568 8217 9571
rect 7745 9531 7803 9537
rect 7852 9540 8217 9568
rect 2590 9500 2596 9512
rect 2551 9472 2596 9500
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4614 9500 4620 9512
rect 4479 9472 4620 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4614 9460 4620 9472
rect 4672 9500 4678 9512
rect 6822 9500 6828 9512
rect 4672 9472 6828 9500
rect 4672 9460 4678 9472
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7282 9500 7288 9512
rect 7243 9472 7288 9500
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7852 9509 7880 9540
rect 8205 9537 8217 9540
rect 8251 9568 8263 9571
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 8251 9540 10701 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 7837 9463 7895 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 10244 9509 10272 9540
rect 10689 9537 10701 9540
rect 10735 9568 10747 9571
rect 15194 9568 15200 9580
rect 10735 9540 15200 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15562 9528 15568 9580
rect 15620 9568 15626 9580
rect 15657 9571 15715 9577
rect 15657 9568 15669 9571
rect 15620 9540 15669 9568
rect 15620 9528 15626 9540
rect 15657 9537 15669 9540
rect 15703 9537 15715 9571
rect 16114 9568 16120 9580
rect 16027 9540 16120 9568
rect 15657 9531 15715 9537
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 16577 9571 16635 9577
rect 16577 9568 16589 9571
rect 16264 9540 16589 9568
rect 16264 9528 16270 9540
rect 16577 9537 16589 9540
rect 16623 9537 16635 9571
rect 16577 9531 16635 9537
rect 21358 9528 21364 9580
rect 21416 9568 21422 9580
rect 21637 9571 21695 9577
rect 21637 9568 21649 9571
rect 21416 9540 21649 9568
rect 21416 9528 21422 9540
rect 21637 9537 21649 9540
rect 21683 9537 21695 9571
rect 21637 9531 21695 9537
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9469 10287 9503
rect 10229 9463 10287 9469
rect 12713 9503 12771 9509
rect 12713 9469 12725 9503
rect 12759 9500 12771 9503
rect 16301 9503 16359 9509
rect 12759 9472 14780 9500
rect 12759 9469 12771 9472
rect 12713 9463 12771 9469
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 8849 9435 8907 9441
rect 8849 9432 8861 9435
rect 8352 9404 8861 9432
rect 8352 9392 8358 9404
rect 8849 9401 8861 9404
rect 8895 9432 8907 9435
rect 12618 9432 12624 9444
rect 8895 9404 10640 9432
rect 12579 9404 12624 9432
rect 8895 9401 8907 9404
rect 8849 9395 8907 9401
rect 4154 9364 4160 9376
rect 4115 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10502 9364 10508 9376
rect 10459 9336 10508 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10612 9364 10640 9404
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 13170 9432 13176 9444
rect 13131 9404 13176 9432
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 14752 9432 14780 9472
rect 16301 9469 16313 9503
rect 16347 9500 16359 9503
rect 16390 9500 16396 9512
rect 16347 9472 16396 9500
rect 16347 9469 16359 9472
rect 16301 9463 16359 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9500 16727 9503
rect 23198 9500 23204 9512
rect 16715 9472 23204 9500
rect 16715 9469 16727 9472
rect 16669 9463 16727 9469
rect 23198 9460 23204 9472
rect 23256 9460 23262 9512
rect 24228 9500 24256 9599
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 26344 9577 26372 9676
rect 26510 9664 26516 9676
rect 26568 9664 26574 9716
rect 26329 9571 26387 9577
rect 26329 9537 26341 9571
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 26605 9571 26663 9577
rect 26605 9537 26617 9571
rect 26651 9568 26663 9571
rect 27890 9568 27896 9580
rect 26651 9540 27896 9568
rect 26651 9537 26663 9540
rect 26605 9531 26663 9537
rect 27890 9528 27896 9540
rect 27948 9528 27954 9580
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 24228 9472 24593 9500
rect 24581 9469 24593 9472
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 16850 9432 16856 9444
rect 14752 9404 16856 9432
rect 16850 9392 16856 9404
rect 16908 9392 16914 9444
rect 12434 9364 12440 9376
rect 10612 9336 12440 9364
rect 12434 9324 12440 9336
rect 12492 9364 12498 9376
rect 13446 9364 13452 9376
rect 12492 9336 13452 9364
rect 12492 9324 12498 9336
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 22278 9364 22284 9376
rect 22239 9336 22284 9364
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 27706 9364 27712 9376
rect 27667 9336 27712 9364
rect 27706 9324 27712 9336
rect 27764 9324 27770 9376
rect 1104 9274 29256 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 29256 9274
rect 1104 9200 29256 9222
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 12676 9132 13737 9160
rect 12676 9120 12682 9132
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 15473 9163 15531 9169
rect 15473 9129 15485 9163
rect 15519 9160 15531 9163
rect 16206 9160 16212 9172
rect 15519 9132 16212 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 27706 9160 27712 9172
rect 16684 9132 27712 9160
rect 11900 9064 12204 9092
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11900 9033 11928 9064
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 10560 8996 11897 9024
rect 10560 8984 10566 8996
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 11422 8956 11428 8968
rect 11383 8928 11428 8956
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 12084 8888 12112 8987
rect 12176 8956 12204 9064
rect 12342 9052 12348 9104
rect 12400 9092 12406 9104
rect 13446 9092 13452 9104
rect 12400 9064 12572 9092
rect 13407 9064 13452 9092
rect 12400 9052 12406 9064
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 12544 9033 12572 9064
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 16574 9092 16580 9104
rect 13648 9064 16580 9092
rect 13648 9033 13676 9064
rect 16574 9052 16580 9064
rect 16632 9052 16638 9104
rect 12437 9027 12495 9033
rect 12437 9024 12449 9027
rect 12308 8996 12449 9024
rect 12308 8984 12314 8996
rect 12437 8993 12449 8996
rect 12483 8993 12495 9027
rect 12437 8987 12495 8993
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 15381 9027 15439 9033
rect 15381 9024 15393 9027
rect 15252 8996 15393 9024
rect 15252 8984 15258 8996
rect 15381 8993 15393 8996
rect 15427 9024 15439 9027
rect 16684 9024 16712 9132
rect 27706 9120 27712 9132
rect 27764 9120 27770 9172
rect 18233 9095 18291 9101
rect 18233 9061 18245 9095
rect 18279 9092 18291 9095
rect 18690 9092 18696 9104
rect 18279 9064 18696 9092
rect 18279 9061 18291 9064
rect 18233 9055 18291 9061
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 15427 8996 15608 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 15580 8956 15608 8996
rect 15948 8996 16712 9024
rect 22281 9027 22339 9033
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 12176 8928 12756 8956
rect 15580 8928 15761 8956
rect 12618 8888 12624 8900
rect 12084 8860 12624 8888
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 12728 8888 12756 8928
rect 15749 8925 15761 8928
rect 15795 8956 15807 8959
rect 15948 8956 15976 8996
rect 22281 8993 22293 9027
rect 22327 9024 22339 9027
rect 24394 9024 24400 9036
rect 22327 8996 24400 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 24394 8984 24400 8996
rect 24452 8984 24458 9036
rect 15795 8928 15976 8956
rect 16577 8959 16635 8965
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 16577 8925 16589 8959
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 18046 8956 18052 8968
rect 16899 8928 18052 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 13354 8888 13360 8900
rect 12728 8860 13360 8888
rect 13354 8848 13360 8860
rect 13412 8848 13418 8900
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 14182 8820 14188 8832
rect 4120 8792 14188 8820
rect 4120 8780 4126 8792
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 16592 8820 16620 8919
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 22833 8959 22891 8965
rect 22833 8956 22845 8959
rect 22756 8928 22845 8956
rect 22756 8832 22784 8928
rect 22833 8925 22845 8928
rect 22879 8925 22891 8959
rect 23106 8956 23112 8968
rect 23067 8928 23112 8956
rect 22833 8919 22891 8925
rect 23106 8916 23112 8928
rect 23164 8916 23170 8968
rect 23198 8916 23204 8968
rect 23256 8956 23262 8968
rect 24213 8959 24271 8965
rect 24213 8956 24225 8959
rect 23256 8928 24225 8956
rect 23256 8916 23262 8928
rect 24213 8925 24225 8928
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 16758 8820 16764 8832
rect 16592 8792 16764 8820
rect 16758 8780 16764 8792
rect 16816 8820 16822 8832
rect 17862 8820 17868 8832
rect 16816 8792 17868 8820
rect 16816 8780 16822 8792
rect 17862 8780 17868 8792
rect 17920 8820 17926 8832
rect 18325 8823 18383 8829
rect 18325 8820 18337 8823
rect 17920 8792 18337 8820
rect 17920 8780 17926 8792
rect 18325 8789 18337 8792
rect 18371 8789 18383 8823
rect 18325 8783 18383 8789
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 22738 8820 22744 8832
rect 22152 8792 22744 8820
rect 22152 8780 22158 8792
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 1104 8730 29256 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 29256 8730
rect 1104 8656 29256 8678
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7524 8588 11284 8616
rect 7524 8576 7530 8588
rect 10962 8548 10968 8560
rect 8496 8520 10968 8548
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3384 8452 3985 8480
rect 3384 8440 3390 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 8496 8480 8524 8520
rect 10962 8508 10968 8520
rect 11020 8508 11026 8560
rect 3973 8443 4031 8449
rect 7392 8452 8524 8480
rect 2590 8412 2596 8424
rect 2503 8384 2596 8412
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 7392 8412 7420 8452
rect 9030 8440 9036 8492
rect 9088 8480 9094 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 9088 8452 9229 8480
rect 9088 8440 9094 8452
rect 9217 8449 9229 8452
rect 9263 8480 9275 8483
rect 11256 8480 11284 8588
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 12713 8619 12771 8625
rect 12713 8616 12725 8619
rect 12584 8588 12725 8616
rect 12584 8576 12590 8588
rect 12713 8585 12725 8588
rect 12759 8585 12771 8619
rect 16482 8616 16488 8628
rect 12713 8579 12771 8585
rect 13372 8588 16488 8616
rect 12342 8480 12348 8492
rect 9263 8452 10732 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 2915 8384 7420 8412
rect 7561 8415 7619 8421
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 7650 8412 7656 8424
rect 7607 8384 7656 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 7837 8415 7895 8421
rect 7837 8381 7849 8415
rect 7883 8412 7895 8415
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 7883 8384 10057 8412
rect 7883 8381 7895 8384
rect 7837 8375 7895 8381
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 10045 8375 10103 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10704 8421 10732 8452
rect 11256 8452 12348 8480
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11256 8421 11284 8452
rect 12342 8440 12348 8452
rect 12400 8480 12406 8492
rect 13372 8480 13400 8588
rect 16482 8576 16488 8588
rect 16540 8616 16546 8628
rect 17126 8616 17132 8628
rect 16540 8588 17132 8616
rect 16540 8576 16546 8588
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 22094 8616 22100 8628
rect 17920 8588 22100 8616
rect 17920 8576 17926 8588
rect 16408 8520 18552 8548
rect 12400 8452 13400 8480
rect 12400 8440 12406 8452
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16408 8489 16436 8520
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 16172 8452 16405 8480
rect 16172 8440 16178 8452
rect 16393 8449 16405 8452
rect 16439 8449 16451 8483
rect 18046 8480 18052 8492
rect 18007 8452 18052 8480
rect 16393 8443 16451 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18524 8489 18552 8520
rect 21100 8489 21128 8588
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 22649 8619 22707 8625
rect 22649 8585 22661 8619
rect 22695 8616 22707 8619
rect 23106 8616 23112 8628
rect 22695 8588 23112 8616
rect 22695 8585 22707 8588
rect 22649 8579 22707 8585
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18969 8483 19027 8489
rect 18969 8449 18981 8483
rect 19015 8449 19027 8483
rect 18969 8443 19027 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 22278 8480 22284 8492
rect 21407 8452 22284 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 11020 8384 11069 8412
rect 11020 8372 11026 8384
rect 11057 8381 11069 8384
rect 11103 8381 11115 8415
rect 11057 8375 11115 8381
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8381 11299 8415
rect 11241 8375 11299 8381
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 12618 8412 12624 8424
rect 12492 8384 12537 8412
rect 12579 8384 12624 8412
rect 12492 8372 12498 8384
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 16574 8412 16580 8424
rect 16535 8384 16580 8412
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 16942 8421 16948 8424
rect 16916 8415 16948 8421
rect 16916 8381 16928 8415
rect 16916 8375 16948 8381
rect 16942 8372 16948 8375
rect 17000 8372 17006 8424
rect 17126 8412 17132 8424
rect 17039 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8412 17190 8424
rect 18690 8412 18696 8424
rect 17184 8384 18184 8412
rect 18651 8384 18696 8412
rect 17184 8372 17190 8384
rect 2608 8276 2636 8372
rect 18156 8344 18184 8384
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 18984 8344 19012 8443
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 19061 8415 19119 8421
rect 19061 8381 19073 8415
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 18156 8316 19012 8344
rect 19076 8344 19104 8375
rect 20530 8344 20536 8356
rect 19076 8316 20536 8344
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 22738 8304 22744 8356
rect 22796 8344 22802 8356
rect 22925 8347 22983 8353
rect 22925 8344 22937 8347
rect 22796 8316 22937 8344
rect 22796 8304 22802 8316
rect 22925 8313 22937 8316
rect 22971 8344 22983 8347
rect 23566 8344 23572 8356
rect 22971 8316 23572 8344
rect 22971 8313 22983 8316
rect 22925 8307 22983 8313
rect 23566 8304 23572 8316
rect 23624 8304 23630 8356
rect 4154 8276 4160 8288
rect 2608 8248 4160 8276
rect 4154 8236 4160 8248
rect 4212 8276 4218 8288
rect 4433 8279 4491 8285
rect 4433 8276 4445 8279
rect 4212 8248 4445 8276
rect 4212 8236 4218 8248
rect 4433 8245 4445 8248
rect 4479 8276 4491 8279
rect 4798 8276 4804 8288
rect 4479 8248 4804 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 9398 8276 9404 8288
rect 9359 8248 9404 8276
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 16206 8276 16212 8288
rect 16167 8248 16212 8276
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 1104 8186 29256 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 29256 8186
rect 1104 8112 29256 8134
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 16724 8044 17509 8072
rect 16724 8032 16730 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 20530 8032 20536 8084
rect 20588 8072 20594 8084
rect 25041 8075 25099 8081
rect 25041 8072 25053 8075
rect 20588 8044 25053 8072
rect 20588 8032 20594 8044
rect 25041 8041 25053 8044
rect 25087 8041 25099 8075
rect 25041 8035 25099 8041
rect 5813 8007 5871 8013
rect 5813 7973 5825 8007
rect 5859 8004 5871 8007
rect 7282 8004 7288 8016
rect 5859 7976 7288 8004
rect 5859 7973 5871 7976
rect 5813 7967 5871 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 12529 8007 12587 8013
rect 12529 7973 12541 8007
rect 12575 8004 12587 8007
rect 12618 8004 12624 8016
rect 12575 7976 12624 8004
rect 12575 7973 12587 7976
rect 12529 7967 12587 7973
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 7006 7936 7012 7948
rect 4120 7908 7012 7936
rect 4120 7896 4126 7908
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7936 11207 7939
rect 11422 7936 11428 7948
rect 11195 7908 11428 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 16264 7908 16405 7936
rect 16264 7896 16270 7908
rect 16393 7905 16405 7908
rect 16439 7905 16451 7939
rect 16393 7899 16451 7905
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7936 22155 7939
rect 22278 7936 22284 7948
rect 22143 7908 22284 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 22278 7896 22284 7908
rect 22336 7896 22342 7948
rect 4154 7868 4160 7880
rect 4115 7840 4160 7868
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4614 7868 4620 7880
rect 4479 7840 4620 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 10870 7868 10876 7880
rect 10831 7840 10876 7868
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16574 7868 16580 7880
rect 16163 7840 16580 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 16574 7828 16580 7840
rect 16632 7868 16638 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 16632 7840 17969 7868
rect 16632 7828 16638 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 23661 7871 23719 7877
rect 23661 7868 23673 7871
rect 17957 7831 18015 7837
rect 23584 7840 23673 7868
rect 23584 7744 23612 7840
rect 23661 7837 23673 7840
rect 23707 7837 23719 7871
rect 23934 7868 23940 7880
rect 23895 7840 23940 7868
rect 23661 7831 23719 7837
rect 23934 7828 23940 7840
rect 23992 7828 23998 7880
rect 5994 7732 6000 7744
rect 5907 7704 6000 7732
rect 5994 7692 6000 7704
rect 6052 7732 6058 7744
rect 6822 7732 6828 7744
rect 6052 7704 6828 7732
rect 6052 7692 6058 7704
rect 6822 7692 6828 7704
rect 6880 7732 6886 7744
rect 7650 7732 7656 7744
rect 6880 7704 7656 7732
rect 6880 7692 6886 7704
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 12713 7735 12771 7741
rect 12713 7701 12725 7735
rect 12759 7732 12771 7735
rect 12802 7732 12808 7744
rect 12759 7704 12808 7732
rect 12759 7701 12771 7704
rect 12713 7695 12771 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 22741 7735 22799 7741
rect 22741 7701 22753 7735
rect 22787 7732 22799 7735
rect 22830 7732 22836 7744
rect 22787 7704 22836 7732
rect 22787 7701 22799 7704
rect 22741 7695 22799 7701
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 23566 7732 23572 7744
rect 23527 7704 23572 7732
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 1104 7642 29256 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 29256 7642
rect 1104 7568 29256 7590
rect 4614 7528 4620 7540
rect 4575 7500 4620 7528
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4856 7500 4905 7528
rect 4856 7488 4862 7500
rect 4893 7497 4905 7500
rect 4939 7528 4951 7531
rect 5994 7528 6000 7540
rect 4939 7500 6000 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 9217 7531 9275 7537
rect 9217 7497 9229 7531
rect 9263 7528 9275 7531
rect 10962 7528 10968 7540
rect 9263 7500 10968 7528
rect 9263 7497 9275 7500
rect 9217 7491 9275 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 15010 7488 15016 7540
rect 15068 7528 15074 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15068 7500 15301 7528
rect 15068 7488 15074 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 9398 7460 9404 7472
rect 9359 7432 9404 7460
rect 9398 7420 9404 7432
rect 9456 7460 9462 7472
rect 9858 7460 9864 7472
rect 9456 7432 9864 7460
rect 9456 7420 9462 7432
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 4798 7392 4804 7404
rect 3099 7364 4804 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 7650 7392 7656 7404
rect 7563 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7392 7714 7404
rect 9416 7392 9444 7420
rect 7708 7364 9444 7392
rect 15304 7392 15332 7491
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15304 7364 15485 7392
rect 7708 7352 7714 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 21729 7395 21787 7401
rect 21729 7361 21741 7395
rect 21775 7392 21787 7395
rect 22830 7392 22836 7404
rect 21775 7364 22836 7392
rect 21775 7361 21787 7364
rect 21729 7355 21787 7361
rect 22830 7352 22836 7364
rect 22888 7352 22894 7404
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 4706 7324 4712 7336
rect 3375 7296 4712 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7324 7987 7327
rect 8386 7324 8392 7336
rect 7975 7296 8392 7324
rect 7975 7293 7987 7296
rect 7929 7287 7987 7293
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 15580 7296 15761 7324
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 15580 7256 15608 7296
rect 15749 7293 15761 7296
rect 15795 7324 15807 7327
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 15795 7296 22385 7324
rect 15795 7293 15807 7296
rect 15749 7287 15807 7293
rect 22373 7293 22385 7296
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 13872 7228 15608 7256
rect 13872 7216 13878 7228
rect 16942 7148 16948 7200
rect 17000 7188 17006 7200
rect 17037 7191 17095 7197
rect 17037 7188 17049 7191
rect 17000 7160 17049 7188
rect 17000 7148 17006 7160
rect 17037 7157 17049 7160
rect 17083 7157 17095 7191
rect 17037 7151 17095 7157
rect 1104 7098 29256 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 29256 7098
rect 1104 7024 29256 7046
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12713 6987 12771 6993
rect 12713 6984 12725 6987
rect 12308 6956 12725 6984
rect 12308 6944 12314 6956
rect 12713 6953 12725 6956
rect 12759 6953 12771 6987
rect 12713 6947 12771 6953
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 12860 6956 13185 6984
rect 12860 6944 12866 6956
rect 13173 6953 13185 6956
rect 13219 6984 13231 6987
rect 15010 6984 15016 6996
rect 13219 6956 15016 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 16684 6956 18429 6984
rect 4706 6848 4712 6860
rect 4667 6820 4712 6848
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10870 6848 10876 6860
rect 9916 6820 10876 6848
rect 9916 6808 9922 6820
rect 10870 6808 10876 6820
rect 10928 6848 10934 6860
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 10928 6820 11345 6848
rect 10928 6808 10934 6820
rect 11333 6817 11345 6820
rect 11379 6848 11391 6851
rect 11698 6848 11704 6860
rect 11379 6820 11704 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 11698 6808 11704 6820
rect 11756 6848 11762 6860
rect 12820 6848 12848 6944
rect 11756 6820 12848 6848
rect 11756 6808 11762 6820
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16684 6857 16712 6956
rect 18417 6953 18429 6956
rect 18463 6953 18475 6987
rect 23934 6984 23940 6996
rect 23895 6956 23940 6984
rect 18417 6947 18475 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16632 6820 16681 6848
rect 16632 6808 16638 6820
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 16669 6811 16727 6817
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 22830 6848 22836 6860
rect 22791 6820 22836 6848
rect 22830 6808 22836 6820
rect 22888 6808 22894 6860
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 10226 6780 10232 6792
rect 6687 6752 10232 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 4080 6712 4108 6743
rect 10226 6740 10232 6752
rect 10284 6780 10290 6792
rect 10962 6780 10968 6792
rect 10284 6752 10968 6780
rect 10284 6740 10290 6752
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11606 6780 11612 6792
rect 11567 6752 11612 6780
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 17034 6740 17040 6792
rect 17092 6780 17098 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17092 6752 18061 6780
rect 17092 6740 17098 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 22465 6783 22523 6789
rect 22465 6749 22477 6783
rect 22511 6780 22523 6783
rect 22557 6783 22615 6789
rect 22557 6780 22569 6783
rect 22511 6752 22569 6780
rect 22511 6749 22523 6752
rect 22465 6743 22523 6749
rect 22557 6749 22569 6752
rect 22603 6780 22615 6783
rect 23566 6780 23572 6792
rect 22603 6752 23572 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 7098 6712 7104 6724
rect 4080 6684 7104 6712
rect 7098 6672 7104 6684
rect 7156 6712 7162 6724
rect 7285 6715 7343 6721
rect 7285 6712 7297 6715
rect 7156 6684 7297 6712
rect 7156 6672 7162 6684
rect 7285 6681 7297 6684
rect 7331 6681 7343 6715
rect 7285 6675 7343 6681
rect 1104 6554 29256 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 29256 6554
rect 1104 6480 29256 6502
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4798 6440 4804 6452
rect 4479 6412 4804 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 11425 6443 11483 6449
rect 11425 6409 11437 6443
rect 11471 6440 11483 6443
rect 11606 6440 11612 6452
rect 11471 6412 11612 6440
rect 11471 6409 11483 6412
rect 11425 6403 11483 6409
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 11756 6412 11801 6440
rect 11756 6400 11762 6412
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 14369 6375 14427 6381
rect 14369 6372 14381 6375
rect 11020 6344 14381 6372
rect 11020 6332 11026 6344
rect 14369 6341 14381 6344
rect 14415 6341 14427 6375
rect 14369 6335 14427 6341
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 7098 6304 7104 6316
rect 2915 6276 6960 6304
rect 7059 6276 7104 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 2590 6236 2596 6248
rect 2551 6208 2596 6236
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 6822 6236 6828 6248
rect 6783 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 3970 6100 3976 6112
rect 3931 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 6932 6100 6960 6276
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 10226 6264 10232 6316
rect 10284 6264 10290 6316
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 13814 6304 13820 6316
rect 13771 6276 13820 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9858 6236 9864 6248
rect 8711 6208 9864 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6236 10195 6239
rect 10244 6236 10272 6264
rect 10183 6208 10272 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 13170 6100 13176 6112
rect 6932 6072 13176 6100
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 1104 6010 29256 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 29256 6010
rect 1104 5936 29256 5958
rect 26789 5763 26847 5769
rect 26789 5760 26801 5763
rect 26252 5732 26801 5760
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 26252 5701 26280 5732
rect 26789 5729 26801 5732
rect 26835 5729 26847 5763
rect 26789 5723 26847 5729
rect 26237 5695 26295 5701
rect 26237 5692 26249 5695
rect 7800 5664 26249 5692
rect 7800 5652 7806 5664
rect 26237 5661 26249 5664
rect 26283 5661 26295 5695
rect 26237 5655 26295 5661
rect 26513 5695 26571 5701
rect 26513 5661 26525 5695
rect 26559 5661 26571 5695
rect 26513 5655 26571 5661
rect 23566 5584 23572 5636
rect 23624 5624 23630 5636
rect 26145 5627 26203 5633
rect 26145 5624 26157 5627
rect 23624 5596 26157 5624
rect 23624 5584 23630 5596
rect 26145 5593 26157 5596
rect 26191 5624 26203 5627
rect 26528 5624 26556 5655
rect 26191 5596 26556 5624
rect 26191 5593 26203 5596
rect 26145 5587 26203 5593
rect 28077 5559 28135 5565
rect 28077 5525 28089 5559
rect 28123 5556 28135 5559
rect 29914 5556 29920 5568
rect 28123 5528 29920 5556
rect 28123 5525 28135 5528
rect 28077 5519 28135 5525
rect 29914 5516 29920 5528
rect 29972 5516 29978 5568
rect 1104 5466 29256 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 29256 5466
rect 1104 5392 29256 5414
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4798 5352 4804 5364
rect 4479 5324 4804 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 2958 5216 2964 5228
rect 2915 5188 2964 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 2590 5148 2596 5160
rect 2503 5120 2596 5148
rect 2590 5108 2596 5120
rect 2648 5148 2654 5160
rect 3234 5148 3240 5160
rect 2648 5120 3240 5148
rect 2648 5108 2654 5120
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 1104 4922 29256 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 29256 4922
rect 1104 4848 29256 4870
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 6546 4808 6552 4820
rect 4120 4780 6552 4808
rect 4120 4768 4126 4780
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 6880 4780 7665 4808
rect 6880 4768 6886 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 7653 4771 7711 4777
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4672 5963 4675
rect 6840 4672 6868 4768
rect 5951 4644 6868 4672
rect 5951 4641 5963 4644
rect 5905 4635 5963 4641
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 8110 4604 8116 4616
rect 6227 4576 8116 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 7285 4471 7343 4477
rect 7285 4468 7297 4471
rect 5132 4440 7297 4468
rect 5132 4428 5138 4440
rect 7285 4437 7297 4440
rect 7331 4437 7343 4471
rect 7285 4431 7343 4437
rect 1104 4378 29256 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 29256 4378
rect 1104 4304 29256 4326
rect 4798 4264 4804 4276
rect 4759 4236 4804 4264
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 3191 4100 4721 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 4709 4097 4721 4100
rect 4755 4128 4767 4131
rect 6178 4128 6184 4140
rect 4755 4100 6184 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 27154 4088 27160 4140
rect 27212 4128 27218 4140
rect 28074 4128 28080 4140
rect 27212 4100 28080 4128
rect 27212 4088 27218 4100
rect 28074 4088 28080 4100
rect 28132 4088 28138 4140
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 3234 4060 3240 4072
rect 2915 4032 3240 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 4062 3952 4068 4004
rect 4120 3992 4126 4004
rect 7558 3992 7564 4004
rect 4120 3964 7564 3992
rect 4120 3952 4126 3964
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4249 3927 4307 3933
rect 4249 3924 4261 3927
rect 4212 3896 4261 3924
rect 4212 3884 4218 3896
rect 4249 3893 4261 3896
rect 4295 3893 4307 3927
rect 4249 3887 4307 3893
rect 1104 3834 29256 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 29256 3834
rect 1104 3760 29256 3782
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 5074 3516 5080 3528
rect 4028 3488 5080 3516
rect 4028 3476 4034 3488
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 56318 3408 56324 3460
rect 56376 3448 56382 3460
rect 84194 3448 84200 3460
rect 56376 3420 84200 3448
rect 56376 3408 56382 3420
rect 84194 3408 84200 3420
rect 84252 3408 84258 3460
rect 1104 3290 29256 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 29256 3290
rect 1104 3216 29256 3238
rect 4982 3136 4988 3188
rect 5040 3176 5046 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 5040 3148 5089 3176
rect 5040 3136 5046 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 5000 3040 5028 3136
rect 3651 3012 5028 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 3292 2944 3341 2972
rect 3292 2932 3298 2944
rect 3329 2941 3341 2944
rect 3375 2972 3387 2975
rect 4798 2972 4804 2984
rect 3375 2944 4804 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 4798 2932 4804 2944
rect 4856 2972 4862 2984
rect 5261 2975 5319 2981
rect 5261 2972 5273 2975
rect 4856 2944 5273 2972
rect 4856 2932 4862 2944
rect 5261 2941 5273 2944
rect 5307 2941 5319 2975
rect 5261 2935 5319 2941
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 2832 2808 4721 2836
rect 2832 2796 2838 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 4709 2799 4767 2805
rect 1104 2746 29256 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 29256 2746
rect 1104 2672 29256 2694
rect 1104 2202 29256 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 29256 2202
rect 1104 2128 29256 2150
<< via1 >>
rect 4068 44140 4120 44192
rect 67272 44140 67324 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 50326 44038 50378 44090
rect 50390 44038 50442 44090
rect 50454 44038 50506 44090
rect 50518 44038 50570 44090
rect 81046 44038 81098 44090
rect 81110 44038 81162 44090
rect 81174 44038 81226 44090
rect 81238 44038 81290 44090
rect 6276 43911 6328 43920
rect 6276 43877 6285 43911
rect 6285 43877 6319 43911
rect 6319 43877 6328 43911
rect 6276 43868 6328 43877
rect 4620 43664 4672 43716
rect 5540 43707 5592 43716
rect 5540 43673 5549 43707
rect 5549 43673 5583 43707
rect 5583 43673 5592 43707
rect 5540 43664 5592 43673
rect 19432 43800 19484 43852
rect 24216 43843 24268 43852
rect 24216 43809 24225 43843
rect 24225 43809 24259 43843
rect 24259 43809 24268 43843
rect 24216 43800 24268 43809
rect 25596 43800 25648 43852
rect 40500 43868 40552 43920
rect 39028 43843 39080 43852
rect 39028 43809 39037 43843
rect 39037 43809 39071 43843
rect 39071 43809 39080 43843
rect 39028 43800 39080 43809
rect 23848 43732 23900 43784
rect 29000 43732 29052 43784
rect 17040 43664 17092 43716
rect 36820 43664 36872 43716
rect 6920 43596 6972 43648
rect 23848 43639 23900 43648
rect 23848 43605 23857 43639
rect 23857 43605 23891 43639
rect 23891 43605 23900 43639
rect 23848 43596 23900 43605
rect 25596 43639 25648 43648
rect 25596 43605 25605 43639
rect 25605 43605 25639 43639
rect 25639 43605 25648 43639
rect 25596 43596 25648 43605
rect 37648 43596 37700 43648
rect 39396 43707 39448 43716
rect 39396 43673 39405 43707
rect 39405 43673 39439 43707
rect 39439 43673 39448 43707
rect 39396 43664 39448 43673
rect 48044 43800 48096 43852
rect 47676 43732 47728 43784
rect 49792 43800 49844 43852
rect 61936 43843 61988 43852
rect 49148 43732 49200 43784
rect 61936 43809 61945 43843
rect 61945 43809 61979 43843
rect 61979 43809 61988 43843
rect 61936 43800 61988 43809
rect 63040 43800 63092 43852
rect 69112 43800 69164 43852
rect 70308 43800 70360 43852
rect 63500 43664 63552 43716
rect 46756 43596 46808 43648
rect 49240 43596 49292 43648
rect 62212 43639 62264 43648
rect 62212 43605 62221 43639
rect 62221 43605 62255 43639
rect 62255 43605 62264 43639
rect 62212 43596 62264 43605
rect 69756 43639 69808 43648
rect 69756 43605 69765 43639
rect 69765 43605 69799 43639
rect 69799 43605 69808 43639
rect 69756 43596 69808 43605
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 65686 43494 65738 43546
rect 65750 43494 65802 43546
rect 65814 43494 65866 43546
rect 65878 43494 65930 43546
rect 96406 43494 96458 43546
rect 96470 43494 96522 43546
rect 96534 43494 96586 43546
rect 96598 43494 96650 43546
rect 19432 43435 19484 43444
rect 19432 43401 19441 43435
rect 19441 43401 19475 43435
rect 19475 43401 19484 43435
rect 19432 43392 19484 43401
rect 36820 43435 36872 43444
rect 36820 43401 36829 43435
rect 36829 43401 36863 43435
rect 36863 43401 36872 43435
rect 36820 43392 36872 43401
rect 4804 43256 4856 43308
rect 18236 43256 18288 43308
rect 5080 43188 5132 43240
rect 6460 43188 6512 43240
rect 4804 43120 4856 43172
rect 6644 43120 6696 43172
rect 9680 43120 9732 43172
rect 10784 43188 10836 43240
rect 18328 43231 18380 43240
rect 12624 43120 12676 43172
rect 5264 43095 5316 43104
rect 5264 43061 5273 43095
rect 5273 43061 5307 43095
rect 5307 43061 5316 43095
rect 5264 43052 5316 43061
rect 6920 43095 6972 43104
rect 6920 43061 6929 43095
rect 6929 43061 6963 43095
rect 6963 43061 6972 43095
rect 6920 43052 6972 43061
rect 8024 43052 8076 43104
rect 11704 43095 11756 43104
rect 11704 43061 11713 43095
rect 11713 43061 11747 43095
rect 11747 43061 11756 43095
rect 11704 43052 11756 43061
rect 17684 43052 17736 43104
rect 18328 43197 18337 43231
rect 18337 43197 18371 43231
rect 18371 43197 18380 43231
rect 18328 43188 18380 43197
rect 29092 43256 29144 43308
rect 30472 43256 30524 43308
rect 45468 43392 45520 43444
rect 70308 43392 70360 43444
rect 48688 43324 48740 43376
rect 66260 43367 66312 43376
rect 66260 43333 66269 43367
rect 66269 43333 66303 43367
rect 66303 43333 66312 43367
rect 66260 43324 66312 43333
rect 46756 43299 46808 43308
rect 24216 43120 24268 43172
rect 26976 43231 27028 43240
rect 26976 43197 26985 43231
rect 26985 43197 27019 43231
rect 27019 43197 27028 43231
rect 26976 43188 27028 43197
rect 46756 43265 46765 43299
rect 46765 43265 46799 43299
rect 46799 43265 46808 43299
rect 46756 43256 46808 43265
rect 61108 43256 61160 43308
rect 29736 43120 29788 43172
rect 19248 43052 19300 43104
rect 23480 43095 23532 43104
rect 23480 43061 23489 43095
rect 23489 43061 23523 43095
rect 23523 43061 23532 43095
rect 23480 43052 23532 43061
rect 25228 43095 25280 43104
rect 25228 43061 25237 43095
rect 25237 43061 25271 43095
rect 25271 43061 25280 43095
rect 25228 43052 25280 43061
rect 26516 43095 26568 43104
rect 26516 43061 26525 43095
rect 26525 43061 26559 43095
rect 26559 43061 26568 43095
rect 26516 43052 26568 43061
rect 34796 43120 34848 43172
rect 39028 43188 39080 43240
rect 40500 43231 40552 43240
rect 40500 43197 40509 43231
rect 40509 43197 40543 43231
rect 40543 43197 40552 43231
rect 40500 43188 40552 43197
rect 38476 43163 38528 43172
rect 38476 43129 38485 43163
rect 38485 43129 38519 43163
rect 38519 43129 38528 43163
rect 38476 43120 38528 43129
rect 38568 43120 38620 43172
rect 43444 43188 43496 43240
rect 48964 43188 49016 43240
rect 49240 43231 49292 43240
rect 34152 43095 34204 43104
rect 34152 43061 34161 43095
rect 34161 43061 34195 43095
rect 34195 43061 34204 43095
rect 34152 43052 34204 43061
rect 39028 43052 39080 43104
rect 43720 43095 43772 43104
rect 43720 43061 43729 43095
rect 43729 43061 43763 43095
rect 43763 43061 43772 43095
rect 43720 43052 43772 43061
rect 47676 43052 47728 43104
rect 47860 43095 47912 43104
rect 47860 43061 47869 43095
rect 47869 43061 47903 43095
rect 47903 43061 47912 43095
rect 47860 43052 47912 43061
rect 49240 43197 49249 43231
rect 49249 43197 49283 43231
rect 49283 43197 49292 43231
rect 49240 43188 49292 43197
rect 49792 43188 49844 43240
rect 50804 43188 50856 43240
rect 55772 43231 55824 43240
rect 55772 43197 55781 43231
rect 55781 43197 55815 43231
rect 55815 43197 55824 43231
rect 55772 43188 55824 43197
rect 56232 43231 56284 43240
rect 49332 43120 49384 43172
rect 55220 43163 55272 43172
rect 55220 43129 55229 43163
rect 55229 43129 55263 43163
rect 55263 43129 55272 43163
rect 55220 43120 55272 43129
rect 56232 43197 56241 43231
rect 56241 43197 56275 43231
rect 56275 43197 56284 43231
rect 56232 43188 56284 43197
rect 59544 43231 59596 43240
rect 59544 43197 59553 43231
rect 59553 43197 59587 43231
rect 59587 43197 59596 43231
rect 59544 43188 59596 43197
rect 66536 43231 66588 43240
rect 56600 43120 56652 43172
rect 57888 43120 57940 43172
rect 66536 43197 66545 43231
rect 66545 43197 66579 43231
rect 66579 43197 66588 43231
rect 66536 43188 66588 43197
rect 66904 43231 66956 43240
rect 66904 43197 66913 43231
rect 66913 43197 66947 43231
rect 66947 43197 66956 43231
rect 66904 43188 66956 43197
rect 69388 43231 69440 43240
rect 49976 43052 50028 43104
rect 60832 43095 60884 43104
rect 60832 43061 60841 43095
rect 60841 43061 60875 43095
rect 60875 43061 60884 43095
rect 60832 43052 60884 43061
rect 61108 43095 61160 43104
rect 61108 43061 61117 43095
rect 61117 43061 61151 43095
rect 61151 43061 61160 43095
rect 61108 43052 61160 43061
rect 66168 43052 66220 43104
rect 69388 43197 69397 43231
rect 69397 43197 69431 43231
rect 69431 43197 69440 43231
rect 69388 43188 69440 43197
rect 69664 43052 69716 43104
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 50326 42950 50378 43002
rect 50390 42950 50442 43002
rect 50454 42950 50506 43002
rect 50518 42950 50570 43002
rect 81046 42950 81098 43002
rect 81110 42950 81162 43002
rect 81174 42950 81226 43002
rect 81238 42950 81290 43002
rect 6644 42891 6696 42900
rect 6644 42857 6653 42891
rect 6653 42857 6687 42891
rect 6687 42857 6696 42891
rect 6644 42848 6696 42857
rect 6460 42823 6512 42832
rect 6460 42789 6469 42823
rect 6469 42789 6503 42823
rect 6503 42789 6512 42823
rect 6460 42780 6512 42789
rect 4804 42755 4856 42764
rect 4804 42721 4813 42755
rect 4813 42721 4847 42755
rect 4847 42721 4856 42755
rect 4804 42712 4856 42721
rect 5540 42712 5592 42764
rect 9680 42712 9732 42764
rect 14096 42712 14148 42764
rect 15660 42755 15712 42764
rect 15660 42721 15669 42755
rect 15669 42721 15703 42755
rect 15703 42721 15712 42755
rect 15660 42712 15712 42721
rect 18420 42848 18472 42900
rect 19984 42848 20036 42900
rect 25228 42848 25280 42900
rect 38568 42848 38620 42900
rect 40500 42848 40552 42900
rect 44916 42848 44968 42900
rect 50804 42891 50856 42900
rect 50804 42857 50813 42891
rect 50813 42857 50847 42891
rect 50847 42857 50856 42891
rect 50804 42848 50856 42857
rect 55772 42848 55824 42900
rect 17040 42780 17092 42832
rect 10692 42687 10744 42696
rect 10692 42653 10701 42687
rect 10701 42653 10735 42687
rect 10735 42653 10744 42687
rect 10692 42644 10744 42653
rect 11704 42644 11756 42696
rect 15016 42644 15068 42696
rect 18328 42712 18380 42764
rect 23112 42712 23164 42764
rect 25596 42780 25648 42832
rect 17040 42687 17092 42696
rect 17040 42653 17049 42687
rect 17049 42653 17083 42687
rect 17083 42653 17092 42687
rect 17040 42644 17092 42653
rect 17684 42687 17736 42696
rect 17684 42653 17693 42687
rect 17693 42653 17727 42687
rect 17727 42653 17736 42687
rect 17684 42644 17736 42653
rect 17960 42687 18012 42696
rect 17960 42653 17969 42687
rect 17969 42653 18003 42687
rect 18003 42653 18012 42687
rect 17960 42644 18012 42653
rect 19340 42687 19392 42696
rect 19340 42653 19349 42687
rect 19349 42653 19383 42687
rect 19383 42653 19392 42687
rect 19340 42644 19392 42653
rect 23388 42644 23440 42696
rect 23848 42687 23900 42696
rect 23848 42653 23857 42687
rect 23857 42653 23891 42687
rect 23891 42653 23900 42687
rect 23848 42644 23900 42653
rect 25228 42712 25280 42764
rect 29000 42755 29052 42764
rect 26976 42644 27028 42696
rect 29000 42721 29009 42755
rect 29009 42721 29043 42755
rect 29043 42721 29052 42755
rect 29000 42712 29052 42721
rect 29092 42712 29144 42764
rect 35440 42712 35492 42764
rect 44088 42712 44140 42764
rect 44364 42712 44416 42764
rect 45284 42755 45336 42764
rect 45284 42721 45293 42755
rect 45293 42721 45327 42755
rect 45327 42721 45336 42755
rect 45284 42712 45336 42721
rect 30380 42687 30432 42696
rect 6920 42508 6972 42560
rect 12164 42508 12216 42560
rect 12256 42508 12308 42560
rect 17592 42508 17644 42560
rect 19248 42508 19300 42560
rect 23296 42551 23348 42560
rect 23296 42517 23305 42551
rect 23305 42517 23339 42551
rect 23339 42517 23348 42551
rect 23296 42508 23348 42517
rect 23572 42508 23624 42560
rect 30380 42653 30389 42687
rect 30389 42653 30423 42687
rect 30423 42653 30432 42687
rect 30380 42644 30432 42653
rect 34152 42644 34204 42696
rect 34428 42644 34480 42696
rect 43444 42687 43496 42696
rect 26516 42508 26568 42560
rect 31576 42508 31628 42560
rect 35532 42576 35584 42628
rect 35348 42508 35400 42560
rect 37832 42551 37884 42560
rect 37832 42517 37841 42551
rect 37841 42517 37875 42551
rect 37875 42517 37884 42551
rect 37832 42508 37884 42517
rect 43444 42653 43453 42687
rect 43453 42653 43487 42687
rect 43487 42653 43496 42687
rect 43444 42644 43496 42653
rect 43904 42644 43956 42696
rect 46756 42712 46808 42764
rect 47676 42755 47728 42764
rect 45836 42687 45888 42696
rect 45836 42653 45845 42687
rect 45845 42653 45879 42687
rect 45879 42653 45888 42687
rect 45836 42644 45888 42653
rect 47676 42721 47685 42755
rect 47685 42721 47719 42755
rect 47719 42721 47728 42755
rect 47676 42712 47728 42721
rect 49332 42780 49384 42832
rect 48688 42644 48740 42696
rect 49056 42712 49108 42764
rect 49332 42644 49384 42696
rect 50620 42712 50672 42764
rect 53748 42644 53800 42696
rect 55220 42644 55272 42696
rect 56232 42712 56284 42764
rect 57888 42712 57940 42764
rect 60832 42712 60884 42764
rect 62212 42712 62264 42764
rect 63500 42712 63552 42764
rect 64604 42712 64656 42764
rect 69204 42755 69256 42764
rect 58532 42644 58584 42696
rect 61108 42644 61160 42696
rect 66076 42687 66128 42696
rect 45468 42576 45520 42628
rect 49148 42576 49200 42628
rect 44548 42508 44600 42560
rect 49976 42508 50028 42560
rect 51080 42508 51132 42560
rect 59452 42576 59504 42628
rect 55956 42508 56008 42560
rect 58532 42551 58584 42560
rect 58532 42517 58541 42551
rect 58541 42517 58575 42551
rect 58575 42517 58584 42551
rect 58532 42508 58584 42517
rect 60372 42551 60424 42560
rect 60372 42517 60381 42551
rect 60381 42517 60415 42551
rect 60415 42517 60424 42551
rect 60372 42508 60424 42517
rect 60832 42508 60884 42560
rect 66076 42653 66085 42687
rect 66085 42653 66119 42687
rect 66119 42653 66128 42687
rect 66076 42644 66128 42653
rect 69204 42721 69213 42755
rect 69213 42721 69247 42755
rect 69247 42721 69256 42755
rect 69204 42712 69256 42721
rect 69296 42755 69348 42764
rect 69296 42721 69305 42755
rect 69305 42721 69339 42755
rect 69339 42721 69348 42755
rect 71412 42755 71464 42764
rect 69296 42712 69348 42721
rect 71412 42721 71421 42755
rect 71421 42721 71455 42755
rect 71455 42721 71464 42755
rect 71412 42712 71464 42721
rect 70400 42644 70452 42696
rect 66812 42576 66864 42628
rect 69664 42576 69716 42628
rect 66996 42508 67048 42560
rect 69388 42508 69440 42560
rect 70032 42508 70084 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 65686 42406 65738 42458
rect 65750 42406 65802 42458
rect 65814 42406 65866 42458
rect 65878 42406 65930 42458
rect 96406 42406 96458 42458
rect 96470 42406 96522 42458
rect 96534 42406 96586 42458
rect 96598 42406 96650 42458
rect 2412 42347 2464 42356
rect 2412 42313 2421 42347
rect 2421 42313 2455 42347
rect 2455 42313 2464 42347
rect 2412 42304 2464 42313
rect 4804 42304 4856 42356
rect 6276 42236 6328 42288
rect 9956 42236 10008 42288
rect 6092 42168 6144 42220
rect 10784 42279 10836 42288
rect 10784 42245 10793 42279
rect 10793 42245 10827 42279
rect 10827 42245 10836 42279
rect 10784 42236 10836 42245
rect 12532 42304 12584 42356
rect 18420 42304 18472 42356
rect 23296 42347 23348 42356
rect 23296 42313 23305 42347
rect 23305 42313 23339 42347
rect 23339 42313 23348 42347
rect 23296 42304 23348 42313
rect 23664 42304 23716 42356
rect 24584 42304 24636 42356
rect 25412 42304 25464 42356
rect 51080 42304 51132 42356
rect 63040 42347 63092 42356
rect 23480 42236 23532 42288
rect 2412 42100 2464 42152
rect 2872 42143 2924 42152
rect 2872 42109 2881 42143
rect 2881 42109 2915 42143
rect 2915 42109 2924 42143
rect 2872 42100 2924 42109
rect 5264 42143 5316 42152
rect 5264 42109 5273 42143
rect 5273 42109 5307 42143
rect 5307 42109 5316 42143
rect 5264 42100 5316 42109
rect 10416 42143 10468 42152
rect 8024 42032 8076 42084
rect 9588 42032 9640 42084
rect 3976 42007 4028 42016
rect 3976 41973 3985 42007
rect 3985 41973 4019 42007
rect 4019 41973 4028 42007
rect 3976 41964 4028 41973
rect 5172 41964 5224 42016
rect 9496 42007 9548 42016
rect 9496 41973 9505 42007
rect 9505 41973 9539 42007
rect 9539 41973 9548 42007
rect 10416 42109 10425 42143
rect 10425 42109 10459 42143
rect 10459 42109 10468 42143
rect 10416 42100 10468 42109
rect 9496 41964 9548 41973
rect 10232 41964 10284 42016
rect 12624 42100 12676 42152
rect 13636 42168 13688 42220
rect 16856 42168 16908 42220
rect 17224 42211 17276 42220
rect 16396 42143 16448 42152
rect 15292 42032 15344 42084
rect 16396 42109 16405 42143
rect 16405 42109 16439 42143
rect 16439 42109 16448 42143
rect 16396 42100 16448 42109
rect 16580 42143 16632 42152
rect 16580 42109 16589 42143
rect 16589 42109 16623 42143
rect 16623 42109 16632 42143
rect 16580 42100 16632 42109
rect 17224 42177 17233 42211
rect 17233 42177 17267 42211
rect 17267 42177 17276 42211
rect 17224 42168 17276 42177
rect 17500 42211 17552 42220
rect 17500 42177 17509 42211
rect 17509 42177 17543 42211
rect 17543 42177 17552 42211
rect 17500 42168 17552 42177
rect 18328 42168 18380 42220
rect 17684 42100 17736 42152
rect 12532 42007 12584 42016
rect 12532 41973 12541 42007
rect 12541 41973 12575 42007
rect 12575 41973 12584 42007
rect 12532 41964 12584 41973
rect 15200 41964 15252 42016
rect 16580 41964 16632 42016
rect 17592 42007 17644 42016
rect 17592 41973 17601 42007
rect 17601 41973 17635 42007
rect 17635 41973 17644 42007
rect 17592 41964 17644 41973
rect 17776 42007 17828 42016
rect 17776 41973 17785 42007
rect 17785 41973 17819 42007
rect 17819 41973 17828 42007
rect 23572 42168 23624 42220
rect 23940 42236 23992 42288
rect 44088 42279 44140 42288
rect 25872 42168 25924 42220
rect 19340 42100 19392 42152
rect 23296 42100 23348 42152
rect 24584 42143 24636 42152
rect 24584 42109 24593 42143
rect 24593 42109 24627 42143
rect 24627 42109 24636 42143
rect 24584 42100 24636 42109
rect 25688 42100 25740 42152
rect 31576 42168 31628 42220
rect 44088 42245 44097 42279
rect 44097 42245 44131 42279
rect 44131 42245 44140 42279
rect 44088 42236 44140 42245
rect 45100 42236 45152 42288
rect 20260 42032 20312 42084
rect 23756 42032 23808 42084
rect 17776 41964 17828 41973
rect 23112 41964 23164 42016
rect 23572 41964 23624 42016
rect 27252 42075 27304 42084
rect 27252 42041 27261 42075
rect 27261 42041 27295 42075
rect 27295 42041 27304 42075
rect 27252 42032 27304 42041
rect 34796 42100 34848 42152
rect 32588 42032 32640 42084
rect 35900 42032 35952 42084
rect 36728 42100 36780 42152
rect 48044 42211 48096 42220
rect 48044 42177 48053 42211
rect 48053 42177 48087 42211
rect 48087 42177 48096 42211
rect 48044 42168 48096 42177
rect 37280 42100 37332 42152
rect 39764 42100 39816 42152
rect 37740 42075 37792 42084
rect 25688 41964 25740 42016
rect 25872 41964 25924 42016
rect 30472 41964 30524 42016
rect 30564 41964 30616 42016
rect 37740 42041 37749 42075
rect 37749 42041 37783 42075
rect 37783 42041 37792 42075
rect 37740 42032 37792 42041
rect 37832 42032 37884 42084
rect 44364 42100 44416 42152
rect 44456 42100 44508 42152
rect 44824 42100 44876 42152
rect 36912 41964 36964 42016
rect 38936 41964 38988 42016
rect 43812 42007 43864 42016
rect 43812 41973 43821 42007
rect 43821 41973 43855 42007
rect 43855 41973 43864 42007
rect 43812 41964 43864 41973
rect 44916 42032 44968 42084
rect 45468 42100 45520 42152
rect 48688 42143 48740 42152
rect 48688 42109 48697 42143
rect 48697 42109 48731 42143
rect 48731 42109 48740 42143
rect 48688 42100 48740 42109
rect 49148 42236 49200 42288
rect 63040 42313 63049 42347
rect 63049 42313 63083 42347
rect 63083 42313 63092 42347
rect 63040 42304 63092 42313
rect 69296 42347 69348 42356
rect 69296 42313 69305 42347
rect 69305 42313 69339 42347
rect 69339 42313 69348 42347
rect 69296 42304 69348 42313
rect 59176 42236 59228 42288
rect 48964 42168 49016 42220
rect 53748 42168 53800 42220
rect 49056 42143 49108 42152
rect 45192 42032 45244 42084
rect 49056 42109 49065 42143
rect 49065 42109 49099 42143
rect 49099 42109 49108 42143
rect 49056 42100 49108 42109
rect 49332 42100 49384 42152
rect 50620 42100 50672 42152
rect 52000 42143 52052 42152
rect 52000 42109 52009 42143
rect 52009 42109 52043 42143
rect 52043 42109 52052 42143
rect 52000 42100 52052 42109
rect 56140 42168 56192 42220
rect 59452 42236 59504 42288
rect 65708 42236 65760 42288
rect 55956 42143 56008 42152
rect 55956 42109 55965 42143
rect 55965 42109 55999 42143
rect 55999 42109 56008 42143
rect 55956 42100 56008 42109
rect 58532 42100 58584 42152
rect 61016 42168 61068 42220
rect 61936 42211 61988 42220
rect 61936 42177 61945 42211
rect 61945 42177 61979 42211
rect 61979 42177 61988 42211
rect 61936 42168 61988 42177
rect 49424 42075 49476 42084
rect 49424 42041 49433 42075
rect 49433 42041 49467 42075
rect 49467 42041 49476 42075
rect 49424 42032 49476 42041
rect 55036 42075 55088 42084
rect 55036 42041 55045 42075
rect 55045 42041 55079 42075
rect 55079 42041 55088 42075
rect 55036 42032 55088 42041
rect 61568 42100 61620 42152
rect 61752 42100 61804 42152
rect 63868 42168 63920 42220
rect 66076 42168 66128 42220
rect 66260 42168 66312 42220
rect 66904 42168 66956 42220
rect 69204 42168 69256 42220
rect 69664 42168 69716 42220
rect 72516 42168 72568 42220
rect 69756 42143 69808 42152
rect 49148 41964 49200 42016
rect 52276 41964 52328 42016
rect 55404 41964 55456 42016
rect 56232 41964 56284 42016
rect 59636 42007 59688 42016
rect 59636 41973 59645 42007
rect 59645 41973 59679 42007
rect 59679 41973 59688 42007
rect 59636 41964 59688 41973
rect 62028 42032 62080 42084
rect 65984 42032 66036 42084
rect 66536 42032 66588 42084
rect 69756 42109 69765 42143
rect 69765 42109 69799 42143
rect 69799 42109 69808 42143
rect 69756 42100 69808 42109
rect 71136 42143 71188 42152
rect 71136 42109 71145 42143
rect 71145 42109 71179 42143
rect 71179 42109 71188 42143
rect 71136 42100 71188 42109
rect 70308 42032 70360 42084
rect 66168 41964 66220 42016
rect 71412 41964 71464 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 50326 41862 50378 41914
rect 50390 41862 50442 41914
rect 50454 41862 50506 41914
rect 50518 41862 50570 41914
rect 81046 41862 81098 41914
rect 81110 41862 81162 41914
rect 81174 41862 81226 41914
rect 81238 41862 81290 41914
rect 5080 41760 5132 41812
rect 10416 41760 10468 41812
rect 10692 41760 10744 41812
rect 10968 41760 11020 41812
rect 12256 41760 12308 41812
rect 4620 41624 4672 41676
rect 8116 41692 8168 41744
rect 9496 41692 9548 41744
rect 5172 41624 5224 41676
rect 8024 41667 8076 41676
rect 8024 41633 8033 41667
rect 8033 41633 8067 41667
rect 8067 41633 8076 41667
rect 8024 41624 8076 41633
rect 8300 41624 8352 41676
rect 8668 41624 8720 41676
rect 9772 41692 9824 41744
rect 5356 41556 5408 41608
rect 9956 41624 10008 41676
rect 10416 41667 10468 41676
rect 10416 41633 10425 41667
rect 10425 41633 10459 41667
rect 10459 41633 10468 41667
rect 10416 41624 10468 41633
rect 10968 41624 11020 41676
rect 11520 41692 11572 41744
rect 14648 41692 14700 41744
rect 13820 41624 13872 41676
rect 15016 41760 15068 41812
rect 16856 41760 16908 41812
rect 17776 41760 17828 41812
rect 17960 41803 18012 41812
rect 17960 41769 17969 41803
rect 17969 41769 18003 41803
rect 18003 41769 18012 41803
rect 17960 41760 18012 41769
rect 18328 41803 18380 41812
rect 18328 41769 18337 41803
rect 18337 41769 18371 41803
rect 18371 41769 18380 41803
rect 18328 41760 18380 41769
rect 20260 41760 20312 41812
rect 23756 41760 23808 41812
rect 23940 41692 23992 41744
rect 8852 41488 8904 41540
rect 9956 41488 10008 41540
rect 14924 41556 14976 41608
rect 17316 41624 17368 41676
rect 17500 41667 17552 41676
rect 17500 41633 17509 41667
rect 17509 41633 17543 41667
rect 17543 41633 17552 41667
rect 17500 41624 17552 41633
rect 17592 41624 17644 41676
rect 17868 41624 17920 41676
rect 23388 41624 23440 41676
rect 23480 41624 23532 41676
rect 24676 41692 24728 41744
rect 25688 41692 25740 41744
rect 30564 41692 30616 41744
rect 31668 41692 31720 41744
rect 35348 41692 35400 41744
rect 23572 41556 23624 41608
rect 24492 41667 24544 41676
rect 24492 41633 24501 41667
rect 24501 41633 24535 41667
rect 24535 41633 24544 41667
rect 24492 41624 24544 41633
rect 25412 41667 25464 41676
rect 25412 41633 25421 41667
rect 25421 41633 25455 41667
rect 25455 41633 25464 41667
rect 25412 41624 25464 41633
rect 26240 41667 26292 41676
rect 26240 41633 26249 41667
rect 26249 41633 26283 41667
rect 26283 41633 26292 41667
rect 26240 41624 26292 41633
rect 29736 41624 29788 41676
rect 30380 41624 30432 41676
rect 30932 41624 30984 41676
rect 35440 41667 35492 41676
rect 35440 41633 35449 41667
rect 35449 41633 35483 41667
rect 35483 41633 35492 41667
rect 35440 41624 35492 41633
rect 35992 41624 36044 41676
rect 37096 41692 37148 41744
rect 37280 41760 37332 41812
rect 37648 41692 37700 41744
rect 36268 41624 36320 41676
rect 38108 41692 38160 41744
rect 38660 41692 38712 41744
rect 43720 41760 43772 41812
rect 44548 41803 44600 41812
rect 44548 41769 44557 41803
rect 44557 41769 44591 41803
rect 44591 41769 44600 41803
rect 44548 41760 44600 41769
rect 45100 41760 45152 41812
rect 49056 41803 49108 41812
rect 44732 41692 44784 41744
rect 49056 41769 49065 41803
rect 49065 41769 49099 41803
rect 49099 41769 49108 41803
rect 49056 41760 49108 41769
rect 51632 41760 51684 41812
rect 52000 41760 52052 41812
rect 58808 41760 58860 41812
rect 59176 41803 59228 41812
rect 59176 41769 59185 41803
rect 59185 41769 59219 41803
rect 59219 41769 59228 41803
rect 59176 41760 59228 41769
rect 63868 41803 63920 41812
rect 51448 41692 51500 41744
rect 43536 41667 43588 41676
rect 43536 41633 43545 41667
rect 43545 41633 43579 41667
rect 43579 41633 43588 41667
rect 43536 41624 43588 41633
rect 43904 41667 43956 41676
rect 43904 41633 43913 41667
rect 43913 41633 43947 41667
rect 43947 41633 43956 41667
rect 43904 41624 43956 41633
rect 9128 41463 9180 41472
rect 9128 41429 9137 41463
rect 9137 41429 9171 41463
rect 9171 41429 9180 41463
rect 9128 41420 9180 41429
rect 10416 41420 10468 41472
rect 11520 41463 11572 41472
rect 11520 41429 11529 41463
rect 11529 41429 11563 41463
rect 11563 41429 11572 41463
rect 11520 41420 11572 41429
rect 13360 41420 13412 41472
rect 13728 41420 13780 41472
rect 14188 41463 14240 41472
rect 14188 41429 14197 41463
rect 14197 41429 14231 41463
rect 14231 41429 14240 41463
rect 14188 41420 14240 41429
rect 15660 41420 15712 41472
rect 18052 41488 18104 41540
rect 23940 41488 23992 41540
rect 26792 41556 26844 41608
rect 31576 41556 31628 41608
rect 37280 41599 37332 41608
rect 26516 41488 26568 41540
rect 37280 41565 37289 41599
rect 37289 41565 37323 41599
rect 37323 41565 37332 41599
rect 37280 41556 37332 41565
rect 45836 41624 45888 41676
rect 45928 41624 45980 41676
rect 47860 41624 47912 41676
rect 51724 41624 51776 41676
rect 53288 41624 53340 41676
rect 17316 41420 17368 41472
rect 17960 41420 18012 41472
rect 18512 41463 18564 41472
rect 18512 41429 18521 41463
rect 18521 41429 18555 41463
rect 18555 41429 18564 41463
rect 18512 41420 18564 41429
rect 23480 41420 23532 41472
rect 24492 41420 24544 41472
rect 25504 41463 25556 41472
rect 25504 41429 25513 41463
rect 25513 41429 25547 41463
rect 25547 41429 25556 41463
rect 25504 41420 25556 41429
rect 25596 41420 25648 41472
rect 37648 41488 37700 41540
rect 37464 41463 37516 41472
rect 37464 41429 37473 41463
rect 37473 41429 37507 41463
rect 37507 41429 37516 41463
rect 38292 41488 38344 41540
rect 37464 41420 37516 41429
rect 38108 41420 38160 41472
rect 44548 41488 44600 41540
rect 51540 41556 51592 41608
rect 52184 41556 52236 41608
rect 54576 41667 54628 41676
rect 54576 41633 54585 41667
rect 54585 41633 54619 41667
rect 54619 41633 54628 41667
rect 54576 41624 54628 41633
rect 57152 41624 57204 41676
rect 59544 41692 59596 41744
rect 59636 41624 59688 41676
rect 61016 41667 61068 41676
rect 61016 41633 61025 41667
rect 61025 41633 61059 41667
rect 61059 41633 61068 41667
rect 61016 41624 61068 41633
rect 63868 41769 63877 41803
rect 63877 41769 63911 41803
rect 63911 41769 63920 41803
rect 63868 41760 63920 41769
rect 69756 41692 69808 41744
rect 50620 41488 50672 41540
rect 60372 41556 60424 41608
rect 63592 41667 63644 41676
rect 63592 41633 63601 41667
rect 63601 41633 63635 41667
rect 63635 41633 63644 41667
rect 63592 41624 63644 41633
rect 62580 41556 62632 41608
rect 62028 41488 62080 41540
rect 65708 41624 65760 41676
rect 66996 41667 67048 41676
rect 66996 41633 67005 41667
rect 67005 41633 67039 41667
rect 67039 41633 67048 41667
rect 66996 41624 67048 41633
rect 68652 41667 68704 41676
rect 68100 41556 68152 41608
rect 68652 41633 68661 41667
rect 68661 41633 68695 41667
rect 68695 41633 68704 41667
rect 68652 41624 68704 41633
rect 69204 41624 69256 41676
rect 69848 41667 69900 41676
rect 69848 41633 69857 41667
rect 69857 41633 69891 41667
rect 69891 41633 69900 41667
rect 69848 41624 69900 41633
rect 70032 41667 70084 41676
rect 70032 41633 70041 41667
rect 70041 41633 70075 41667
rect 70075 41633 70084 41667
rect 70032 41624 70084 41633
rect 71412 41667 71464 41676
rect 71412 41633 71421 41667
rect 71421 41633 71455 41667
rect 71455 41633 71464 41667
rect 71412 41624 71464 41633
rect 70308 41599 70360 41608
rect 70308 41565 70317 41599
rect 70317 41565 70351 41599
rect 70351 41565 70360 41599
rect 70308 41556 70360 41565
rect 78220 41599 78272 41608
rect 64512 41488 64564 41540
rect 78220 41565 78229 41599
rect 78229 41565 78263 41599
rect 78263 41565 78272 41599
rect 78220 41556 78272 41565
rect 45008 41420 45060 41472
rect 46756 41420 46808 41472
rect 52184 41420 52236 41472
rect 52552 41420 52604 41472
rect 54668 41420 54720 41472
rect 55404 41420 55456 41472
rect 55496 41463 55548 41472
rect 55496 41429 55505 41463
rect 55505 41429 55539 41463
rect 55539 41429 55548 41463
rect 55496 41420 55548 41429
rect 63040 41420 63092 41472
rect 65984 41463 66036 41472
rect 65984 41429 65993 41463
rect 65993 41429 66027 41463
rect 66027 41429 66036 41463
rect 65984 41420 66036 41429
rect 69020 41420 69072 41472
rect 70032 41420 70084 41472
rect 71596 41463 71648 41472
rect 71596 41429 71605 41463
rect 71605 41429 71639 41463
rect 71639 41429 71648 41463
rect 71596 41420 71648 41429
rect 72516 41420 72568 41472
rect 77944 41420 77996 41472
rect 79784 41420 79836 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 65686 41318 65738 41370
rect 65750 41318 65802 41370
rect 65814 41318 65866 41370
rect 65878 41318 65930 41370
rect 96406 41318 96458 41370
rect 96470 41318 96522 41370
rect 96534 41318 96586 41370
rect 96598 41318 96650 41370
rect 10232 41259 10284 41268
rect 10232 41225 10241 41259
rect 10241 41225 10275 41259
rect 10275 41225 10284 41259
rect 10232 41216 10284 41225
rect 3608 41012 3660 41064
rect 3884 41055 3936 41064
rect 3884 41021 3893 41055
rect 3893 41021 3927 41055
rect 3927 41021 3936 41055
rect 3884 41012 3936 41021
rect 5448 41055 5500 41064
rect 4620 40944 4672 40996
rect 5448 41021 5457 41055
rect 5457 41021 5491 41055
rect 5491 41021 5500 41055
rect 5448 41012 5500 41021
rect 8300 41012 8352 41064
rect 9128 41012 9180 41064
rect 7288 40944 7340 40996
rect 8852 40987 8904 40996
rect 8852 40953 8861 40987
rect 8861 40953 8895 40987
rect 8895 40953 8904 40987
rect 8852 40944 8904 40953
rect 3884 40876 3936 40928
rect 8024 40876 8076 40928
rect 9956 41012 10008 41064
rect 10968 41148 11020 41200
rect 13084 41216 13136 41268
rect 15200 41216 15252 41268
rect 17500 41216 17552 41268
rect 18236 41259 18288 41268
rect 18236 41225 18245 41259
rect 18245 41225 18279 41259
rect 18279 41225 18288 41259
rect 18236 41216 18288 41225
rect 18512 41216 18564 41268
rect 23388 41216 23440 41268
rect 17960 41148 18012 41200
rect 23940 41216 23992 41268
rect 29828 41259 29880 41268
rect 29828 41225 29837 41259
rect 29837 41225 29871 41259
rect 29871 41225 29880 41259
rect 29828 41216 29880 41225
rect 12808 41080 12860 41132
rect 26240 41148 26292 41200
rect 12716 41055 12768 41064
rect 12716 41021 12725 41055
rect 12725 41021 12759 41055
rect 12759 41021 12768 41055
rect 12716 41012 12768 41021
rect 10508 40919 10560 40928
rect 10508 40885 10517 40919
rect 10517 40885 10551 40919
rect 10551 40885 10560 40919
rect 10508 40876 10560 40885
rect 13636 40876 13688 40928
rect 14004 40919 14056 40928
rect 14004 40885 14013 40919
rect 14013 40885 14047 40919
rect 14047 40885 14056 40919
rect 14004 40876 14056 40885
rect 16948 41012 17000 41064
rect 20904 41012 20956 41064
rect 23664 41012 23716 41064
rect 24124 41055 24176 41064
rect 24124 41021 24133 41055
rect 24133 41021 24167 41055
rect 24167 41021 24176 41055
rect 24124 41012 24176 41021
rect 25504 41080 25556 41132
rect 27344 41080 27396 41132
rect 24676 41055 24728 41064
rect 24676 41021 24685 41055
rect 24685 41021 24719 41055
rect 24719 41021 24728 41055
rect 24676 41012 24728 41021
rect 26240 41012 26292 41064
rect 31576 41216 31628 41268
rect 44640 41216 44692 41268
rect 44732 41216 44784 41268
rect 45468 41216 45520 41268
rect 51816 41216 51868 41268
rect 53104 41216 53156 41268
rect 54576 41216 54628 41268
rect 63500 41216 63552 41268
rect 64696 41216 64748 41268
rect 68100 41259 68152 41268
rect 68100 41225 68109 41259
rect 68109 41225 68143 41259
rect 68143 41225 68152 41259
rect 68100 41216 68152 41225
rect 68652 41216 68704 41268
rect 69020 41216 69072 41268
rect 27620 41080 27672 41132
rect 16396 40876 16448 40928
rect 21732 40876 21784 40928
rect 30012 40944 30064 40996
rect 30656 41055 30708 41064
rect 24124 40876 24176 40928
rect 24584 40876 24636 40928
rect 25228 40876 25280 40928
rect 25688 40876 25740 40928
rect 25872 40876 25924 40928
rect 30656 41021 30665 41055
rect 30665 41021 30699 41055
rect 30699 41021 30708 41055
rect 30656 41012 30708 41021
rect 36176 41148 36228 41200
rect 38568 41148 38620 41200
rect 60648 41148 60700 41200
rect 62028 41148 62080 41200
rect 63040 41191 63092 41200
rect 63040 41157 63049 41191
rect 63049 41157 63083 41191
rect 63083 41157 63092 41191
rect 63040 41148 63092 41157
rect 63132 41148 63184 41200
rect 34796 41080 34848 41132
rect 35992 41080 36044 41132
rect 38476 41123 38528 41132
rect 38476 41089 38485 41123
rect 38485 41089 38519 41123
rect 38519 41089 38528 41123
rect 38476 41080 38528 41089
rect 32680 40944 32732 40996
rect 36268 41012 36320 41064
rect 36452 41012 36504 41064
rect 36636 41055 36688 41064
rect 36636 41021 36645 41055
rect 36645 41021 36679 41055
rect 36679 41021 36688 41055
rect 36636 41012 36688 41021
rect 37740 41012 37792 41064
rect 38660 41080 38712 41132
rect 39028 41080 39080 41132
rect 43720 41012 43772 41064
rect 43812 41012 43864 41064
rect 44824 41055 44876 41064
rect 44824 41021 44833 41055
rect 44833 41021 44867 41055
rect 44867 41021 44876 41055
rect 44824 41012 44876 41021
rect 52460 41012 52512 41064
rect 52920 41055 52972 41064
rect 39948 40944 40000 40996
rect 40040 40944 40092 40996
rect 42892 40944 42944 40996
rect 45100 40944 45152 40996
rect 49424 40944 49476 40996
rect 52920 41021 52929 41055
rect 52929 41021 52963 41055
rect 52963 41021 52972 41055
rect 52920 41012 52972 41021
rect 53104 41055 53156 41064
rect 53104 41021 53113 41055
rect 53113 41021 53147 41055
rect 53147 41021 53156 41055
rect 53104 41012 53156 41021
rect 54484 41055 54536 41064
rect 54484 41021 54493 41055
rect 54493 41021 54527 41055
rect 54527 41021 54536 41055
rect 54484 41012 54536 41021
rect 55496 41055 55548 41064
rect 55496 41021 55505 41055
rect 55505 41021 55539 41055
rect 55539 41021 55548 41055
rect 55496 41012 55548 41021
rect 60832 41012 60884 41064
rect 61568 41012 61620 41064
rect 63040 41012 63092 41064
rect 64236 41012 64288 41064
rect 31576 40876 31628 40928
rect 36544 40876 36596 40928
rect 36636 40876 36688 40928
rect 37096 40876 37148 40928
rect 39028 40876 39080 40928
rect 39120 40876 39172 40928
rect 42800 40876 42852 40928
rect 42984 40876 43036 40928
rect 43812 40876 43864 40928
rect 53472 40944 53524 40996
rect 55128 40944 55180 40996
rect 53380 40876 53432 40928
rect 56600 40944 56652 40996
rect 57060 40944 57112 40996
rect 57152 40944 57204 40996
rect 55956 40919 56008 40928
rect 55956 40885 55965 40919
rect 55965 40885 55999 40919
rect 55999 40885 56008 40919
rect 55956 40876 56008 40885
rect 61568 40919 61620 40928
rect 61568 40885 61577 40919
rect 61577 40885 61611 40919
rect 61611 40885 61620 40919
rect 61568 40876 61620 40885
rect 61844 40919 61896 40928
rect 61844 40885 61853 40919
rect 61853 40885 61887 40919
rect 61887 40885 61896 40919
rect 61844 40876 61896 40885
rect 62580 40876 62632 40928
rect 63316 40876 63368 40928
rect 68100 41012 68152 41064
rect 69388 41080 69440 41132
rect 70400 41123 70452 41132
rect 70400 41089 70409 41123
rect 70409 41089 70443 41123
rect 70443 41089 70452 41123
rect 71688 41148 71740 41200
rect 71136 41123 71188 41132
rect 70400 41080 70452 41089
rect 71136 41089 71145 41123
rect 71145 41089 71179 41123
rect 71179 41089 71188 41123
rect 71136 41080 71188 41089
rect 70492 41012 70544 41064
rect 78128 41080 78180 41132
rect 64420 40944 64472 40996
rect 70308 40944 70360 40996
rect 71964 40987 72016 40996
rect 71964 40953 71973 40987
rect 71973 40953 72007 40987
rect 72007 40953 72016 40987
rect 71964 40944 72016 40953
rect 64328 40919 64380 40928
rect 64328 40885 64337 40919
rect 64337 40885 64371 40919
rect 64371 40885 64380 40919
rect 64328 40876 64380 40885
rect 66720 40876 66772 40928
rect 68376 40919 68428 40928
rect 68376 40885 68385 40919
rect 68385 40885 68419 40919
rect 68419 40885 68428 40919
rect 68376 40876 68428 40885
rect 69020 40876 69072 40928
rect 71596 40876 71648 40928
rect 74264 40876 74316 40928
rect 76840 40876 76892 40928
rect 77852 41012 77904 41064
rect 79784 41055 79836 41064
rect 79784 41021 79793 41055
rect 79793 41021 79827 41055
rect 79827 41021 79836 41055
rect 79784 41012 79836 41021
rect 77576 40876 77628 40928
rect 79876 40919 79928 40928
rect 79876 40885 79885 40919
rect 79885 40885 79919 40919
rect 79919 40885 79928 40919
rect 79876 40876 79928 40885
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 50326 40774 50378 40826
rect 50390 40774 50442 40826
rect 50454 40774 50506 40826
rect 50518 40774 50570 40826
rect 81046 40774 81098 40826
rect 81110 40774 81162 40826
rect 81174 40774 81226 40826
rect 81238 40774 81290 40826
rect 9956 40672 10008 40724
rect 10508 40672 10560 40724
rect 4712 40536 4764 40588
rect 12808 40672 12860 40724
rect 14004 40672 14056 40724
rect 28632 40672 28684 40724
rect 36176 40715 36228 40724
rect 36176 40681 36185 40715
rect 36185 40681 36219 40715
rect 36219 40681 36228 40715
rect 36176 40672 36228 40681
rect 36268 40672 36320 40724
rect 23664 40604 23716 40656
rect 16488 40536 16540 40588
rect 5540 40468 5592 40520
rect 11152 40511 11204 40520
rect 11152 40477 11161 40511
rect 11161 40477 11195 40511
rect 11195 40477 11204 40511
rect 11152 40468 11204 40477
rect 12900 40468 12952 40520
rect 16396 40468 16448 40520
rect 5724 40332 5776 40384
rect 12624 40332 12676 40384
rect 18236 40375 18288 40384
rect 18236 40341 18245 40375
rect 18245 40341 18279 40375
rect 18279 40341 18288 40375
rect 18236 40332 18288 40341
rect 18420 40375 18472 40384
rect 18420 40341 18429 40375
rect 18429 40341 18463 40375
rect 18463 40341 18472 40375
rect 18420 40332 18472 40341
rect 24584 40579 24636 40588
rect 24584 40545 24593 40579
rect 24593 40545 24627 40579
rect 24627 40545 24636 40579
rect 25688 40604 25740 40656
rect 27252 40604 27304 40656
rect 34612 40647 34664 40656
rect 24584 40536 24636 40545
rect 25228 40536 25280 40588
rect 27620 40536 27672 40588
rect 30012 40579 30064 40588
rect 28724 40468 28776 40520
rect 28816 40468 28868 40520
rect 29000 40468 29052 40520
rect 25688 40400 25740 40452
rect 23940 40332 23992 40384
rect 25044 40332 25096 40384
rect 26608 40332 26660 40384
rect 28264 40375 28316 40384
rect 28264 40341 28273 40375
rect 28273 40341 28307 40375
rect 28307 40341 28316 40375
rect 28264 40332 28316 40341
rect 28356 40332 28408 40384
rect 30012 40545 30021 40579
rect 30021 40545 30055 40579
rect 30055 40545 30064 40579
rect 30012 40536 30064 40545
rect 34612 40613 34621 40647
rect 34621 40613 34655 40647
rect 34655 40613 34664 40647
rect 34612 40604 34664 40613
rect 32956 40468 33008 40520
rect 35348 40536 35400 40588
rect 35624 40579 35676 40588
rect 35624 40545 35633 40579
rect 35633 40545 35667 40579
rect 35667 40545 35676 40579
rect 35624 40536 35676 40545
rect 35716 40579 35768 40588
rect 35716 40545 35725 40579
rect 35725 40545 35759 40579
rect 35759 40545 35768 40579
rect 35716 40536 35768 40545
rect 36544 40604 36596 40656
rect 37464 40604 37516 40656
rect 37924 40604 37976 40656
rect 38292 40647 38344 40656
rect 38292 40613 38301 40647
rect 38301 40613 38335 40647
rect 38335 40613 38344 40647
rect 38292 40604 38344 40613
rect 39120 40672 39172 40724
rect 40040 40604 40092 40656
rect 36636 40536 36688 40588
rect 42616 40604 42668 40656
rect 42892 40604 42944 40656
rect 43536 40604 43588 40656
rect 44456 40604 44508 40656
rect 45192 40604 45244 40656
rect 45376 40647 45428 40656
rect 45376 40613 45385 40647
rect 45385 40613 45419 40647
rect 45419 40613 45428 40647
rect 45376 40604 45428 40613
rect 46296 40672 46348 40724
rect 72516 40715 72568 40724
rect 55772 40604 55824 40656
rect 57060 40647 57112 40656
rect 57060 40613 57069 40647
rect 57069 40613 57103 40647
rect 57103 40613 57112 40647
rect 57060 40604 57112 40613
rect 60740 40647 60792 40656
rect 60740 40613 60749 40647
rect 60749 40613 60783 40647
rect 60783 40613 60792 40647
rect 60740 40604 60792 40613
rect 41236 40536 41288 40588
rect 38476 40468 38528 40520
rect 39396 40468 39448 40520
rect 40960 40468 41012 40520
rect 43352 40536 43404 40588
rect 45008 40579 45060 40588
rect 45008 40545 45017 40579
rect 45017 40545 45051 40579
rect 45051 40545 45060 40579
rect 45008 40536 45060 40545
rect 52276 40579 52328 40588
rect 52276 40545 52285 40579
rect 52285 40545 52319 40579
rect 52319 40545 52328 40579
rect 52276 40536 52328 40545
rect 53104 40536 53156 40588
rect 52920 40468 52972 40520
rect 54760 40536 54812 40588
rect 55128 40536 55180 40588
rect 55864 40579 55916 40588
rect 55864 40545 55873 40579
rect 55873 40545 55907 40579
rect 55907 40545 55916 40579
rect 55864 40536 55916 40545
rect 62304 40579 62356 40588
rect 62304 40545 62313 40579
rect 62313 40545 62347 40579
rect 62347 40545 62356 40579
rect 62304 40536 62356 40545
rect 62948 40604 63000 40656
rect 63868 40647 63920 40656
rect 63868 40613 63877 40647
rect 63877 40613 63911 40647
rect 63911 40613 63920 40647
rect 63868 40604 63920 40613
rect 64604 40647 64656 40656
rect 64604 40613 64613 40647
rect 64613 40613 64647 40647
rect 64647 40613 64656 40647
rect 64604 40604 64656 40613
rect 64696 40604 64748 40656
rect 70124 40604 70176 40656
rect 57244 40468 57296 40520
rect 62580 40536 62632 40588
rect 62764 40468 62816 40520
rect 63776 40536 63828 40588
rect 64420 40579 64472 40588
rect 64420 40545 64429 40579
rect 64429 40545 64463 40579
rect 64463 40545 64472 40579
rect 64420 40536 64472 40545
rect 66720 40579 66772 40588
rect 66720 40545 66729 40579
rect 66729 40545 66763 40579
rect 66763 40545 66772 40579
rect 66720 40536 66772 40545
rect 68468 40579 68520 40588
rect 68468 40545 68477 40579
rect 68477 40545 68511 40579
rect 68511 40545 68520 40579
rect 68468 40536 68520 40545
rect 69388 40536 69440 40588
rect 69848 40536 69900 40588
rect 70400 40468 70452 40520
rect 72516 40681 72525 40715
rect 72525 40681 72559 40715
rect 72559 40681 72568 40715
rect 72516 40672 72568 40681
rect 77944 40672 77996 40724
rect 78220 40604 78272 40656
rect 75828 40536 75880 40588
rect 77576 40579 77628 40588
rect 77576 40545 77585 40579
rect 77585 40545 77619 40579
rect 77619 40545 77628 40579
rect 77576 40536 77628 40545
rect 77668 40536 77720 40588
rect 77852 40579 77904 40588
rect 77852 40545 77861 40579
rect 77861 40545 77895 40579
rect 77895 40545 77904 40579
rect 77852 40536 77904 40545
rect 78128 40579 78180 40588
rect 78128 40545 78137 40579
rect 78137 40545 78171 40579
rect 78171 40545 78180 40579
rect 78128 40536 78180 40545
rect 74448 40468 74500 40520
rect 80796 40468 80848 40520
rect 83648 40511 83700 40520
rect 83648 40477 83657 40511
rect 83657 40477 83691 40511
rect 83691 40477 83700 40511
rect 83648 40468 83700 40477
rect 62672 40400 62724 40452
rect 66812 40400 66864 40452
rect 34796 40375 34848 40384
rect 34796 40341 34805 40375
rect 34805 40341 34839 40375
rect 34839 40341 34848 40375
rect 34796 40332 34848 40341
rect 35716 40332 35768 40384
rect 36820 40332 36872 40384
rect 37648 40332 37700 40384
rect 38568 40375 38620 40384
rect 38568 40341 38577 40375
rect 38577 40341 38611 40375
rect 38611 40341 38620 40375
rect 38568 40332 38620 40341
rect 38660 40332 38712 40384
rect 42708 40332 42760 40384
rect 42800 40332 42852 40384
rect 43628 40332 43680 40384
rect 53288 40375 53340 40384
rect 53288 40341 53297 40375
rect 53297 40341 53331 40375
rect 53331 40341 53340 40375
rect 53288 40332 53340 40341
rect 56876 40375 56928 40384
rect 56876 40341 56885 40375
rect 56885 40341 56919 40375
rect 56919 40341 56928 40375
rect 56876 40332 56928 40341
rect 57336 40375 57388 40384
rect 57336 40341 57345 40375
rect 57345 40341 57379 40375
rect 57379 40341 57388 40375
rect 57336 40332 57388 40341
rect 57796 40375 57848 40384
rect 57796 40341 57805 40375
rect 57805 40341 57839 40375
rect 57839 40341 57848 40375
rect 57796 40332 57848 40341
rect 62948 40332 63000 40384
rect 68652 40375 68704 40384
rect 68652 40341 68661 40375
rect 68661 40341 68695 40375
rect 68695 40341 68704 40375
rect 68652 40332 68704 40341
rect 69388 40375 69440 40384
rect 69388 40341 69397 40375
rect 69397 40341 69431 40375
rect 69431 40341 69440 40375
rect 69388 40332 69440 40341
rect 69848 40375 69900 40384
rect 69848 40341 69857 40375
rect 69857 40341 69891 40375
rect 69891 40341 69900 40375
rect 69848 40332 69900 40341
rect 70032 40332 70084 40384
rect 71964 40332 72016 40384
rect 73988 40375 74040 40384
rect 73988 40341 73997 40375
rect 73997 40341 74031 40375
rect 74031 40341 74040 40375
rect 73988 40332 74040 40341
rect 75828 40332 75880 40384
rect 78036 40332 78088 40384
rect 80244 40375 80296 40384
rect 80244 40341 80253 40375
rect 80253 40341 80287 40375
rect 80287 40341 80296 40375
rect 80244 40332 80296 40341
rect 84752 40375 84804 40384
rect 84752 40341 84761 40375
rect 84761 40341 84795 40375
rect 84795 40341 84804 40375
rect 84752 40332 84804 40341
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 65686 40230 65738 40282
rect 65750 40230 65802 40282
rect 65814 40230 65866 40282
rect 65878 40230 65930 40282
rect 96406 40230 96458 40282
rect 96470 40230 96522 40282
rect 96534 40230 96586 40282
rect 96598 40230 96650 40282
rect 5448 40128 5500 40180
rect 6920 40171 6972 40180
rect 6920 40137 6929 40171
rect 6929 40137 6963 40171
rect 6963 40137 6972 40171
rect 6920 40128 6972 40137
rect 11152 40171 11204 40180
rect 11152 40137 11161 40171
rect 11161 40137 11195 40171
rect 11195 40137 11204 40171
rect 11152 40128 11204 40137
rect 12900 40128 12952 40180
rect 31576 40128 31628 40180
rect 4712 40103 4764 40112
rect 4712 40069 4721 40103
rect 4721 40069 4755 40103
rect 4755 40069 4764 40103
rect 4712 40060 4764 40069
rect 4620 39992 4672 40044
rect 9772 39992 9824 40044
rect 5724 39967 5776 39976
rect 5724 39933 5733 39967
rect 5733 39933 5767 39967
rect 5767 39933 5776 39967
rect 5724 39924 5776 39933
rect 7104 39967 7156 39976
rect 7104 39933 7105 39967
rect 7105 39933 7139 39967
rect 7139 39933 7156 39967
rect 7104 39924 7156 39933
rect 7288 39924 7340 39976
rect 10692 40060 10744 40112
rect 14188 40060 14240 40112
rect 16856 40060 16908 40112
rect 17684 40035 17736 40044
rect 17684 40001 17693 40035
rect 17693 40001 17727 40035
rect 17727 40001 17736 40035
rect 17684 39992 17736 40001
rect 10692 39967 10744 39976
rect 10692 39933 10701 39967
rect 10701 39933 10735 39967
rect 10735 39933 10744 39967
rect 10692 39924 10744 39933
rect 10876 39967 10928 39976
rect 10876 39933 10885 39967
rect 10885 39933 10919 39967
rect 10919 39933 10928 39967
rect 10876 39924 10928 39933
rect 12992 39924 13044 39976
rect 13360 39924 13412 39976
rect 4068 39856 4120 39908
rect 19984 40060 20036 40112
rect 23388 40060 23440 40112
rect 23572 39992 23624 40044
rect 25504 40060 25556 40112
rect 25688 40060 25740 40112
rect 26516 40060 26568 40112
rect 27528 40060 27580 40112
rect 19340 39924 19392 39976
rect 23480 39924 23532 39976
rect 24860 39992 24912 40044
rect 5816 39831 5868 39840
rect 5816 39797 5825 39831
rect 5825 39797 5859 39831
rect 5859 39797 5868 39831
rect 5816 39788 5868 39797
rect 7840 39788 7892 39840
rect 9772 39831 9824 39840
rect 9772 39797 9781 39831
rect 9781 39797 9815 39831
rect 9815 39797 9824 39831
rect 9772 39788 9824 39797
rect 11704 39788 11756 39840
rect 13268 39831 13320 39840
rect 13268 39797 13277 39831
rect 13277 39797 13311 39831
rect 13311 39797 13320 39831
rect 13268 39788 13320 39797
rect 13360 39788 13412 39840
rect 14648 39788 14700 39840
rect 19984 39856 20036 39908
rect 23572 39856 23624 39908
rect 24584 39924 24636 39976
rect 26516 39967 26568 39976
rect 20444 39788 20496 39840
rect 23296 39788 23348 39840
rect 24860 39856 24912 39908
rect 26516 39933 26525 39967
rect 26525 39933 26559 39967
rect 26559 39933 26568 39967
rect 26516 39924 26568 39933
rect 26608 39967 26660 39976
rect 26608 39933 26617 39967
rect 26617 39933 26651 39967
rect 26651 39933 26660 39967
rect 28356 40060 28408 40112
rect 28632 40060 28684 40112
rect 35900 40128 35952 40180
rect 32220 39992 32272 40044
rect 32680 39992 32732 40044
rect 32956 40035 33008 40044
rect 32956 40001 32965 40035
rect 32965 40001 32999 40035
rect 32999 40001 33008 40035
rect 32956 39992 33008 40001
rect 30564 39967 30616 39976
rect 26608 39924 26660 39933
rect 30564 39933 30573 39967
rect 30573 39933 30607 39967
rect 30607 39933 30616 39967
rect 30564 39924 30616 39933
rect 30748 39924 30800 39976
rect 30932 39924 30984 39976
rect 31116 39967 31168 39976
rect 31116 39933 31125 39967
rect 31125 39933 31159 39967
rect 31159 39933 31168 39967
rect 32588 39967 32640 39976
rect 31116 39924 31168 39933
rect 32128 39856 32180 39908
rect 32588 39933 32597 39967
rect 32597 39933 32631 39967
rect 32631 39933 32640 39967
rect 32588 39924 32640 39933
rect 33416 39924 33468 39976
rect 34796 40060 34848 40112
rect 35624 40060 35676 40112
rect 34060 39992 34112 40044
rect 35348 39992 35400 40044
rect 35716 39924 35768 39976
rect 38660 40128 38712 40180
rect 54852 40128 54904 40180
rect 55772 40128 55824 40180
rect 61568 40171 61620 40180
rect 61568 40137 61577 40171
rect 61577 40137 61611 40171
rect 61611 40137 61620 40171
rect 61568 40128 61620 40137
rect 62672 40128 62724 40180
rect 69112 40128 69164 40180
rect 70124 40128 70176 40180
rect 70308 40128 70360 40180
rect 70492 40128 70544 40180
rect 36820 40060 36872 40112
rect 37924 40103 37976 40112
rect 37924 40069 37933 40103
rect 37933 40069 37967 40103
rect 37967 40069 37976 40103
rect 37924 40060 37976 40069
rect 36912 39924 36964 39976
rect 38200 39967 38252 39976
rect 38200 39933 38209 39967
rect 38209 39933 38243 39967
rect 38243 39933 38252 39967
rect 38200 39924 38252 39933
rect 38384 39967 38436 39976
rect 38384 39933 38393 39967
rect 38393 39933 38427 39967
rect 38427 39933 38436 39967
rect 38384 39924 38436 39933
rect 38936 39967 38988 39976
rect 38936 39933 38945 39967
rect 38945 39933 38979 39967
rect 38979 39933 38988 39967
rect 38936 39924 38988 39933
rect 40040 39924 40092 39976
rect 41512 39967 41564 39976
rect 41512 39933 41521 39967
rect 41521 39933 41555 39967
rect 41555 39933 41564 39967
rect 41512 39924 41564 39933
rect 42248 40060 42300 40112
rect 44640 40060 44692 40112
rect 42708 40035 42760 40044
rect 42708 40001 42717 40035
rect 42717 40001 42751 40035
rect 42751 40001 42760 40035
rect 42708 39992 42760 40001
rect 56876 40060 56928 40112
rect 57796 40060 57848 40112
rect 66168 40060 66220 40112
rect 74264 40060 74316 40112
rect 26148 39788 26200 39840
rect 26516 39788 26568 39840
rect 31116 39788 31168 39840
rect 31760 39788 31812 39840
rect 38108 39856 38160 39908
rect 35532 39788 35584 39840
rect 35808 39788 35860 39840
rect 38200 39788 38252 39840
rect 38384 39788 38436 39840
rect 41052 39788 41104 39840
rect 41512 39788 41564 39840
rect 42248 39967 42300 39976
rect 42248 39933 42257 39967
rect 42257 39933 42291 39967
rect 42291 39933 42300 39967
rect 42248 39924 42300 39933
rect 43536 39924 43588 39976
rect 43996 39924 44048 39976
rect 48872 39992 48924 40044
rect 47676 39967 47728 39976
rect 47676 39933 47685 39967
rect 47685 39933 47719 39967
rect 47719 39933 47728 39967
rect 47676 39924 47728 39933
rect 43720 39899 43772 39908
rect 42248 39788 42300 39840
rect 43076 39831 43128 39840
rect 43076 39797 43085 39831
rect 43085 39797 43119 39831
rect 43119 39797 43128 39831
rect 43076 39788 43128 39797
rect 43720 39865 43729 39899
rect 43729 39865 43763 39899
rect 43763 39865 43772 39899
rect 43720 39856 43772 39865
rect 48136 39967 48188 39976
rect 48136 39933 48145 39967
rect 48145 39933 48179 39967
rect 48179 39933 48188 39967
rect 49148 39967 49200 39976
rect 48136 39924 48188 39933
rect 49148 39933 49157 39967
rect 49157 39933 49191 39967
rect 49191 39933 49200 39967
rect 49148 39924 49200 39933
rect 52460 39924 52512 39976
rect 52552 39967 52604 39976
rect 52552 39933 52561 39967
rect 52561 39933 52595 39967
rect 52595 39933 52604 39967
rect 53748 39967 53800 39976
rect 52552 39924 52604 39933
rect 53748 39933 53757 39967
rect 53757 39933 53791 39967
rect 53791 39933 53800 39967
rect 53748 39924 53800 39933
rect 54024 39967 54076 39976
rect 54024 39933 54033 39967
rect 54033 39933 54067 39967
rect 54067 39933 54076 39967
rect 54024 39924 54076 39933
rect 54116 39924 54168 39976
rect 55496 39967 55548 39976
rect 55496 39933 55505 39967
rect 55505 39933 55539 39967
rect 55539 39933 55548 39967
rect 55496 39924 55548 39933
rect 44272 39788 44324 39840
rect 44548 39788 44600 39840
rect 52184 39856 52236 39908
rect 48596 39831 48648 39840
rect 48596 39797 48605 39831
rect 48605 39797 48639 39831
rect 48639 39797 48648 39831
rect 48596 39788 48648 39797
rect 48688 39788 48740 39840
rect 52276 39788 52328 39840
rect 52552 39788 52604 39840
rect 56048 39992 56100 40044
rect 61936 40035 61988 40044
rect 61936 40001 61945 40035
rect 61945 40001 61979 40035
rect 61979 40001 61988 40035
rect 61936 39992 61988 40001
rect 64420 39992 64472 40044
rect 60740 39924 60792 39976
rect 66812 39992 66864 40044
rect 67272 40035 67324 40044
rect 67272 40001 67281 40035
rect 67281 40001 67315 40035
rect 67315 40001 67324 40035
rect 67272 39992 67324 40001
rect 67732 39992 67784 40044
rect 68376 39992 68428 40044
rect 69388 39992 69440 40044
rect 69940 40035 69992 40044
rect 69940 40001 69949 40035
rect 69949 40001 69983 40035
rect 69983 40001 69992 40035
rect 69940 39992 69992 40001
rect 70308 39992 70360 40044
rect 68468 39924 68520 39976
rect 70032 39967 70084 39976
rect 70032 39933 70041 39967
rect 70041 39933 70075 39967
rect 70075 39933 70084 39967
rect 70032 39924 70084 39933
rect 70400 39967 70452 39976
rect 70400 39933 70409 39967
rect 70409 39933 70443 39967
rect 70443 39933 70452 39967
rect 71412 39967 71464 39976
rect 70400 39924 70452 39933
rect 71412 39933 71421 39967
rect 71421 39933 71455 39967
rect 71455 39933 71464 39967
rect 71412 39924 71464 39933
rect 71872 39924 71924 39976
rect 68560 39856 68612 39908
rect 69388 39899 69440 39908
rect 69388 39865 69397 39899
rect 69397 39865 69431 39899
rect 69431 39865 69440 39899
rect 69388 39856 69440 39865
rect 64788 39788 64840 39840
rect 67180 39788 67232 39840
rect 69664 39788 69716 39840
rect 70952 39831 71004 39840
rect 70952 39797 70961 39831
rect 70961 39797 70995 39831
rect 70995 39797 71004 39831
rect 70952 39788 71004 39797
rect 71688 39788 71740 39840
rect 74540 39992 74592 40044
rect 77668 39992 77720 40044
rect 75184 39924 75236 39976
rect 75828 39967 75880 39976
rect 75828 39933 75837 39967
rect 75837 39933 75871 39967
rect 75871 39933 75880 39967
rect 75828 39924 75880 39933
rect 76196 39856 76248 39908
rect 78128 40128 78180 40180
rect 83648 40128 83700 40180
rect 78036 40060 78088 40112
rect 84752 40060 84804 40112
rect 79876 39924 79928 39976
rect 80244 39924 80296 39976
rect 83740 39924 83792 39976
rect 85212 39924 85264 39976
rect 77392 39899 77444 39908
rect 75828 39788 75880 39840
rect 76656 39831 76708 39840
rect 76656 39797 76665 39831
rect 76665 39797 76699 39831
rect 76699 39797 76708 39831
rect 76656 39788 76708 39797
rect 77392 39865 77401 39899
rect 77401 39865 77435 39899
rect 77435 39865 77444 39899
rect 77392 39856 77444 39865
rect 85396 39899 85448 39908
rect 85396 39865 85405 39899
rect 85405 39865 85439 39899
rect 85439 39865 85448 39899
rect 85396 39856 85448 39865
rect 85948 39899 86000 39908
rect 85948 39865 85957 39899
rect 85957 39865 85991 39899
rect 85991 39865 86000 39899
rect 85948 39856 86000 39865
rect 77024 39788 77076 39840
rect 79600 39788 79652 39840
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 50326 39686 50378 39738
rect 50390 39686 50442 39738
rect 50454 39686 50506 39738
rect 50518 39686 50570 39738
rect 81046 39686 81098 39738
rect 81110 39686 81162 39738
rect 81174 39686 81226 39738
rect 81238 39686 81290 39738
rect 5540 39584 5592 39636
rect 8024 39584 8076 39636
rect 5816 39448 5868 39500
rect 11704 39516 11756 39568
rect 12716 39516 12768 39568
rect 12992 39559 13044 39568
rect 12992 39525 13001 39559
rect 13001 39525 13035 39559
rect 13035 39525 13044 39559
rect 12992 39516 13044 39525
rect 17408 39516 17460 39568
rect 26516 39559 26568 39568
rect 3608 39244 3660 39296
rect 12624 39448 12676 39500
rect 12900 39491 12952 39500
rect 12900 39457 12909 39491
rect 12909 39457 12943 39491
rect 12943 39457 12952 39491
rect 12900 39448 12952 39457
rect 16396 39491 16448 39500
rect 16396 39457 16405 39491
rect 16405 39457 16439 39491
rect 16439 39457 16448 39491
rect 16396 39448 16448 39457
rect 9772 39380 9824 39432
rect 15752 39380 15804 39432
rect 16672 39423 16724 39432
rect 16672 39389 16681 39423
rect 16681 39389 16715 39423
rect 16715 39389 16724 39423
rect 16672 39380 16724 39389
rect 18236 39448 18288 39500
rect 23296 39448 23348 39500
rect 23572 39491 23624 39500
rect 23572 39457 23581 39491
rect 23581 39457 23615 39491
rect 23615 39457 23624 39491
rect 23572 39448 23624 39457
rect 23940 39491 23992 39500
rect 23940 39457 23949 39491
rect 23949 39457 23983 39491
rect 23983 39457 23992 39491
rect 23940 39448 23992 39457
rect 19340 39380 19392 39432
rect 22928 39380 22980 39432
rect 24860 39491 24912 39500
rect 24860 39457 24869 39491
rect 24869 39457 24903 39491
rect 24903 39457 24912 39491
rect 25044 39491 25096 39500
rect 24860 39448 24912 39457
rect 25044 39457 25053 39491
rect 25053 39457 25087 39491
rect 25087 39457 25096 39491
rect 25044 39448 25096 39457
rect 26516 39525 26525 39559
rect 26525 39525 26559 39559
rect 26559 39525 26568 39559
rect 26516 39516 26568 39525
rect 29828 39584 29880 39636
rect 30564 39584 30616 39636
rect 31024 39516 31076 39568
rect 31392 39584 31444 39636
rect 26976 39448 27028 39500
rect 29828 39491 29880 39500
rect 29828 39457 29837 39491
rect 29837 39457 29871 39491
rect 29871 39457 29880 39491
rect 29828 39448 29880 39457
rect 29920 39448 29972 39500
rect 31116 39448 31168 39500
rect 32220 39448 32272 39500
rect 36176 39584 36228 39636
rect 36820 39627 36872 39636
rect 36820 39593 36829 39627
rect 36829 39593 36863 39627
rect 36863 39593 36872 39627
rect 36820 39584 36872 39593
rect 38476 39584 38528 39636
rect 35532 39516 35584 39568
rect 35348 39491 35400 39500
rect 35348 39457 35357 39491
rect 35357 39457 35391 39491
rect 35391 39457 35400 39491
rect 35348 39448 35400 39457
rect 35808 39491 35860 39500
rect 26884 39423 26936 39432
rect 26884 39389 26893 39423
rect 26893 39389 26927 39423
rect 26927 39389 26936 39423
rect 26884 39380 26936 39389
rect 27252 39423 27304 39432
rect 27252 39389 27261 39423
rect 27261 39389 27295 39423
rect 27295 39389 27304 39423
rect 27252 39380 27304 39389
rect 29736 39423 29788 39432
rect 29736 39389 29745 39423
rect 29745 39389 29779 39423
rect 29779 39389 29788 39423
rect 29736 39380 29788 39389
rect 31760 39380 31812 39432
rect 34152 39380 34204 39432
rect 35808 39457 35817 39491
rect 35817 39457 35851 39491
rect 35851 39457 35860 39491
rect 35808 39448 35860 39457
rect 36084 39448 36136 39500
rect 38568 39516 38620 39568
rect 43720 39516 43772 39568
rect 43812 39516 43864 39568
rect 44640 39559 44692 39568
rect 40868 39448 40920 39500
rect 41696 39491 41748 39500
rect 36636 39423 36688 39432
rect 8760 39312 8812 39364
rect 10600 39312 10652 39364
rect 10876 39312 10928 39364
rect 34612 39312 34664 39364
rect 18052 39244 18104 39296
rect 18420 39244 18472 39296
rect 18972 39244 19024 39296
rect 23756 39244 23808 39296
rect 23940 39244 23992 39296
rect 25780 39244 25832 39296
rect 26332 39244 26384 39296
rect 26792 39287 26844 39296
rect 26792 39253 26801 39287
rect 26801 39253 26835 39287
rect 26835 39253 26844 39287
rect 26792 39244 26844 39253
rect 30840 39287 30892 39296
rect 30840 39253 30849 39287
rect 30849 39253 30883 39287
rect 30883 39253 30892 39287
rect 30840 39244 30892 39253
rect 34704 39244 34756 39296
rect 36636 39389 36645 39423
rect 36645 39389 36679 39423
rect 36679 39389 36688 39423
rect 36636 39380 36688 39389
rect 37740 39380 37792 39432
rect 40960 39380 41012 39432
rect 35072 39312 35124 39364
rect 41696 39457 41705 39491
rect 41705 39457 41739 39491
rect 41739 39457 41748 39491
rect 41696 39448 41748 39457
rect 42432 39448 42484 39500
rect 42248 39380 42300 39432
rect 43260 39380 43312 39432
rect 43536 39491 43588 39500
rect 43536 39457 43545 39491
rect 43545 39457 43579 39491
rect 43579 39457 43588 39491
rect 44088 39491 44140 39500
rect 43536 39448 43588 39457
rect 44088 39457 44097 39491
rect 44097 39457 44131 39491
rect 44131 39457 44140 39491
rect 44088 39448 44140 39457
rect 44180 39448 44232 39500
rect 44640 39525 44649 39559
rect 44649 39525 44683 39559
rect 44683 39525 44692 39559
rect 44640 39516 44692 39525
rect 48688 39516 48740 39568
rect 49976 39516 50028 39568
rect 52000 39516 52052 39568
rect 44824 39448 44876 39500
rect 48780 39448 48832 39500
rect 48964 39491 49016 39500
rect 48964 39457 48973 39491
rect 48973 39457 49007 39491
rect 49007 39457 49016 39491
rect 48964 39448 49016 39457
rect 50988 39448 51040 39500
rect 51724 39448 51776 39500
rect 52552 39448 52604 39500
rect 52828 39448 52880 39500
rect 53196 39516 53248 39568
rect 54024 39516 54076 39568
rect 55404 39516 55456 39568
rect 56048 39516 56100 39568
rect 61660 39559 61712 39568
rect 61660 39525 61669 39559
rect 61669 39525 61703 39559
rect 61703 39525 61712 39559
rect 61660 39516 61712 39525
rect 66536 39516 66588 39568
rect 69664 39584 69716 39636
rect 53472 39448 53524 39500
rect 54760 39491 54812 39500
rect 54760 39457 54769 39491
rect 54769 39457 54803 39491
rect 54803 39457 54812 39491
rect 54760 39448 54812 39457
rect 54852 39491 54904 39500
rect 54852 39457 54861 39491
rect 54861 39457 54895 39491
rect 54895 39457 54904 39491
rect 54852 39448 54904 39457
rect 43720 39380 43772 39432
rect 44640 39380 44692 39432
rect 48688 39380 48740 39432
rect 49240 39423 49292 39432
rect 49240 39389 49249 39423
rect 49249 39389 49283 39423
rect 49283 39389 49292 39423
rect 49240 39380 49292 39389
rect 49332 39380 49384 39432
rect 35348 39244 35400 39296
rect 36636 39244 36688 39296
rect 36912 39244 36964 39296
rect 40960 39244 41012 39296
rect 41604 39312 41656 39364
rect 43168 39312 43220 39364
rect 43996 39312 44048 39364
rect 44088 39312 44140 39364
rect 44824 39312 44876 39364
rect 41880 39244 41932 39296
rect 42524 39287 42576 39296
rect 42524 39253 42533 39287
rect 42533 39253 42567 39287
rect 42567 39253 42576 39287
rect 42892 39287 42944 39296
rect 42524 39244 42576 39253
rect 42892 39253 42901 39287
rect 42901 39253 42935 39287
rect 42935 39253 42944 39287
rect 42892 39244 42944 39253
rect 43076 39287 43128 39296
rect 43076 39253 43085 39287
rect 43085 39253 43119 39287
rect 43119 39253 43128 39287
rect 43076 39244 43128 39253
rect 44456 39244 44508 39296
rect 55864 39312 55916 39364
rect 50160 39244 50212 39296
rect 54576 39287 54628 39296
rect 54576 39253 54585 39287
rect 54585 39253 54619 39287
rect 54619 39253 54628 39287
rect 54576 39244 54628 39253
rect 55404 39244 55456 39296
rect 55496 39244 55548 39296
rect 57336 39448 57388 39500
rect 61844 39491 61896 39500
rect 61844 39457 61853 39491
rect 61853 39457 61887 39491
rect 61887 39457 61896 39491
rect 61844 39448 61896 39457
rect 62212 39491 62264 39500
rect 62212 39457 62221 39491
rect 62221 39457 62255 39491
rect 62255 39457 62264 39491
rect 62212 39448 62264 39457
rect 63040 39491 63092 39500
rect 63040 39457 63049 39491
rect 63049 39457 63083 39491
rect 63083 39457 63092 39491
rect 63040 39448 63092 39457
rect 63500 39448 63552 39500
rect 64604 39448 64656 39500
rect 66720 39491 66772 39500
rect 66720 39457 66729 39491
rect 66729 39457 66763 39491
rect 66763 39457 66772 39491
rect 66720 39448 66772 39457
rect 67640 39491 67692 39500
rect 67640 39457 67649 39491
rect 67649 39457 67683 39491
rect 67683 39457 67692 39491
rect 67640 39448 67692 39457
rect 65524 39380 65576 39432
rect 63224 39312 63276 39364
rect 66536 39355 66588 39364
rect 66536 39321 66545 39355
rect 66545 39321 66579 39355
rect 66579 39321 66588 39355
rect 66536 39312 66588 39321
rect 69020 39448 69072 39500
rect 69388 39448 69440 39500
rect 56048 39244 56100 39296
rect 61660 39244 61712 39296
rect 62764 39244 62816 39296
rect 63500 39244 63552 39296
rect 64696 39244 64748 39296
rect 67732 39287 67784 39296
rect 67732 39253 67741 39287
rect 67741 39253 67775 39287
rect 67775 39253 67784 39287
rect 67732 39244 67784 39253
rect 69940 39312 69992 39364
rect 70952 39312 71004 39364
rect 75828 39491 75880 39500
rect 75828 39457 75837 39491
rect 75837 39457 75871 39491
rect 75871 39457 75880 39491
rect 75828 39448 75880 39457
rect 76196 39584 76248 39636
rect 80796 39627 80848 39636
rect 80796 39593 80805 39627
rect 80805 39593 80839 39627
rect 80839 39593 80848 39627
rect 80796 39584 80848 39593
rect 76472 39516 76524 39568
rect 83464 39516 83516 39568
rect 83740 39559 83792 39568
rect 83740 39525 83749 39559
rect 83749 39525 83783 39559
rect 83783 39525 83792 39559
rect 83740 39516 83792 39525
rect 85396 39584 85448 39636
rect 78036 39491 78088 39500
rect 78036 39457 78045 39491
rect 78045 39457 78079 39491
rect 78079 39457 78088 39491
rect 78036 39448 78088 39457
rect 79140 39491 79192 39500
rect 79140 39457 79149 39491
rect 79149 39457 79183 39491
rect 79183 39457 79192 39491
rect 79140 39448 79192 39457
rect 79416 39491 79468 39500
rect 79416 39457 79425 39491
rect 79425 39457 79459 39491
rect 79459 39457 79468 39491
rect 79416 39448 79468 39457
rect 80704 39491 80756 39500
rect 80704 39457 80713 39491
rect 80713 39457 80747 39491
rect 80747 39457 80756 39491
rect 80704 39448 80756 39457
rect 84384 39491 84436 39500
rect 84384 39457 84393 39491
rect 84393 39457 84427 39491
rect 84427 39457 84436 39491
rect 84384 39448 84436 39457
rect 76472 39312 76524 39364
rect 76380 39244 76432 39296
rect 77300 39244 77352 39296
rect 82912 39244 82964 39296
rect 84016 39312 84068 39364
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 65686 39142 65738 39194
rect 65750 39142 65802 39194
rect 65814 39142 65866 39194
rect 65878 39142 65930 39194
rect 96406 39142 96458 39194
rect 96470 39142 96522 39194
rect 96534 39142 96586 39194
rect 96598 39142 96650 39194
rect 3792 39040 3844 39092
rect 9772 39040 9824 39092
rect 11520 39040 11572 39092
rect 4068 38972 4120 39024
rect 15016 38972 15068 39024
rect 16672 39040 16724 39092
rect 2596 38836 2648 38888
rect 5264 38879 5316 38888
rect 5264 38845 5273 38879
rect 5273 38845 5307 38879
rect 5307 38845 5316 38879
rect 5264 38836 5316 38845
rect 14648 38904 14700 38956
rect 10968 38879 11020 38888
rect 4160 38700 4212 38752
rect 4436 38743 4488 38752
rect 4436 38709 4445 38743
rect 4445 38709 4479 38743
rect 4479 38709 4488 38743
rect 4436 38700 4488 38709
rect 9772 38768 9824 38820
rect 10968 38845 10977 38879
rect 10977 38845 11011 38879
rect 11011 38845 11020 38879
rect 10968 38836 11020 38845
rect 11244 38836 11296 38888
rect 11520 38879 11572 38888
rect 11520 38845 11529 38879
rect 11529 38845 11563 38879
rect 11563 38845 11572 38879
rect 11520 38836 11572 38845
rect 13268 38836 13320 38888
rect 14832 38836 14884 38888
rect 15016 38879 15068 38888
rect 15016 38845 15025 38879
rect 15025 38845 15059 38879
rect 15059 38845 15068 38879
rect 15016 38836 15068 38845
rect 14004 38768 14056 38820
rect 20444 38972 20496 39024
rect 23848 38972 23900 39024
rect 25964 38972 26016 39024
rect 19340 38904 19392 38956
rect 16672 38836 16724 38888
rect 16948 38879 17000 38888
rect 16948 38845 16957 38879
rect 16957 38845 16991 38879
rect 16991 38845 17000 38879
rect 16948 38836 17000 38845
rect 18052 38879 18104 38888
rect 18052 38845 18061 38879
rect 18061 38845 18095 38879
rect 18095 38845 18104 38879
rect 18052 38836 18104 38845
rect 18972 38836 19024 38888
rect 21180 38904 21232 38956
rect 26240 38947 26292 38956
rect 26240 38913 26249 38947
rect 26249 38913 26283 38947
rect 26283 38913 26292 38947
rect 27436 39040 27488 39092
rect 29736 39083 29788 39092
rect 29736 39049 29745 39083
rect 29745 39049 29779 39083
rect 29779 39049 29788 39083
rect 29736 39040 29788 39049
rect 29828 39040 29880 39092
rect 31392 39040 31444 39092
rect 34612 39040 34664 39092
rect 26976 38972 27028 39024
rect 34704 38972 34756 39024
rect 26240 38904 26292 38913
rect 34796 38904 34848 38956
rect 23848 38879 23900 38888
rect 23848 38845 23857 38879
rect 23857 38845 23891 38879
rect 23891 38845 23900 38879
rect 23848 38836 23900 38845
rect 24400 38879 24452 38888
rect 24400 38845 24409 38879
rect 24409 38845 24443 38879
rect 24443 38845 24452 38879
rect 24400 38836 24452 38845
rect 23572 38768 23624 38820
rect 24768 38836 24820 38888
rect 25228 38879 25280 38888
rect 25228 38845 25237 38879
rect 25237 38845 25271 38879
rect 25271 38845 25280 38879
rect 25228 38836 25280 38845
rect 25780 38836 25832 38888
rect 26148 38836 26200 38888
rect 26792 38836 26844 38888
rect 29460 38836 29512 38888
rect 29644 38879 29696 38888
rect 29644 38845 29653 38879
rect 29653 38845 29687 38879
rect 29687 38845 29696 38879
rect 37648 38972 37700 39024
rect 37740 38947 37792 38956
rect 37740 38913 37749 38947
rect 37749 38913 37783 38947
rect 37783 38913 37792 38947
rect 37740 38904 37792 38913
rect 37924 39040 37976 39092
rect 39488 39040 39540 39092
rect 49332 39040 49384 39092
rect 53380 39040 53432 39092
rect 62120 39040 62172 39092
rect 41144 38904 41196 38956
rect 29644 38836 29696 38845
rect 37096 38879 37148 38888
rect 37096 38845 37105 38879
rect 37105 38845 37139 38879
rect 37139 38845 37148 38879
rect 37096 38836 37148 38845
rect 38476 38836 38528 38888
rect 41604 38836 41656 38888
rect 41880 38972 41932 39024
rect 43536 39015 43588 39024
rect 43536 38981 43545 39015
rect 43545 38981 43579 39015
rect 43579 38981 43588 39015
rect 43536 38972 43588 38981
rect 43628 38972 43680 39024
rect 43996 39015 44048 39024
rect 43996 38981 44005 39015
rect 44005 38981 44039 39015
rect 44039 38981 44048 39015
rect 43996 38972 44048 38981
rect 44548 38972 44600 39024
rect 48872 39015 48924 39024
rect 42708 38947 42760 38956
rect 42708 38913 42717 38947
rect 42717 38913 42751 38947
rect 42751 38913 42760 38947
rect 42708 38904 42760 38913
rect 42248 38879 42300 38888
rect 42248 38845 42257 38879
rect 42257 38845 42291 38879
rect 42291 38845 42300 38879
rect 43168 38904 43220 38956
rect 44272 38904 44324 38956
rect 47400 38947 47452 38956
rect 47400 38913 47409 38947
rect 47409 38913 47443 38947
rect 47443 38913 47452 38947
rect 47400 38904 47452 38913
rect 42248 38836 42300 38845
rect 43536 38836 43588 38888
rect 48872 38981 48881 39015
rect 48881 38981 48915 39015
rect 48915 38981 48924 39015
rect 48872 38972 48924 38981
rect 49148 38972 49200 39024
rect 47584 38836 47636 38888
rect 48044 38879 48096 38888
rect 48044 38845 48053 38879
rect 48053 38845 48087 38879
rect 48087 38845 48096 38879
rect 48044 38836 48096 38845
rect 26056 38768 26108 38820
rect 26608 38811 26660 38820
rect 26608 38777 26617 38811
rect 26617 38777 26651 38811
rect 26651 38777 26660 38811
rect 26608 38768 26660 38777
rect 26700 38768 26752 38820
rect 47860 38768 47912 38820
rect 52552 38768 52604 38820
rect 52828 38879 52880 38888
rect 52828 38845 52837 38879
rect 52837 38845 52871 38879
rect 52871 38845 52880 38879
rect 53288 38879 53340 38888
rect 52828 38836 52880 38845
rect 53288 38845 53297 38879
rect 53297 38845 53331 38879
rect 53331 38845 53340 38879
rect 53288 38836 53340 38845
rect 53380 38879 53432 38888
rect 53380 38845 53389 38879
rect 53389 38845 53423 38879
rect 53423 38845 53432 38879
rect 53380 38836 53432 38845
rect 53564 38768 53616 38820
rect 16580 38700 16632 38752
rect 16856 38700 16908 38752
rect 20812 38743 20864 38752
rect 20812 38709 20821 38743
rect 20821 38709 20855 38743
rect 20855 38709 20864 38743
rect 20812 38700 20864 38709
rect 21180 38743 21232 38752
rect 21180 38709 21189 38743
rect 21189 38709 21223 38743
rect 21223 38709 21232 38743
rect 21180 38700 21232 38709
rect 24400 38700 24452 38752
rect 25412 38743 25464 38752
rect 25412 38709 25421 38743
rect 25421 38709 25455 38743
rect 25455 38709 25464 38743
rect 25412 38700 25464 38709
rect 34060 38700 34112 38752
rect 34152 38700 34204 38752
rect 36912 38700 36964 38752
rect 38476 38700 38528 38752
rect 39580 38700 39632 38752
rect 41696 38700 41748 38752
rect 42524 38700 42576 38752
rect 42892 38700 42944 38752
rect 43260 38743 43312 38752
rect 43260 38709 43269 38743
rect 43269 38709 43303 38743
rect 43303 38709 43312 38743
rect 43260 38700 43312 38709
rect 47584 38700 47636 38752
rect 48136 38700 48188 38752
rect 48412 38700 48464 38752
rect 48504 38743 48556 38752
rect 48504 38709 48513 38743
rect 48513 38709 48547 38743
rect 48547 38709 48556 38743
rect 48504 38700 48556 38709
rect 53748 38700 53800 38752
rect 56232 38972 56284 39024
rect 67640 39040 67692 39092
rect 69112 39040 69164 39092
rect 70952 39083 71004 39092
rect 70952 39049 70961 39083
rect 70961 39049 70995 39083
rect 70995 39049 71004 39083
rect 70952 39040 71004 39049
rect 56140 38904 56192 38956
rect 68744 38972 68796 39024
rect 72608 39083 72660 39092
rect 72608 39049 72617 39083
rect 72617 39049 72651 39083
rect 72651 39049 72660 39083
rect 72608 39040 72660 39049
rect 73988 39040 74040 39092
rect 75184 39083 75236 39092
rect 75184 39049 75193 39083
rect 75193 39049 75227 39083
rect 75227 39049 75236 39083
rect 75184 39040 75236 39049
rect 78956 39040 79008 39092
rect 63776 38947 63828 38956
rect 63776 38913 63785 38947
rect 63785 38913 63819 38947
rect 63819 38913 63828 38947
rect 63776 38904 63828 38913
rect 64052 38904 64104 38956
rect 64512 38904 64564 38956
rect 65524 38904 65576 38956
rect 55680 38879 55732 38888
rect 55680 38845 55689 38879
rect 55689 38845 55723 38879
rect 55723 38845 55732 38879
rect 55680 38836 55732 38845
rect 55772 38879 55824 38888
rect 55772 38845 55781 38879
rect 55781 38845 55815 38879
rect 55815 38845 55824 38879
rect 55772 38836 55824 38845
rect 56048 38879 56100 38888
rect 56048 38845 56057 38879
rect 56057 38845 56091 38879
rect 56091 38845 56100 38879
rect 56048 38836 56100 38845
rect 62304 38836 62356 38888
rect 63224 38879 63276 38888
rect 63224 38845 63233 38879
rect 63233 38845 63267 38879
rect 63267 38845 63276 38879
rect 63224 38836 63276 38845
rect 63684 38836 63736 38888
rect 64788 38836 64840 38888
rect 68560 38879 68612 38888
rect 68560 38845 68569 38879
rect 68569 38845 68603 38879
rect 68603 38845 68612 38879
rect 68560 38836 68612 38845
rect 55864 38768 55916 38820
rect 60832 38700 60884 38752
rect 62120 38768 62172 38820
rect 69480 38811 69532 38820
rect 69480 38777 69489 38811
rect 69489 38777 69523 38811
rect 69523 38777 69532 38811
rect 71412 38836 71464 38888
rect 72608 38836 72660 38888
rect 75736 38904 75788 38956
rect 77576 38904 77628 38956
rect 79784 38972 79836 39024
rect 82728 39040 82780 39092
rect 83464 39083 83516 39092
rect 83464 39049 83473 39083
rect 83473 39049 83507 39083
rect 83507 39049 83516 39083
rect 83464 39040 83516 39049
rect 84384 39040 84436 39092
rect 85304 39040 85356 39092
rect 80244 38972 80296 39024
rect 76380 38836 76432 38888
rect 77760 38879 77812 38888
rect 77760 38845 77769 38879
rect 77769 38845 77803 38879
rect 77803 38845 77812 38879
rect 77760 38836 77812 38845
rect 69480 38768 69532 38777
rect 76104 38768 76156 38820
rect 77024 38768 77076 38820
rect 79600 38904 79652 38956
rect 80336 38904 80388 38956
rect 83740 38947 83792 38956
rect 83740 38913 83749 38947
rect 83749 38913 83783 38947
rect 83783 38913 83792 38947
rect 83740 38904 83792 38913
rect 79784 38811 79836 38820
rect 79784 38777 79793 38811
rect 79793 38777 79827 38811
rect 79827 38777 79836 38811
rect 79784 38768 79836 38777
rect 83648 38879 83700 38888
rect 83648 38845 83662 38879
rect 83662 38845 83696 38879
rect 83696 38845 83700 38879
rect 83648 38836 83700 38845
rect 80244 38768 80296 38820
rect 65984 38700 66036 38752
rect 67272 38700 67324 38752
rect 68468 38700 68520 38752
rect 68744 38743 68796 38752
rect 68744 38709 68753 38743
rect 68753 38709 68787 38743
rect 68787 38709 68796 38743
rect 68744 38700 68796 38709
rect 69756 38700 69808 38752
rect 70308 38700 70360 38752
rect 76288 38700 76340 38752
rect 76656 38700 76708 38752
rect 77576 38700 77628 38752
rect 78220 38700 78272 38752
rect 83464 38768 83516 38820
rect 85212 38836 85264 38888
rect 85396 38879 85448 38888
rect 85396 38845 85405 38879
rect 85405 38845 85439 38879
rect 85439 38845 85448 38879
rect 85396 38836 85448 38845
rect 86776 38879 86828 38888
rect 86776 38845 86785 38879
rect 86785 38845 86819 38879
rect 86819 38845 86828 38879
rect 86776 38836 86828 38845
rect 80520 38700 80572 38752
rect 86408 38743 86460 38752
rect 86408 38709 86417 38743
rect 86417 38709 86451 38743
rect 86451 38709 86460 38743
rect 86408 38700 86460 38709
rect 87880 38743 87932 38752
rect 87880 38709 87889 38743
rect 87889 38709 87923 38743
rect 87923 38709 87932 38743
rect 87880 38700 87932 38709
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 50326 38598 50378 38650
rect 50390 38598 50442 38650
rect 50454 38598 50506 38650
rect 50518 38598 50570 38650
rect 81046 38598 81098 38650
rect 81110 38598 81162 38650
rect 81174 38598 81226 38650
rect 81238 38598 81290 38650
rect 3700 38496 3752 38548
rect 8116 38496 8168 38548
rect 9956 38539 10008 38548
rect 9956 38505 9965 38539
rect 9965 38505 9999 38539
rect 9999 38505 10008 38539
rect 9956 38496 10008 38505
rect 11244 38496 11296 38548
rect 13084 38539 13136 38548
rect 10416 38428 10468 38480
rect 10968 38428 11020 38480
rect 4436 38360 4488 38412
rect 5080 38360 5132 38412
rect 8024 38403 8076 38412
rect 8024 38369 8033 38403
rect 8033 38369 8067 38403
rect 8067 38369 8076 38403
rect 8024 38360 8076 38369
rect 8760 38403 8812 38412
rect 4620 38335 4672 38344
rect 4620 38301 4629 38335
rect 4629 38301 4663 38335
rect 4663 38301 4672 38335
rect 4620 38292 4672 38301
rect 5448 38292 5500 38344
rect 8760 38369 8769 38403
rect 8769 38369 8803 38403
rect 8803 38369 8812 38403
rect 8760 38360 8812 38369
rect 10784 38360 10836 38412
rect 11244 38360 11296 38412
rect 13084 38505 13093 38539
rect 13093 38505 13127 38539
rect 13127 38505 13136 38539
rect 13084 38496 13136 38505
rect 14188 38496 14240 38548
rect 16488 38539 16540 38548
rect 16488 38505 16497 38539
rect 16497 38505 16531 38539
rect 16531 38505 16540 38539
rect 16488 38496 16540 38505
rect 16580 38496 16632 38548
rect 17408 38496 17460 38548
rect 14464 38428 14516 38480
rect 19248 38496 19300 38548
rect 25412 38539 25464 38548
rect 25412 38505 25421 38539
rect 25421 38505 25455 38539
rect 25455 38505 25464 38539
rect 25412 38496 25464 38505
rect 27528 38496 27580 38548
rect 29644 38539 29696 38548
rect 22284 38428 22336 38480
rect 23940 38428 23992 38480
rect 26884 38428 26936 38480
rect 29644 38505 29653 38539
rect 29653 38505 29687 38539
rect 29687 38505 29696 38539
rect 29644 38496 29696 38505
rect 46020 38496 46072 38548
rect 46112 38496 46164 38548
rect 52552 38496 52604 38548
rect 51816 38428 51868 38480
rect 11980 38360 12032 38412
rect 10876 38292 10928 38344
rect 12164 38360 12216 38412
rect 14004 38360 14056 38412
rect 14832 38360 14884 38412
rect 10048 38224 10100 38276
rect 15384 38292 15436 38344
rect 15936 38360 15988 38412
rect 16580 38360 16632 38412
rect 20536 38360 20588 38412
rect 23848 38403 23900 38412
rect 23848 38369 23857 38403
rect 23857 38369 23891 38403
rect 23891 38369 23900 38403
rect 23848 38360 23900 38369
rect 24400 38403 24452 38412
rect 24400 38369 24407 38403
rect 24407 38369 24441 38403
rect 24441 38369 24452 38403
rect 24400 38360 24452 38369
rect 24584 38403 24636 38412
rect 24584 38369 24593 38403
rect 24593 38369 24627 38403
rect 24627 38369 24636 38403
rect 24584 38360 24636 38369
rect 26608 38360 26660 38412
rect 30656 38403 30708 38412
rect 25228 38335 25280 38344
rect 15200 38224 15252 38276
rect 25228 38301 25237 38335
rect 25237 38301 25271 38335
rect 25271 38301 25280 38335
rect 25228 38292 25280 38301
rect 25872 38292 25924 38344
rect 28356 38335 28408 38344
rect 28356 38301 28365 38335
rect 28365 38301 28399 38335
rect 28399 38301 28408 38335
rect 28356 38292 28408 38301
rect 30656 38369 30665 38403
rect 30665 38369 30699 38403
rect 30699 38369 30708 38403
rect 30656 38360 30708 38369
rect 31484 38360 31536 38412
rect 36544 38403 36596 38412
rect 36544 38369 36553 38403
rect 36553 38369 36587 38403
rect 36587 38369 36596 38403
rect 36544 38360 36596 38369
rect 37740 38403 37792 38412
rect 37740 38369 37749 38403
rect 37749 38369 37783 38403
rect 37783 38369 37792 38403
rect 37740 38360 37792 38369
rect 37924 38403 37976 38412
rect 37924 38369 37933 38403
rect 37933 38369 37967 38403
rect 37967 38369 37976 38403
rect 37924 38360 37976 38369
rect 38016 38360 38068 38412
rect 38476 38403 38528 38412
rect 38476 38369 38485 38403
rect 38485 38369 38519 38403
rect 38519 38369 38528 38403
rect 38476 38360 38528 38369
rect 38660 38360 38712 38412
rect 40868 38403 40920 38412
rect 40868 38369 40877 38403
rect 40877 38369 40911 38403
rect 40911 38369 40920 38403
rect 40868 38360 40920 38369
rect 32864 38292 32916 38344
rect 36452 38292 36504 38344
rect 43904 38360 43956 38412
rect 47676 38360 47728 38412
rect 50160 38360 50212 38412
rect 51724 38360 51776 38412
rect 41236 38335 41288 38344
rect 41236 38301 41245 38335
rect 41245 38301 41279 38335
rect 41279 38301 41288 38335
rect 41236 38292 41288 38301
rect 51540 38292 51592 38344
rect 51816 38335 51868 38344
rect 51816 38301 51825 38335
rect 51825 38301 51859 38335
rect 51859 38301 51868 38335
rect 51816 38292 51868 38301
rect 4712 38156 4764 38208
rect 14832 38156 14884 38208
rect 16948 38224 17000 38276
rect 18420 38156 18472 38208
rect 24124 38156 24176 38208
rect 26884 38156 26936 38208
rect 29092 38224 29144 38276
rect 38844 38224 38896 38276
rect 30748 38199 30800 38208
rect 30748 38165 30757 38199
rect 30757 38165 30791 38199
rect 30791 38165 30800 38199
rect 30748 38156 30800 38165
rect 33140 38156 33192 38208
rect 33232 38156 33284 38208
rect 40868 38224 40920 38276
rect 39488 38199 39540 38208
rect 39488 38165 39497 38199
rect 39497 38165 39531 38199
rect 39531 38165 39540 38199
rect 39488 38156 39540 38165
rect 39948 38156 40000 38208
rect 41512 38156 41564 38208
rect 42064 38156 42116 38208
rect 49700 38224 49752 38276
rect 50160 38224 50212 38276
rect 53380 38496 53432 38548
rect 57796 38496 57848 38548
rect 65524 38496 65576 38548
rect 68652 38496 68704 38548
rect 67640 38428 67692 38480
rect 59820 38360 59872 38412
rect 77760 38496 77812 38548
rect 83648 38496 83700 38548
rect 84016 38539 84068 38548
rect 84016 38505 84025 38539
rect 84025 38505 84059 38539
rect 84059 38505 84068 38539
rect 84016 38496 84068 38505
rect 70124 38403 70176 38412
rect 60280 38292 60332 38344
rect 61844 38224 61896 38276
rect 64420 38335 64472 38344
rect 64420 38301 64429 38335
rect 64429 38301 64463 38335
rect 64463 38301 64472 38335
rect 64420 38292 64472 38301
rect 70124 38369 70133 38403
rect 70133 38369 70167 38403
rect 70167 38369 70176 38403
rect 70124 38360 70176 38369
rect 70400 38360 70452 38412
rect 71872 38360 71924 38412
rect 76932 38428 76984 38480
rect 77024 38471 77076 38480
rect 77024 38437 77033 38471
rect 77033 38437 77067 38471
rect 77067 38437 77076 38471
rect 77024 38428 77076 38437
rect 77208 38428 77260 38480
rect 77392 38428 77444 38480
rect 82728 38428 82780 38480
rect 75736 38403 75788 38412
rect 75736 38369 75745 38403
rect 75745 38369 75779 38403
rect 75779 38369 75788 38403
rect 75736 38360 75788 38369
rect 65156 38292 65208 38344
rect 70308 38335 70360 38344
rect 70032 38224 70084 38276
rect 70308 38301 70317 38335
rect 70317 38301 70351 38335
rect 70351 38301 70360 38335
rect 70308 38292 70360 38301
rect 76104 38335 76156 38344
rect 76104 38301 76113 38335
rect 76113 38301 76147 38335
rect 76147 38301 76156 38335
rect 76104 38292 76156 38301
rect 77300 38360 77352 38412
rect 78404 38360 78456 38412
rect 83556 38403 83608 38412
rect 83556 38369 83565 38403
rect 83565 38369 83599 38403
rect 83599 38369 83608 38403
rect 83556 38360 83608 38369
rect 86316 38428 86368 38480
rect 86776 38428 86828 38480
rect 85856 38403 85908 38412
rect 77668 38335 77720 38344
rect 77668 38301 77677 38335
rect 77677 38301 77711 38335
rect 77711 38301 77720 38335
rect 77668 38292 77720 38301
rect 85856 38369 85865 38403
rect 85865 38369 85899 38403
rect 85899 38369 85908 38403
rect 85856 38360 85908 38369
rect 85948 38403 86000 38412
rect 85948 38369 85957 38403
rect 85957 38369 85991 38403
rect 85991 38369 86000 38403
rect 85948 38360 86000 38369
rect 75644 38224 75696 38276
rect 76380 38267 76432 38276
rect 76380 38233 76389 38267
rect 76389 38233 76423 38267
rect 76423 38233 76432 38267
rect 76380 38224 76432 38233
rect 77484 38224 77536 38276
rect 46296 38199 46348 38208
rect 46296 38165 46305 38199
rect 46305 38165 46339 38199
rect 46339 38165 46348 38199
rect 47676 38199 47728 38208
rect 46296 38156 46348 38165
rect 47676 38165 47685 38199
rect 47685 38165 47719 38199
rect 47719 38165 47728 38199
rect 47676 38156 47728 38165
rect 47768 38156 47820 38208
rect 52828 38156 52880 38208
rect 53104 38156 53156 38208
rect 53380 38199 53432 38208
rect 53380 38165 53389 38199
rect 53389 38165 53423 38199
rect 53423 38165 53432 38199
rect 53380 38156 53432 38165
rect 64512 38156 64564 38208
rect 64880 38199 64932 38208
rect 64880 38165 64889 38199
rect 64889 38165 64923 38199
rect 64923 38165 64932 38199
rect 64880 38156 64932 38165
rect 67640 38156 67692 38208
rect 68928 38156 68980 38208
rect 76288 38156 76340 38208
rect 78404 38199 78456 38208
rect 78404 38165 78413 38199
rect 78413 38165 78447 38199
rect 78447 38165 78456 38199
rect 78404 38156 78456 38165
rect 82820 38156 82872 38208
rect 84752 38156 84804 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 65686 38054 65738 38106
rect 65750 38054 65802 38106
rect 65814 38054 65866 38106
rect 65878 38054 65930 38106
rect 96406 38054 96458 38106
rect 96470 38054 96522 38106
rect 96534 38054 96586 38106
rect 96598 38054 96650 38106
rect 3976 37995 4028 38004
rect 3976 37961 3985 37995
rect 3985 37961 4019 37995
rect 4019 37961 4028 37995
rect 3976 37952 4028 37961
rect 6092 37995 6144 38004
rect 6092 37961 6101 37995
rect 6101 37961 6135 37995
rect 6135 37961 6144 37995
rect 6092 37952 6144 37961
rect 9864 37952 9916 38004
rect 12164 37952 12216 38004
rect 14188 37995 14240 38004
rect 14188 37961 14197 37995
rect 14197 37961 14231 37995
rect 14231 37961 14240 37995
rect 14188 37952 14240 37961
rect 14280 37952 14332 38004
rect 16396 37952 16448 38004
rect 16488 37952 16540 38004
rect 20536 37995 20588 38004
rect 3884 37884 3936 37936
rect 2596 37859 2648 37868
rect 2596 37825 2605 37859
rect 2605 37825 2639 37859
rect 2639 37825 2648 37859
rect 2596 37816 2648 37825
rect 4528 37816 4580 37868
rect 5080 37816 5132 37868
rect 5264 37791 5316 37800
rect 5264 37757 5273 37791
rect 5273 37757 5307 37791
rect 5307 37757 5316 37791
rect 5264 37748 5316 37757
rect 6092 37748 6144 37800
rect 10048 37816 10100 37868
rect 10600 37791 10652 37800
rect 5908 37680 5960 37732
rect 10140 37723 10192 37732
rect 10140 37689 10149 37723
rect 10149 37689 10183 37723
rect 10183 37689 10192 37723
rect 10140 37680 10192 37689
rect 10600 37757 10609 37791
rect 10609 37757 10643 37791
rect 10643 37757 10652 37791
rect 10600 37748 10652 37757
rect 10968 37816 11020 37868
rect 11428 37884 11480 37936
rect 18420 37884 18472 37936
rect 20536 37961 20545 37995
rect 20545 37961 20579 37995
rect 20579 37961 20588 37995
rect 20536 37952 20588 37961
rect 21180 37884 21232 37936
rect 29092 37884 29144 37936
rect 30656 37927 30708 37936
rect 30656 37893 30665 37927
rect 30665 37893 30699 37927
rect 30699 37893 30708 37927
rect 30656 37884 30708 37893
rect 31576 37884 31628 37936
rect 32680 37884 32732 37936
rect 33232 37884 33284 37936
rect 34428 37884 34480 37936
rect 36636 37952 36688 38004
rect 47768 37952 47820 38004
rect 51632 37952 51684 38004
rect 14464 37816 14516 37868
rect 15200 37816 15252 37868
rect 10876 37748 10928 37800
rect 12624 37748 12676 37800
rect 14280 37748 14332 37800
rect 15292 37680 15344 37732
rect 15936 37791 15988 37800
rect 15936 37757 15945 37791
rect 15945 37757 15979 37791
rect 15979 37757 15988 37791
rect 15936 37748 15988 37757
rect 16304 37748 16356 37800
rect 16580 37748 16632 37800
rect 16856 37748 16908 37800
rect 17684 37748 17736 37800
rect 18972 37791 19024 37800
rect 18972 37757 18981 37791
rect 18981 37757 19015 37791
rect 19015 37757 19024 37791
rect 18972 37748 19024 37757
rect 19248 37791 19300 37800
rect 19248 37757 19257 37791
rect 19257 37757 19291 37791
rect 19291 37757 19300 37791
rect 19248 37748 19300 37757
rect 26148 37816 26200 37868
rect 32128 37859 32180 37868
rect 32128 37825 32137 37859
rect 32137 37825 32171 37859
rect 32171 37825 32180 37859
rect 32128 37816 32180 37825
rect 42064 37884 42116 37936
rect 35992 37816 36044 37868
rect 36176 37816 36228 37868
rect 41420 37816 41472 37868
rect 46020 37884 46072 37936
rect 49240 37884 49292 37936
rect 53564 37952 53616 38004
rect 25504 37748 25556 37800
rect 26056 37791 26108 37800
rect 26056 37757 26065 37791
rect 26065 37757 26099 37791
rect 26099 37757 26108 37791
rect 26056 37748 26108 37757
rect 25412 37680 25464 37732
rect 26884 37748 26936 37800
rect 29092 37748 29144 37800
rect 29276 37791 29328 37800
rect 29276 37757 29292 37791
rect 29292 37757 29326 37791
rect 29326 37757 29328 37791
rect 29276 37748 29328 37757
rect 27068 37680 27120 37732
rect 30748 37748 30800 37800
rect 36636 37748 36688 37800
rect 38016 37791 38068 37800
rect 38016 37757 38025 37791
rect 38025 37757 38059 37791
rect 38059 37757 38068 37791
rect 38016 37748 38068 37757
rect 40592 37748 40644 37800
rect 41880 37748 41932 37800
rect 4528 37655 4580 37664
rect 4528 37621 4537 37655
rect 4537 37621 4571 37655
rect 4571 37621 4580 37655
rect 4528 37612 4580 37621
rect 4620 37612 4672 37664
rect 6920 37655 6972 37664
rect 6920 37621 6929 37655
rect 6929 37621 6963 37655
rect 6963 37621 6972 37655
rect 6920 37612 6972 37621
rect 15568 37655 15620 37664
rect 15568 37621 15577 37655
rect 15577 37621 15611 37655
rect 15611 37621 15620 37655
rect 15568 37612 15620 37621
rect 16304 37612 16356 37664
rect 25504 37655 25556 37664
rect 25504 37621 25513 37655
rect 25513 37621 25547 37655
rect 25547 37621 25556 37655
rect 25504 37612 25556 37621
rect 26056 37612 26108 37664
rect 26700 37612 26752 37664
rect 30380 37680 30432 37732
rect 33416 37680 33468 37732
rect 36544 37680 36596 37732
rect 30288 37612 30340 37664
rect 31576 37655 31628 37664
rect 31576 37621 31585 37655
rect 31585 37621 31619 37655
rect 31619 37621 31628 37655
rect 31576 37612 31628 37621
rect 38200 37612 38252 37664
rect 41420 37612 41472 37664
rect 41604 37612 41656 37664
rect 42616 37748 42668 37800
rect 51816 37816 51868 37868
rect 53380 37816 53432 37868
rect 54024 37859 54076 37868
rect 54024 37825 54033 37859
rect 54033 37825 54067 37859
rect 54067 37825 54076 37859
rect 54024 37816 54076 37825
rect 44180 37680 44232 37732
rect 46112 37680 46164 37732
rect 46296 37680 46348 37732
rect 47676 37748 47728 37800
rect 48688 37748 48740 37800
rect 52000 37748 52052 37800
rect 51908 37680 51960 37732
rect 52644 37748 52696 37800
rect 53656 37748 53708 37800
rect 53932 37791 53984 37800
rect 53932 37757 53941 37791
rect 53941 37757 53975 37791
rect 53975 37757 53984 37791
rect 53932 37748 53984 37757
rect 58716 37952 58768 38004
rect 57704 37859 57756 37868
rect 57704 37825 57713 37859
rect 57713 37825 57747 37859
rect 57747 37825 57756 37859
rect 57704 37816 57756 37825
rect 61752 37952 61804 38004
rect 64420 37952 64472 38004
rect 65156 37995 65208 38004
rect 65156 37961 65165 37995
rect 65165 37961 65199 37995
rect 65199 37961 65208 37995
rect 65156 37952 65208 37961
rect 69020 37952 69072 38004
rect 70308 37952 70360 38004
rect 76104 37952 76156 38004
rect 77116 37952 77168 38004
rect 83740 37952 83792 38004
rect 86316 37952 86368 38004
rect 64512 37859 64564 37868
rect 64512 37825 64521 37859
rect 64521 37825 64555 37859
rect 64555 37825 64564 37859
rect 75736 37859 75788 37868
rect 64512 37816 64564 37825
rect 58624 37791 58676 37800
rect 58624 37757 58633 37791
rect 58633 37757 58667 37791
rect 58667 37757 58676 37791
rect 58624 37748 58676 37757
rect 60280 37791 60332 37800
rect 60280 37757 60289 37791
rect 60289 37757 60323 37791
rect 60323 37757 60332 37791
rect 60280 37748 60332 37757
rect 61844 37748 61896 37800
rect 43444 37612 43496 37664
rect 47032 37612 47084 37664
rect 52092 37655 52144 37664
rect 52092 37621 52101 37655
rect 52101 37621 52135 37655
rect 52135 37621 52144 37655
rect 52092 37612 52144 37621
rect 52184 37612 52236 37664
rect 62120 37680 62172 37732
rect 65156 37748 65208 37800
rect 64880 37680 64932 37732
rect 75736 37825 75745 37859
rect 75745 37825 75779 37859
rect 75779 37825 75788 37859
rect 75736 37816 75788 37825
rect 69020 37748 69072 37800
rect 69572 37791 69624 37800
rect 69572 37757 69581 37791
rect 69581 37757 69615 37791
rect 69615 37757 69624 37791
rect 69572 37748 69624 37757
rect 57152 37612 57204 37664
rect 67456 37612 67508 37664
rect 70676 37655 70728 37664
rect 70676 37621 70685 37655
rect 70685 37621 70719 37655
rect 70719 37621 70728 37655
rect 70676 37612 70728 37621
rect 71136 37612 71188 37664
rect 75644 37791 75696 37800
rect 75644 37757 75653 37791
rect 75653 37757 75687 37791
rect 75687 37757 75696 37791
rect 78404 37816 78456 37868
rect 80336 37816 80388 37868
rect 84752 37816 84804 37868
rect 85856 37859 85908 37868
rect 85856 37825 85865 37859
rect 85865 37825 85899 37859
rect 85899 37825 85908 37859
rect 85856 37816 85908 37825
rect 75644 37748 75696 37757
rect 76932 37791 76984 37800
rect 71688 37680 71740 37732
rect 76932 37757 76941 37791
rect 76941 37757 76975 37791
rect 76975 37757 76984 37791
rect 76932 37748 76984 37757
rect 82728 37791 82780 37800
rect 82728 37757 82737 37791
rect 82737 37757 82771 37791
rect 82771 37757 82780 37791
rect 82728 37748 82780 37757
rect 82636 37680 82688 37732
rect 85304 37748 85356 37800
rect 87880 37816 87932 37868
rect 86776 37791 86828 37800
rect 86776 37757 86785 37791
rect 86785 37757 86819 37791
rect 86819 37757 86828 37791
rect 86776 37748 86828 37757
rect 77944 37612 77996 37664
rect 80152 37612 80204 37664
rect 82820 37655 82872 37664
rect 82820 37621 82829 37655
rect 82829 37621 82863 37655
rect 82863 37621 82872 37655
rect 82820 37612 82872 37621
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 81046 37510 81098 37562
rect 81110 37510 81162 37562
rect 81174 37510 81226 37562
rect 81238 37510 81290 37562
rect 4804 37272 4856 37324
rect 10048 37451 10100 37460
rect 10048 37417 10057 37451
rect 10057 37417 10091 37451
rect 10091 37417 10100 37451
rect 10048 37408 10100 37417
rect 8300 37340 8352 37392
rect 10968 37340 11020 37392
rect 6920 37272 6972 37324
rect 9864 37315 9916 37324
rect 9864 37281 9873 37315
rect 9873 37281 9907 37315
rect 9907 37281 9916 37315
rect 9864 37272 9916 37281
rect 11428 37315 11480 37324
rect 11428 37281 11437 37315
rect 11437 37281 11471 37315
rect 11471 37281 11480 37315
rect 11428 37272 11480 37281
rect 13544 37340 13596 37392
rect 11980 37315 12032 37324
rect 11980 37281 11989 37315
rect 11989 37281 12023 37315
rect 12023 37281 12032 37315
rect 11980 37272 12032 37281
rect 15568 37408 15620 37460
rect 16488 37451 16540 37460
rect 16488 37417 16497 37451
rect 16497 37417 16531 37451
rect 16531 37417 16540 37451
rect 16488 37408 16540 37417
rect 16580 37408 16632 37460
rect 21088 37451 21140 37460
rect 21088 37417 21097 37451
rect 21097 37417 21131 37451
rect 21131 37417 21140 37451
rect 21088 37408 21140 37417
rect 25412 37408 25464 37460
rect 26056 37451 26108 37460
rect 26056 37417 26065 37451
rect 26065 37417 26099 37451
rect 26099 37417 26108 37451
rect 26056 37408 26108 37417
rect 26148 37408 26200 37460
rect 52092 37408 52144 37460
rect 52828 37408 52880 37460
rect 15384 37340 15436 37392
rect 3516 37204 3568 37256
rect 4896 37204 4948 37256
rect 4068 37136 4120 37188
rect 4712 37136 4764 37188
rect 15476 37315 15528 37324
rect 15476 37281 15485 37315
rect 15485 37281 15519 37315
rect 15519 37281 15528 37315
rect 17776 37340 17828 37392
rect 15476 37272 15528 37281
rect 16948 37272 17000 37324
rect 17684 37315 17736 37324
rect 17684 37281 17693 37315
rect 17693 37281 17727 37315
rect 17727 37281 17736 37315
rect 17684 37272 17736 37281
rect 18420 37315 18472 37324
rect 18420 37281 18429 37315
rect 18429 37281 18463 37315
rect 18463 37281 18472 37315
rect 18420 37272 18472 37281
rect 19248 37340 19300 37392
rect 20812 37272 20864 37324
rect 20904 37315 20956 37324
rect 20904 37281 20913 37315
rect 20913 37281 20947 37315
rect 20947 37281 20956 37315
rect 20904 37272 20956 37281
rect 21824 37272 21876 37324
rect 16488 37136 16540 37188
rect 6368 37111 6420 37120
rect 6368 37077 6377 37111
rect 6377 37077 6411 37111
rect 6411 37077 6420 37111
rect 6368 37068 6420 37077
rect 14924 37068 14976 37120
rect 24768 37136 24820 37188
rect 26700 37315 26752 37324
rect 26700 37281 26709 37315
rect 26709 37281 26743 37315
rect 26743 37281 26752 37315
rect 26700 37272 26752 37281
rect 27252 37315 27304 37324
rect 27252 37281 27261 37315
rect 27261 37281 27295 37315
rect 27295 37281 27304 37315
rect 27252 37272 27304 37281
rect 27436 37315 27488 37324
rect 27436 37281 27445 37315
rect 27445 37281 27479 37315
rect 27479 37281 27488 37315
rect 27436 37272 27488 37281
rect 28356 37340 28408 37392
rect 29000 37340 29052 37392
rect 30380 37340 30432 37392
rect 30840 37272 30892 37324
rect 31668 37315 31720 37324
rect 31668 37281 31677 37315
rect 31677 37281 31711 37315
rect 31711 37281 31720 37315
rect 31668 37272 31720 37281
rect 34428 37272 34480 37324
rect 37096 37340 37148 37392
rect 39764 37340 39816 37392
rect 38200 37272 38252 37324
rect 38292 37272 38344 37324
rect 26056 37204 26108 37256
rect 35440 37247 35492 37256
rect 21364 37068 21416 37120
rect 30564 37136 30616 37188
rect 30472 37111 30524 37120
rect 30472 37077 30481 37111
rect 30481 37077 30515 37111
rect 30515 37077 30524 37111
rect 30472 37068 30524 37077
rect 31484 37111 31536 37120
rect 31484 37077 31493 37111
rect 31493 37077 31527 37111
rect 31527 37077 31536 37111
rect 31484 37068 31536 37077
rect 34612 37068 34664 37120
rect 35440 37213 35449 37247
rect 35449 37213 35483 37247
rect 35483 37213 35492 37247
rect 35440 37204 35492 37213
rect 40592 37315 40644 37324
rect 40592 37281 40601 37315
rect 40601 37281 40635 37315
rect 40635 37281 40644 37315
rect 40592 37272 40644 37281
rect 42616 37340 42668 37392
rect 48688 37340 48740 37392
rect 49700 37383 49752 37392
rect 49700 37349 49709 37383
rect 49709 37349 49743 37383
rect 49743 37349 49752 37383
rect 49700 37340 49752 37349
rect 41880 37272 41932 37324
rect 43352 37272 43404 37324
rect 47216 37272 47268 37324
rect 51724 37340 51776 37392
rect 50988 37272 51040 37324
rect 52000 37272 52052 37324
rect 53012 37315 53064 37324
rect 53012 37281 53021 37315
rect 53021 37281 53055 37315
rect 53055 37281 53064 37315
rect 53012 37272 53064 37281
rect 53104 37315 53156 37324
rect 53104 37281 53113 37315
rect 53113 37281 53147 37315
rect 53147 37281 53156 37315
rect 53104 37272 53156 37281
rect 53472 37315 53524 37324
rect 53472 37281 53481 37315
rect 53481 37281 53515 37315
rect 53515 37281 53524 37315
rect 53472 37272 53524 37281
rect 53656 37272 53708 37324
rect 57060 37408 57112 37460
rect 57244 37451 57296 37460
rect 57244 37417 57253 37451
rect 57253 37417 57287 37451
rect 57287 37417 57296 37451
rect 57244 37408 57296 37417
rect 57704 37451 57756 37460
rect 55312 37315 55364 37324
rect 55312 37281 55321 37315
rect 55321 37281 55355 37315
rect 55355 37281 55364 37315
rect 55312 37272 55364 37281
rect 57704 37417 57713 37451
rect 57713 37417 57747 37451
rect 57747 37417 57756 37451
rect 57704 37408 57756 37417
rect 57796 37408 57848 37460
rect 60556 37408 60608 37460
rect 61844 37451 61896 37460
rect 61844 37417 61853 37451
rect 61853 37417 61887 37451
rect 61887 37417 61896 37451
rect 61844 37408 61896 37417
rect 64788 37408 64840 37460
rect 67180 37451 67232 37460
rect 67180 37417 67189 37451
rect 67189 37417 67223 37451
rect 67223 37417 67232 37451
rect 67180 37408 67232 37417
rect 64052 37340 64104 37392
rect 58716 37315 58768 37324
rect 58716 37281 58725 37315
rect 58725 37281 58759 37315
rect 58759 37281 58768 37315
rect 58716 37272 58768 37281
rect 61752 37315 61804 37324
rect 50344 37204 50396 37256
rect 57704 37204 57756 37256
rect 59820 37204 59872 37256
rect 61752 37281 61761 37315
rect 61761 37281 61795 37315
rect 61795 37281 61804 37315
rect 61752 37272 61804 37281
rect 62580 37315 62632 37324
rect 62580 37281 62589 37315
rect 62589 37281 62623 37315
rect 62623 37281 62632 37315
rect 62580 37272 62632 37281
rect 63592 37272 63644 37324
rect 63684 37272 63736 37324
rect 64328 37272 64380 37324
rect 66260 37315 66312 37324
rect 66260 37281 66269 37315
rect 66269 37281 66303 37315
rect 66303 37281 66312 37315
rect 66260 37272 66312 37281
rect 66444 37315 66496 37324
rect 66444 37281 66453 37315
rect 66453 37281 66487 37315
rect 66487 37281 66496 37315
rect 66444 37272 66496 37281
rect 66628 37272 66680 37324
rect 82636 37408 82688 37460
rect 82728 37408 82780 37460
rect 69572 37340 69624 37392
rect 71136 37383 71188 37392
rect 67456 37272 67508 37324
rect 69112 37272 69164 37324
rect 71136 37349 71145 37383
rect 71145 37349 71179 37383
rect 71179 37349 71188 37383
rect 71136 37340 71188 37349
rect 70032 37315 70084 37324
rect 70032 37281 70041 37315
rect 70041 37281 70075 37315
rect 70075 37281 70084 37315
rect 70032 37272 70084 37281
rect 70124 37272 70176 37324
rect 70308 37315 70360 37324
rect 70308 37281 70317 37315
rect 70317 37281 70351 37315
rect 70351 37281 70360 37315
rect 70308 37272 70360 37281
rect 71688 37315 71740 37324
rect 71688 37281 71697 37315
rect 71697 37281 71731 37315
rect 71731 37281 71740 37315
rect 71688 37272 71740 37281
rect 76932 37340 76984 37392
rect 72056 37272 72108 37324
rect 77208 37315 77260 37324
rect 77208 37281 77217 37315
rect 77217 37281 77251 37315
rect 77251 37281 77260 37315
rect 77208 37272 77260 37281
rect 77484 37272 77536 37324
rect 66168 37204 66220 37256
rect 66720 37247 66772 37256
rect 66720 37213 66729 37247
rect 66729 37213 66763 37247
rect 66763 37213 66772 37247
rect 66720 37204 66772 37213
rect 75184 37204 75236 37256
rect 80336 37340 80388 37392
rect 78680 37272 78732 37324
rect 83188 37340 83240 37392
rect 40868 37068 40920 37120
rect 46112 37068 46164 37120
rect 50988 37068 51040 37120
rect 52460 37111 52512 37120
rect 52460 37077 52469 37111
rect 52469 37077 52503 37111
rect 52503 37077 52512 37111
rect 52460 37068 52512 37077
rect 54392 37068 54444 37120
rect 54852 37068 54904 37120
rect 69940 37136 69992 37188
rect 77944 37204 77996 37256
rect 86408 37340 86460 37392
rect 86868 37340 86920 37392
rect 84752 37272 84804 37324
rect 85948 37272 86000 37324
rect 86224 37315 86276 37324
rect 86224 37281 86233 37315
rect 86233 37281 86267 37315
rect 86267 37281 86276 37315
rect 86224 37272 86276 37281
rect 87420 37272 87472 37324
rect 65984 37068 66036 37120
rect 66168 37068 66220 37120
rect 67732 37068 67784 37120
rect 68652 37068 68704 37120
rect 70676 37068 70728 37120
rect 77024 37068 77076 37120
rect 80428 37068 80480 37120
rect 83556 37068 83608 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 65686 36966 65738 37018
rect 65750 36966 65802 37018
rect 65814 36966 65866 37018
rect 65878 36966 65930 37018
rect 96406 36966 96458 37018
rect 96470 36966 96522 37018
rect 96534 36966 96586 37018
rect 96598 36966 96650 37018
rect 10876 36864 10928 36916
rect 18236 36864 18288 36916
rect 5540 36796 5592 36848
rect 26608 36864 26660 36916
rect 30472 36864 30524 36916
rect 41328 36864 41380 36916
rect 41512 36907 41564 36916
rect 41512 36873 41521 36907
rect 41521 36873 41555 36907
rect 41555 36873 41564 36907
rect 41512 36864 41564 36873
rect 43996 36864 44048 36916
rect 46848 36864 46900 36916
rect 51632 36864 51684 36916
rect 51816 36907 51868 36916
rect 51816 36873 51825 36907
rect 51825 36873 51859 36907
rect 51859 36873 51868 36907
rect 51816 36864 51868 36873
rect 54392 36864 54444 36916
rect 54484 36864 54536 36916
rect 60648 36864 60700 36916
rect 60740 36864 60792 36916
rect 5264 36703 5316 36712
rect 5264 36669 5273 36703
rect 5273 36669 5307 36703
rect 5307 36669 5316 36703
rect 5264 36660 5316 36669
rect 8852 36660 8904 36712
rect 10784 36703 10836 36712
rect 10784 36669 10793 36703
rect 10793 36669 10827 36703
rect 10827 36669 10836 36703
rect 10784 36660 10836 36669
rect 15476 36728 15528 36780
rect 18420 36728 18472 36780
rect 16488 36660 16540 36712
rect 17224 36660 17276 36712
rect 21364 36796 21416 36848
rect 25412 36796 25464 36848
rect 19892 36660 19944 36712
rect 20168 36703 20220 36712
rect 20168 36669 20177 36703
rect 20177 36669 20211 36703
rect 20211 36669 20220 36703
rect 20168 36660 20220 36669
rect 21088 36660 21140 36712
rect 21732 36703 21784 36712
rect 21732 36669 21741 36703
rect 21741 36669 21775 36703
rect 21775 36669 21784 36703
rect 21732 36660 21784 36669
rect 25412 36660 25464 36712
rect 25596 36703 25648 36712
rect 25596 36669 25605 36703
rect 25605 36669 25639 36703
rect 25639 36669 25648 36703
rect 25596 36660 25648 36669
rect 33140 36796 33192 36848
rect 35992 36839 36044 36848
rect 27160 36728 27212 36780
rect 27436 36728 27488 36780
rect 34612 36728 34664 36780
rect 35992 36805 36001 36839
rect 36001 36805 36035 36839
rect 36035 36805 36044 36839
rect 35992 36796 36044 36805
rect 39764 36796 39816 36848
rect 41420 36796 41472 36848
rect 39488 36728 39540 36780
rect 41696 36728 41748 36780
rect 46940 36796 46992 36848
rect 47216 36839 47268 36848
rect 47216 36805 47225 36839
rect 47225 36805 47259 36839
rect 47259 36805 47268 36839
rect 47216 36796 47268 36805
rect 47308 36796 47360 36848
rect 50712 36796 50764 36848
rect 53472 36796 53524 36848
rect 70952 36864 71004 36916
rect 71136 36907 71188 36916
rect 71136 36873 71145 36907
rect 71145 36873 71179 36907
rect 71179 36873 71188 36907
rect 71136 36864 71188 36873
rect 77024 36864 77076 36916
rect 82912 36907 82964 36916
rect 82912 36873 82921 36907
rect 82921 36873 82955 36907
rect 82955 36873 82964 36907
rect 82912 36864 82964 36873
rect 83188 36864 83240 36916
rect 5172 36567 5224 36576
rect 5172 36533 5181 36567
rect 5181 36533 5215 36567
rect 5215 36533 5224 36567
rect 5172 36524 5224 36533
rect 14924 36567 14976 36576
rect 14924 36533 14933 36567
rect 14933 36533 14967 36567
rect 14967 36533 14976 36567
rect 14924 36524 14976 36533
rect 19340 36524 19392 36576
rect 20168 36524 20220 36576
rect 24860 36592 24912 36644
rect 32404 36592 32456 36644
rect 20720 36567 20772 36576
rect 20720 36533 20729 36567
rect 20729 36533 20763 36567
rect 20763 36533 20772 36567
rect 20720 36524 20772 36533
rect 21548 36524 21600 36576
rect 25412 36524 25464 36576
rect 25596 36524 25648 36576
rect 35624 36703 35676 36712
rect 35624 36669 35633 36703
rect 35633 36669 35667 36703
rect 35667 36669 35676 36703
rect 35624 36660 35676 36669
rect 35808 36703 35860 36712
rect 35808 36669 35817 36703
rect 35817 36669 35851 36703
rect 35851 36669 35860 36703
rect 35808 36660 35860 36669
rect 35992 36660 36044 36712
rect 41328 36660 41380 36712
rect 40868 36635 40920 36644
rect 40868 36601 40877 36635
rect 40877 36601 40911 36635
rect 40911 36601 40920 36635
rect 40868 36592 40920 36601
rect 36544 36524 36596 36576
rect 36636 36524 36688 36576
rect 43996 36660 44048 36712
rect 44180 36703 44232 36712
rect 44180 36669 44189 36703
rect 44189 36669 44223 36703
rect 44223 36669 44232 36703
rect 44180 36660 44232 36669
rect 44548 36703 44600 36712
rect 44548 36669 44562 36703
rect 44562 36669 44600 36703
rect 44548 36660 44600 36669
rect 46112 36703 46164 36712
rect 46112 36669 46121 36703
rect 46121 36669 46155 36703
rect 46155 36669 46164 36703
rect 46112 36660 46164 36669
rect 49240 36728 49292 36780
rect 53748 36771 53800 36780
rect 53748 36737 53757 36771
rect 53757 36737 53791 36771
rect 53791 36737 53800 36771
rect 53748 36728 53800 36737
rect 71504 36839 71556 36848
rect 71504 36805 71513 36839
rect 71513 36805 71547 36839
rect 71547 36805 71556 36839
rect 71504 36796 71556 36805
rect 75184 36796 75236 36848
rect 80152 36796 80204 36848
rect 83924 36864 83976 36916
rect 86960 36907 87012 36916
rect 86960 36873 86969 36907
rect 86969 36873 87003 36907
rect 87003 36873 87012 36907
rect 86960 36864 87012 36873
rect 54300 36728 54352 36780
rect 46848 36703 46900 36712
rect 46848 36669 46857 36703
rect 46857 36669 46891 36703
rect 46891 36669 46900 36703
rect 46848 36660 46900 36669
rect 47032 36703 47084 36712
rect 47032 36669 47041 36703
rect 47041 36669 47075 36703
rect 47075 36669 47084 36703
rect 47032 36660 47084 36669
rect 48412 36660 48464 36712
rect 49700 36703 49752 36712
rect 49700 36669 49709 36703
rect 49709 36669 49743 36703
rect 49743 36669 49752 36703
rect 49700 36660 49752 36669
rect 50804 36660 50856 36712
rect 51724 36703 51776 36712
rect 51724 36669 51733 36703
rect 51733 36669 51767 36703
rect 51767 36669 51776 36703
rect 51724 36660 51776 36669
rect 53656 36703 53708 36712
rect 53656 36669 53665 36703
rect 53665 36669 53699 36703
rect 53699 36669 53708 36703
rect 53656 36660 53708 36669
rect 53932 36660 53984 36712
rect 54208 36660 54260 36712
rect 61108 36660 61160 36712
rect 66628 36771 66680 36780
rect 41512 36524 41564 36576
rect 42524 36567 42576 36576
rect 42524 36533 42533 36567
rect 42533 36533 42567 36567
rect 42567 36533 42576 36567
rect 42524 36524 42576 36533
rect 54852 36592 54904 36644
rect 62120 36592 62172 36644
rect 51632 36524 51684 36576
rect 55036 36524 55088 36576
rect 56600 36524 56652 36576
rect 63592 36660 63644 36712
rect 63776 36660 63828 36712
rect 64512 36660 64564 36712
rect 65432 36660 65484 36712
rect 66628 36737 66637 36771
rect 66637 36737 66671 36771
rect 66671 36737 66680 36771
rect 66628 36728 66680 36737
rect 71136 36728 71188 36780
rect 71596 36771 71648 36780
rect 71596 36737 71605 36771
rect 71605 36737 71639 36771
rect 71639 36737 71648 36771
rect 71596 36728 71648 36737
rect 71964 36728 72016 36780
rect 66168 36703 66220 36712
rect 66168 36669 66177 36703
rect 66177 36669 66211 36703
rect 66211 36669 66220 36703
rect 66444 36703 66496 36712
rect 66168 36660 66220 36669
rect 66444 36669 66453 36703
rect 66453 36669 66487 36703
rect 66487 36669 66496 36703
rect 66444 36660 66496 36669
rect 68652 36703 68704 36712
rect 68652 36669 68661 36703
rect 68661 36669 68695 36703
rect 68695 36669 68704 36703
rect 68652 36660 68704 36669
rect 69756 36703 69808 36712
rect 69756 36669 69765 36703
rect 69765 36669 69799 36703
rect 69799 36669 69808 36703
rect 69756 36660 69808 36669
rect 69940 36703 69992 36712
rect 69940 36669 69949 36703
rect 69949 36669 69983 36703
rect 69983 36669 69992 36703
rect 69940 36660 69992 36669
rect 72608 36660 72660 36712
rect 72792 36703 72844 36712
rect 72792 36669 72801 36703
rect 72801 36669 72835 36703
rect 72835 36669 72844 36703
rect 72792 36660 72844 36669
rect 76840 36660 76892 36712
rect 78220 36703 78272 36712
rect 64604 36524 64656 36576
rect 70308 36592 70360 36644
rect 70584 36592 70636 36644
rect 70124 36524 70176 36576
rect 74448 36592 74500 36644
rect 78220 36669 78229 36703
rect 78229 36669 78263 36703
rect 78263 36669 78272 36703
rect 78220 36660 78272 36669
rect 83556 36728 83608 36780
rect 85948 36771 86000 36780
rect 85948 36737 85957 36771
rect 85957 36737 85991 36771
rect 85991 36737 86000 36771
rect 85948 36728 86000 36737
rect 87420 36771 87472 36780
rect 87420 36737 87429 36771
rect 87429 36737 87463 36771
rect 87463 36737 87472 36771
rect 87420 36728 87472 36737
rect 82176 36703 82228 36712
rect 82176 36669 82185 36703
rect 82185 36669 82219 36703
rect 82219 36669 82228 36703
rect 82176 36660 82228 36669
rect 83924 36703 83976 36712
rect 83924 36669 83933 36703
rect 83933 36669 83967 36703
rect 83967 36669 83976 36703
rect 84200 36703 84252 36712
rect 83924 36660 83976 36669
rect 84200 36669 84209 36703
rect 84209 36669 84243 36703
rect 84243 36669 84252 36703
rect 84200 36660 84252 36669
rect 77208 36567 77260 36576
rect 77208 36533 77217 36567
rect 77217 36533 77251 36567
rect 77251 36533 77260 36567
rect 77208 36524 77260 36533
rect 77852 36524 77904 36576
rect 83004 36567 83056 36576
rect 83004 36533 83013 36567
rect 83013 36533 83047 36567
rect 83047 36533 83056 36567
rect 83004 36524 83056 36533
rect 86960 36660 87012 36712
rect 86776 36592 86828 36644
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 81046 36422 81098 36474
rect 81110 36422 81162 36474
rect 81174 36422 81226 36474
rect 81238 36422 81290 36474
rect 4988 36363 5040 36372
rect 4988 36329 4997 36363
rect 4997 36329 5031 36363
rect 5031 36329 5040 36363
rect 4988 36320 5040 36329
rect 15476 36363 15528 36372
rect 15476 36329 15485 36363
rect 15485 36329 15519 36363
rect 15519 36329 15528 36363
rect 15476 36320 15528 36329
rect 17224 36363 17276 36372
rect 17224 36329 17233 36363
rect 17233 36329 17267 36363
rect 17267 36329 17276 36363
rect 17224 36320 17276 36329
rect 26608 36363 26660 36372
rect 9864 36252 9916 36304
rect 10600 36295 10652 36304
rect 10600 36261 10609 36295
rect 10609 36261 10643 36295
rect 10643 36261 10652 36295
rect 10600 36252 10652 36261
rect 5356 36227 5408 36236
rect 5356 36193 5365 36227
rect 5365 36193 5399 36227
rect 5399 36193 5408 36227
rect 5356 36184 5408 36193
rect 8208 36184 8260 36236
rect 16764 36252 16816 36304
rect 16488 36227 16540 36236
rect 5264 36116 5316 36168
rect 11060 36159 11112 36168
rect 11060 36125 11069 36159
rect 11069 36125 11103 36159
rect 11103 36125 11112 36159
rect 11060 36116 11112 36125
rect 16488 36193 16497 36227
rect 16497 36193 16531 36227
rect 16531 36193 16540 36227
rect 16488 36184 16540 36193
rect 26608 36329 26617 36363
rect 26617 36329 26651 36363
rect 26651 36329 26660 36363
rect 26608 36320 26660 36329
rect 25504 36252 25556 36304
rect 33692 36320 33744 36372
rect 35440 36320 35492 36372
rect 36544 36320 36596 36372
rect 41328 36320 41380 36372
rect 41696 36363 41748 36372
rect 41696 36329 41705 36363
rect 41705 36329 41739 36363
rect 41739 36329 41748 36363
rect 41696 36320 41748 36329
rect 41788 36320 41840 36372
rect 44548 36363 44600 36372
rect 16764 36116 16816 36168
rect 24860 36184 24912 36236
rect 24952 36184 25004 36236
rect 26148 36227 26200 36236
rect 26148 36193 26157 36227
rect 26157 36193 26191 36227
rect 26191 36193 26200 36227
rect 32220 36252 32272 36304
rect 36636 36252 36688 36304
rect 44548 36329 44557 36363
rect 44557 36329 44591 36363
rect 44591 36329 44600 36363
rect 44548 36320 44600 36329
rect 26148 36184 26200 36193
rect 20996 36159 21048 36168
rect 20996 36125 21005 36159
rect 21005 36125 21039 36159
rect 21039 36125 21048 36159
rect 20996 36116 21048 36125
rect 21272 36159 21324 36168
rect 21272 36125 21281 36159
rect 21281 36125 21315 36159
rect 21315 36125 21324 36159
rect 21272 36116 21324 36125
rect 27068 36159 27120 36168
rect 27068 36125 27077 36159
rect 27077 36125 27111 36159
rect 27111 36125 27120 36159
rect 27068 36116 27120 36125
rect 27436 36159 27488 36168
rect 27436 36125 27445 36159
rect 27445 36125 27479 36159
rect 27479 36125 27488 36159
rect 27436 36116 27488 36125
rect 31484 36184 31536 36236
rect 32404 36227 32456 36236
rect 32404 36193 32413 36227
rect 32413 36193 32447 36227
rect 32447 36193 32456 36227
rect 32404 36184 32456 36193
rect 34152 36227 34204 36236
rect 34152 36193 34161 36227
rect 34161 36193 34195 36227
rect 34195 36193 34204 36227
rect 34152 36184 34204 36193
rect 35348 36227 35400 36236
rect 35348 36193 35357 36227
rect 35357 36193 35391 36227
rect 35391 36193 35400 36227
rect 35348 36184 35400 36193
rect 35992 36184 36044 36236
rect 36452 36184 36504 36236
rect 39120 36184 39172 36236
rect 40684 36227 40736 36236
rect 40684 36193 40693 36227
rect 40693 36193 40727 36227
rect 40727 36193 40736 36227
rect 40684 36184 40736 36193
rect 41788 36184 41840 36236
rect 42248 36184 42300 36236
rect 43536 36227 43588 36236
rect 43536 36193 43545 36227
rect 43545 36193 43579 36227
rect 43579 36193 43588 36227
rect 43536 36184 43588 36193
rect 16488 35980 16540 36032
rect 16764 36023 16816 36032
rect 16764 35989 16773 36023
rect 16773 35989 16807 36023
rect 16807 35989 16816 36023
rect 16764 35980 16816 35989
rect 20996 35980 21048 36032
rect 22008 35980 22060 36032
rect 25320 36048 25372 36100
rect 25872 36048 25924 36100
rect 27528 36048 27580 36100
rect 29184 36048 29236 36100
rect 30288 36116 30340 36168
rect 35900 36116 35952 36168
rect 37556 36116 37608 36168
rect 40224 36116 40276 36168
rect 43720 36184 43772 36236
rect 43996 36227 44048 36236
rect 43996 36193 44005 36227
rect 44005 36193 44039 36227
rect 44039 36193 44048 36227
rect 43996 36184 44048 36193
rect 49976 36320 50028 36372
rect 46020 36227 46072 36236
rect 46020 36193 46029 36227
rect 46029 36193 46063 36227
rect 46063 36193 46072 36227
rect 46020 36184 46072 36193
rect 44916 36159 44968 36168
rect 44916 36125 44925 36159
rect 44925 36125 44959 36159
rect 44959 36125 44968 36159
rect 44916 36116 44968 36125
rect 45836 36159 45888 36168
rect 45836 36125 45845 36159
rect 45845 36125 45879 36159
rect 45879 36125 45888 36159
rect 46940 36252 46992 36304
rect 45836 36116 45888 36125
rect 35256 36048 35308 36100
rect 46940 36116 46992 36168
rect 47676 36184 47728 36236
rect 49056 36184 49108 36236
rect 49792 36116 49844 36168
rect 54484 36320 54536 36372
rect 61108 36320 61160 36372
rect 68652 36320 68704 36372
rect 72792 36320 72844 36372
rect 50160 36184 50212 36236
rect 51172 36252 51224 36304
rect 51540 36252 51592 36304
rect 50712 36184 50764 36236
rect 52460 36252 52512 36304
rect 51172 36116 51224 36168
rect 54300 36184 54352 36236
rect 58624 36252 58676 36304
rect 64788 36252 64840 36304
rect 23664 35980 23716 36032
rect 26240 36023 26292 36032
rect 26240 35989 26249 36023
rect 26249 35989 26283 36023
rect 26283 35989 26292 36023
rect 26240 35980 26292 35989
rect 27160 35980 27212 36032
rect 27436 35980 27488 36032
rect 34612 35980 34664 36032
rect 38752 35980 38804 36032
rect 39580 36023 39632 36032
rect 39580 35989 39589 36023
rect 39589 35989 39623 36023
rect 39623 35989 39632 36023
rect 39580 35980 39632 35989
rect 39948 35980 40000 36032
rect 40224 35980 40276 36032
rect 49148 35980 49200 36032
rect 49516 35980 49568 36032
rect 51264 36048 51316 36100
rect 56600 36116 56652 36168
rect 56876 36159 56928 36168
rect 56876 36125 56885 36159
rect 56885 36125 56919 36159
rect 56919 36125 56928 36159
rect 56876 36116 56928 36125
rect 54852 36048 54904 36100
rect 55956 36048 56008 36100
rect 53288 35980 53340 36032
rect 55036 35980 55088 36032
rect 58716 36184 58768 36236
rect 62212 36184 62264 36236
rect 65984 36184 66036 36236
rect 71504 36252 71556 36304
rect 77944 36320 77996 36372
rect 78680 36363 78732 36372
rect 78680 36329 78689 36363
rect 78689 36329 78723 36363
rect 78723 36329 78732 36363
rect 78680 36320 78732 36329
rect 82176 36320 82228 36372
rect 86960 36363 87012 36372
rect 81348 36252 81400 36304
rect 83556 36252 83608 36304
rect 86960 36329 86969 36363
rect 86969 36329 87003 36363
rect 87003 36329 87012 36363
rect 86960 36320 87012 36329
rect 86224 36252 86276 36304
rect 69572 36184 69624 36236
rect 62120 36116 62172 36168
rect 65524 36116 65576 36168
rect 71688 36184 71740 36236
rect 77300 36227 77352 36236
rect 60556 36048 60608 36100
rect 71596 36116 71648 36168
rect 62212 36023 62264 36032
rect 62212 35989 62221 36023
rect 62221 35989 62255 36023
rect 62255 35989 62264 36023
rect 62212 35980 62264 35989
rect 64512 35980 64564 36032
rect 69020 35980 69072 36032
rect 70124 35980 70176 36032
rect 77300 36193 77309 36227
rect 77309 36193 77343 36227
rect 77343 36193 77352 36227
rect 77300 36184 77352 36193
rect 79968 36227 80020 36236
rect 79968 36193 79977 36227
rect 79977 36193 80011 36227
rect 80011 36193 80020 36227
rect 79968 36184 80020 36193
rect 82820 36227 82872 36236
rect 82820 36193 82829 36227
rect 82829 36193 82863 36227
rect 82863 36193 82872 36227
rect 82820 36184 82872 36193
rect 72516 36159 72568 36168
rect 72516 36125 72525 36159
rect 72525 36125 72559 36159
rect 72559 36125 72568 36159
rect 72516 36116 72568 36125
rect 77576 36159 77628 36168
rect 77576 36125 77585 36159
rect 77585 36125 77619 36159
rect 77619 36125 77628 36159
rect 77576 36116 77628 36125
rect 79692 36048 79744 36100
rect 83004 36091 83056 36100
rect 83004 36057 83013 36091
rect 83013 36057 83047 36091
rect 83047 36057 83056 36091
rect 84200 36184 84252 36236
rect 86316 36184 86368 36236
rect 86776 36227 86828 36236
rect 86776 36193 86785 36227
rect 86785 36193 86819 36227
rect 86819 36193 86828 36227
rect 86776 36184 86828 36193
rect 83004 36048 83056 36057
rect 78220 35980 78272 36032
rect 80244 35980 80296 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 65686 35878 65738 35930
rect 65750 35878 65802 35930
rect 65814 35878 65866 35930
rect 65878 35878 65930 35930
rect 96406 35878 96458 35930
rect 96470 35878 96522 35930
rect 96534 35878 96586 35930
rect 96598 35878 96650 35930
rect 4068 35776 4120 35828
rect 6368 35776 6420 35828
rect 26148 35776 26200 35828
rect 21732 35751 21784 35760
rect 21732 35717 21741 35751
rect 21741 35717 21775 35751
rect 21775 35717 21784 35751
rect 21732 35708 21784 35717
rect 22468 35708 22520 35760
rect 30840 35776 30892 35828
rect 30932 35776 30984 35828
rect 31668 35776 31720 35828
rect 32220 35776 32272 35828
rect 32312 35776 32364 35828
rect 35256 35776 35308 35828
rect 35348 35776 35400 35828
rect 38384 35776 38436 35828
rect 38476 35776 38528 35828
rect 40776 35776 40828 35828
rect 40868 35776 40920 35828
rect 5172 35640 5224 35692
rect 5632 35640 5684 35692
rect 14924 35640 14976 35692
rect 20720 35640 20772 35692
rect 3700 35572 3752 35624
rect 6276 35572 6328 35624
rect 10140 35572 10192 35624
rect 4804 35504 4856 35556
rect 10324 35547 10376 35556
rect 10324 35513 10333 35547
rect 10333 35513 10367 35547
rect 10367 35513 10376 35547
rect 10324 35504 10376 35513
rect 4160 35436 4212 35488
rect 6092 35436 6144 35488
rect 10232 35479 10284 35488
rect 10232 35445 10241 35479
rect 10241 35445 10275 35479
rect 10275 35445 10284 35479
rect 10968 35572 11020 35624
rect 13636 35615 13688 35624
rect 11520 35479 11572 35488
rect 10232 35436 10284 35445
rect 11520 35445 11529 35479
rect 11529 35445 11563 35479
rect 11563 35445 11572 35479
rect 11520 35436 11572 35445
rect 13636 35581 13645 35615
rect 13645 35581 13679 35615
rect 13679 35581 13688 35615
rect 13636 35572 13688 35581
rect 14556 35572 14608 35624
rect 20996 35572 21048 35624
rect 15016 35547 15068 35556
rect 15016 35513 15025 35547
rect 15025 35513 15059 35547
rect 15059 35513 15068 35547
rect 15016 35504 15068 35513
rect 13452 35436 13504 35488
rect 22928 35572 22980 35624
rect 25412 35615 25464 35624
rect 25412 35581 25421 35615
rect 25421 35581 25455 35615
rect 25455 35581 25464 35615
rect 25412 35572 25464 35581
rect 27528 35708 27580 35760
rect 31392 35708 31444 35760
rect 30564 35683 30616 35692
rect 21364 35504 21416 35556
rect 27252 35572 27304 35624
rect 28632 35572 28684 35624
rect 29460 35615 29512 35624
rect 29460 35581 29469 35615
rect 29469 35581 29503 35615
rect 29503 35581 29512 35615
rect 29460 35572 29512 35581
rect 30564 35649 30573 35683
rect 30573 35649 30607 35683
rect 30607 35649 30616 35683
rect 30564 35640 30616 35649
rect 30012 35615 30064 35624
rect 30012 35581 30021 35615
rect 30021 35581 30055 35615
rect 30055 35581 30064 35615
rect 30932 35640 30984 35692
rect 30012 35572 30064 35581
rect 31024 35572 31076 35624
rect 31576 35572 31628 35624
rect 32680 35751 32732 35760
rect 32680 35717 32689 35751
rect 32689 35717 32723 35751
rect 32723 35717 32732 35751
rect 32680 35708 32732 35717
rect 32220 35615 32272 35624
rect 32220 35581 32229 35615
rect 32229 35581 32263 35615
rect 32263 35581 32272 35615
rect 41328 35708 41380 35760
rect 41972 35708 42024 35760
rect 48964 35776 49016 35828
rect 49700 35776 49752 35828
rect 50804 35776 50856 35828
rect 52000 35751 52052 35760
rect 52000 35717 52009 35751
rect 52009 35717 52043 35751
rect 52043 35717 52052 35751
rect 52000 35708 52052 35717
rect 53656 35776 53708 35828
rect 54852 35819 54904 35828
rect 54852 35785 54861 35819
rect 54861 35785 54895 35819
rect 54895 35785 54904 35819
rect 54852 35776 54904 35785
rect 55036 35819 55088 35828
rect 55036 35785 55045 35819
rect 55045 35785 55079 35819
rect 55079 35785 55088 35819
rect 55036 35776 55088 35785
rect 55680 35776 55732 35828
rect 58256 35776 58308 35828
rect 35716 35640 35768 35692
rect 35992 35640 36044 35692
rect 32220 35572 32272 35581
rect 33416 35504 33468 35556
rect 33508 35504 33560 35556
rect 35256 35504 35308 35556
rect 38568 35640 38620 35692
rect 39488 35683 39540 35692
rect 39488 35649 39497 35683
rect 39497 35649 39531 35683
rect 39531 35649 39540 35683
rect 39488 35640 39540 35649
rect 22008 35436 22060 35488
rect 26516 35436 26568 35488
rect 28632 35436 28684 35488
rect 29460 35436 29512 35488
rect 30012 35436 30064 35488
rect 31024 35436 31076 35488
rect 31392 35436 31444 35488
rect 38476 35572 38528 35624
rect 40776 35615 40828 35624
rect 39948 35504 40000 35556
rect 37832 35479 37884 35488
rect 37832 35445 37841 35479
rect 37841 35445 37875 35479
rect 37875 35445 37884 35479
rect 37832 35436 37884 35445
rect 38016 35479 38068 35488
rect 38016 35445 38025 35479
rect 38025 35445 38059 35479
rect 38059 35445 38068 35479
rect 38016 35436 38068 35445
rect 38384 35436 38436 35488
rect 38476 35436 38528 35488
rect 40776 35581 40785 35615
rect 40785 35581 40819 35615
rect 40819 35581 40828 35615
rect 40776 35572 40828 35581
rect 43628 35640 43680 35692
rect 49056 35640 49108 35692
rect 41236 35615 41288 35624
rect 41236 35581 41245 35615
rect 41245 35581 41279 35615
rect 41279 35581 41288 35615
rect 41236 35572 41288 35581
rect 42708 35547 42760 35556
rect 42708 35513 42717 35547
rect 42717 35513 42751 35547
rect 42751 35513 42760 35547
rect 42708 35504 42760 35513
rect 48964 35504 49016 35556
rect 49424 35615 49476 35624
rect 49424 35581 49433 35615
rect 49433 35581 49467 35615
rect 49467 35581 49476 35615
rect 49424 35572 49476 35581
rect 49700 35572 49752 35624
rect 53196 35640 53248 35692
rect 51448 35572 51500 35624
rect 53012 35572 53064 35624
rect 53288 35615 53340 35624
rect 53288 35581 53297 35615
rect 53297 35581 53331 35615
rect 53331 35581 53340 35615
rect 53288 35572 53340 35581
rect 43352 35479 43404 35488
rect 43352 35445 43361 35479
rect 43361 35445 43395 35479
rect 43395 35445 43404 35479
rect 43352 35436 43404 35445
rect 49056 35479 49108 35488
rect 49056 35445 49065 35479
rect 49065 35445 49099 35479
rect 49099 35445 49108 35479
rect 49056 35436 49108 35445
rect 49240 35479 49292 35488
rect 49240 35445 49249 35479
rect 49249 35445 49283 35479
rect 49283 35445 49292 35479
rect 49240 35436 49292 35445
rect 49516 35436 49568 35488
rect 50160 35436 50212 35488
rect 50988 35504 51040 35556
rect 55036 35572 55088 35624
rect 55220 35547 55272 35556
rect 55220 35513 55229 35547
rect 55229 35513 55263 35547
rect 55263 35513 55272 35547
rect 55220 35504 55272 35513
rect 55680 35615 55732 35624
rect 55680 35581 55689 35615
rect 55689 35581 55723 35615
rect 55723 35581 55732 35615
rect 55680 35572 55732 35581
rect 55956 35572 56008 35624
rect 56600 35615 56652 35624
rect 56600 35581 56609 35615
rect 56609 35581 56643 35615
rect 56643 35581 56652 35615
rect 56600 35572 56652 35581
rect 59544 35708 59596 35760
rect 60280 35708 60332 35760
rect 62120 35708 62172 35760
rect 62948 35708 63000 35760
rect 63776 35708 63828 35760
rect 68928 35708 68980 35760
rect 70124 35751 70176 35760
rect 70124 35717 70133 35751
rect 70133 35717 70167 35751
rect 70167 35717 70176 35751
rect 70124 35708 70176 35717
rect 71320 35708 71372 35760
rect 74448 35776 74500 35828
rect 77208 35708 77260 35760
rect 58348 35504 58400 35556
rect 62948 35572 63000 35624
rect 66168 35572 66220 35624
rect 68928 35615 68980 35624
rect 68928 35581 68937 35615
rect 68937 35581 68971 35615
rect 68971 35581 68980 35615
rect 68928 35572 68980 35581
rect 69020 35615 69072 35624
rect 69020 35581 69029 35615
rect 69029 35581 69063 35615
rect 69063 35581 69072 35615
rect 69020 35572 69072 35581
rect 70124 35572 70176 35624
rect 70216 35572 70268 35624
rect 70584 35615 70636 35624
rect 70584 35581 70593 35615
rect 70593 35581 70627 35615
rect 70627 35581 70636 35615
rect 70584 35572 70636 35581
rect 70676 35572 70728 35624
rect 72792 35615 72844 35624
rect 69572 35547 69624 35556
rect 69572 35513 69581 35547
rect 69581 35513 69615 35547
rect 69615 35513 69624 35547
rect 69572 35504 69624 35513
rect 72792 35581 72801 35615
rect 72801 35581 72835 35615
rect 72835 35581 72844 35615
rect 72792 35572 72844 35581
rect 77576 35640 77628 35692
rect 77852 35683 77904 35692
rect 77852 35649 77861 35683
rect 77861 35649 77895 35683
rect 77895 35649 77904 35683
rect 77852 35640 77904 35649
rect 80428 35819 80480 35828
rect 80428 35785 80437 35819
rect 80437 35785 80471 35819
rect 80471 35785 80480 35819
rect 80428 35776 80480 35785
rect 82820 35776 82872 35828
rect 78128 35615 78180 35624
rect 78128 35581 78137 35615
rect 78137 35581 78171 35615
rect 78171 35581 78180 35615
rect 78128 35572 78180 35581
rect 83096 35751 83148 35760
rect 83096 35717 83105 35751
rect 83105 35717 83139 35751
rect 83139 35717 83148 35751
rect 83096 35708 83148 35717
rect 79968 35683 80020 35692
rect 79968 35649 79974 35683
rect 79974 35649 80020 35683
rect 79968 35640 80020 35649
rect 80152 35683 80204 35692
rect 80152 35649 80161 35683
rect 80161 35649 80195 35683
rect 80195 35649 80204 35683
rect 80152 35640 80204 35649
rect 82912 35640 82964 35692
rect 84200 35640 84252 35692
rect 79692 35504 79744 35556
rect 82728 35572 82780 35624
rect 83924 35615 83976 35624
rect 83004 35504 83056 35556
rect 83924 35581 83933 35615
rect 83933 35581 83967 35615
rect 83967 35581 83976 35615
rect 83924 35572 83976 35581
rect 84384 35615 84436 35624
rect 84384 35581 84393 35615
rect 84393 35581 84427 35615
rect 84427 35581 84436 35615
rect 86500 35776 86552 35828
rect 86868 35776 86920 35828
rect 84384 35572 84436 35581
rect 86868 35572 86920 35624
rect 88340 35572 88392 35624
rect 53840 35436 53892 35488
rect 63776 35436 63828 35488
rect 65432 35436 65484 35488
rect 69848 35436 69900 35488
rect 70860 35436 70912 35488
rect 77024 35436 77076 35488
rect 80152 35436 80204 35488
rect 82728 35436 82780 35488
rect 83924 35436 83976 35488
rect 85028 35436 85080 35488
rect 88248 35436 88300 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 81046 35334 81098 35386
rect 81110 35334 81162 35386
rect 81174 35334 81226 35386
rect 81238 35334 81290 35386
rect 4712 35275 4764 35284
rect 4712 35241 4721 35275
rect 4721 35241 4755 35275
rect 4755 35241 4764 35275
rect 4712 35232 4764 35241
rect 5356 35096 5408 35148
rect 6276 35139 6328 35148
rect 6276 35105 6285 35139
rect 6285 35105 6319 35139
rect 6319 35105 6328 35139
rect 6276 35096 6328 35105
rect 9772 35164 9824 35216
rect 8300 35096 8352 35148
rect 11060 35164 11112 35216
rect 2872 34960 2924 35012
rect 8208 35028 8260 35080
rect 10324 35096 10376 35148
rect 12348 35232 12400 35284
rect 15016 35096 15068 35148
rect 21364 35232 21416 35284
rect 11520 35028 11572 35080
rect 22468 35164 22520 35216
rect 32772 35232 32824 35284
rect 16396 35139 16448 35148
rect 16396 35105 16405 35139
rect 16405 35105 16439 35139
rect 16439 35105 16448 35139
rect 16396 35096 16448 35105
rect 16488 35028 16540 35080
rect 21732 35096 21784 35148
rect 21824 35096 21876 35148
rect 23664 35139 23716 35148
rect 23664 35105 23673 35139
rect 23673 35105 23707 35139
rect 23707 35105 23716 35139
rect 23664 35096 23716 35105
rect 25136 35096 25188 35148
rect 20720 35028 20772 35080
rect 22008 35028 22060 35080
rect 9128 34960 9180 35012
rect 10968 34960 11020 35012
rect 26240 34960 26292 35012
rect 13912 34935 13964 34944
rect 13912 34901 13921 34935
rect 13921 34901 13955 34935
rect 13955 34901 13964 34935
rect 13912 34892 13964 34901
rect 16580 34935 16632 34944
rect 16580 34901 16589 34935
rect 16589 34901 16623 34935
rect 16623 34901 16632 34935
rect 16580 34892 16632 34901
rect 25872 34892 25924 34944
rect 26700 35139 26752 35148
rect 26700 35105 26709 35139
rect 26709 35105 26743 35139
rect 26743 35105 26752 35139
rect 27896 35164 27948 35216
rect 26700 35096 26752 35105
rect 28172 35096 28224 35148
rect 28908 35139 28960 35148
rect 28908 35105 28917 35139
rect 28917 35105 28951 35139
rect 28951 35105 28960 35139
rect 30380 35139 30432 35148
rect 28908 35096 28960 35105
rect 30380 35105 30389 35139
rect 30389 35105 30423 35139
rect 30423 35105 30432 35139
rect 30380 35096 30432 35105
rect 41236 35232 41288 35284
rect 41328 35232 41380 35284
rect 61292 35232 61344 35284
rect 39120 35164 39172 35216
rect 27804 35071 27856 35080
rect 27804 35037 27813 35071
rect 27813 35037 27847 35071
rect 27847 35037 27856 35071
rect 27804 35028 27856 35037
rect 33232 35096 33284 35148
rect 33416 35139 33468 35148
rect 33416 35105 33425 35139
rect 33425 35105 33459 35139
rect 33459 35105 33468 35139
rect 33416 35096 33468 35105
rect 39396 35139 39448 35148
rect 38108 35028 38160 35080
rect 38476 35071 38528 35080
rect 38476 35037 38485 35071
rect 38485 35037 38519 35071
rect 38519 35037 38528 35071
rect 38476 35028 38528 35037
rect 35624 34960 35676 35012
rect 38568 34960 38620 35012
rect 39396 35105 39405 35139
rect 39405 35105 39439 35139
rect 39439 35105 39448 35139
rect 39396 35096 39448 35105
rect 39764 35071 39816 35080
rect 39764 35037 39773 35071
rect 39773 35037 39807 35071
rect 39807 35037 39816 35071
rect 39764 35028 39816 35037
rect 40224 35028 40276 35080
rect 40960 35028 41012 35080
rect 40868 34960 40920 35012
rect 41512 35164 41564 35216
rect 41972 35207 42024 35216
rect 41236 35096 41288 35148
rect 41420 35139 41472 35148
rect 41420 35105 41429 35139
rect 41429 35105 41463 35139
rect 41463 35105 41472 35139
rect 41972 35173 41981 35207
rect 41981 35173 42015 35207
rect 42015 35173 42024 35207
rect 41972 35164 42024 35173
rect 43720 35164 43772 35216
rect 42248 35139 42300 35148
rect 41420 35096 41472 35105
rect 42248 35105 42257 35139
rect 42257 35105 42291 35139
rect 42291 35105 42300 35139
rect 42248 35096 42300 35105
rect 49884 35139 49936 35148
rect 49884 35105 49893 35139
rect 49893 35105 49927 35139
rect 49927 35105 49936 35139
rect 49884 35096 49936 35105
rect 52000 35164 52052 35216
rect 53196 35207 53248 35216
rect 53196 35173 53205 35207
rect 53205 35173 53239 35207
rect 53239 35173 53248 35207
rect 53196 35164 53248 35173
rect 50436 35139 50488 35148
rect 50436 35105 50445 35139
rect 50445 35105 50479 35139
rect 50479 35105 50488 35139
rect 50436 35096 50488 35105
rect 51172 35096 51224 35148
rect 51816 35096 51868 35148
rect 52092 35139 52144 35148
rect 52092 35105 52101 35139
rect 52101 35105 52135 35139
rect 52135 35105 52144 35139
rect 52092 35096 52144 35105
rect 42524 35028 42576 35080
rect 49424 35028 49476 35080
rect 49700 35071 49752 35080
rect 49700 35037 49709 35071
rect 49709 35037 49743 35071
rect 49743 35037 49752 35071
rect 49700 35028 49752 35037
rect 51724 35028 51776 35080
rect 52644 35139 52696 35148
rect 52644 35105 52653 35139
rect 52653 35105 52687 35139
rect 52687 35105 52696 35139
rect 56140 35164 56192 35216
rect 57060 35164 57112 35216
rect 58348 35164 58400 35216
rect 58808 35164 58860 35216
rect 70584 35232 70636 35284
rect 70860 35232 70912 35284
rect 63040 35164 63092 35216
rect 82820 35232 82872 35284
rect 83004 35275 83056 35284
rect 83004 35241 83013 35275
rect 83013 35241 83047 35275
rect 83047 35241 83056 35275
rect 83004 35232 83056 35241
rect 83096 35232 83148 35284
rect 83280 35232 83332 35284
rect 86500 35275 86552 35284
rect 72516 35164 72568 35216
rect 52644 35096 52696 35105
rect 58716 35139 58768 35148
rect 43352 34960 43404 35012
rect 51448 34960 51500 35012
rect 38108 34935 38160 34944
rect 38108 34901 38117 34935
rect 38117 34901 38151 34935
rect 38151 34901 38160 34935
rect 38108 34892 38160 34901
rect 38292 34935 38344 34944
rect 38292 34901 38301 34935
rect 38301 34901 38335 34935
rect 38335 34901 38344 34935
rect 38292 34892 38344 34901
rect 39396 34892 39448 34944
rect 40408 34892 40460 34944
rect 48872 34892 48924 34944
rect 49332 34935 49384 34944
rect 49332 34901 49341 34935
rect 49341 34901 49375 34935
rect 49375 34901 49384 34935
rect 49332 34892 49384 34901
rect 49516 34892 49568 34944
rect 49700 34892 49752 34944
rect 49884 34892 49936 34944
rect 51172 34892 51224 34944
rect 51264 34935 51316 34944
rect 51264 34901 51273 34935
rect 51273 34901 51307 34935
rect 51307 34901 51316 34935
rect 51540 34935 51592 34944
rect 51264 34892 51316 34901
rect 51540 34901 51549 34935
rect 51549 34901 51583 34935
rect 51583 34901 51592 34935
rect 51724 34935 51776 34944
rect 51540 34892 51592 34901
rect 51724 34901 51733 34935
rect 51733 34901 51767 34935
rect 51767 34901 51776 34935
rect 51724 34892 51776 34901
rect 51816 34892 51868 34944
rect 55956 35028 56008 35080
rect 56048 35071 56100 35080
rect 56048 35037 56057 35071
rect 56057 35037 56091 35071
rect 56091 35037 56100 35071
rect 56324 35071 56376 35080
rect 56048 35028 56100 35037
rect 56324 35037 56333 35071
rect 56333 35037 56367 35071
rect 56367 35037 56376 35071
rect 56324 35028 56376 35037
rect 56416 35028 56468 35080
rect 58440 35028 58492 35080
rect 58716 35105 58725 35139
rect 58725 35105 58759 35139
rect 58759 35105 58768 35139
rect 58716 35096 58768 35105
rect 62028 35139 62080 35148
rect 62028 35105 62037 35139
rect 62037 35105 62071 35139
rect 62071 35105 62080 35139
rect 62028 35096 62080 35105
rect 64512 35139 64564 35148
rect 64512 35105 64521 35139
rect 64521 35105 64555 35139
rect 64555 35105 64564 35139
rect 64512 35096 64564 35105
rect 66720 35096 66772 35148
rect 69296 35139 69348 35148
rect 69296 35105 69305 35139
rect 69305 35105 69339 35139
rect 69339 35105 69348 35139
rect 69296 35096 69348 35105
rect 69848 35096 69900 35148
rect 70032 35096 70084 35148
rect 71412 35096 71464 35148
rect 71688 35096 71740 35148
rect 53472 35003 53524 35012
rect 53472 34969 53481 35003
rect 53481 34969 53515 35003
rect 53515 34969 53524 35003
rect 59636 35028 59688 35080
rect 62304 35071 62356 35080
rect 62304 35037 62313 35071
rect 62313 35037 62347 35071
rect 62347 35037 62356 35071
rect 62304 35028 62356 35037
rect 53472 34960 53524 34969
rect 55588 34935 55640 34944
rect 55588 34901 55597 34935
rect 55597 34901 55631 34935
rect 55631 34901 55640 34935
rect 55588 34892 55640 34901
rect 57428 34935 57480 34944
rect 57428 34901 57437 34935
rect 57437 34901 57471 34935
rect 57471 34901 57480 34935
rect 57428 34892 57480 34901
rect 62028 34960 62080 35012
rect 58808 34935 58860 34944
rect 58808 34901 58817 34935
rect 58817 34901 58851 34935
rect 58851 34901 58860 34935
rect 58808 34892 58860 34901
rect 58900 34892 58952 34944
rect 59084 34892 59136 34944
rect 59728 34892 59780 34944
rect 61292 34892 61344 34944
rect 69112 34960 69164 35012
rect 64604 34935 64656 34944
rect 64604 34901 64613 34935
rect 64613 34901 64647 34935
rect 64647 34901 64656 34935
rect 64604 34892 64656 34901
rect 64696 34892 64748 34944
rect 66260 34892 66312 34944
rect 71596 35028 71648 35080
rect 72240 35096 72292 35148
rect 80060 35164 80112 35216
rect 80244 35207 80296 35216
rect 80244 35173 80253 35207
rect 80253 35173 80287 35207
rect 80287 35173 80296 35207
rect 80244 35164 80296 35173
rect 84384 35164 84436 35216
rect 84936 35207 84988 35216
rect 84936 35173 84945 35207
rect 84945 35173 84979 35207
rect 84979 35173 84988 35207
rect 84936 35164 84988 35173
rect 86500 35241 86509 35275
rect 86509 35241 86543 35275
rect 86543 35241 86552 35275
rect 86500 35232 86552 35241
rect 77024 35139 77076 35148
rect 72148 35028 72200 35080
rect 77024 35105 77033 35139
rect 77033 35105 77067 35139
rect 77067 35105 77076 35139
rect 77024 35096 77076 35105
rect 78588 35139 78640 35148
rect 78588 35105 78597 35139
rect 78597 35105 78631 35139
rect 78631 35105 78640 35139
rect 78588 35096 78640 35105
rect 78956 35096 79008 35148
rect 80152 35139 80204 35148
rect 80152 35105 80161 35139
rect 80161 35105 80195 35139
rect 80195 35105 80204 35139
rect 80152 35096 80204 35105
rect 77760 35028 77812 35080
rect 83096 35096 83148 35148
rect 84752 35139 84804 35148
rect 84752 35105 84761 35139
rect 84761 35105 84795 35139
rect 84795 35105 84804 35139
rect 84752 35096 84804 35105
rect 85028 35139 85080 35148
rect 85028 35105 85037 35139
rect 85037 35105 85071 35139
rect 85071 35105 85080 35139
rect 85028 35096 85080 35105
rect 82176 35028 82228 35080
rect 86868 35096 86920 35148
rect 87328 35096 87380 35148
rect 88248 35139 88300 35148
rect 88248 35105 88257 35139
rect 88257 35105 88291 35139
rect 88291 35105 88300 35139
rect 88248 35096 88300 35105
rect 85488 35071 85540 35080
rect 85488 35037 85497 35071
rect 85497 35037 85531 35071
rect 85531 35037 85540 35071
rect 85488 35028 85540 35037
rect 87236 35028 87288 35080
rect 78680 34960 78732 35012
rect 84200 34960 84252 35012
rect 88248 34960 88300 35012
rect 71596 34892 71648 34944
rect 71872 34892 71924 34944
rect 76012 34935 76064 34944
rect 76012 34901 76021 34935
rect 76021 34901 76055 34935
rect 76055 34901 76064 34935
rect 76012 34892 76064 34901
rect 77208 34935 77260 34944
rect 77208 34901 77217 34935
rect 77217 34901 77251 34935
rect 77251 34901 77260 34935
rect 77208 34892 77260 34901
rect 80520 34935 80572 34944
rect 80520 34901 80529 34935
rect 80529 34901 80563 34935
rect 80563 34901 80572 34935
rect 80520 34892 80572 34901
rect 83280 34892 83332 34944
rect 85948 34935 86000 34944
rect 85948 34901 85957 34935
rect 85957 34901 85991 34935
rect 85991 34901 86000 34935
rect 85948 34892 86000 34901
rect 86132 34935 86184 34944
rect 86132 34901 86141 34935
rect 86141 34901 86175 34935
rect 86175 34901 86184 34935
rect 86132 34892 86184 34901
rect 86684 34935 86736 34944
rect 86684 34901 86693 34935
rect 86693 34901 86727 34935
rect 86727 34901 86736 34935
rect 86684 34892 86736 34901
rect 87512 34892 87564 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 65686 34790 65738 34842
rect 65750 34790 65802 34842
rect 65814 34790 65866 34842
rect 65878 34790 65930 34842
rect 96406 34790 96458 34842
rect 96470 34790 96522 34842
rect 96534 34790 96586 34842
rect 96598 34790 96650 34842
rect 4988 34552 5040 34604
rect 5632 34595 5684 34604
rect 5632 34561 5641 34595
rect 5641 34561 5675 34595
rect 5675 34561 5684 34595
rect 5632 34552 5684 34561
rect 3700 34484 3752 34536
rect 4804 34484 4856 34536
rect 5356 34527 5408 34536
rect 5356 34493 5365 34527
rect 5365 34493 5399 34527
rect 5399 34493 5408 34527
rect 5356 34484 5408 34493
rect 10416 34620 10468 34672
rect 10600 34620 10652 34672
rect 25136 34688 25188 34740
rect 25504 34731 25556 34740
rect 25504 34697 25513 34731
rect 25513 34697 25547 34731
rect 25547 34697 25556 34731
rect 25504 34688 25556 34697
rect 25872 34688 25924 34740
rect 9864 34552 9916 34604
rect 9404 34484 9456 34536
rect 15752 34620 15804 34672
rect 11152 34484 11204 34536
rect 26424 34620 26476 34672
rect 26976 34620 27028 34672
rect 30380 34688 30432 34740
rect 30748 34688 30800 34740
rect 37832 34731 37884 34740
rect 37832 34697 37841 34731
rect 37841 34697 37875 34731
rect 37875 34697 37884 34731
rect 37832 34688 37884 34697
rect 38568 34688 38620 34740
rect 39304 34688 39356 34740
rect 42708 34688 42760 34740
rect 43628 34731 43680 34740
rect 43628 34697 43637 34731
rect 43637 34697 43671 34731
rect 43671 34697 43680 34731
rect 43628 34688 43680 34697
rect 46756 34688 46808 34740
rect 48412 34731 48464 34740
rect 48412 34697 48421 34731
rect 48421 34697 48455 34731
rect 48455 34697 48464 34731
rect 48412 34688 48464 34697
rect 48872 34688 48924 34740
rect 13452 34484 13504 34536
rect 14280 34527 14332 34536
rect 14280 34493 14289 34527
rect 14289 34493 14323 34527
rect 14323 34493 14332 34527
rect 14280 34484 14332 34493
rect 19984 34527 20036 34536
rect 19984 34493 19993 34527
rect 19993 34493 20027 34527
rect 20027 34493 20036 34527
rect 19984 34484 20036 34493
rect 20628 34527 20680 34536
rect 20628 34493 20637 34527
rect 20637 34493 20671 34527
rect 20671 34493 20680 34527
rect 20628 34484 20680 34493
rect 21364 34484 21416 34536
rect 21732 34484 21784 34536
rect 21272 34459 21324 34468
rect 3976 34391 4028 34400
rect 3976 34357 3985 34391
rect 3985 34357 4019 34391
rect 4019 34357 4028 34391
rect 3976 34348 4028 34357
rect 21272 34425 21281 34459
rect 21281 34425 21315 34459
rect 21315 34425 21324 34459
rect 21272 34416 21324 34425
rect 14556 34348 14608 34400
rect 19340 34348 19392 34400
rect 20260 34348 20312 34400
rect 21824 34348 21876 34400
rect 24676 34348 24728 34400
rect 25872 34527 25924 34536
rect 25872 34493 25881 34527
rect 25881 34493 25915 34527
rect 25915 34493 25924 34527
rect 25872 34484 25924 34493
rect 27344 34552 27396 34604
rect 30748 34552 30800 34604
rect 30840 34552 30892 34604
rect 26424 34484 26476 34536
rect 28908 34416 28960 34468
rect 26792 34391 26844 34400
rect 26792 34357 26801 34391
rect 26801 34357 26835 34391
rect 26835 34357 26844 34391
rect 26792 34348 26844 34357
rect 29184 34484 29236 34536
rect 29552 34527 29604 34536
rect 29552 34493 29561 34527
rect 29561 34493 29595 34527
rect 29595 34493 29604 34527
rect 29552 34484 29604 34493
rect 34152 34484 34204 34536
rect 38384 34620 38436 34672
rect 40408 34620 40460 34672
rect 39396 34552 39448 34604
rect 49792 34620 49844 34672
rect 50252 34731 50304 34740
rect 50252 34697 50261 34731
rect 50261 34697 50295 34731
rect 50295 34697 50304 34731
rect 50252 34688 50304 34697
rect 52092 34688 52144 34740
rect 53196 34688 53248 34740
rect 46664 34595 46716 34604
rect 38568 34484 38620 34536
rect 39948 34484 40000 34536
rect 42064 34527 42116 34536
rect 42064 34493 42073 34527
rect 42073 34493 42107 34527
rect 42107 34493 42116 34527
rect 42064 34484 42116 34493
rect 46664 34561 46673 34595
rect 46673 34561 46707 34595
rect 46707 34561 46716 34595
rect 46664 34552 46716 34561
rect 30288 34416 30340 34468
rect 48964 34552 49016 34604
rect 56324 34688 56376 34740
rect 57428 34688 57480 34740
rect 62028 34688 62080 34740
rect 71412 34731 71464 34740
rect 61936 34663 61988 34672
rect 53840 34595 53892 34604
rect 53840 34561 53849 34595
rect 53849 34561 53883 34595
rect 53883 34561 53892 34595
rect 53840 34552 53892 34561
rect 56784 34595 56836 34604
rect 56784 34561 56793 34595
rect 56793 34561 56827 34595
rect 56827 34561 56836 34595
rect 56784 34552 56836 34561
rect 58624 34595 58676 34604
rect 30380 34348 30432 34400
rect 37832 34348 37884 34400
rect 38568 34348 38620 34400
rect 48872 34527 48924 34536
rect 48872 34493 48881 34527
rect 48881 34493 48915 34527
rect 48915 34493 48924 34527
rect 48872 34484 48924 34493
rect 49424 34527 49476 34536
rect 49424 34493 49433 34527
rect 49433 34493 49467 34527
rect 49467 34493 49476 34527
rect 49424 34484 49476 34493
rect 50620 34484 50672 34536
rect 48320 34348 48372 34400
rect 48504 34391 48556 34400
rect 48504 34357 48513 34391
rect 48513 34357 48547 34391
rect 48547 34357 48556 34391
rect 48504 34348 48556 34357
rect 48596 34348 48648 34400
rect 55312 34484 55364 34536
rect 56140 34484 56192 34536
rect 56600 34527 56652 34536
rect 53932 34348 53984 34400
rect 55588 34416 55640 34468
rect 55128 34391 55180 34400
rect 55128 34357 55137 34391
rect 55137 34357 55171 34391
rect 55171 34357 55180 34391
rect 55128 34348 55180 34357
rect 56600 34493 56609 34527
rect 56609 34493 56643 34527
rect 56643 34493 56652 34527
rect 58624 34561 58633 34595
rect 58633 34561 58667 34595
rect 58667 34561 58676 34595
rect 58624 34552 58676 34561
rect 59452 34552 59504 34604
rect 61936 34629 61945 34663
rect 61945 34629 61979 34663
rect 61979 34629 61988 34663
rect 61936 34620 61988 34629
rect 62580 34620 62632 34672
rect 64328 34663 64380 34672
rect 64328 34629 64337 34663
rect 64337 34629 64371 34663
rect 64371 34629 64380 34663
rect 64328 34620 64380 34629
rect 69940 34663 69992 34672
rect 69940 34629 69949 34663
rect 69949 34629 69983 34663
rect 69983 34629 69992 34663
rect 69940 34620 69992 34629
rect 71412 34697 71421 34731
rect 71421 34697 71455 34731
rect 71455 34697 71464 34731
rect 71412 34688 71464 34697
rect 72608 34731 72660 34740
rect 72240 34620 72292 34672
rect 72148 34552 72200 34604
rect 56600 34484 56652 34493
rect 58256 34527 58308 34536
rect 58256 34493 58265 34527
rect 58265 34493 58299 34527
rect 58299 34493 58308 34527
rect 58992 34527 59044 34536
rect 58256 34484 58308 34493
rect 58992 34493 59001 34527
rect 59001 34493 59035 34527
rect 59035 34493 59044 34527
rect 58992 34484 59044 34493
rect 59176 34527 59228 34536
rect 59176 34493 59185 34527
rect 59185 34493 59219 34527
rect 59219 34493 59228 34527
rect 59176 34484 59228 34493
rect 59360 34527 59412 34536
rect 59360 34493 59369 34527
rect 59369 34493 59403 34527
rect 59403 34493 59412 34527
rect 59360 34484 59412 34493
rect 59636 34484 59688 34536
rect 61752 34484 61804 34536
rect 62948 34527 63000 34536
rect 59544 34391 59596 34400
rect 59544 34357 59553 34391
rect 59553 34357 59587 34391
rect 59587 34357 59596 34391
rect 59544 34348 59596 34357
rect 59636 34348 59688 34400
rect 62948 34493 62957 34527
rect 62957 34493 62991 34527
rect 62991 34493 63000 34527
rect 62948 34484 63000 34493
rect 62672 34459 62724 34468
rect 62672 34425 62681 34459
rect 62681 34425 62715 34459
rect 62715 34425 62724 34459
rect 62672 34416 62724 34425
rect 64328 34484 64380 34536
rect 69940 34484 69992 34536
rect 70124 34484 70176 34536
rect 72608 34697 72617 34731
rect 72617 34697 72651 34731
rect 72651 34697 72660 34731
rect 72608 34688 72660 34697
rect 77300 34688 77352 34740
rect 77760 34731 77812 34740
rect 77760 34697 77769 34731
rect 77769 34697 77803 34731
rect 77803 34697 77812 34731
rect 77760 34688 77812 34697
rect 79968 34688 80020 34740
rect 83924 34688 83976 34740
rect 85764 34688 85816 34740
rect 86776 34688 86828 34740
rect 86868 34688 86920 34740
rect 88340 34731 88392 34740
rect 88340 34697 88349 34731
rect 88349 34697 88383 34731
rect 88383 34697 88392 34731
rect 88340 34688 88392 34697
rect 87052 34620 87104 34672
rect 80520 34552 80572 34604
rect 78956 34484 79008 34536
rect 81348 34484 81400 34536
rect 82176 34527 82228 34536
rect 82176 34493 82185 34527
rect 82185 34493 82219 34527
rect 82219 34493 82228 34527
rect 82176 34484 82228 34493
rect 83280 34484 83332 34536
rect 85488 34552 85540 34604
rect 87420 34552 87472 34604
rect 85764 34527 85816 34536
rect 85764 34493 85773 34527
rect 85773 34493 85807 34527
rect 85807 34493 85816 34527
rect 85764 34484 85816 34493
rect 86960 34484 87012 34536
rect 87880 34527 87932 34536
rect 87880 34493 87889 34527
rect 87889 34493 87923 34527
rect 87923 34493 87932 34527
rect 87880 34484 87932 34493
rect 88248 34527 88300 34536
rect 88248 34493 88257 34527
rect 88257 34493 88291 34527
rect 88291 34493 88300 34527
rect 88248 34484 88300 34493
rect 78588 34348 78640 34400
rect 84936 34348 84988 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 81046 34246 81098 34298
rect 81110 34246 81162 34298
rect 81174 34246 81226 34298
rect 81238 34246 81290 34298
rect 4068 34144 4120 34196
rect 13544 34144 13596 34196
rect 5356 34076 5408 34128
rect 14280 34119 14332 34128
rect 5448 34008 5500 34060
rect 3700 33940 3752 33992
rect 5448 33872 5500 33924
rect 9036 33940 9088 33992
rect 10232 33983 10284 33992
rect 10232 33949 10241 33983
rect 10241 33949 10275 33983
rect 10275 33949 10284 33983
rect 10232 33940 10284 33949
rect 9496 33847 9548 33856
rect 9496 33813 9505 33847
rect 9505 33813 9539 33847
rect 9539 33813 9548 33847
rect 10600 34008 10652 34060
rect 13176 34051 13228 34060
rect 13176 34017 13185 34051
rect 13185 34017 13219 34051
rect 13219 34017 13228 34051
rect 13176 34008 13228 34017
rect 14280 34085 14289 34119
rect 14289 34085 14323 34119
rect 14323 34085 14332 34119
rect 14280 34076 14332 34085
rect 12808 33940 12860 33992
rect 15752 34144 15804 34196
rect 18880 34008 18932 34060
rect 18696 33940 18748 33992
rect 19708 34008 19760 34060
rect 20168 34008 20220 34060
rect 20628 33940 20680 33992
rect 21548 34008 21600 34060
rect 21824 34144 21876 34196
rect 30288 34144 30340 34196
rect 28172 34119 28224 34128
rect 28172 34085 28181 34119
rect 28181 34085 28215 34119
rect 28215 34085 28224 34119
rect 28172 34076 28224 34085
rect 28356 34076 28408 34128
rect 51540 34144 51592 34196
rect 62672 34144 62724 34196
rect 26792 34051 26844 34060
rect 26516 33983 26568 33992
rect 26516 33949 26525 33983
rect 26525 33949 26559 33983
rect 26559 33949 26568 33983
rect 26516 33940 26568 33949
rect 26792 34017 26801 34051
rect 26801 34017 26835 34051
rect 26835 34017 26844 34051
rect 26792 34008 26844 34017
rect 27988 34008 28040 34060
rect 42064 34076 42116 34128
rect 70032 34008 70084 34060
rect 12808 33847 12860 33856
rect 9496 33804 9548 33813
rect 12808 33813 12817 33847
rect 12817 33813 12851 33847
rect 12851 33813 12860 33847
rect 12808 33804 12860 33813
rect 20168 33847 20220 33856
rect 20168 33813 20177 33847
rect 20177 33813 20211 33847
rect 20211 33813 20220 33847
rect 20168 33804 20220 33813
rect 20628 33847 20680 33856
rect 20628 33813 20637 33847
rect 20637 33813 20671 33847
rect 20671 33813 20680 33847
rect 20628 33804 20680 33813
rect 28264 33847 28316 33856
rect 28264 33813 28273 33847
rect 28273 33813 28307 33847
rect 28307 33813 28316 33847
rect 28264 33804 28316 33813
rect 29184 33804 29236 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 5356 33600 5408 33652
rect 13636 33643 13688 33652
rect 13636 33609 13645 33643
rect 13645 33609 13679 33643
rect 13679 33609 13688 33643
rect 13636 33600 13688 33609
rect 14556 33643 14608 33652
rect 14556 33609 14565 33643
rect 14565 33609 14599 33643
rect 14599 33609 14608 33643
rect 14556 33600 14608 33609
rect 18696 33600 18748 33652
rect 19340 33643 19392 33652
rect 19340 33609 19349 33643
rect 19349 33609 19383 33643
rect 19383 33609 19392 33643
rect 19340 33600 19392 33609
rect 20168 33600 20220 33652
rect 4712 33464 4764 33516
rect 9036 33507 9088 33516
rect 9036 33473 9045 33507
rect 9045 33473 9079 33507
rect 9079 33473 9088 33507
rect 9036 33464 9088 33473
rect 4344 33396 4396 33448
rect 8208 33439 8260 33448
rect 8208 33405 8217 33439
rect 8217 33405 8251 33439
rect 8251 33405 8260 33439
rect 8208 33396 8260 33405
rect 12532 33396 12584 33448
rect 4160 33303 4212 33312
rect 4160 33269 4169 33303
rect 4169 33269 4203 33303
rect 4203 33269 4212 33303
rect 4160 33260 4212 33269
rect 10876 33328 10928 33380
rect 4620 33260 4672 33312
rect 4896 33260 4948 33312
rect 8300 33260 8352 33312
rect 10968 33260 11020 33312
rect 12808 33396 12860 33448
rect 13912 33396 13964 33448
rect 14556 33396 14608 33448
rect 19340 33396 19392 33448
rect 14740 33328 14792 33380
rect 20076 33396 20128 33448
rect 26056 33600 26108 33652
rect 26700 33600 26752 33652
rect 27252 33600 27304 33652
rect 28264 33600 28316 33652
rect 61936 33600 61988 33652
rect 62212 33532 62264 33584
rect 24400 33396 24452 33448
rect 25044 33464 25096 33516
rect 25964 33507 26016 33516
rect 25964 33473 25973 33507
rect 25973 33473 26007 33507
rect 26007 33473 26016 33507
rect 25964 33464 26016 33473
rect 26056 33464 26108 33516
rect 64604 33464 64656 33516
rect 25228 33396 25280 33448
rect 14832 33303 14884 33312
rect 14832 33269 14841 33303
rect 14841 33269 14875 33303
rect 14875 33269 14884 33303
rect 14832 33260 14884 33269
rect 19340 33260 19392 33312
rect 20628 33328 20680 33380
rect 25872 33396 25924 33448
rect 23572 33260 23624 33312
rect 26056 33328 26108 33380
rect 69296 33328 69348 33380
rect 25044 33260 25096 33312
rect 25780 33260 25832 33312
rect 76012 33260 76064 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 3240 33056 3292 33108
rect 14004 33056 14056 33108
rect 16672 33056 16724 33108
rect 25780 33099 25832 33108
rect 25780 33065 25789 33099
rect 25789 33065 25823 33099
rect 25823 33065 25832 33099
rect 25780 33056 25832 33065
rect 25964 33056 26016 33108
rect 34612 33056 34664 33108
rect 4344 32963 4396 32972
rect 4344 32929 4353 32963
rect 4353 32929 4387 32963
rect 4387 32929 4396 32963
rect 4344 32920 4396 32929
rect 9404 32988 9456 33040
rect 8208 32963 8260 32972
rect 8208 32929 8217 32963
rect 8217 32929 8251 32963
rect 8251 32929 8260 32963
rect 8208 32920 8260 32929
rect 12900 32988 12952 33040
rect 13360 32988 13412 33040
rect 17224 32988 17276 33040
rect 55128 32988 55180 33040
rect 5356 32852 5408 32904
rect 6000 32895 6052 32904
rect 4896 32716 4948 32768
rect 6000 32861 6009 32895
rect 6009 32861 6043 32895
rect 6043 32861 6052 32895
rect 6000 32852 6052 32861
rect 8944 32852 8996 32904
rect 7380 32716 7432 32768
rect 12348 32784 12400 32836
rect 18052 32852 18104 32904
rect 18696 32920 18748 32972
rect 19248 32963 19300 32972
rect 19248 32929 19257 32963
rect 19257 32929 19291 32963
rect 19291 32929 19300 32963
rect 19248 32920 19300 32929
rect 19432 32920 19484 32972
rect 21364 32963 21416 32972
rect 18604 32852 18656 32904
rect 20168 32852 20220 32904
rect 21364 32929 21373 32963
rect 21373 32929 21407 32963
rect 21407 32929 21416 32963
rect 21364 32920 21416 32929
rect 21548 32963 21600 32972
rect 21548 32929 21557 32963
rect 21557 32929 21591 32963
rect 21591 32929 21600 32963
rect 21548 32920 21600 32929
rect 22008 32963 22060 32972
rect 22008 32929 22017 32963
rect 22017 32929 22051 32963
rect 22051 32929 22060 32963
rect 22008 32920 22060 32929
rect 24400 32963 24452 32972
rect 24400 32929 24409 32963
rect 24409 32929 24443 32963
rect 24443 32929 24452 32963
rect 24400 32920 24452 32929
rect 24492 32920 24544 32972
rect 26056 32963 26108 32972
rect 26056 32929 26065 32963
rect 26065 32929 26099 32963
rect 26099 32929 26108 32963
rect 26056 32920 26108 32929
rect 27160 32920 27212 32972
rect 38292 32920 38344 32972
rect 84016 32920 84068 32972
rect 86684 32920 86736 32972
rect 23848 32852 23900 32904
rect 24216 32895 24268 32904
rect 24216 32861 24225 32895
rect 24225 32861 24259 32895
rect 24259 32861 24268 32895
rect 24216 32852 24268 32861
rect 26332 32852 26384 32904
rect 28816 32852 28868 32904
rect 49332 32852 49384 32904
rect 56600 32784 56652 32836
rect 7748 32716 7800 32768
rect 8668 32716 8720 32768
rect 10048 32716 10100 32768
rect 12532 32716 12584 32768
rect 13912 32759 13964 32768
rect 13912 32725 13921 32759
rect 13921 32725 13955 32759
rect 13955 32725 13964 32759
rect 13912 32716 13964 32725
rect 18052 32716 18104 32768
rect 19248 32716 19300 32768
rect 20352 32716 20404 32768
rect 24216 32716 24268 32768
rect 27804 32716 27856 32768
rect 28264 32716 28316 32768
rect 49240 32716 49292 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 32772 32580 32824 32632
rect 49056 32580 49108 32632
rect 4804 32512 4856 32564
rect 5632 32376 5684 32428
rect 7932 32512 7984 32564
rect 8208 32555 8260 32564
rect 8208 32521 8217 32555
rect 8217 32521 8251 32555
rect 8251 32521 8260 32555
rect 8208 32512 8260 32521
rect 8760 32512 8812 32564
rect 17224 32512 17276 32564
rect 20076 32512 20128 32564
rect 22744 32512 22796 32564
rect 26976 32512 27028 32564
rect 27068 32512 27120 32564
rect 55220 32512 55272 32564
rect 10048 32444 10100 32496
rect 14740 32444 14792 32496
rect 18420 32444 18472 32496
rect 18972 32444 19024 32496
rect 19432 32444 19484 32496
rect 5816 32240 5868 32292
rect 6276 32240 6328 32292
rect 6552 32240 6604 32292
rect 8116 32376 8168 32428
rect 8024 32308 8076 32360
rect 7932 32240 7984 32292
rect 3976 32215 4028 32224
rect 3976 32181 3985 32215
rect 3985 32181 4019 32215
rect 4019 32181 4028 32215
rect 3976 32172 4028 32181
rect 4988 32172 5040 32224
rect 8208 32172 8260 32224
rect 8668 32172 8720 32224
rect 12992 32240 13044 32292
rect 12072 32172 12124 32224
rect 12808 32172 12860 32224
rect 13544 32308 13596 32360
rect 23756 32376 23808 32428
rect 23940 32376 23992 32428
rect 24492 32376 24544 32428
rect 15200 32308 15252 32360
rect 18604 32308 18656 32360
rect 13728 32240 13780 32292
rect 19432 32351 19484 32360
rect 19432 32317 19441 32351
rect 19441 32317 19475 32351
rect 19475 32317 19484 32351
rect 19432 32308 19484 32317
rect 19708 32351 19760 32360
rect 19708 32317 19717 32351
rect 19717 32317 19751 32351
rect 19751 32317 19760 32351
rect 19708 32308 19760 32317
rect 21732 32308 21784 32360
rect 46112 32444 46164 32496
rect 55128 32444 55180 32496
rect 24860 32376 24912 32428
rect 69020 32376 69072 32428
rect 24768 32351 24820 32360
rect 24768 32317 24777 32351
rect 24777 32317 24811 32351
rect 24811 32317 24820 32351
rect 24768 32308 24820 32317
rect 25228 32308 25280 32360
rect 25596 32308 25648 32360
rect 26976 32308 27028 32360
rect 38016 32308 38068 32360
rect 14832 32172 14884 32224
rect 18788 32172 18840 32224
rect 19524 32240 19576 32292
rect 40040 32240 40092 32292
rect 20996 32215 21048 32224
rect 20996 32181 21005 32215
rect 21005 32181 21039 32215
rect 21039 32181 21048 32215
rect 20996 32172 21048 32181
rect 24676 32172 24728 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 84016 32104 84068 32156
rect 4620 31968 4672 32020
rect 6000 31968 6052 32020
rect 8116 32011 8168 32020
rect 8116 31977 8125 32011
rect 8125 31977 8159 32011
rect 8159 31977 8168 32011
rect 8116 31968 8168 31977
rect 8208 31968 8260 32020
rect 16672 31968 16724 32020
rect 18052 32011 18104 32020
rect 18052 31977 18061 32011
rect 18061 31977 18095 32011
rect 18095 31977 18104 32011
rect 18052 31968 18104 31977
rect 4620 31832 4672 31884
rect 5816 31875 5868 31884
rect 5816 31841 5825 31875
rect 5825 31841 5859 31875
rect 5859 31841 5868 31875
rect 5816 31832 5868 31841
rect 6552 31875 6604 31884
rect 6552 31841 6561 31875
rect 6561 31841 6595 31875
rect 6595 31841 6604 31875
rect 6552 31832 6604 31841
rect 7380 31832 7432 31884
rect 3516 31696 3568 31748
rect 12716 31900 12768 31952
rect 12992 31900 13044 31952
rect 19708 31900 19760 31952
rect 11244 31832 11296 31884
rect 12072 31832 12124 31884
rect 12808 31875 12860 31884
rect 12808 31841 12817 31875
rect 12817 31841 12851 31875
rect 12851 31841 12860 31875
rect 12808 31832 12860 31841
rect 8852 31764 8904 31816
rect 12716 31807 12768 31816
rect 12716 31773 12725 31807
rect 12725 31773 12759 31807
rect 12759 31773 12768 31807
rect 12716 31764 12768 31773
rect 12992 31764 13044 31816
rect 18512 31832 18564 31884
rect 19156 31875 19208 31884
rect 19156 31841 19165 31875
rect 19165 31841 19199 31875
rect 19199 31841 19208 31875
rect 23480 31968 23532 32020
rect 24952 32011 25004 32020
rect 24952 31977 24961 32011
rect 24961 31977 24995 32011
rect 24995 31977 25004 32011
rect 24952 31968 25004 31977
rect 27528 31968 27580 32020
rect 20352 31900 20404 31952
rect 22284 31900 22336 31952
rect 27804 31943 27856 31952
rect 27804 31909 27813 31943
rect 27813 31909 27847 31943
rect 27847 31909 27856 31943
rect 27804 31900 27856 31909
rect 48504 31968 48556 32020
rect 20996 31875 21048 31884
rect 19156 31832 19208 31841
rect 20996 31841 21005 31875
rect 21005 31841 21039 31875
rect 21039 31841 21048 31875
rect 20996 31832 21048 31841
rect 21548 31832 21600 31884
rect 24952 31832 25004 31884
rect 13820 31764 13872 31816
rect 18052 31764 18104 31816
rect 20536 31764 20588 31816
rect 27344 31764 27396 31816
rect 27620 31832 27672 31884
rect 27712 31764 27764 31816
rect 43076 31764 43128 31816
rect 13636 31696 13688 31748
rect 15200 31696 15252 31748
rect 16488 31696 16540 31748
rect 19892 31696 19944 31748
rect 8576 31628 8628 31680
rect 8852 31628 8904 31680
rect 12992 31628 13044 31680
rect 13728 31628 13780 31680
rect 16212 31628 16264 31680
rect 24584 31628 24636 31680
rect 26792 31628 26844 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 2872 31331 2924 31340
rect 2872 31297 2881 31331
rect 2881 31297 2915 31331
rect 2915 31297 2924 31331
rect 2872 31288 2924 31297
rect 4896 31424 4948 31476
rect 8024 31467 8076 31476
rect 8024 31433 8033 31467
rect 8033 31433 8067 31467
rect 8067 31433 8076 31467
rect 8024 31424 8076 31433
rect 7472 31356 7524 31408
rect 7656 31356 7708 31408
rect 6276 31288 6328 31340
rect 7656 31220 7708 31272
rect 8668 31424 8720 31476
rect 9772 31424 9824 31476
rect 19248 31424 19300 31476
rect 33508 31424 33560 31476
rect 5080 31152 5132 31204
rect 12900 31356 12952 31408
rect 13176 31356 13228 31408
rect 18052 31288 18104 31340
rect 19432 31288 19484 31340
rect 20168 31331 20220 31340
rect 20168 31297 20177 31331
rect 20177 31297 20211 31331
rect 20211 31297 20220 31331
rect 20168 31288 20220 31297
rect 21548 31331 21600 31340
rect 21548 31297 21557 31331
rect 21557 31297 21591 31331
rect 21591 31297 21600 31331
rect 21548 31288 21600 31297
rect 10048 31263 10100 31272
rect 9588 31195 9640 31204
rect 9588 31161 9597 31195
rect 9597 31161 9631 31195
rect 9631 31161 9640 31195
rect 9588 31152 9640 31161
rect 4160 31127 4212 31136
rect 4160 31093 4169 31127
rect 4169 31093 4203 31127
rect 4203 31093 4212 31127
rect 4160 31084 4212 31093
rect 9680 31127 9732 31136
rect 9680 31093 9689 31127
rect 9689 31093 9723 31127
rect 9723 31093 9732 31127
rect 10048 31229 10057 31263
rect 10057 31229 10091 31263
rect 10091 31229 10100 31263
rect 10048 31220 10100 31229
rect 11152 31195 11204 31204
rect 11152 31161 11161 31195
rect 11161 31161 11195 31195
rect 11195 31161 11204 31195
rect 11152 31152 11204 31161
rect 13728 31220 13780 31272
rect 12992 31152 13044 31204
rect 16488 31220 16540 31272
rect 20628 31220 20680 31272
rect 23756 31220 23808 31272
rect 27344 31356 27396 31408
rect 27528 31399 27580 31408
rect 27528 31365 27537 31399
rect 27537 31365 27571 31399
rect 27571 31365 27580 31399
rect 27528 31356 27580 31365
rect 32036 31356 32088 31408
rect 59728 31560 59780 31612
rect 87144 31560 87196 31612
rect 87880 31560 87932 31612
rect 59360 31492 59412 31544
rect 24032 31288 24084 31340
rect 24676 31220 24728 31272
rect 24952 31220 25004 31272
rect 26792 31220 26844 31272
rect 32404 31288 32456 31340
rect 16396 31152 16448 31204
rect 19432 31152 19484 31204
rect 9680 31084 9732 31093
rect 20996 31152 21048 31204
rect 28356 31152 28408 31204
rect 21548 31084 21600 31136
rect 23940 31127 23992 31136
rect 23940 31093 23949 31127
rect 23949 31093 23983 31127
rect 23983 31093 23992 31127
rect 23940 31084 23992 31093
rect 26792 31084 26844 31136
rect 27344 31084 27396 31136
rect 41604 31220 41656 31272
rect 56600 31220 56652 31272
rect 32680 31152 32732 31204
rect 87236 31152 87288 31204
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 2964 30880 3016 30932
rect 2780 30744 2832 30796
rect 3976 30744 4028 30796
rect 20352 30880 20404 30932
rect 20444 30880 20496 30932
rect 25964 30880 26016 30932
rect 27712 30880 27764 30932
rect 9588 30812 9640 30864
rect 12164 30812 12216 30864
rect 4712 30719 4764 30728
rect 4712 30685 4721 30719
rect 4721 30685 4755 30719
rect 4755 30685 4764 30719
rect 4712 30676 4764 30685
rect 7748 30744 7800 30796
rect 11060 30744 11112 30796
rect 13360 30744 13412 30796
rect 13728 30787 13780 30796
rect 5724 30608 5776 30660
rect 4620 30540 4672 30592
rect 4896 30540 4948 30592
rect 12900 30676 12952 30728
rect 13728 30753 13737 30787
rect 13737 30753 13771 30787
rect 13771 30753 13780 30787
rect 13728 30744 13780 30753
rect 15016 30676 15068 30728
rect 17776 30812 17828 30864
rect 18052 30855 18104 30864
rect 18052 30821 18061 30855
rect 18061 30821 18095 30855
rect 18095 30821 18104 30855
rect 18052 30812 18104 30821
rect 18972 30812 19024 30864
rect 16304 30744 16356 30796
rect 16764 30744 16816 30796
rect 18880 30744 18932 30796
rect 19156 30812 19208 30864
rect 21640 30812 21692 30864
rect 22652 30812 22704 30864
rect 24032 30812 24084 30864
rect 25596 30855 25648 30864
rect 25596 30821 25605 30855
rect 25605 30821 25639 30855
rect 25639 30821 25648 30855
rect 25596 30812 25648 30821
rect 27528 30812 27580 30864
rect 86868 31084 86920 31136
rect 87420 31084 87472 31136
rect 32496 31016 32548 31068
rect 86132 31016 86184 31068
rect 86960 31016 87012 31068
rect 32588 30948 32640 31000
rect 108304 31016 108356 31068
rect 87052 30880 87104 30932
rect 86224 30812 86276 30864
rect 25228 30744 25280 30796
rect 26792 30787 26844 30796
rect 26792 30753 26801 30787
rect 26801 30753 26835 30787
rect 26835 30753 26844 30787
rect 26792 30744 26844 30753
rect 23480 30676 23532 30728
rect 19064 30608 19116 30660
rect 9220 30540 9272 30592
rect 12164 30540 12216 30592
rect 13360 30540 13412 30592
rect 15200 30540 15252 30592
rect 16672 30540 16724 30592
rect 26976 30540 27028 30592
rect 27252 30540 27304 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 4620 30336 4672 30388
rect 5724 30379 5776 30388
rect 3148 30268 3200 30320
rect 3976 30200 4028 30252
rect 2688 30175 2740 30184
rect 2688 30141 2697 30175
rect 2697 30141 2731 30175
rect 2731 30141 2740 30175
rect 2688 30132 2740 30141
rect 4528 30175 4580 30184
rect 4528 30141 4537 30175
rect 4537 30141 4571 30175
rect 4571 30141 4580 30175
rect 4528 30132 4580 30141
rect 5724 30345 5733 30379
rect 5733 30345 5767 30379
rect 5767 30345 5776 30379
rect 5724 30336 5776 30345
rect 7656 30336 7708 30388
rect 10600 30336 10652 30388
rect 13176 30336 13228 30388
rect 11060 30311 11112 30320
rect 11060 30277 11069 30311
rect 11069 30277 11103 30311
rect 11103 30277 11112 30311
rect 11060 30268 11112 30277
rect 13820 30336 13872 30388
rect 16304 30336 16356 30388
rect 5172 30132 5224 30184
rect 9680 30132 9732 30184
rect 10600 30175 10652 30184
rect 10600 30141 10609 30175
rect 10609 30141 10643 30175
rect 10643 30141 10652 30175
rect 10600 30132 10652 30141
rect 11520 30200 11572 30252
rect 12072 30132 12124 30184
rect 12900 30132 12952 30184
rect 3792 30064 3844 30116
rect 14464 30064 14516 30116
rect 15292 30132 15344 30184
rect 17224 30268 17276 30320
rect 19432 30336 19484 30388
rect 19340 30268 19392 30320
rect 25044 30336 25096 30388
rect 21088 30268 21140 30320
rect 16764 30200 16816 30252
rect 17500 30200 17552 30252
rect 18236 30243 18288 30252
rect 18236 30209 18242 30243
rect 18242 30209 18288 30243
rect 18236 30200 18288 30209
rect 18420 30243 18472 30252
rect 18420 30209 18429 30243
rect 18429 30209 18463 30243
rect 18463 30209 18472 30243
rect 18420 30200 18472 30209
rect 21640 30200 21692 30252
rect 23480 30200 23532 30252
rect 24492 30268 24544 30320
rect 28816 30268 28868 30320
rect 19340 30132 19392 30184
rect 21548 30175 21600 30184
rect 21548 30141 21557 30175
rect 21557 30141 21591 30175
rect 21591 30141 21600 30175
rect 21548 30132 21600 30141
rect 22744 30132 22796 30184
rect 24492 30175 24544 30184
rect 17224 30107 17276 30116
rect 17224 30073 17233 30107
rect 17233 30073 17267 30107
rect 17267 30073 17276 30107
rect 17224 30064 17276 30073
rect 4528 29996 4580 30048
rect 5540 29996 5592 30048
rect 9772 30039 9824 30048
rect 9772 30005 9781 30039
rect 9781 30005 9815 30039
rect 9815 30005 9824 30039
rect 9772 29996 9824 30005
rect 12992 29996 13044 30048
rect 15016 30039 15068 30048
rect 15016 30005 15025 30039
rect 15025 30005 15059 30039
rect 15059 30005 15068 30039
rect 15016 29996 15068 30005
rect 15384 30039 15436 30048
rect 15384 30005 15393 30039
rect 15393 30005 15427 30039
rect 15427 30005 15436 30039
rect 15384 29996 15436 30005
rect 16672 29996 16724 30048
rect 18052 30107 18104 30116
rect 18052 30073 18061 30107
rect 18061 30073 18095 30107
rect 18095 30073 18104 30107
rect 18052 30064 18104 30073
rect 18328 30064 18380 30116
rect 24492 30141 24501 30175
rect 24501 30141 24535 30175
rect 24535 30141 24544 30175
rect 24492 30132 24544 30141
rect 24584 30175 24636 30184
rect 24584 30141 24593 30175
rect 24593 30141 24627 30175
rect 24627 30141 24636 30175
rect 24584 30132 24636 30141
rect 58440 30132 58492 30184
rect 58900 30132 58952 30184
rect 17500 30039 17552 30048
rect 17500 30005 17509 30039
rect 17509 30005 17543 30039
rect 17543 30005 17552 30039
rect 17500 29996 17552 30005
rect 18696 30039 18748 30048
rect 18696 30005 18705 30039
rect 18705 30005 18739 30039
rect 18739 30005 18748 30039
rect 18696 29996 18748 30005
rect 22744 29996 22796 30048
rect 27068 30064 27120 30116
rect 25044 30039 25096 30048
rect 25044 30005 25053 30039
rect 25053 30005 25087 30039
rect 25087 30005 25096 30039
rect 25044 29996 25096 30005
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 3332 29835 3384 29844
rect 3332 29801 3341 29835
rect 3341 29801 3375 29835
rect 3375 29801 3384 29835
rect 3332 29792 3384 29801
rect 4988 29835 5040 29844
rect 4988 29801 4997 29835
rect 4997 29801 5031 29835
rect 5031 29801 5040 29835
rect 4988 29792 5040 29801
rect 12072 29835 12124 29844
rect 12072 29801 12081 29835
rect 12081 29801 12115 29835
rect 12115 29801 12124 29835
rect 12072 29792 12124 29801
rect 14096 29835 14148 29844
rect 14096 29801 14105 29835
rect 14105 29801 14139 29835
rect 14139 29801 14148 29835
rect 14096 29792 14148 29801
rect 17500 29792 17552 29844
rect 2688 29699 2740 29708
rect 2688 29665 2697 29699
rect 2697 29665 2731 29699
rect 2731 29665 2740 29699
rect 2688 29656 2740 29665
rect 3700 29656 3752 29708
rect 3884 29656 3936 29708
rect 16580 29724 16632 29776
rect 6092 29699 6144 29708
rect 6092 29665 6101 29699
rect 6101 29665 6135 29699
rect 6135 29665 6144 29699
rect 6092 29656 6144 29665
rect 11152 29656 11204 29708
rect 13912 29699 13964 29708
rect 13912 29665 13921 29699
rect 13921 29665 13955 29699
rect 13955 29665 13964 29699
rect 13912 29656 13964 29665
rect 18052 29724 18104 29776
rect 18880 29724 18932 29776
rect 17316 29699 17368 29708
rect 17316 29665 17325 29699
rect 17325 29665 17359 29699
rect 17359 29665 17368 29699
rect 17316 29656 17368 29665
rect 18144 29656 18196 29708
rect 19708 29724 19760 29776
rect 24860 29792 24912 29844
rect 58440 29792 58492 29844
rect 59084 29792 59136 29844
rect 19892 29724 19944 29776
rect 2964 29631 3016 29640
rect 2964 29597 2973 29631
rect 2973 29597 3007 29631
rect 3007 29597 3016 29631
rect 2964 29588 3016 29597
rect 4068 29588 4120 29640
rect 3056 29520 3108 29572
rect 4804 29588 4856 29640
rect 7932 29588 7984 29640
rect 17500 29520 17552 29572
rect 4988 29452 5040 29504
rect 16580 29452 16632 29504
rect 17316 29452 17368 29504
rect 18420 29452 18472 29504
rect 20628 29452 20680 29504
rect 25044 29656 25096 29708
rect 25872 29588 25924 29640
rect 86224 29520 86276 29572
rect 87236 29520 87288 29572
rect 24676 29495 24728 29504
rect 24676 29461 24685 29495
rect 24685 29461 24719 29495
rect 24719 29461 24728 29495
rect 24676 29452 24728 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 3976 29248 4028 29300
rect 11520 29248 11572 29300
rect 18144 29291 18196 29300
rect 18144 29257 18153 29291
rect 18153 29257 18187 29291
rect 18187 29257 18196 29291
rect 18144 29248 18196 29257
rect 20260 29248 20312 29300
rect 24492 29248 24544 29300
rect 26700 29291 26752 29300
rect 5264 29180 5316 29232
rect 18696 29180 18748 29232
rect 26700 29257 26709 29291
rect 26709 29257 26743 29291
rect 26743 29257 26752 29291
rect 26700 29248 26752 29257
rect 29000 29248 29052 29300
rect 31484 29180 31536 29232
rect 4160 29044 4212 29096
rect 8576 29112 8628 29164
rect 13360 29112 13412 29164
rect 5172 29044 5224 29096
rect 13544 29044 13596 29096
rect 16764 29112 16816 29164
rect 26976 29112 27028 29164
rect 15016 29044 15068 29096
rect 14188 29019 14240 29028
rect 14188 28985 14197 29019
rect 14197 28985 14231 29019
rect 14231 28985 14240 29019
rect 14188 28976 14240 28985
rect 19340 29044 19392 29096
rect 25412 29087 25464 29096
rect 25412 29053 25421 29087
rect 25421 29053 25455 29087
rect 25455 29053 25464 29087
rect 25412 29044 25464 29053
rect 24676 28976 24728 29028
rect 3884 28951 3936 28960
rect 3884 28917 3893 28951
rect 3893 28917 3927 28951
rect 3927 28917 3936 28951
rect 3884 28908 3936 28917
rect 5172 28908 5224 28960
rect 9036 28908 9088 28960
rect 15016 28951 15068 28960
rect 15016 28917 15025 28951
rect 15025 28917 15059 28951
rect 15059 28917 15068 28951
rect 15016 28908 15068 28917
rect 17132 28908 17184 28960
rect 18420 28951 18472 28960
rect 18420 28917 18429 28951
rect 18429 28917 18463 28951
rect 18463 28917 18472 28951
rect 18420 28908 18472 28917
rect 26976 28951 27028 28960
rect 26976 28917 26985 28951
rect 26985 28917 27019 28951
rect 27019 28917 27028 28951
rect 26976 28908 27028 28917
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 4068 28704 4120 28756
rect 4988 28704 5040 28756
rect 4160 28636 4212 28688
rect 5264 28636 5316 28688
rect 5448 28568 5500 28620
rect 13912 28704 13964 28756
rect 13176 28636 13228 28688
rect 4620 28543 4672 28552
rect 4620 28509 4629 28543
rect 4629 28509 4663 28543
rect 4663 28509 4672 28543
rect 4620 28500 4672 28509
rect 5908 28364 5960 28416
rect 6828 28364 6880 28416
rect 13728 28611 13780 28620
rect 13728 28577 13737 28611
rect 13737 28577 13771 28611
rect 13771 28577 13780 28611
rect 13728 28568 13780 28577
rect 12992 28500 13044 28552
rect 16580 28500 16632 28552
rect 11704 28432 11756 28484
rect 12624 28475 12676 28484
rect 12624 28441 12633 28475
rect 12633 28441 12667 28475
rect 12667 28441 12676 28475
rect 12624 28432 12676 28441
rect 13912 28475 13964 28484
rect 13912 28441 13921 28475
rect 13921 28441 13955 28475
rect 13955 28441 13964 28475
rect 13912 28432 13964 28441
rect 17500 28611 17552 28620
rect 17500 28577 17509 28611
rect 17509 28577 17543 28611
rect 17543 28577 17552 28611
rect 17500 28568 17552 28577
rect 20260 28704 20312 28756
rect 26700 28568 26752 28620
rect 28080 28568 28132 28620
rect 28632 28500 28684 28552
rect 8484 28407 8536 28416
rect 8484 28373 8493 28407
rect 8493 28373 8527 28407
rect 8527 28373 8536 28407
rect 8484 28364 8536 28373
rect 17132 28407 17184 28416
rect 17132 28373 17141 28407
rect 17141 28373 17175 28407
rect 17175 28373 17184 28407
rect 17132 28364 17184 28373
rect 18420 28364 18472 28416
rect 19892 28407 19944 28416
rect 19892 28373 19901 28407
rect 19901 28373 19935 28407
rect 19935 28373 19944 28407
rect 19892 28364 19944 28373
rect 25228 28364 25280 28416
rect 27436 28407 27488 28416
rect 27436 28373 27445 28407
rect 27445 28373 27479 28407
rect 27479 28373 27488 28407
rect 27436 28364 27488 28373
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 8484 28160 8536 28212
rect 3608 28024 3660 28076
rect 18328 28160 18380 28212
rect 20720 28160 20772 28212
rect 20996 28160 21048 28212
rect 28080 28203 28132 28212
rect 28080 28169 28089 28203
rect 28089 28169 28123 28203
rect 28123 28169 28132 28203
rect 28080 28160 28132 28169
rect 28908 28160 28960 28212
rect 86224 28160 86276 28212
rect 87052 28160 87104 28212
rect 9864 28135 9916 28144
rect 9864 28101 9873 28135
rect 9873 28101 9907 28135
rect 9907 28101 9916 28135
rect 9864 28092 9916 28101
rect 11336 28135 11388 28144
rect 11336 28101 11345 28135
rect 11345 28101 11379 28135
rect 11379 28101 11388 28135
rect 11336 28092 11388 28101
rect 2596 27999 2648 28008
rect 2596 27965 2605 27999
rect 2605 27965 2639 27999
rect 2639 27965 2648 27999
rect 2596 27956 2648 27965
rect 5264 27999 5316 28008
rect 5264 27965 5273 27999
rect 5273 27965 5307 27999
rect 5307 27965 5316 27999
rect 5264 27956 5316 27965
rect 8484 27956 8536 28008
rect 3608 27888 3660 27940
rect 8760 27931 8812 27940
rect 4160 27863 4212 27872
rect 4160 27829 4169 27863
rect 4169 27829 4203 27863
rect 4203 27829 4212 27863
rect 4160 27820 4212 27829
rect 4804 27820 4856 27872
rect 8760 27897 8769 27931
rect 8769 27897 8803 27931
rect 8803 27897 8812 27931
rect 8760 27888 8812 27897
rect 9404 27956 9456 28008
rect 9680 27956 9732 28008
rect 11244 27888 11296 27940
rect 7656 27863 7708 27872
rect 7656 27829 7665 27863
rect 7665 27829 7699 27863
rect 7699 27829 7708 27863
rect 7656 27820 7708 27829
rect 11152 27863 11204 27872
rect 11152 27829 11161 27863
rect 11161 27829 11195 27863
rect 11195 27829 11204 27863
rect 16672 28092 16724 28144
rect 25412 28135 25464 28144
rect 25412 28101 25421 28135
rect 25421 28101 25455 28135
rect 25455 28101 25464 28135
rect 25412 28092 25464 28101
rect 13636 28067 13688 28076
rect 13636 28033 13645 28067
rect 13645 28033 13679 28067
rect 13679 28033 13688 28067
rect 13636 28024 13688 28033
rect 19432 28024 19484 28076
rect 26976 28024 27028 28076
rect 58440 28024 58492 28076
rect 59544 28024 59596 28076
rect 13084 27999 13136 28008
rect 13084 27965 13093 27999
rect 13093 27965 13127 27999
rect 13127 27965 13136 27999
rect 13084 27956 13136 27965
rect 13912 27956 13964 28008
rect 16396 27956 16448 28008
rect 19892 27999 19944 28008
rect 19892 27965 19901 27999
rect 19901 27965 19935 27999
rect 19935 27965 19944 27999
rect 19892 27956 19944 27965
rect 23940 27956 23992 28008
rect 16580 27888 16632 27940
rect 20996 27931 21048 27940
rect 11152 27820 11204 27829
rect 12992 27820 13044 27872
rect 13084 27820 13136 27872
rect 15016 27820 15068 27872
rect 19432 27820 19484 27872
rect 20996 27897 21005 27931
rect 21005 27897 21039 27931
rect 21039 27897 21048 27931
rect 20996 27888 21048 27897
rect 25228 27999 25280 28008
rect 25228 27965 25237 27999
rect 25237 27965 25271 27999
rect 25271 27965 25280 27999
rect 25228 27956 25280 27965
rect 27804 27956 27856 28008
rect 26608 27888 26660 27940
rect 59544 27931 59596 27940
rect 59544 27897 59553 27931
rect 59553 27897 59587 27931
rect 59587 27897 59596 27931
rect 59544 27888 59596 27897
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 8484 27659 8536 27668
rect 8484 27625 8493 27659
rect 8493 27625 8527 27659
rect 8527 27625 8536 27659
rect 8484 27616 8536 27625
rect 5264 27548 5316 27600
rect 5080 27480 5132 27532
rect 8760 27548 8812 27600
rect 9312 27616 9364 27668
rect 11152 27616 11204 27668
rect 12072 27616 12124 27668
rect 13728 27616 13780 27668
rect 26608 27616 26660 27668
rect 29000 27616 29052 27668
rect 59360 27616 59412 27668
rect 17316 27591 17368 27600
rect 9128 27523 9180 27532
rect 9128 27489 9137 27523
rect 9137 27489 9171 27523
rect 9171 27489 9180 27523
rect 9128 27480 9180 27489
rect 10600 27523 10652 27532
rect 10600 27489 10609 27523
rect 10609 27489 10643 27523
rect 10643 27489 10652 27523
rect 10600 27480 10652 27489
rect 12624 27480 12676 27532
rect 17316 27557 17325 27591
rect 17325 27557 17359 27591
rect 17359 27557 17368 27591
rect 17316 27548 17368 27557
rect 24860 27548 24912 27600
rect 25136 27548 25188 27600
rect 27804 27591 27856 27600
rect 27804 27557 27813 27591
rect 27813 27557 27847 27591
rect 27847 27557 27856 27591
rect 27804 27548 27856 27557
rect 15936 27523 15988 27532
rect 15936 27489 15945 27523
rect 15945 27489 15979 27523
rect 15979 27489 15988 27523
rect 16396 27523 16448 27532
rect 15936 27480 15988 27489
rect 16396 27489 16405 27523
rect 16405 27489 16439 27523
rect 16439 27489 16448 27523
rect 16396 27480 16448 27489
rect 2872 27412 2924 27464
rect 3516 27344 3568 27396
rect 10968 27344 11020 27396
rect 9588 27276 9640 27328
rect 11704 27412 11756 27464
rect 20996 27480 21048 27532
rect 24124 27480 24176 27532
rect 26700 27523 26752 27532
rect 26700 27489 26709 27523
rect 26709 27489 26743 27523
rect 26743 27489 26752 27523
rect 26700 27480 26752 27489
rect 27436 27523 27488 27532
rect 27436 27489 27445 27523
rect 27445 27489 27479 27523
rect 27479 27489 27488 27523
rect 27436 27480 27488 27489
rect 17132 27412 17184 27464
rect 20628 27412 20680 27464
rect 22284 27412 22336 27464
rect 23756 27412 23808 27464
rect 13084 27319 13136 27328
rect 13084 27285 13093 27319
rect 13093 27285 13127 27319
rect 13127 27285 13136 27319
rect 13084 27276 13136 27285
rect 16856 27319 16908 27328
rect 16856 27285 16865 27319
rect 16865 27285 16899 27319
rect 16899 27285 16908 27319
rect 16856 27276 16908 27285
rect 16948 27276 17000 27328
rect 17868 27276 17920 27328
rect 23572 27319 23624 27328
rect 23572 27285 23581 27319
rect 23581 27285 23615 27319
rect 23615 27285 23624 27319
rect 23572 27276 23624 27285
rect 26240 27319 26292 27328
rect 26240 27285 26249 27319
rect 26249 27285 26283 27319
rect 26283 27285 26292 27319
rect 26240 27276 26292 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 2596 26979 2648 26988
rect 2596 26945 2605 26979
rect 2605 26945 2639 26979
rect 2639 26945 2648 26979
rect 2596 26936 2648 26945
rect 2872 26979 2924 26988
rect 2872 26945 2881 26979
rect 2881 26945 2915 26979
rect 2915 26945 2924 26979
rect 2872 26936 2924 26945
rect 9404 26936 9456 26988
rect 4252 26868 4304 26920
rect 4804 26868 4856 26920
rect 8576 26911 8628 26920
rect 8576 26877 8585 26911
rect 8585 26877 8619 26911
rect 8619 26877 8628 26911
rect 9220 26911 9272 26920
rect 8576 26868 8628 26877
rect 9220 26877 9229 26911
rect 9229 26877 9263 26911
rect 9263 26877 9272 26911
rect 9220 26868 9272 26877
rect 11336 27072 11388 27124
rect 13176 27115 13228 27124
rect 13176 27081 13185 27115
rect 13185 27081 13219 27115
rect 13219 27081 13228 27115
rect 13176 27072 13228 27081
rect 15936 27072 15988 27124
rect 26240 27072 26292 27124
rect 26608 27115 26660 27124
rect 26608 27081 26617 27115
rect 26617 27081 26651 27115
rect 26651 27081 26660 27115
rect 26608 27072 26660 27081
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 16856 26936 16908 26988
rect 13084 26911 13136 26920
rect 8392 26800 8444 26852
rect 13084 26877 13093 26911
rect 13093 26877 13127 26911
rect 13127 26877 13136 26911
rect 13084 26868 13136 26877
rect 12348 26800 12400 26852
rect 20812 26868 20864 26920
rect 22192 26936 22244 26988
rect 31024 26936 31076 26988
rect 87052 26936 87104 26988
rect 87328 26936 87380 26988
rect 21088 26868 21140 26920
rect 21548 26868 21600 26920
rect 4160 26775 4212 26784
rect 4160 26741 4169 26775
rect 4169 26741 4203 26775
rect 4203 26741 4212 26775
rect 4160 26732 4212 26741
rect 7564 26775 7616 26784
rect 7564 26741 7573 26775
rect 7573 26741 7607 26775
rect 7607 26741 7616 26775
rect 7564 26732 7616 26741
rect 11796 26732 11848 26784
rect 15660 26775 15712 26784
rect 15660 26741 15669 26775
rect 15669 26741 15703 26775
rect 15703 26741 15712 26775
rect 15660 26732 15712 26741
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 21548 26732 21600 26784
rect 25320 26911 25372 26920
rect 22376 26732 22428 26784
rect 25320 26877 25329 26911
rect 25329 26877 25363 26911
rect 25363 26877 25372 26911
rect 25320 26868 25372 26877
rect 58440 26800 58492 26852
rect 59360 26800 59412 26852
rect 25136 26732 25188 26784
rect 86224 26732 86276 26784
rect 87236 26732 87288 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 58440 26596 58492 26648
rect 59452 26596 59504 26648
rect 5908 26528 5960 26580
rect 6828 26528 6880 26580
rect 16856 26528 16908 26580
rect 22192 26528 22244 26580
rect 22376 26528 22428 26580
rect 27160 26528 27212 26580
rect 17592 26460 17644 26512
rect 17868 26503 17920 26512
rect 17868 26469 17877 26503
rect 17877 26469 17911 26503
rect 17911 26469 17920 26503
rect 17868 26460 17920 26469
rect 4620 26392 4672 26444
rect 7656 26392 7708 26444
rect 17132 26392 17184 26444
rect 21548 26435 21600 26444
rect 4252 26324 4304 26376
rect 9588 26324 9640 26376
rect 16672 26324 16724 26376
rect 21548 26401 21557 26435
rect 21557 26401 21591 26435
rect 21591 26401 21600 26435
rect 21548 26392 21600 26401
rect 26608 26392 26660 26444
rect 27804 26392 27856 26444
rect 17776 26256 17828 26308
rect 3516 26188 3568 26240
rect 25504 26231 25556 26240
rect 25504 26197 25513 26231
rect 25513 26197 25547 26231
rect 25547 26197 25556 26231
rect 25504 26188 25556 26197
rect 26792 26231 26844 26240
rect 26792 26197 26801 26231
rect 26801 26197 26835 26231
rect 26835 26197 26844 26231
rect 26792 26188 26844 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 3976 25984 4028 26036
rect 6276 25984 6328 26036
rect 8576 25984 8628 26036
rect 9312 26027 9364 26036
rect 9312 25993 9321 26027
rect 9321 25993 9355 26027
rect 9355 25993 9364 26027
rect 9312 25984 9364 25993
rect 8116 25916 8168 25968
rect 8668 25916 8720 25968
rect 11980 25916 12032 25968
rect 16672 25959 16724 25968
rect 7288 25848 7340 25900
rect 16672 25925 16681 25959
rect 16681 25925 16715 25959
rect 16715 25925 16724 25959
rect 16672 25916 16724 25925
rect 2596 25823 2648 25832
rect 2596 25789 2605 25823
rect 2605 25789 2639 25823
rect 2639 25789 2648 25823
rect 2596 25780 2648 25789
rect 7012 25780 7064 25832
rect 8392 25823 8444 25832
rect 8392 25789 8401 25823
rect 8401 25789 8435 25823
rect 8435 25789 8444 25823
rect 8392 25780 8444 25789
rect 8668 25823 8720 25832
rect 8668 25789 8677 25823
rect 8677 25789 8711 25823
rect 8711 25789 8720 25823
rect 8668 25780 8720 25789
rect 9312 25780 9364 25832
rect 4160 25687 4212 25696
rect 4160 25653 4169 25687
rect 4169 25653 4203 25687
rect 4203 25653 4212 25687
rect 4160 25644 4212 25653
rect 5448 25644 5500 25696
rect 7748 25644 7800 25696
rect 9956 25644 10008 25696
rect 10600 25644 10652 25696
rect 16304 25823 16356 25832
rect 16304 25789 16313 25823
rect 16313 25789 16347 25823
rect 16347 25789 16356 25823
rect 16304 25780 16356 25789
rect 23572 25984 23624 26036
rect 25320 25984 25372 26036
rect 27804 26027 27856 26036
rect 27804 25993 27813 26027
rect 27813 25993 27847 26027
rect 27847 25993 27856 26027
rect 27804 25984 27856 25993
rect 28908 25984 28960 26036
rect 17960 25780 18012 25832
rect 24124 25823 24176 25832
rect 19432 25712 19484 25764
rect 24124 25789 24133 25823
rect 24133 25789 24167 25823
rect 24167 25789 24176 25823
rect 24124 25780 24176 25789
rect 25504 25780 25556 25832
rect 15384 25644 15436 25696
rect 15936 25644 15988 25696
rect 18144 25687 18196 25696
rect 18144 25653 18153 25687
rect 18153 25653 18187 25687
rect 18187 25653 18196 25687
rect 18144 25644 18196 25653
rect 25228 25644 25280 25696
rect 26516 25823 26568 25832
rect 26516 25789 26525 25823
rect 26525 25789 26559 25823
rect 26559 25789 26568 25823
rect 26516 25780 26568 25789
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 86224 25576 86276 25628
rect 87144 25576 87196 25628
rect 11060 25440 11112 25492
rect 11980 25483 12032 25492
rect 11980 25449 11989 25483
rect 11989 25449 12023 25483
rect 12023 25449 12032 25483
rect 11980 25440 12032 25449
rect 7012 25304 7064 25356
rect 7748 25347 7800 25356
rect 7748 25313 7757 25347
rect 7757 25313 7791 25347
rect 7791 25313 7800 25347
rect 7748 25304 7800 25313
rect 11980 25304 12032 25356
rect 16304 25304 16356 25356
rect 20812 25440 20864 25492
rect 26516 25440 26568 25492
rect 18144 25372 18196 25424
rect 28264 25372 28316 25424
rect 17868 25304 17920 25356
rect 23572 25304 23624 25356
rect 24124 25304 24176 25356
rect 26792 25304 26844 25356
rect 16488 25279 16540 25288
rect 16488 25245 16497 25279
rect 16497 25245 16531 25279
rect 16531 25245 16540 25279
rect 16488 25236 16540 25245
rect 5448 25100 5500 25152
rect 8300 25100 8352 25152
rect 18328 25100 18380 25152
rect 24032 25143 24084 25152
rect 24032 25109 24041 25143
rect 24041 25109 24075 25143
rect 24075 25109 24084 25143
rect 24032 25100 24084 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 13176 24939 13228 24948
rect 13176 24905 13185 24939
rect 13185 24905 13219 24939
rect 13219 24905 13228 24939
rect 13176 24896 13228 24905
rect 14188 24896 14240 24948
rect 3608 24760 3660 24812
rect 12348 24828 12400 24880
rect 13360 24871 13412 24880
rect 13360 24837 13369 24871
rect 13369 24837 13403 24871
rect 13403 24837 13412 24871
rect 13360 24828 13412 24837
rect 2596 24735 2648 24744
rect 2596 24701 2605 24735
rect 2605 24701 2639 24735
rect 2639 24701 2648 24735
rect 2596 24692 2648 24701
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 7840 24735 7892 24744
rect 4620 24624 4672 24676
rect 5724 24624 5776 24676
rect 7840 24701 7849 24735
rect 7849 24701 7883 24735
rect 7883 24701 7892 24735
rect 7840 24692 7892 24701
rect 8024 24735 8076 24744
rect 8024 24701 8033 24735
rect 8033 24701 8067 24735
rect 8067 24701 8076 24735
rect 8024 24692 8076 24701
rect 8668 24692 8720 24744
rect 9956 24692 10008 24744
rect 8208 24624 8260 24676
rect 13544 24760 13596 24812
rect 15660 24760 15712 24812
rect 18328 24803 18380 24812
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 19432 24760 19484 24812
rect 20536 24760 20588 24812
rect 29000 24828 29052 24880
rect 11060 24624 11112 24676
rect 5448 24556 5500 24608
rect 9588 24556 9640 24608
rect 9956 24556 10008 24608
rect 11704 24692 11756 24744
rect 14188 24735 14240 24744
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 14280 24735 14332 24744
rect 14280 24701 14289 24735
rect 14289 24701 14323 24735
rect 14323 24701 14332 24735
rect 14280 24692 14332 24701
rect 16028 24735 16080 24744
rect 16028 24701 16037 24735
rect 16037 24701 16071 24735
rect 16071 24701 16080 24735
rect 16028 24692 16080 24701
rect 16396 24624 16448 24676
rect 16948 24692 17000 24744
rect 18144 24624 18196 24676
rect 13084 24556 13136 24608
rect 13728 24556 13780 24608
rect 14188 24556 14240 24608
rect 16028 24556 16080 24608
rect 16856 24556 16908 24608
rect 20720 24556 20772 24608
rect 24492 24692 24544 24744
rect 25228 24556 25280 24608
rect 25320 24556 25372 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 3976 24352 4028 24404
rect 9772 24352 9824 24404
rect 13544 24352 13596 24404
rect 16028 24352 16080 24404
rect 16488 24352 16540 24404
rect 24492 24395 24544 24404
rect 14004 24284 14056 24336
rect 5448 24216 5500 24268
rect 9956 24259 10008 24268
rect 9956 24225 9965 24259
rect 9965 24225 9999 24259
rect 9999 24225 10008 24259
rect 9956 24216 10008 24225
rect 15844 24216 15896 24268
rect 16856 24259 16908 24268
rect 16856 24225 16865 24259
rect 16865 24225 16899 24259
rect 16899 24225 16908 24259
rect 16856 24216 16908 24225
rect 20996 24284 21048 24336
rect 5816 24148 5868 24200
rect 8300 24148 8352 24200
rect 9588 24148 9640 24200
rect 15752 24148 15804 24200
rect 16764 24148 16816 24200
rect 17776 24148 17828 24200
rect 20720 24148 20772 24200
rect 6920 24055 6972 24064
rect 6920 24021 6929 24055
rect 6929 24021 6963 24055
rect 6963 24021 6972 24055
rect 6920 24012 6972 24021
rect 11152 24012 11204 24064
rect 11704 24012 11756 24064
rect 15844 24055 15896 24064
rect 15844 24021 15853 24055
rect 15853 24021 15887 24055
rect 15887 24021 15896 24055
rect 15844 24012 15896 24021
rect 15936 24012 15988 24064
rect 24492 24361 24501 24395
rect 24501 24361 24535 24395
rect 24535 24361 24544 24395
rect 24492 24352 24544 24361
rect 28724 24352 28776 24404
rect 23572 24216 23624 24268
rect 24124 24216 24176 24268
rect 25320 24216 25372 24268
rect 26516 24259 26568 24268
rect 26516 24225 26525 24259
rect 26525 24225 26559 24259
rect 26559 24225 26568 24259
rect 26516 24216 26568 24225
rect 22468 24080 22520 24132
rect 17960 24055 18012 24064
rect 17960 24021 17969 24055
rect 17969 24021 18003 24055
rect 18003 24021 18012 24055
rect 17960 24012 18012 24021
rect 26240 24148 26292 24200
rect 86224 24216 86276 24268
rect 86960 24216 87012 24268
rect 29000 24148 29052 24200
rect 25044 24080 25096 24132
rect 26700 24055 26752 24064
rect 26700 24021 26709 24055
rect 26709 24021 26743 24055
rect 26743 24021 26752 24055
rect 26700 24012 26752 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 5448 23808 5500 23860
rect 5816 23851 5868 23860
rect 5816 23817 5825 23851
rect 5825 23817 5859 23851
rect 5859 23817 5868 23851
rect 5816 23808 5868 23817
rect 12348 23808 12400 23860
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 16948 23808 17000 23860
rect 18052 23808 18104 23860
rect 19432 23808 19484 23860
rect 26240 23851 26292 23860
rect 9588 23740 9640 23792
rect 16028 23740 16080 23792
rect 24032 23740 24084 23792
rect 26240 23817 26249 23851
rect 26249 23817 26283 23851
rect 26283 23817 26292 23851
rect 26240 23808 26292 23817
rect 28724 23808 28776 23860
rect 26516 23740 26568 23792
rect 3884 23672 3936 23724
rect 7472 23715 7524 23724
rect 7472 23681 7481 23715
rect 7481 23681 7515 23715
rect 7515 23681 7524 23715
rect 7472 23672 7524 23681
rect 13084 23672 13136 23724
rect 26884 23672 26936 23724
rect 2596 23647 2648 23656
rect 2596 23613 2605 23647
rect 2605 23613 2639 23647
rect 2639 23613 2648 23647
rect 2596 23604 2648 23613
rect 5724 23647 5776 23656
rect 5724 23613 5733 23647
rect 5733 23613 5767 23647
rect 5767 23613 5776 23647
rect 5724 23604 5776 23613
rect 6920 23604 6972 23656
rect 7932 23604 7984 23656
rect 8852 23647 8904 23656
rect 8852 23613 8861 23647
rect 8861 23613 8895 23647
rect 8895 23613 8904 23647
rect 8852 23604 8904 23613
rect 10232 23579 10284 23588
rect 10232 23545 10241 23579
rect 10241 23545 10275 23579
rect 10275 23545 10284 23579
rect 10232 23536 10284 23545
rect 14096 23604 14148 23656
rect 14832 23604 14884 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 11336 23536 11388 23588
rect 15844 23579 15896 23588
rect 15844 23545 15853 23579
rect 15853 23545 15887 23579
rect 15887 23545 15896 23579
rect 15844 23536 15896 23545
rect 3976 23511 4028 23520
rect 3976 23477 3985 23511
rect 3985 23477 4019 23511
rect 4019 23477 4028 23511
rect 3976 23468 4028 23477
rect 7748 23511 7800 23520
rect 7748 23477 7757 23511
rect 7757 23477 7791 23511
rect 7791 23477 7800 23511
rect 7748 23468 7800 23477
rect 17868 23468 17920 23520
rect 21916 23511 21968 23520
rect 21916 23477 21925 23511
rect 21925 23477 21959 23511
rect 21959 23477 21968 23511
rect 21916 23468 21968 23477
rect 22468 23604 22520 23656
rect 22560 23468 22612 23520
rect 24216 23511 24268 23520
rect 24216 23477 24225 23511
rect 24225 23477 24259 23511
rect 24259 23477 24268 23511
rect 24216 23468 24268 23477
rect 25412 23604 25464 23656
rect 58440 23604 58492 23656
rect 58992 23604 59044 23656
rect 27160 23579 27212 23588
rect 27160 23545 27169 23579
rect 27169 23545 27203 23579
rect 27203 23545 27212 23579
rect 27160 23536 27212 23545
rect 25228 23468 25280 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 10232 23264 10284 23316
rect 32036 23264 32088 23316
rect 10692 23196 10744 23248
rect 11980 23239 12032 23248
rect 11980 23205 11989 23239
rect 11989 23205 12023 23239
rect 12023 23205 12032 23239
rect 11980 23196 12032 23205
rect 15200 23196 15252 23248
rect 20720 23239 20772 23248
rect 3332 23060 3384 23112
rect 4620 23060 4672 23112
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 12164 23128 12216 23180
rect 20720 23205 20729 23239
rect 20729 23205 20763 23239
rect 20763 23205 20772 23239
rect 22560 23239 22612 23248
rect 20720 23196 20772 23205
rect 9680 22924 9732 22976
rect 12164 22967 12216 22976
rect 12164 22933 12173 22967
rect 12173 22933 12207 22967
rect 12207 22933 12216 22967
rect 12164 22924 12216 22933
rect 13728 22924 13780 22976
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 14740 22924 14792 22976
rect 17868 23128 17920 23180
rect 22560 23205 22569 23239
rect 22569 23205 22603 23239
rect 22603 23205 22612 23239
rect 22560 23196 22612 23205
rect 24124 23196 24176 23248
rect 25412 23239 25464 23248
rect 25044 23171 25096 23180
rect 25044 23137 25053 23171
rect 25053 23137 25087 23171
rect 25087 23137 25096 23171
rect 25044 23128 25096 23137
rect 25412 23205 25421 23239
rect 25421 23205 25455 23239
rect 25455 23205 25464 23239
rect 25412 23196 25464 23205
rect 26700 23171 26752 23180
rect 26700 23137 26709 23171
rect 26709 23137 26743 23171
rect 26743 23137 26752 23171
rect 26700 23128 26752 23137
rect 27712 23128 27764 23180
rect 15752 23103 15804 23112
rect 15752 23069 15761 23103
rect 15761 23069 15795 23103
rect 15795 23069 15804 23103
rect 15752 23060 15804 23069
rect 21180 23103 21232 23112
rect 21180 23069 21189 23103
rect 21189 23069 21223 23103
rect 21223 23069 21232 23103
rect 21180 23060 21232 23069
rect 15476 22924 15528 22976
rect 21088 22924 21140 22976
rect 22652 22924 22704 22976
rect 26792 22924 26844 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 4068 22720 4120 22772
rect 25320 22720 25372 22772
rect 27620 22720 27672 22772
rect 29092 22720 29144 22772
rect 4804 22652 4856 22704
rect 5448 22652 5500 22704
rect 9588 22652 9640 22704
rect 14832 22695 14884 22704
rect 14832 22661 14841 22695
rect 14841 22661 14875 22695
rect 14875 22661 14884 22695
rect 14832 22652 14884 22661
rect 21180 22695 21232 22704
rect 21180 22661 21189 22695
rect 21189 22661 21223 22695
rect 21223 22661 21232 22695
rect 21180 22652 21232 22661
rect 5172 22584 5224 22636
rect 5356 22584 5408 22636
rect 5724 22584 5776 22636
rect 2596 22559 2648 22568
rect 2596 22525 2605 22559
rect 2605 22525 2639 22559
rect 2639 22525 2648 22559
rect 2596 22516 2648 22525
rect 8576 22559 8628 22568
rect 8576 22525 8585 22559
rect 8585 22525 8619 22559
rect 8619 22525 8628 22559
rect 8576 22516 8628 22525
rect 13728 22516 13780 22568
rect 9956 22491 10008 22500
rect 9956 22457 9965 22491
rect 9965 22457 9999 22491
rect 9999 22457 10008 22491
rect 9956 22448 10008 22457
rect 14004 22559 14056 22568
rect 14004 22525 14013 22559
rect 14013 22525 14047 22559
rect 14047 22525 14056 22559
rect 14004 22516 14056 22525
rect 14372 22516 14424 22568
rect 15752 22516 15804 22568
rect 2872 22380 2924 22432
rect 16672 22380 16724 22432
rect 25228 22584 25280 22636
rect 26792 22627 26844 22636
rect 26792 22593 26801 22627
rect 26801 22593 26835 22627
rect 26835 22593 26844 22627
rect 26792 22584 26844 22593
rect 20812 22559 20864 22568
rect 18696 22448 18748 22500
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 20812 22516 20864 22525
rect 21640 22516 21692 22568
rect 21916 22516 21968 22568
rect 21088 22448 21140 22500
rect 18604 22380 18656 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 8576 22219 8628 22228
rect 8576 22185 8585 22219
rect 8585 22185 8619 22219
rect 8619 22185 8628 22219
rect 8576 22176 8628 22185
rect 18604 22151 18656 22160
rect 18604 22117 18613 22151
rect 18613 22117 18647 22151
rect 18647 22117 18656 22151
rect 18604 22108 18656 22117
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 7288 21972 7340 22024
rect 10232 22040 10284 22092
rect 11336 22040 11388 22092
rect 11980 22040 12032 22092
rect 16764 22083 16816 22092
rect 16764 22049 16773 22083
rect 16773 22049 16807 22083
rect 16807 22049 16816 22083
rect 22376 22108 22428 22160
rect 16764 22040 16816 22049
rect 9772 21972 9824 22024
rect 17224 22015 17276 22024
rect 17224 21981 17233 22015
rect 17233 21981 17267 22015
rect 17267 21981 17276 22015
rect 17224 21972 17276 21981
rect 4068 21904 4120 21956
rect 27620 22083 27672 22092
rect 20720 21972 20772 22024
rect 21088 21972 21140 22024
rect 21640 22015 21692 22024
rect 21640 21981 21649 22015
rect 21649 21981 21683 22015
rect 21683 21981 21692 22015
rect 21640 21972 21692 21981
rect 27620 22049 27629 22083
rect 27629 22049 27663 22083
rect 27663 22049 27672 22083
rect 27620 22040 27672 22049
rect 27712 22083 27764 22092
rect 27712 22049 27721 22083
rect 27721 22049 27755 22083
rect 27755 22049 27764 22083
rect 27712 22040 27764 22049
rect 59360 22040 59412 22092
rect 59544 22040 59596 22092
rect 6920 21836 6972 21888
rect 7288 21836 7340 21888
rect 9036 21836 9088 21888
rect 11980 21879 12032 21888
rect 11980 21845 11989 21879
rect 11989 21845 12023 21879
rect 12023 21845 12032 21879
rect 11980 21836 12032 21845
rect 12164 21836 12216 21888
rect 21180 21904 21232 21956
rect 19800 21836 19852 21888
rect 21088 21836 21140 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 3608 21632 3660 21684
rect 4804 21632 4856 21684
rect 2596 21471 2648 21480
rect 2596 21437 2605 21471
rect 2605 21437 2639 21471
rect 2639 21437 2648 21471
rect 2596 21428 2648 21437
rect 8852 21564 8904 21616
rect 9680 21632 9732 21684
rect 11244 21564 11296 21616
rect 8208 21496 8260 21548
rect 7104 21292 7156 21344
rect 8116 21471 8168 21480
rect 8116 21437 8125 21471
rect 8125 21437 8159 21471
rect 8159 21437 8168 21471
rect 8116 21428 8168 21437
rect 9036 21428 9088 21480
rect 10876 21428 10928 21480
rect 11888 21496 11940 21548
rect 14096 21632 14148 21684
rect 17224 21632 17276 21684
rect 19340 21675 19392 21684
rect 19340 21641 19349 21675
rect 19349 21641 19383 21675
rect 19383 21641 19392 21675
rect 19340 21632 19392 21641
rect 22652 21564 22704 21616
rect 21272 21539 21324 21548
rect 21272 21505 21281 21539
rect 21281 21505 21315 21539
rect 21315 21505 21324 21539
rect 21272 21496 21324 21505
rect 13084 21471 13136 21480
rect 13084 21437 13093 21471
rect 13093 21437 13127 21471
rect 13127 21437 13136 21471
rect 13084 21428 13136 21437
rect 13176 21428 13228 21480
rect 16672 21471 16724 21480
rect 14464 21403 14516 21412
rect 14464 21369 14473 21403
rect 14473 21369 14507 21403
rect 14507 21369 14516 21403
rect 14464 21360 14516 21369
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 18788 21428 18840 21480
rect 20812 21428 20864 21480
rect 22008 21471 22060 21480
rect 22008 21437 22017 21471
rect 22017 21437 22051 21471
rect 22051 21437 22060 21471
rect 22008 21428 22060 21437
rect 22100 21428 22152 21480
rect 16764 21360 16816 21412
rect 22652 21360 22704 21412
rect 12440 21292 12492 21344
rect 21272 21292 21324 21344
rect 23940 21335 23992 21344
rect 23940 21301 23949 21335
rect 23949 21301 23983 21335
rect 23983 21301 23992 21335
rect 23940 21292 23992 21301
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 9956 21131 10008 21140
rect 9956 21097 9965 21131
rect 9965 21097 9999 21131
rect 9999 21097 10008 21131
rect 9956 21088 10008 21097
rect 11612 21131 11664 21140
rect 11612 21097 11621 21131
rect 11621 21097 11655 21131
rect 11655 21097 11664 21131
rect 11612 21088 11664 21097
rect 14464 21088 14516 21140
rect 13084 21020 13136 21072
rect 26148 21088 26200 21140
rect 27988 21088 28040 21140
rect 10692 20995 10744 21004
rect 10692 20961 10701 20995
rect 10701 20961 10735 20995
rect 10735 20961 10744 20995
rect 10692 20952 10744 20961
rect 11612 20952 11664 21004
rect 11888 20995 11940 21004
rect 11888 20961 11897 20995
rect 11897 20961 11931 20995
rect 11931 20961 11940 20995
rect 11888 20952 11940 20961
rect 12440 20995 12492 21004
rect 12440 20961 12449 20995
rect 12449 20961 12483 20995
rect 12483 20961 12492 20995
rect 12440 20952 12492 20961
rect 12900 20952 12952 21004
rect 14464 20952 14516 21004
rect 4068 20884 4120 20936
rect 11060 20816 11112 20868
rect 15016 20952 15068 21004
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 10968 20748 11020 20800
rect 11980 20748 12032 20800
rect 15200 20816 15252 20868
rect 16672 20952 16724 21004
rect 16764 20952 16816 21004
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 14740 20748 14792 20800
rect 21088 20884 21140 20936
rect 22008 20748 22060 20800
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 26240 20859 26292 20868
rect 26240 20825 26249 20859
rect 26249 20825 26283 20859
rect 26283 20825 26292 20859
rect 26240 20816 26292 20825
rect 23940 20791 23992 20800
rect 23940 20757 23949 20791
rect 23949 20757 23983 20791
rect 23983 20757 23992 20791
rect 23940 20748 23992 20757
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 2596 20544 2648 20596
rect 4804 20544 4856 20596
rect 11888 20544 11940 20596
rect 16764 20544 16816 20596
rect 20628 20544 20680 20596
rect 21180 20587 21232 20596
rect 21180 20553 21189 20587
rect 21189 20553 21223 20587
rect 21223 20553 21232 20587
rect 21180 20544 21232 20553
rect 22744 20544 22796 20596
rect 26240 20544 26292 20596
rect 27528 20544 27580 20596
rect 27896 20544 27948 20596
rect 18788 20476 18840 20528
rect 3148 20340 3200 20392
rect 10692 20383 10744 20392
rect 10692 20349 10701 20383
rect 10701 20349 10735 20383
rect 10735 20349 10744 20383
rect 10692 20340 10744 20349
rect 10876 20383 10928 20392
rect 10876 20349 10885 20383
rect 10885 20349 10919 20383
rect 10919 20349 10928 20383
rect 10876 20340 10928 20349
rect 12716 20340 12768 20392
rect 15292 20340 15344 20392
rect 16948 20272 17000 20324
rect 18788 20272 18840 20324
rect 3332 20204 3384 20256
rect 14832 20247 14884 20256
rect 14832 20213 14841 20247
rect 14841 20213 14875 20247
rect 14875 20213 14884 20247
rect 14832 20204 14884 20213
rect 18144 20204 18196 20256
rect 20168 20383 20220 20392
rect 19432 20272 19484 20324
rect 19156 20247 19208 20256
rect 19156 20213 19165 20247
rect 19165 20213 19199 20247
rect 19199 20213 19208 20247
rect 20168 20349 20177 20383
rect 20177 20349 20211 20383
rect 20211 20349 20220 20383
rect 20168 20340 20220 20349
rect 21088 20476 21140 20528
rect 22008 20476 22060 20528
rect 25320 20476 25372 20528
rect 21180 20340 21232 20392
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22100 20408 22152 20417
rect 25412 20408 25464 20460
rect 19984 20272 20036 20324
rect 22744 20383 22796 20392
rect 22744 20349 22753 20383
rect 22753 20349 22787 20383
rect 22787 20349 22796 20383
rect 22744 20340 22796 20349
rect 26240 20340 26292 20392
rect 58440 20272 58492 20324
rect 59176 20272 59228 20324
rect 19156 20204 19208 20213
rect 23756 20204 23808 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 2780 20043 2832 20052
rect 2780 20009 2789 20043
rect 2789 20009 2823 20043
rect 2823 20009 2832 20043
rect 2780 20000 2832 20009
rect 11060 19932 11112 19984
rect 13728 20000 13780 20052
rect 16764 20000 16816 20052
rect 21364 20000 21416 20052
rect 25412 20043 25464 20052
rect 25412 20009 25421 20043
rect 25421 20009 25455 20043
rect 25455 20009 25464 20043
rect 25412 20000 25464 20009
rect 27528 20043 27580 20052
rect 27528 20009 27537 20043
rect 27537 20009 27571 20043
rect 27571 20009 27580 20043
rect 27528 20000 27580 20009
rect 4620 19907 4672 19916
rect 4620 19873 4629 19907
rect 4629 19873 4663 19907
rect 4663 19873 4672 19907
rect 4620 19864 4672 19873
rect 5816 19907 5868 19916
rect 5816 19873 5825 19907
rect 5825 19873 5859 19907
rect 5859 19873 5868 19907
rect 5816 19864 5868 19873
rect 9496 19907 9548 19916
rect 9496 19873 9505 19907
rect 9505 19873 9539 19907
rect 9539 19873 9548 19907
rect 9496 19864 9548 19873
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 10048 19907 10100 19916
rect 10048 19873 10057 19907
rect 10057 19873 10091 19907
rect 10091 19873 10100 19907
rect 10048 19864 10100 19873
rect 10508 19907 10560 19916
rect 10508 19873 10517 19907
rect 10517 19873 10551 19907
rect 10551 19873 10560 19907
rect 10508 19864 10560 19873
rect 14740 19932 14792 19984
rect 12716 19907 12768 19916
rect 12716 19873 12725 19907
rect 12725 19873 12759 19907
rect 12759 19873 12768 19907
rect 12716 19864 12768 19873
rect 11244 19796 11296 19848
rect 15568 19839 15620 19848
rect 9772 19728 9824 19780
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 17040 19864 17092 19916
rect 24860 19864 24912 19916
rect 25780 19932 25832 19984
rect 25412 19864 25464 19916
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 16948 19839 17000 19848
rect 16948 19805 16957 19839
rect 16957 19805 16991 19839
rect 16991 19805 17000 19839
rect 16948 19796 17000 19805
rect 18144 19728 18196 19780
rect 24768 19728 24820 19780
rect 27988 19796 28040 19848
rect 4068 19660 4120 19712
rect 10048 19660 10100 19712
rect 10324 19660 10376 19712
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 14372 19660 14424 19712
rect 14924 19660 14976 19712
rect 26700 19703 26752 19712
rect 26700 19669 26709 19703
rect 26709 19669 26743 19703
rect 26743 19669 26752 19703
rect 26700 19660 26752 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 10324 19499 10376 19508
rect 10324 19465 10333 19499
rect 10333 19465 10367 19499
rect 10367 19465 10376 19499
rect 10324 19456 10376 19465
rect 11244 19456 11296 19508
rect 16764 19499 16816 19508
rect 16764 19465 16773 19499
rect 16773 19465 16807 19499
rect 16807 19465 16816 19499
rect 16764 19456 16816 19465
rect 20628 19456 20680 19508
rect 20904 19456 20956 19508
rect 7932 19363 7984 19372
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 9036 19320 9088 19372
rect 10140 19363 10192 19372
rect 2596 19295 2648 19304
rect 2596 19261 2605 19295
rect 2605 19261 2639 19295
rect 2639 19261 2648 19295
rect 2596 19252 2648 19261
rect 2964 19252 3016 19304
rect 5908 19252 5960 19304
rect 10140 19329 10149 19363
rect 10149 19329 10183 19363
rect 10183 19329 10192 19363
rect 10140 19320 10192 19329
rect 9680 19252 9732 19304
rect 10508 19252 10560 19304
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 11060 19252 11112 19304
rect 15568 19320 15620 19372
rect 2596 19116 2648 19168
rect 4896 19184 4948 19236
rect 5632 19227 5684 19236
rect 5632 19193 5641 19227
rect 5641 19193 5675 19227
rect 5675 19193 5684 19227
rect 5632 19184 5684 19193
rect 7196 19227 7248 19236
rect 7196 19193 7205 19227
rect 7205 19193 7239 19227
rect 7239 19193 7248 19227
rect 7196 19184 7248 19193
rect 7564 19227 7616 19236
rect 7564 19193 7573 19227
rect 7573 19193 7607 19227
rect 7607 19193 7616 19227
rect 7564 19184 7616 19193
rect 3976 19159 4028 19168
rect 3976 19125 3985 19159
rect 3985 19125 4019 19159
rect 4019 19125 4028 19159
rect 3976 19116 4028 19125
rect 7380 19159 7432 19168
rect 7380 19125 7389 19159
rect 7389 19125 7423 19159
rect 7423 19125 7432 19159
rect 7380 19116 7432 19125
rect 8576 19116 8628 19168
rect 17592 19252 17644 19304
rect 17868 19116 17920 19168
rect 19432 19252 19484 19304
rect 25688 19295 25740 19304
rect 24860 19184 24912 19236
rect 24952 19159 25004 19168
rect 24952 19125 24961 19159
rect 24961 19125 24995 19159
rect 24995 19125 25004 19159
rect 25688 19261 25697 19295
rect 25697 19261 25731 19295
rect 25731 19261 25740 19295
rect 25688 19252 25740 19261
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 26792 19184 26844 19236
rect 24952 19116 25004 19125
rect 25688 19116 25740 19168
rect 26700 19116 26752 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 4160 18955 4212 18964
rect 4160 18921 4169 18955
rect 4169 18921 4203 18955
rect 4203 18921 4212 18955
rect 4160 18912 4212 18921
rect 5632 18844 5684 18896
rect 9680 18844 9732 18896
rect 11060 18912 11112 18964
rect 11336 18912 11388 18964
rect 10416 18887 10468 18896
rect 10416 18853 10425 18887
rect 10425 18853 10459 18887
rect 10459 18853 10468 18887
rect 10416 18844 10468 18853
rect 10968 18844 11020 18896
rect 12164 18844 12216 18896
rect 18420 18912 18472 18964
rect 23756 18912 23808 18964
rect 18144 18887 18196 18896
rect 5080 18776 5132 18828
rect 8576 18776 8628 18828
rect 11336 18776 11388 18828
rect 6368 18708 6420 18760
rect 7196 18708 7248 18760
rect 8852 18708 8904 18760
rect 3424 18640 3476 18692
rect 4988 18572 5040 18624
rect 9220 18640 9272 18692
rect 10416 18640 10468 18692
rect 10784 18640 10836 18692
rect 18144 18853 18153 18887
rect 18153 18853 18187 18887
rect 18187 18853 18196 18887
rect 18144 18844 18196 18853
rect 14280 18708 14332 18760
rect 16396 18776 16448 18828
rect 18972 18819 19024 18828
rect 18972 18785 18981 18819
rect 18981 18785 19015 18819
rect 19015 18785 19024 18819
rect 18972 18776 19024 18785
rect 20168 18844 20220 18896
rect 19432 18819 19484 18828
rect 19432 18785 19441 18819
rect 19441 18785 19475 18819
rect 19475 18785 19484 18819
rect 19432 18776 19484 18785
rect 21180 18776 21232 18828
rect 24032 18776 24084 18828
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 18788 18708 18840 18760
rect 24216 18751 24268 18760
rect 24216 18717 24225 18751
rect 24225 18717 24259 18751
rect 24259 18717 24268 18751
rect 24216 18708 24268 18717
rect 24124 18640 24176 18692
rect 25044 18708 25096 18760
rect 25780 18640 25832 18692
rect 14464 18572 14516 18624
rect 15752 18615 15804 18624
rect 15752 18581 15761 18615
rect 15761 18581 15795 18615
rect 15795 18581 15804 18615
rect 15752 18572 15804 18581
rect 17040 18615 17092 18624
rect 17040 18581 17049 18615
rect 17049 18581 17083 18615
rect 17083 18581 17092 18615
rect 17040 18572 17092 18581
rect 17132 18572 17184 18624
rect 21732 18572 21784 18624
rect 24032 18615 24084 18624
rect 24032 18581 24041 18615
rect 24041 18581 24075 18615
rect 24075 18581 24084 18615
rect 24032 18572 24084 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 5080 18368 5132 18420
rect 7196 18300 7248 18352
rect 7288 18300 7340 18352
rect 12440 18300 12492 18352
rect 13544 18300 13596 18352
rect 13636 18300 13688 18352
rect 14832 18368 14884 18420
rect 15200 18368 15252 18420
rect 24032 18368 24084 18420
rect 25320 18368 25372 18420
rect 25872 18368 25924 18420
rect 27712 18411 27764 18420
rect 27712 18377 27721 18411
rect 27721 18377 27755 18411
rect 27755 18377 27764 18411
rect 27712 18368 27764 18377
rect 21180 18343 21232 18352
rect 21180 18309 21189 18343
rect 21189 18309 21223 18343
rect 21223 18309 21232 18343
rect 21180 18300 21232 18309
rect 25780 18300 25832 18352
rect 5816 18275 5868 18284
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 5816 18232 5868 18241
rect 8852 18232 8904 18284
rect 18512 18232 18564 18284
rect 3148 18096 3200 18148
rect 2964 18028 3016 18080
rect 5172 18207 5224 18216
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 5172 18164 5224 18173
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 6276 18164 6328 18216
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 8576 18164 8628 18216
rect 11152 18164 11204 18216
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 13452 18207 13504 18216
rect 13452 18173 13461 18207
rect 13461 18173 13495 18207
rect 13495 18173 13504 18207
rect 13452 18164 13504 18173
rect 13544 18164 13596 18216
rect 15016 18207 15068 18216
rect 15016 18173 15022 18207
rect 15022 18173 15068 18207
rect 15016 18164 15068 18173
rect 16396 18207 16448 18216
rect 8116 18071 8168 18080
rect 3424 18028 3476 18037
rect 8116 18037 8125 18071
rect 8125 18037 8159 18071
rect 8159 18037 8168 18071
rect 8116 18028 8168 18037
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 10048 18096 10100 18148
rect 13176 18096 13228 18148
rect 16396 18173 16405 18207
rect 16405 18173 16439 18207
rect 16439 18173 16448 18207
rect 16396 18164 16448 18173
rect 24768 18164 24820 18216
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 25780 18207 25832 18216
rect 25780 18173 25789 18207
rect 25789 18173 25823 18207
rect 25823 18173 25832 18207
rect 25780 18164 25832 18173
rect 25872 18207 25924 18216
rect 25872 18173 25881 18207
rect 25881 18173 25915 18207
rect 25915 18173 25924 18207
rect 25872 18164 25924 18173
rect 15752 18096 15804 18148
rect 18972 18096 19024 18148
rect 10876 18028 10928 18080
rect 11796 18028 11848 18080
rect 13452 18028 13504 18080
rect 15200 18028 15252 18080
rect 16672 18028 16724 18080
rect 17868 18028 17920 18080
rect 21180 18096 21232 18148
rect 32772 18232 32824 18284
rect 27712 18164 27764 18216
rect 26424 18139 26476 18148
rect 26424 18105 26433 18139
rect 26433 18105 26467 18139
rect 26467 18105 26476 18139
rect 26424 18096 26476 18105
rect 21548 18028 21600 18080
rect 24768 18028 24820 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 4620 17824 4672 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 9220 17824 9272 17876
rect 10784 17824 10836 17876
rect 5172 17756 5224 17808
rect 2964 17731 3016 17740
rect 2964 17697 2973 17731
rect 2973 17697 3007 17731
rect 3007 17697 3016 17731
rect 2964 17688 3016 17697
rect 4620 17688 4672 17740
rect 6000 17731 6052 17740
rect 5080 17620 5132 17672
rect 2964 17484 3016 17536
rect 3148 17484 3200 17536
rect 3700 17484 3752 17536
rect 6000 17697 6009 17731
rect 6009 17697 6043 17731
rect 6043 17697 6052 17731
rect 6000 17688 6052 17697
rect 6276 17731 6328 17740
rect 6276 17697 6285 17731
rect 6285 17697 6319 17731
rect 6319 17697 6328 17731
rect 6276 17688 6328 17697
rect 7932 17756 7984 17808
rect 10508 17799 10560 17808
rect 9036 17688 9088 17740
rect 10508 17765 10517 17799
rect 10517 17765 10551 17799
rect 10551 17765 10560 17799
rect 10508 17756 10560 17765
rect 10876 17756 10928 17808
rect 12716 17824 12768 17876
rect 11060 17756 11112 17808
rect 12164 17799 12216 17808
rect 12164 17765 12173 17799
rect 12173 17765 12207 17799
rect 12207 17765 12216 17799
rect 12164 17756 12216 17765
rect 5356 17552 5408 17604
rect 9680 17688 9732 17740
rect 10416 17688 10468 17740
rect 11244 17688 11296 17740
rect 11336 17688 11388 17740
rect 18696 17756 18748 17808
rect 10876 17620 10928 17672
rect 12624 17620 12676 17672
rect 9680 17552 9732 17604
rect 16488 17620 16540 17672
rect 10508 17484 10560 17536
rect 15108 17484 15160 17536
rect 17960 17688 18012 17740
rect 20720 17688 20772 17740
rect 20904 17731 20956 17740
rect 20904 17697 20913 17731
rect 20913 17697 20947 17731
rect 20947 17697 20956 17731
rect 20904 17688 20956 17697
rect 22376 17731 22428 17740
rect 17040 17620 17092 17672
rect 19432 17620 19484 17672
rect 22376 17697 22385 17731
rect 22385 17697 22419 17731
rect 22419 17697 22428 17731
rect 22376 17688 22428 17697
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 23848 17824 23900 17876
rect 24032 17824 24084 17876
rect 26240 17867 26292 17876
rect 23756 17756 23808 17808
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 27712 17824 27764 17876
rect 26332 17688 26384 17740
rect 26424 17688 26476 17740
rect 23664 17620 23716 17672
rect 25688 17620 25740 17672
rect 26240 17620 26292 17672
rect 17500 17552 17552 17604
rect 22192 17552 22244 17604
rect 20904 17484 20956 17536
rect 22100 17484 22152 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 3424 17280 3476 17332
rect 3424 17076 3476 17128
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 4252 17119 4304 17128
rect 4252 17085 4261 17119
rect 4261 17085 4295 17119
rect 4295 17085 4304 17119
rect 4252 17076 4304 17085
rect 4620 17076 4672 17128
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 6276 17280 6328 17332
rect 9588 17280 9640 17332
rect 8852 17212 8904 17264
rect 9404 17212 9456 17264
rect 4896 17076 4948 17085
rect 5172 17008 5224 17060
rect 9036 17119 9088 17128
rect 9036 17085 9045 17119
rect 9045 17085 9079 17119
rect 9079 17085 9088 17119
rect 9036 17076 9088 17085
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 7288 17008 7340 17060
rect 9864 17008 9916 17060
rect 10416 17008 10468 17060
rect 16856 17323 16908 17332
rect 16856 17289 16865 17323
rect 16865 17289 16899 17323
rect 16899 17289 16908 17323
rect 16856 17280 16908 17289
rect 21180 17280 21232 17332
rect 21824 17323 21876 17332
rect 14096 17119 14148 17128
rect 14096 17085 14105 17119
rect 14105 17085 14139 17119
rect 14139 17085 14148 17119
rect 14096 17076 14148 17085
rect 15016 17144 15068 17196
rect 16764 17212 16816 17264
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 14372 17076 14424 17128
rect 15476 17119 15528 17128
rect 15476 17085 15485 17119
rect 15485 17085 15519 17119
rect 15519 17085 15528 17119
rect 15476 17076 15528 17085
rect 16672 17119 16724 17128
rect 16672 17085 16681 17119
rect 16681 17085 16715 17119
rect 16715 17085 16724 17119
rect 24952 17144 25004 17196
rect 25228 17144 25280 17196
rect 16672 17076 16724 17085
rect 15200 17008 15252 17060
rect 3056 16940 3108 16992
rect 4068 16940 4120 16992
rect 8944 16940 8996 16992
rect 12532 16983 12584 16992
rect 12532 16949 12541 16983
rect 12541 16949 12575 16983
rect 12575 16949 12584 16983
rect 12532 16940 12584 16949
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 15568 16940 15620 16949
rect 22376 17076 22428 17128
rect 25320 17076 25372 17128
rect 26332 17119 26384 17128
rect 26332 17085 26341 17119
rect 26341 17085 26375 17119
rect 26375 17085 26384 17119
rect 26332 17076 26384 17085
rect 27252 17076 27304 17128
rect 21088 17008 21140 17060
rect 24676 17008 24728 17060
rect 26792 17008 26844 17060
rect 21732 16940 21784 16992
rect 22560 16940 22612 16992
rect 25228 16983 25280 16992
rect 25228 16949 25237 16983
rect 25237 16949 25271 16983
rect 25271 16949 25280 16983
rect 25228 16940 25280 16949
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 4160 16736 4212 16788
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 5356 16779 5408 16788
rect 4252 16736 4304 16745
rect 5356 16745 5365 16779
rect 5365 16745 5399 16779
rect 5399 16745 5408 16779
rect 5356 16736 5408 16745
rect 7380 16668 7432 16720
rect 9220 16668 9272 16720
rect 9496 16711 9548 16720
rect 9496 16677 9505 16711
rect 9505 16677 9539 16711
rect 9539 16677 9548 16711
rect 9496 16668 9548 16677
rect 3700 16600 3752 16652
rect 5264 16600 5316 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 10048 16643 10100 16652
rect 10048 16609 10057 16643
rect 10057 16609 10091 16643
rect 10091 16609 10100 16643
rect 10048 16600 10100 16609
rect 10140 16600 10192 16652
rect 10508 16643 10560 16652
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 10692 16600 10744 16652
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 11428 16600 11480 16652
rect 15108 16736 15160 16788
rect 17500 16779 17552 16788
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 14372 16668 14424 16720
rect 15200 16668 15252 16720
rect 16488 16668 16540 16720
rect 12348 16532 12400 16584
rect 16396 16643 16448 16652
rect 16396 16609 16405 16643
rect 16405 16609 16439 16643
rect 16439 16609 16448 16643
rect 16396 16600 16448 16609
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 17960 16736 18012 16788
rect 21916 16736 21968 16788
rect 22560 16779 22612 16788
rect 22560 16745 22569 16779
rect 22569 16745 22603 16779
rect 22603 16745 22612 16779
rect 22560 16736 22612 16745
rect 16764 16600 16816 16652
rect 13820 16575 13872 16584
rect 13820 16541 13829 16575
rect 13829 16541 13863 16575
rect 13863 16541 13872 16575
rect 13820 16532 13872 16541
rect 14096 16532 14148 16584
rect 14280 16532 14332 16584
rect 16948 16532 17000 16584
rect 19984 16668 20036 16720
rect 20812 16600 20864 16652
rect 20904 16643 20956 16652
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 21088 16643 21140 16652
rect 20904 16600 20956 16609
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 21180 16600 21232 16652
rect 21732 16643 21784 16652
rect 21732 16609 21741 16643
rect 21741 16609 21775 16643
rect 21775 16609 21784 16643
rect 21732 16600 21784 16609
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 24216 16600 24268 16652
rect 3884 16464 3936 16516
rect 16304 16464 16356 16516
rect 2964 16396 3016 16448
rect 12256 16396 12308 16448
rect 13268 16396 13320 16448
rect 32680 16532 32732 16584
rect 17776 16464 17828 16516
rect 32496 16464 32548 16516
rect 20628 16396 20680 16448
rect 23296 16439 23348 16448
rect 23296 16405 23305 16439
rect 23305 16405 23339 16439
rect 23339 16405 23348 16439
rect 23296 16396 23348 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 6000 16192 6052 16244
rect 13176 16235 13228 16244
rect 13176 16201 13185 16235
rect 13185 16201 13219 16235
rect 13219 16201 13228 16235
rect 13176 16192 13228 16201
rect 16028 16192 16080 16244
rect 21180 16192 21232 16244
rect 21640 16192 21692 16244
rect 27252 16235 27304 16244
rect 27252 16201 27261 16235
rect 27261 16201 27295 16235
rect 27295 16201 27304 16235
rect 27252 16192 27304 16201
rect 16304 16124 16356 16176
rect 20076 16124 20128 16176
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 2872 16099 2924 16108
rect 2872 16065 2881 16099
rect 2881 16065 2915 16099
rect 2915 16065 2924 16099
rect 2872 16056 2924 16065
rect 12348 16056 12400 16108
rect 12532 16056 12584 16108
rect 13912 16056 13964 16108
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 9312 15988 9364 16040
rect 9772 16031 9824 16040
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 7288 15920 7340 15972
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 4252 15852 4304 15904
rect 6736 15852 6788 15904
rect 8760 15852 8812 15904
rect 10600 15988 10652 16040
rect 12716 15988 12768 16040
rect 14096 16031 14148 16040
rect 14096 15997 14105 16031
rect 14105 15997 14139 16031
rect 14139 15997 14148 16031
rect 14096 15988 14148 15997
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 15200 16031 15252 16040
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15200 15988 15252 15997
rect 11336 15920 11388 15972
rect 17132 15920 17184 15972
rect 32588 16124 32640 16176
rect 20812 16056 20864 16108
rect 20996 16031 21048 16040
rect 20996 15997 21005 16031
rect 21005 15997 21039 16031
rect 21039 15997 21048 16031
rect 20996 15988 21048 15997
rect 22008 16056 22060 16108
rect 21640 15988 21692 16040
rect 21916 16031 21968 16040
rect 21916 15997 21925 16031
rect 21925 15997 21959 16031
rect 21959 15997 21968 16031
rect 21916 15988 21968 15997
rect 20536 15963 20588 15972
rect 20536 15929 20545 15963
rect 20545 15929 20579 15963
rect 20579 15929 20588 15963
rect 20536 15920 20588 15929
rect 22008 15920 22060 15972
rect 22560 15988 22612 16040
rect 23664 16031 23716 16040
rect 23664 15997 23673 16031
rect 23673 15997 23707 16031
rect 23707 15997 23716 16031
rect 23664 15988 23716 15997
rect 20812 15895 20864 15904
rect 20812 15861 20821 15895
rect 20821 15861 20855 15895
rect 20855 15861 20864 15895
rect 20812 15852 20864 15861
rect 22100 15852 22152 15904
rect 22928 15852 22980 15904
rect 27528 15895 27580 15904
rect 27528 15861 27537 15895
rect 27537 15861 27571 15895
rect 27571 15861 27580 15895
rect 27528 15852 27580 15861
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 4068 15648 4120 15700
rect 5540 15648 5592 15700
rect 6368 15691 6420 15700
rect 6368 15657 6377 15691
rect 6377 15657 6411 15691
rect 6411 15657 6420 15691
rect 8760 15691 8812 15700
rect 6368 15648 6420 15657
rect 4712 15512 4764 15564
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 6736 15623 6788 15632
rect 6736 15589 6745 15623
rect 6745 15589 6779 15623
rect 6779 15589 6788 15623
rect 6736 15580 6788 15589
rect 2596 15444 2648 15496
rect 4252 15444 4304 15496
rect 4528 15444 4580 15496
rect 9864 15512 9916 15564
rect 11428 15648 11480 15700
rect 12716 15691 12768 15700
rect 12716 15657 12725 15691
rect 12725 15657 12759 15691
rect 12759 15657 12768 15691
rect 12716 15648 12768 15657
rect 14372 15648 14424 15700
rect 13636 15623 13688 15632
rect 13636 15589 13645 15623
rect 13645 15589 13679 15623
rect 13679 15589 13688 15623
rect 13636 15580 13688 15589
rect 12440 15512 12492 15564
rect 13820 15555 13872 15564
rect 13820 15521 13826 15555
rect 13826 15521 13872 15555
rect 13820 15512 13872 15521
rect 6184 15376 6236 15428
rect 11336 15376 11388 15428
rect 13544 15444 13596 15496
rect 14464 15444 14516 15496
rect 15568 15512 15620 15564
rect 16856 15580 16908 15632
rect 16028 15555 16080 15564
rect 16028 15521 16037 15555
rect 16037 15521 16071 15555
rect 16071 15521 16080 15555
rect 16028 15512 16080 15521
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 17132 15648 17184 15700
rect 21088 15648 21140 15700
rect 22008 15648 22060 15700
rect 24124 15648 24176 15700
rect 26240 15691 26292 15700
rect 21640 15580 21692 15632
rect 17960 15512 18012 15564
rect 21824 15555 21876 15564
rect 21824 15521 21833 15555
rect 21833 15521 21867 15555
rect 21867 15521 21876 15555
rect 21824 15512 21876 15521
rect 22560 15555 22612 15564
rect 22560 15521 22569 15555
rect 22569 15521 22603 15555
rect 22603 15521 22612 15555
rect 22560 15512 22612 15521
rect 23296 15444 23348 15496
rect 15200 15376 15252 15428
rect 26240 15657 26249 15691
rect 26249 15657 26283 15691
rect 26283 15657 26292 15691
rect 26240 15648 26292 15657
rect 27528 15580 27580 15632
rect 32404 15580 32456 15632
rect 26792 15555 26844 15564
rect 26792 15521 26801 15555
rect 26801 15521 26835 15555
rect 26835 15521 26844 15555
rect 26792 15512 26844 15521
rect 24860 15376 24912 15428
rect 7932 15308 7984 15360
rect 14188 15308 14240 15360
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 25688 15308 25740 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 58440 15172 58492 15224
rect 59360 15172 59412 15224
rect 4896 15104 4948 15156
rect 25504 15104 25556 15156
rect 3792 15036 3844 15088
rect 4620 15079 4672 15088
rect 4620 15045 4629 15079
rect 4629 15045 4663 15079
rect 4663 15045 4672 15079
rect 4620 15036 4672 15045
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 8760 15036 8812 15088
rect 19340 14968 19392 15020
rect 20720 14968 20772 15020
rect 21732 14968 21784 15020
rect 24768 14968 24820 15020
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 12992 14900 13044 14952
rect 13912 14900 13964 14952
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 15660 14900 15712 14952
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 10968 14764 11020 14816
rect 12716 14764 12768 14816
rect 13544 14764 13596 14816
rect 14188 14764 14240 14816
rect 14924 14764 14976 14816
rect 15016 14764 15068 14816
rect 16672 14764 16724 14816
rect 17868 14764 17920 14816
rect 25688 14943 25740 14952
rect 25688 14909 25697 14943
rect 25697 14909 25731 14943
rect 25731 14909 25740 14943
rect 25688 14900 25740 14909
rect 29092 14900 29144 14952
rect 26792 14875 26844 14884
rect 26792 14841 26801 14875
rect 26801 14841 26835 14875
rect 26835 14841 26844 14875
rect 26792 14832 26844 14841
rect 86224 14832 86276 14884
rect 87144 14832 87196 14884
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 9496 14560 9548 14612
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 14372 14560 14424 14612
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 12624 14424 12676 14476
rect 13912 14467 13964 14476
rect 13912 14433 13921 14467
rect 13921 14433 13955 14467
rect 13955 14433 13964 14467
rect 13912 14424 13964 14433
rect 14464 14424 14516 14476
rect 16212 14560 16264 14612
rect 20720 14560 20772 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 26240 14603 26292 14612
rect 26240 14569 26249 14603
rect 26249 14569 26283 14603
rect 26283 14569 26292 14603
rect 26240 14560 26292 14569
rect 22928 14492 22980 14544
rect 29092 14492 29144 14544
rect 13820 14399 13872 14408
rect 13820 14365 13829 14399
rect 13829 14365 13863 14399
rect 13863 14365 13872 14399
rect 13820 14356 13872 14365
rect 21456 14356 21508 14408
rect 22008 14356 22060 14408
rect 8116 14331 8168 14340
rect 8116 14297 8125 14331
rect 8125 14297 8159 14331
rect 8159 14297 8168 14331
rect 8116 14288 8168 14297
rect 16948 14288 17000 14340
rect 7012 14220 7064 14272
rect 12532 14220 12584 14272
rect 19064 14220 19116 14272
rect 26792 14467 26844 14476
rect 26792 14433 26801 14467
rect 26801 14433 26835 14467
rect 26835 14433 26844 14467
rect 26792 14424 26844 14433
rect 24032 14220 24084 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 4804 14016 4856 14068
rect 8208 14016 8260 14068
rect 16948 14016 17000 14068
rect 19340 14059 19392 14068
rect 19340 14025 19349 14059
rect 19349 14025 19383 14059
rect 19383 14025 19392 14059
rect 19340 14016 19392 14025
rect 4620 13991 4672 14000
rect 4620 13957 4629 13991
rect 4629 13957 4663 13991
rect 4663 13957 4672 13991
rect 4620 13948 4672 13957
rect 12716 13948 12768 14000
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 15016 13923 15068 13932
rect 10968 13812 11020 13864
rect 15016 13889 15025 13923
rect 15025 13889 15059 13923
rect 15059 13889 15068 13923
rect 15016 13880 15068 13889
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 18788 13948 18840 14000
rect 17776 13812 17828 13821
rect 19064 13855 19116 13864
rect 16672 13744 16724 13796
rect 16764 13744 16816 13796
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19064 13812 19116 13821
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 4068 13676 4120 13728
rect 19156 13676 19208 13728
rect 21364 13855 21416 13864
rect 21364 13821 21373 13855
rect 21373 13821 21407 13855
rect 21407 13821 21416 13855
rect 21364 13812 21416 13821
rect 24032 13923 24084 13932
rect 24032 13889 24041 13923
rect 24041 13889 24075 13923
rect 24075 13889 24084 13923
rect 24032 13880 24084 13889
rect 22008 13744 22060 13796
rect 28080 13812 28132 13864
rect 29000 13812 29052 13864
rect 22652 13787 22704 13796
rect 22652 13753 22661 13787
rect 22661 13753 22695 13787
rect 22695 13753 22704 13787
rect 22652 13744 22704 13753
rect 27712 13719 27764 13728
rect 27712 13685 27721 13719
rect 27721 13685 27755 13719
rect 27755 13685 27764 13719
rect 27712 13676 27764 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 7840 13472 7892 13524
rect 6828 13404 6880 13456
rect 11612 13472 11664 13524
rect 12992 13472 13044 13524
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 5724 13336 5776 13345
rect 7196 13336 7248 13388
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 7932 13336 7984 13388
rect 10968 13379 11020 13388
rect 10968 13345 10977 13379
rect 10977 13345 11011 13379
rect 11011 13345 11020 13379
rect 10968 13336 11020 13345
rect 20812 13472 20864 13524
rect 21364 13472 21416 13524
rect 25228 13472 25280 13524
rect 16672 13447 16724 13456
rect 16672 13413 16681 13447
rect 16681 13413 16715 13447
rect 16715 13413 16724 13447
rect 16672 13404 16724 13413
rect 19340 13404 19392 13456
rect 20536 13404 20588 13456
rect 24032 13447 24084 13456
rect 24032 13413 24041 13447
rect 24041 13413 24075 13447
rect 24075 13413 24084 13447
rect 24032 13404 24084 13413
rect 22652 13379 22704 13388
rect 22652 13345 22661 13379
rect 22661 13345 22695 13379
rect 22695 13345 22704 13379
rect 22652 13336 22704 13345
rect 25136 13336 25188 13388
rect 25688 13336 25740 13388
rect 27712 13336 27764 13388
rect 3700 13132 3752 13184
rect 6920 13268 6972 13320
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 14280 13268 14332 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 22376 13311 22428 13320
rect 22376 13277 22385 13311
rect 22385 13277 22419 13311
rect 22419 13277 22428 13311
rect 22376 13268 22428 13277
rect 23388 13268 23440 13320
rect 26240 13200 26292 13252
rect 8852 13132 8904 13184
rect 12256 13132 12308 13184
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 26792 13132 26844 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 5448 12928 5500 12980
rect 6552 12792 6604 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 5724 12724 5776 12776
rect 7472 12860 7524 12912
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 8852 12724 8904 12776
rect 11244 12903 11296 12912
rect 11244 12869 11253 12903
rect 11253 12869 11287 12903
rect 11287 12869 11296 12903
rect 11244 12860 11296 12869
rect 10876 12767 10928 12776
rect 10876 12733 10885 12767
rect 10885 12733 10919 12767
rect 10919 12733 10928 12767
rect 10876 12724 10928 12733
rect 11980 12724 12032 12776
rect 12532 12724 12584 12776
rect 19340 12928 19392 12980
rect 21180 12792 21232 12844
rect 21548 12928 21600 12980
rect 24860 12928 24912 12980
rect 26240 12928 26292 12980
rect 28080 12971 28132 12980
rect 28080 12937 28089 12971
rect 28089 12937 28123 12971
rect 28123 12937 28132 12971
rect 28080 12928 28132 12937
rect 26516 12835 26568 12844
rect 26516 12801 26525 12835
rect 26525 12801 26559 12835
rect 26559 12801 26568 12835
rect 26516 12792 26568 12801
rect 26792 12835 26844 12844
rect 26792 12801 26801 12835
rect 26801 12801 26835 12835
rect 26835 12801 26844 12835
rect 26792 12792 26844 12801
rect 22284 12767 22336 12776
rect 12900 12656 12952 12708
rect 22008 12656 22060 12708
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 23388 12724 23440 12776
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 4160 12588 4212 12597
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 8024 12631 8076 12640
rect 8024 12597 8033 12631
rect 8033 12597 8067 12631
rect 8067 12597 8076 12631
rect 8024 12588 8076 12597
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 10876 12588 10928 12640
rect 12532 12588 12584 12640
rect 17040 12588 17092 12640
rect 18144 12631 18196 12640
rect 18144 12597 18153 12631
rect 18153 12597 18187 12631
rect 18187 12597 18196 12631
rect 18144 12588 18196 12597
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 8852 12384 8904 12436
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 4068 12248 4120 12300
rect 12624 12316 12676 12368
rect 17132 12384 17184 12436
rect 22284 12384 22336 12436
rect 21180 12316 21232 12368
rect 12992 12248 13044 12300
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 14372 12248 14424 12300
rect 16672 12248 16724 12300
rect 17040 12291 17092 12300
rect 17040 12257 17049 12291
rect 17049 12257 17083 12291
rect 17083 12257 17092 12291
rect 17040 12248 17092 12257
rect 18144 12248 18196 12300
rect 24860 12384 24912 12436
rect 4620 12044 4672 12096
rect 8024 12180 8076 12232
rect 12532 12180 12584 12232
rect 12624 12112 12676 12164
rect 22100 12112 22152 12164
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 12900 12044 12952 12053
rect 13452 12044 13504 12096
rect 21272 12044 21324 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 6920 11840 6972 11892
rect 8208 11840 8260 11892
rect 3976 11772 4028 11824
rect 12532 11840 12584 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 12900 11840 12952 11892
rect 15016 11840 15068 11892
rect 20720 11840 20772 11892
rect 21732 11840 21784 11892
rect 29644 11840 29696 11892
rect 2596 11679 2648 11688
rect 2596 11645 2605 11679
rect 2605 11645 2639 11679
rect 2639 11645 2648 11679
rect 2596 11636 2648 11645
rect 6920 11679 6972 11688
rect 6920 11645 6929 11679
rect 6929 11645 6963 11679
rect 6963 11645 6972 11679
rect 6920 11636 6972 11645
rect 7932 11636 7984 11688
rect 10600 11636 10652 11688
rect 15384 11636 15436 11688
rect 20720 11636 20772 11688
rect 22376 11636 22428 11688
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 24400 11636 24452 11688
rect 8116 11568 8168 11620
rect 14096 11568 14148 11620
rect 14556 11611 14608 11620
rect 14556 11577 14565 11611
rect 14565 11577 14599 11611
rect 14599 11577 14608 11611
rect 14556 11568 14608 11577
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 4620 11500 4672 11552
rect 5540 11500 5592 11552
rect 11336 11500 11388 11552
rect 18604 11500 18656 11552
rect 26240 11543 26292 11552
rect 26240 11509 26249 11543
rect 26249 11509 26283 11543
rect 26283 11509 26292 11543
rect 26240 11500 26292 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 5540 11296 5592 11348
rect 10692 11296 10744 11348
rect 12716 11296 12768 11348
rect 13820 11296 13872 11348
rect 14464 11296 14516 11348
rect 15384 11339 15436 11348
rect 15384 11305 15393 11339
rect 15393 11305 15427 11339
rect 15427 11305 15436 11339
rect 15384 11296 15436 11305
rect 21088 11296 21140 11348
rect 9128 11228 9180 11280
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 12624 11160 12676 11212
rect 14556 11160 14608 11212
rect 18604 11203 18656 11212
rect 2964 11024 3016 11076
rect 8024 11092 8076 11144
rect 13820 11092 13872 11144
rect 16212 11135 16264 11144
rect 15292 11024 15344 11076
rect 16212 11101 16221 11135
rect 16221 11101 16255 11135
rect 16255 11101 16264 11135
rect 16212 11092 16264 11101
rect 17960 11092 18012 11144
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 21088 11092 21140 11144
rect 22284 11135 22336 11144
rect 22284 11101 22293 11135
rect 22293 11101 22327 11135
rect 22327 11101 22336 11135
rect 22284 11092 22336 11101
rect 6828 10956 6880 11008
rect 17776 10956 17828 11008
rect 23572 10999 23624 11008
rect 23572 10965 23581 10999
rect 23581 10965 23615 10999
rect 23615 10965 23624 10999
rect 23572 10956 23624 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 3976 10752 4028 10804
rect 6828 10752 6880 10804
rect 7932 10752 7984 10804
rect 2596 10591 2648 10600
rect 2596 10557 2605 10591
rect 2605 10557 2639 10591
rect 2639 10557 2648 10591
rect 2596 10548 2648 10557
rect 15200 10752 15252 10804
rect 22284 10752 22336 10804
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 7564 10523 7616 10532
rect 7564 10489 7573 10523
rect 7573 10489 7607 10523
rect 7607 10489 7616 10523
rect 7564 10480 7616 10489
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 4620 10412 4672 10464
rect 23572 10616 23624 10668
rect 26240 10616 26292 10668
rect 16212 10548 16264 10600
rect 21088 10591 21140 10600
rect 21088 10557 21097 10591
rect 21097 10557 21131 10591
rect 21131 10557 21140 10591
rect 21088 10548 21140 10557
rect 21364 10591 21416 10600
rect 21364 10557 21373 10591
rect 21373 10557 21407 10591
rect 21407 10557 21416 10591
rect 21364 10548 21416 10557
rect 26516 10548 26568 10600
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 16488 10412 16540 10464
rect 26792 10412 26844 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 7564 10208 7616 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 6828 10072 6880 10124
rect 8300 10072 8352 10124
rect 15016 10251 15068 10260
rect 6920 10004 6972 10056
rect 12532 10004 12584 10056
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 16396 10208 16448 10260
rect 21364 10208 21416 10260
rect 21732 10251 21784 10260
rect 21732 10217 21741 10251
rect 21741 10217 21775 10251
rect 21775 10217 21784 10251
rect 21732 10208 21784 10217
rect 20628 10140 20680 10192
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 7380 9868 7432 9920
rect 11060 9868 11112 9920
rect 27896 9911 27948 9920
rect 27896 9877 27905 9911
rect 27905 9877 27939 9911
rect 27939 9877 27948 9911
rect 27896 9868 27948 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 9128 9707 9180 9716
rect 9128 9673 9137 9707
rect 9137 9673 9171 9707
rect 9171 9673 9180 9707
rect 9128 9664 9180 9673
rect 11336 9664 11388 9716
rect 8024 9596 8076 9648
rect 13360 9596 13412 9648
rect 20812 9596 20864 9648
rect 24400 9639 24452 9648
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7380 9528 7432 9580
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 4620 9460 4672 9512
rect 6828 9460 6880 9512
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 15200 9528 15252 9580
rect 15568 9528 15620 9580
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 16212 9528 16264 9580
rect 21364 9528 21416 9580
rect 8300 9392 8352 9444
rect 12624 9435 12676 9444
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 10508 9324 10560 9376
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 16396 9460 16448 9512
rect 23204 9460 23256 9512
rect 24400 9605 24409 9639
rect 24409 9605 24443 9639
rect 24443 9605 24452 9639
rect 24400 9596 24452 9605
rect 26516 9664 26568 9716
rect 27896 9528 27948 9580
rect 16856 9392 16908 9444
rect 12440 9324 12492 9376
rect 13452 9324 13504 9376
rect 22284 9367 22336 9376
rect 22284 9333 22293 9367
rect 22293 9333 22327 9367
rect 22327 9333 22336 9367
rect 22284 9324 22336 9333
rect 27712 9367 27764 9376
rect 27712 9333 27721 9367
rect 27721 9333 27755 9367
rect 27755 9333 27764 9367
rect 27712 9324 27764 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 12624 9120 12676 9172
rect 16212 9120 16264 9172
rect 10508 8984 10560 9036
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 12348 9052 12400 9104
rect 13452 9095 13504 9104
rect 12256 8984 12308 9036
rect 13452 9061 13461 9095
rect 13461 9061 13495 9095
rect 13495 9061 13504 9095
rect 13452 9052 13504 9061
rect 16580 9052 16632 9104
rect 15200 8984 15252 9036
rect 27712 9120 27764 9172
rect 18696 9052 18748 9104
rect 12624 8848 12676 8900
rect 24400 8984 24452 9036
rect 13360 8848 13412 8900
rect 4068 8780 4120 8832
rect 14188 8780 14240 8832
rect 18052 8916 18104 8968
rect 23112 8959 23164 8968
rect 23112 8925 23121 8959
rect 23121 8925 23155 8959
rect 23155 8925 23164 8959
rect 23112 8916 23164 8925
rect 23204 8916 23256 8968
rect 16764 8780 16816 8832
rect 17868 8780 17920 8832
rect 22100 8823 22152 8832
rect 22100 8789 22109 8823
rect 22109 8789 22143 8823
rect 22143 8789 22152 8823
rect 22744 8823 22796 8832
rect 22100 8780 22152 8789
rect 22744 8789 22753 8823
rect 22753 8789 22787 8823
rect 22787 8789 22796 8823
rect 22744 8780 22796 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 7472 8576 7524 8628
rect 3332 8440 3384 8492
rect 10968 8508 11020 8560
rect 2596 8415 2648 8424
rect 2596 8381 2605 8415
rect 2605 8381 2639 8415
rect 2639 8381 2648 8415
rect 2596 8372 2648 8381
rect 9036 8440 9088 8492
rect 12532 8576 12584 8628
rect 7656 8372 7708 8424
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 10968 8372 11020 8424
rect 12348 8440 12400 8492
rect 16488 8576 16540 8628
rect 17132 8576 17184 8628
rect 17868 8576 17920 8628
rect 16120 8440 16172 8492
rect 18052 8483 18104 8492
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 22100 8576 22152 8628
rect 23112 8576 23164 8628
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12624 8415 12676 8424
rect 12440 8372 12492 8381
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 16580 8415 16632 8424
rect 16580 8381 16589 8415
rect 16589 8381 16623 8415
rect 16623 8381 16632 8415
rect 16580 8372 16632 8381
rect 16948 8415 17000 8424
rect 16948 8381 16962 8415
rect 16962 8381 17000 8415
rect 16948 8372 17000 8381
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 18696 8415 18748 8424
rect 17132 8372 17184 8381
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 22284 8440 22336 8492
rect 20536 8304 20588 8356
rect 22744 8304 22796 8356
rect 23572 8304 23624 8356
rect 4160 8236 4212 8288
rect 4804 8236 4856 8288
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 16672 8032 16724 8084
rect 20536 8032 20588 8084
rect 7288 7964 7340 8016
rect 12624 7964 12676 8016
rect 4068 7896 4120 7948
rect 7012 7896 7064 7948
rect 11428 7896 11480 7948
rect 16212 7896 16264 7948
rect 22284 7896 22336 7948
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4620 7828 4672 7880
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 16580 7828 16632 7880
rect 23940 7871 23992 7880
rect 23940 7837 23949 7871
rect 23949 7837 23983 7871
rect 23983 7837 23992 7871
rect 23940 7828 23992 7837
rect 6000 7735 6052 7744
rect 6000 7701 6009 7735
rect 6009 7701 6043 7735
rect 6043 7701 6052 7735
rect 6000 7692 6052 7701
rect 6828 7692 6880 7744
rect 7656 7692 7708 7744
rect 12808 7692 12860 7744
rect 22836 7692 22888 7744
rect 23572 7735 23624 7744
rect 23572 7701 23581 7735
rect 23581 7701 23615 7735
rect 23615 7701 23624 7735
rect 23572 7692 23624 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 4620 7531 4672 7540
rect 4620 7497 4629 7531
rect 4629 7497 4663 7531
rect 4663 7497 4672 7531
rect 4620 7488 4672 7497
rect 4804 7488 4856 7540
rect 6000 7488 6052 7540
rect 10968 7488 11020 7540
rect 15016 7488 15068 7540
rect 9404 7463 9456 7472
rect 9404 7429 9413 7463
rect 9413 7429 9447 7463
rect 9447 7429 9456 7463
rect 9404 7420 9456 7429
rect 9864 7420 9916 7472
rect 4804 7352 4856 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 22836 7352 22888 7404
rect 4712 7284 4764 7336
rect 8392 7284 8444 7336
rect 13820 7216 13872 7268
rect 16948 7148 17000 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 12256 6944 12308 6996
rect 12808 6944 12860 6996
rect 15016 6944 15068 6996
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 9864 6808 9916 6860
rect 10876 6808 10928 6860
rect 11704 6808 11756 6860
rect 16580 6808 16632 6860
rect 23940 6987 23992 6996
rect 23940 6953 23949 6987
rect 23949 6953 23983 6987
rect 23983 6953 23992 6987
rect 23940 6944 23992 6953
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 22836 6851 22888 6860
rect 22836 6817 22845 6851
rect 22845 6817 22879 6851
rect 22879 6817 22888 6851
rect 22836 6808 22888 6817
rect 10232 6740 10284 6792
rect 10968 6740 11020 6792
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 17040 6740 17092 6792
rect 23572 6740 23624 6792
rect 7104 6672 7156 6724
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 4804 6400 4856 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 11612 6400 11664 6452
rect 11704 6443 11756 6452
rect 11704 6409 11713 6443
rect 11713 6409 11747 6443
rect 11747 6409 11756 6443
rect 11704 6400 11756 6409
rect 10968 6332 11020 6384
rect 7104 6307 7156 6316
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 10232 6264 10284 6316
rect 13820 6264 13872 6316
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 13176 6060 13228 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 7748 5652 7800 5704
rect 23572 5584 23624 5636
rect 29920 5516 29972 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 4804 5312 4856 5364
rect 2964 5176 3016 5228
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 3240 5108 3292 5160
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 4068 4768 4120 4820
rect 6552 4768 6604 4820
rect 6828 4768 6880 4820
rect 8116 4564 8168 4616
rect 5080 4428 5132 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 4804 4267 4856 4276
rect 4804 4233 4813 4267
rect 4813 4233 4847 4267
rect 4847 4233 4856 4267
rect 4804 4224 4856 4233
rect 6184 4088 6236 4140
rect 27160 4088 27212 4140
rect 28080 4088 28132 4140
rect 3240 4020 3292 4072
rect 4068 3952 4120 4004
rect 7564 3952 7616 4004
rect 4160 3884 4212 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 3976 3476 4028 3528
rect 5080 3476 5132 3528
rect 56324 3408 56376 3460
rect 84200 3408 84252 3460
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 4988 3136 5040 3188
rect 3240 2932 3292 2984
rect 4804 2932 4856 2984
rect 2780 2796 2832 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
<< metal2 >>
rect 4066 45928 4122 45937
rect 4066 45863 4122 45872
rect 2410 45384 2466 45393
rect 2410 45319 2466 45328
rect 2424 42362 2452 45319
rect 4080 44198 4108 45863
rect 56138 45440 56194 46240
rect 7654 44704 7710 44713
rect 7654 44639 7710 44648
rect 4068 44192 4120 44198
rect 4068 44134 4120 44140
rect 6276 43920 6328 43926
rect 6276 43862 6328 43868
rect 4620 43716 4672 43722
rect 4620 43658 4672 43664
rect 5540 43716 5592 43722
rect 5540 43658 5592 43664
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 2412 42356 2464 42362
rect 2412 42298 2464 42304
rect 2424 42158 2452 42298
rect 2412 42152 2464 42158
rect 2412 42094 2464 42100
rect 2872 42152 2924 42158
rect 2872 42094 2924 42100
rect 2596 38888 2648 38894
rect 2596 38830 2648 38836
rect 2608 37874 2636 38830
rect 2884 38706 2912 42094
rect 3976 42016 4028 42022
rect 3976 41958 4028 41964
rect 3988 41721 4016 41958
rect 3974 41712 4030 41721
rect 4632 41682 4660 43658
rect 4804 43308 4856 43314
rect 4804 43250 4856 43256
rect 4816 43178 4844 43250
rect 5080 43240 5132 43246
rect 5080 43182 5132 43188
rect 4804 43172 4856 43178
rect 4804 43114 4856 43120
rect 4816 42770 4844 43114
rect 4804 42764 4856 42770
rect 4804 42706 4856 42712
rect 4816 42362 4844 42706
rect 4804 42356 4856 42362
rect 4804 42298 4856 42304
rect 5092 41818 5120 43182
rect 5264 43104 5316 43110
rect 5264 43046 5316 43052
rect 5276 42158 5304 43046
rect 5552 42770 5580 43658
rect 5540 42764 5592 42770
rect 5540 42706 5592 42712
rect 6288 42294 6316 43862
rect 6920 43648 6972 43654
rect 6920 43590 6972 43596
rect 6460 43240 6512 43246
rect 6460 43182 6512 43188
rect 6472 42838 6500 43182
rect 6644 43172 6696 43178
rect 6644 43114 6696 43120
rect 6656 42906 6684 43114
rect 6932 43110 6960 43590
rect 6920 43104 6972 43110
rect 6920 43046 6972 43052
rect 6644 42900 6696 42906
rect 6644 42842 6696 42848
rect 6460 42832 6512 42838
rect 6460 42774 6512 42780
rect 6920 42560 6972 42566
rect 6920 42502 6972 42508
rect 6276 42288 6328 42294
rect 6276 42230 6328 42236
rect 6092 42220 6144 42226
rect 6092 42162 6144 42168
rect 5264 42152 5316 42158
rect 5264 42094 5316 42100
rect 5172 42016 5224 42022
rect 5172 41958 5224 41964
rect 5080 41812 5132 41818
rect 5080 41754 5132 41760
rect 5184 41682 5212 41958
rect 3974 41647 4030 41656
rect 4620 41676 4672 41682
rect 4620 41618 4672 41624
rect 5172 41676 5224 41682
rect 5172 41618 5224 41624
rect 4632 41562 4660 41618
rect 5356 41608 5408 41614
rect 4632 41534 4936 41562
rect 5356 41550 5408 41556
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 3608 41064 3660 41070
rect 3608 41006 3660 41012
rect 3884 41064 3936 41070
rect 3884 41006 3936 41012
rect 3422 40488 3478 40497
rect 3422 40423 3478 40432
rect 2884 38678 3004 38706
rect 2596 37868 2648 37874
rect 2596 37810 2648 37816
rect 2872 35012 2924 35018
rect 2872 34954 2924 34960
rect 2884 31346 2912 34954
rect 2872 31340 2924 31346
rect 2872 31282 2924 31288
rect 2976 30938 3004 38678
rect 3330 36136 3386 36145
rect 3330 36071 3386 36080
rect 3240 33108 3292 33114
rect 3240 33050 3292 33056
rect 3252 32745 3280 33050
rect 3238 32736 3294 32745
rect 3238 32671 3294 32680
rect 2964 30932 3016 30938
rect 2964 30874 3016 30880
rect 2780 30796 2832 30802
rect 2780 30738 2832 30744
rect 2688 30184 2740 30190
rect 2688 30126 2740 30132
rect 2700 29714 2728 30126
rect 2688 29708 2740 29714
rect 2688 29650 2740 29656
rect 2596 28008 2648 28014
rect 2596 27950 2648 27956
rect 2608 26994 2636 27950
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2792 26330 2820 30738
rect 3148 30320 3200 30326
rect 3148 30262 3200 30268
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 2872 27464 2924 27470
rect 2872 27406 2924 27412
rect 2884 26994 2912 27406
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2700 26302 2820 26330
rect 2700 25922 2728 26302
rect 2700 25894 2820 25922
rect 2596 25832 2648 25838
rect 2596 25774 2648 25780
rect 2608 24750 2636 25774
rect 2596 24744 2648 24750
rect 2596 24686 2648 24692
rect 2608 23662 2636 24686
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2608 22574 2636 23598
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2608 21486 2636 22510
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 2608 20602 2636 21422
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2792 20058 2820 25894
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2884 20097 2912 22374
rect 2870 20088 2926 20097
rect 2780 20052 2832 20058
rect 2870 20023 2926 20032
rect 2780 19994 2832 20000
rect 2976 19394 3004 29582
rect 3056 29572 3108 29578
rect 3056 29514 3108 29520
rect 2884 19366 3004 19394
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2608 19174 2636 19246
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2608 16114 2636 19110
rect 2884 16114 2912 19366
rect 2964 19304 3016 19310
rect 3068 19292 3096 29514
rect 3160 20398 3188 30262
rect 3344 29850 3372 36071
rect 3332 29844 3384 29850
rect 3332 29786 3384 29792
rect 3436 24698 3464 40423
rect 3620 39302 3648 41006
rect 3896 40934 3924 41006
rect 4620 40996 4672 41002
rect 4620 40938 4672 40944
rect 3884 40928 3936 40934
rect 3884 40870 3936 40876
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4632 40050 4660 40938
rect 4712 40588 4764 40594
rect 4712 40530 4764 40536
rect 4724 40118 4752 40530
rect 4712 40112 4764 40118
rect 4712 40054 4764 40060
rect 4620 40044 4672 40050
rect 4620 39986 4672 39992
rect 4066 39944 4122 39953
rect 4066 39879 4068 39888
rect 4120 39879 4122 39888
rect 4068 39850 4120 39856
rect 3974 39400 4030 39409
rect 3974 39335 4030 39344
rect 3608 39296 3660 39302
rect 3608 39238 3660 39244
rect 3516 37256 3568 37262
rect 3516 37198 3568 37204
rect 3528 36281 3556 37198
rect 3514 36272 3570 36281
rect 3514 36207 3570 36216
rect 3516 31748 3568 31754
rect 3516 31690 3568 31696
rect 3528 27985 3556 31690
rect 3620 30297 3648 39238
rect 3792 39092 3844 39098
rect 3792 39034 3844 39040
rect 3700 38548 3752 38554
rect 3700 38490 3752 38496
rect 3712 37505 3740 38490
rect 3698 37496 3754 37505
rect 3698 37431 3754 37440
rect 3700 35624 3752 35630
rect 3700 35566 3752 35572
rect 3712 34542 3740 35566
rect 3700 34536 3752 34542
rect 3700 34478 3752 34484
rect 3700 33992 3752 33998
rect 3700 33934 3752 33940
rect 3606 30288 3662 30297
rect 3606 30223 3662 30232
rect 3712 29866 3740 33934
rect 3804 31521 3832 39034
rect 3988 38010 4016 39335
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4068 39024 4120 39030
rect 4068 38966 4120 38972
rect 4080 38729 4108 38966
rect 4160 38752 4212 38758
rect 4066 38720 4122 38729
rect 4160 38694 4212 38700
rect 4436 38752 4488 38758
rect 4436 38694 4488 38700
rect 4066 38655 4122 38664
rect 4172 38196 4200 38694
rect 4448 38418 4476 38694
rect 4436 38412 4488 38418
rect 4436 38354 4488 38360
rect 4620 38344 4672 38350
rect 4620 38286 4672 38292
rect 4080 38185 4200 38196
rect 4066 38176 4200 38185
rect 4122 38168 4200 38176
rect 4066 38111 4122 38120
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 3976 38004 4028 38010
rect 3976 37946 4028 37952
rect 3884 37936 3936 37942
rect 3884 37878 3936 37884
rect 3790 31512 3846 31521
rect 3790 31447 3846 31456
rect 3792 30116 3844 30122
rect 3792 30058 3844 30064
rect 3620 29838 3740 29866
rect 3620 28082 3648 29838
rect 3700 29708 3752 29714
rect 3700 29650 3752 29656
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3514 27976 3570 27985
rect 3514 27911 3570 27920
rect 3608 27940 3660 27946
rect 3608 27882 3660 27888
rect 3516 27396 3568 27402
rect 3516 27338 3568 27344
rect 3528 26761 3556 27338
rect 3514 26752 3570 26761
rect 3514 26687 3570 26696
rect 3516 26240 3568 26246
rect 3516 26182 3568 26188
rect 3528 26081 3556 26182
rect 3514 26072 3570 26081
rect 3514 26007 3570 26016
rect 3620 24818 3648 27882
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 3436 24670 3648 24698
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3344 22545 3372 23054
rect 3330 22536 3386 22545
rect 3330 22471 3386 22480
rect 3620 21690 3648 24670
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3016 19264 3096 19292
rect 2964 19246 3016 19252
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2976 17746 3004 18022
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2976 17542 3004 17682
rect 3160 17542 3188 18090
rect 3344 17785 3372 20198
rect 3712 19553 3740 29650
rect 3698 19544 3754 19553
rect 3698 19479 3754 19488
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3436 18329 3464 18634
rect 3422 18320 3478 18329
rect 3422 18255 3478 18264
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3330 17776 3386 17785
rect 3330 17711 3386 17720
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2976 16454 3004 17478
rect 3436 17338 3464 18022
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3436 17134 3464 17274
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2608 15502 2636 16050
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 15026 2636 15438
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2608 13938 2636 14962
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2608 11694 2636 12718
rect 2976 12322 3004 16390
rect 2884 12294 3004 12322
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 10606 2636 11630
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2608 9518 2636 10542
rect 2884 9636 2912 12294
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2700 9608 2912 9636
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 8430 2636 9454
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2608 5166 2636 6190
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2700 2689 2728 9608
rect 2976 5234 3004 11018
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2686 2680 2742 2689
rect 2686 2615 2742 2624
rect 2792 921 2820 2790
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 3068 377 3096 16934
rect 3712 16658 3740 17478
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3712 14906 3740 16594
rect 3804 15094 3832 30058
rect 3896 29714 3924 37878
rect 4528 37868 4580 37874
rect 4528 37810 4580 37816
rect 4540 37670 4568 37810
rect 4632 37670 4660 38286
rect 4712 38208 4764 38214
rect 4712 38150 4764 38156
rect 4528 37664 4580 37670
rect 4528 37606 4580 37612
rect 4620 37664 4672 37670
rect 4620 37606 4672 37612
rect 4540 37210 4568 37606
rect 4068 37188 4120 37194
rect 4540 37182 4660 37210
rect 4724 37194 4752 38150
rect 4804 37324 4856 37330
rect 4804 37266 4856 37272
rect 4068 37130 4120 37136
rect 4080 36961 4108 37130
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4066 36952 4122 36961
rect 4220 36944 4516 36964
rect 4066 36887 4122 36896
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4068 35828 4120 35834
rect 4068 35770 4120 35776
rect 4080 35737 4108 35770
rect 4066 35728 4122 35737
rect 4066 35663 4122 35672
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4172 35034 4200 35430
rect 4080 35006 4200 35034
rect 4080 34513 4108 35006
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4066 34504 4122 34513
rect 4066 34439 4122 34448
rect 3976 34400 4028 34406
rect 3976 34342 4028 34348
rect 3988 33289 4016 34342
rect 4068 34196 4120 34202
rect 4068 34138 4120 34144
rect 4080 33969 4108 34138
rect 4066 33960 4122 33969
rect 4066 33895 4122 33904
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4344 33448 4396 33454
rect 4344 33390 4396 33396
rect 4160 33312 4212 33318
rect 3974 33280 4030 33289
rect 4160 33254 4212 33260
rect 3974 33215 4030 33224
rect 4172 32756 4200 33254
rect 4356 32978 4384 33390
rect 4632 33318 4660 37182
rect 4712 37188 4764 37194
rect 4712 37130 4764 37136
rect 4816 35562 4844 37266
rect 4908 37262 4936 41534
rect 5264 38888 5316 38894
rect 5264 38830 5316 38836
rect 5080 38412 5132 38418
rect 5080 38354 5132 38360
rect 5092 37874 5120 38354
rect 5080 37868 5132 37874
rect 5080 37810 5132 37816
rect 5276 37806 5304 38830
rect 5264 37800 5316 37806
rect 5264 37742 5316 37748
rect 4896 37256 4948 37262
rect 4896 37198 4948 37204
rect 5276 36718 5304 37742
rect 5264 36712 5316 36718
rect 5264 36654 5316 36660
rect 5172 36576 5224 36582
rect 5172 36518 5224 36524
rect 4988 36372 5040 36378
rect 4988 36314 5040 36320
rect 4804 35556 4856 35562
rect 4804 35498 4856 35504
rect 4712 35284 4764 35290
rect 4712 35226 4764 35232
rect 4724 33522 4752 35226
rect 4816 34542 4844 35498
rect 5000 34610 5028 36314
rect 5184 35698 5212 36518
rect 5276 36174 5304 36654
rect 5368 36242 5396 41550
rect 5448 41064 5500 41070
rect 5448 41006 5500 41012
rect 5460 40186 5488 41006
rect 5540 40520 5592 40526
rect 5540 40462 5592 40468
rect 5448 40180 5500 40186
rect 5448 40122 5500 40128
rect 5552 39642 5580 40462
rect 5724 40384 5776 40390
rect 5724 40326 5776 40332
rect 5736 39982 5764 40326
rect 5724 39976 5776 39982
rect 5724 39918 5776 39924
rect 5816 39840 5868 39846
rect 5816 39782 5868 39788
rect 5540 39636 5592 39642
rect 5540 39578 5592 39584
rect 5828 39506 5856 39782
rect 5816 39500 5868 39506
rect 5816 39442 5868 39448
rect 5448 38344 5500 38350
rect 5448 38286 5500 38292
rect 5356 36236 5408 36242
rect 5356 36178 5408 36184
rect 5264 36168 5316 36174
rect 5264 36110 5316 36116
rect 5172 35692 5224 35698
rect 5172 35634 5224 35640
rect 5356 35148 5408 35154
rect 5356 35090 5408 35096
rect 4988 34604 5040 34610
rect 4988 34546 5040 34552
rect 5368 34542 5396 35090
rect 4804 34536 4856 34542
rect 4804 34478 4856 34484
rect 5356 34536 5408 34542
rect 5356 34478 5408 34484
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4344 32972 4396 32978
rect 4344 32914 4396 32920
rect 4080 32728 4200 32756
rect 4356 32756 4384 32914
rect 4356 32728 4660 32756
rect 3976 32224 4028 32230
rect 4080 32201 4108 32728
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 3976 32166 4028 32172
rect 4066 32192 4122 32201
rect 3988 30977 4016 32166
rect 4066 32127 4122 32136
rect 4632 32026 4660 32728
rect 4816 32570 4844 34478
rect 5368 34134 5396 34478
rect 5356 34128 5408 34134
rect 5356 34070 5408 34076
rect 5368 33658 5396 34070
rect 5460 34066 5488 38286
rect 6104 38010 6132 42162
rect 6932 41177 6960 42502
rect 6918 41168 6974 41177
rect 6918 41103 6974 41112
rect 6932 40186 6960 41103
rect 7288 40996 7340 41002
rect 7288 40938 7340 40944
rect 6920 40180 6972 40186
rect 6920 40122 6972 40128
rect 6932 39964 6960 40122
rect 7300 39982 7328 40938
rect 7104 39976 7156 39982
rect 6932 39936 7104 39964
rect 7104 39918 7156 39924
rect 7288 39976 7340 39982
rect 7288 39918 7340 39924
rect 6092 38004 6144 38010
rect 6092 37946 6144 37952
rect 6104 37806 6132 37946
rect 6092 37800 6144 37806
rect 6092 37742 6144 37748
rect 5908 37732 5960 37738
rect 5908 37674 5960 37680
rect 5540 36848 5592 36854
rect 5540 36790 5592 36796
rect 5448 34060 5500 34066
rect 5448 34002 5500 34008
rect 5448 33924 5500 33930
rect 5448 33866 5500 33872
rect 5356 33652 5408 33658
rect 5356 33594 5408 33600
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 4908 32774 4936 33254
rect 5356 32904 5408 32910
rect 5356 32846 5408 32852
rect 4896 32768 4948 32774
rect 4896 32710 4948 32716
rect 4804 32564 4856 32570
rect 4804 32506 4856 32512
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4160 31136 4212 31142
rect 4160 31078 4212 31084
rect 3974 30968 4030 30977
rect 3974 30903 4030 30912
rect 3976 30796 4028 30802
rect 3976 30738 4028 30744
rect 3988 30258 4016 30738
rect 4172 30682 4200 31078
rect 4080 30654 4200 30682
rect 3976 30252 4028 30258
rect 3976 30194 4028 30200
rect 4080 29753 4108 30654
rect 4632 30598 4660 31826
rect 4908 31482 4936 32710
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 4896 31476 4948 31482
rect 4896 31418 4948 31424
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4632 30394 4660 30534
rect 4620 30388 4672 30394
rect 4620 30330 4672 30336
rect 4528 30184 4580 30190
rect 4528 30126 4580 30132
rect 4540 30054 4568 30126
rect 4528 30048 4580 30054
rect 4528 29990 4580 29996
rect 4066 29744 4122 29753
rect 3884 29708 3936 29714
rect 4066 29679 4122 29688
rect 3884 29650 3936 29656
rect 4068 29640 4120 29646
rect 4068 29582 4120 29588
rect 3976 29300 4028 29306
rect 3976 29242 4028 29248
rect 3988 29073 4016 29242
rect 4080 29186 4108 29582
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4080 29158 4200 29186
rect 4172 29102 4200 29158
rect 4160 29096 4212 29102
rect 3974 29064 4030 29073
rect 4160 29038 4212 29044
rect 3974 28999 4030 29008
rect 3884 28960 3936 28966
rect 3884 28902 3936 28908
rect 3896 23730 3924 28902
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 4080 28529 4108 28698
rect 4172 28694 4200 29038
rect 4160 28688 4212 28694
rect 4160 28630 4212 28636
rect 4620 28552 4672 28558
rect 4066 28520 4122 28529
rect 4620 28494 4672 28500
rect 4066 28455 4122 28464
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4160 27872 4212 27878
rect 4160 27814 4212 27820
rect 4172 27418 4200 27814
rect 4080 27390 4200 27418
rect 4080 27305 4108 27390
rect 4066 27296 4122 27305
rect 4066 27231 4122 27240
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4252 26920 4304 26926
rect 4252 26862 4304 26868
rect 4160 26784 4212 26790
rect 4160 26726 4212 26732
rect 4172 26330 4200 26726
rect 4264 26382 4292 26862
rect 4632 26450 4660 28494
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 4080 26302 4200 26330
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3988 25537 4016 25978
rect 3974 25528 4030 25537
rect 3974 25463 4030 25472
rect 4080 25378 4108 26302
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4160 25696 4212 25702
rect 4160 25638 4212 25644
rect 3988 25350 4108 25378
rect 3988 24993 4016 25350
rect 4172 25242 4200 25638
rect 4080 25214 4200 25242
rect 3974 24984 4030 24993
rect 3974 24919 4030 24928
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3988 24313 4016 24346
rect 3974 24304 4030 24313
rect 3974 24239 4030 24248
rect 4080 23769 4108 25214
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4066 23760 4122 23769
rect 3884 23724 3936 23730
rect 4066 23695 4122 23704
rect 3884 23666 3936 23672
rect 3976 23520 4028 23526
rect 3976 23462 4028 23468
rect 3988 21321 4016 23462
rect 4632 23118 4660 24618
rect 4620 23112 4672 23118
rect 4066 23080 4122 23089
rect 4620 23054 4672 23060
rect 4066 23015 4122 23024
rect 4080 22778 4108 23015
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4068 21956 4120 21962
rect 4068 21898 4120 21904
rect 4080 21865 4108 21898
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 3974 21312 4030 21321
rect 3974 21247 4030 21256
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4080 20777 4108 20878
rect 4066 20768 4122 20777
rect 4066 20703 4122 20712
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4724 20210 4752 30670
rect 4896 30592 4948 30598
rect 4896 30534 4948 30540
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4816 27878 4844 29582
rect 4804 27872 4856 27878
rect 4804 27814 4856 27820
rect 4816 26926 4844 27814
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4816 21690 4844 22646
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4816 20602 4844 21626
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 4724 20182 4844 20210
rect 4816 19938 4844 20182
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 4724 19910 4844 19938
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3988 18873 4016 19110
rect 4080 18986 4108 19654
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4080 18970 4200 18986
rect 4080 18964 4212 18970
rect 4080 18958 4160 18964
rect 4160 18906 4212 18912
rect 3974 18864 4030 18873
rect 3974 18799 4030 18808
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4632 17882 4660 19858
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4632 17134 4660 17682
rect 4160 17128 4212 17134
rect 4066 17096 4122 17105
rect 4160 17070 4212 17076
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4066 17031 4122 17040
rect 4080 16998 4108 17031
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4172 16794 4200 17070
rect 4264 16794 4292 17070
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4066 16552 4122 16561
rect 3884 16516 3936 16522
rect 4066 16487 4122 16496
rect 3884 16458 3936 16464
rect 3896 15881 3924 16458
rect 3976 15904 4028 15910
rect 3882 15872 3938 15881
rect 3976 15846 4028 15852
rect 3882 15807 3938 15816
rect 3988 15337 4016 15846
rect 4080 15706 4108 16487
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4264 15502 4292 15846
rect 4724 15570 4752 19910
rect 4908 19802 4936 30534
rect 5000 29850 5028 32166
rect 5080 31204 5132 31210
rect 5080 31146 5132 31152
rect 4988 29844 5040 29850
rect 4988 29786 5040 29792
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 5000 28762 5028 29446
rect 4988 28756 5040 28762
rect 4988 28698 5040 28704
rect 5092 27538 5120 31146
rect 5172 30184 5224 30190
rect 5172 30126 5224 30132
rect 5184 29102 5212 30126
rect 5264 29232 5316 29238
rect 5264 29174 5316 29180
rect 5172 29096 5224 29102
rect 5172 29038 5224 29044
rect 5172 28960 5224 28966
rect 5172 28902 5224 28908
rect 5080 27532 5132 27538
rect 5080 27474 5132 27480
rect 5184 22642 5212 28902
rect 5276 28694 5304 29174
rect 5264 28688 5316 28694
rect 5264 28630 5316 28636
rect 5276 28014 5304 28630
rect 5264 28008 5316 28014
rect 5264 27950 5316 27956
rect 5276 27606 5304 27950
rect 5264 27600 5316 27606
rect 5264 27542 5316 27548
rect 5368 22642 5396 32846
rect 5460 28626 5488 33866
rect 5552 30054 5580 36790
rect 5632 35692 5684 35698
rect 5632 35634 5684 35640
rect 5644 35193 5672 35634
rect 5630 35184 5686 35193
rect 5630 35119 5686 35128
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5644 32434 5672 34546
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 5816 32292 5868 32298
rect 5816 32234 5868 32240
rect 5828 31890 5856 32234
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5724 30660 5776 30666
rect 5724 30602 5776 30608
rect 5736 30394 5764 30602
rect 5724 30388 5776 30394
rect 5724 30330 5776 30336
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5448 28620 5500 28626
rect 5448 28562 5500 28568
rect 5920 28422 5948 37674
rect 6920 37664 6972 37670
rect 6920 37606 6972 37612
rect 6932 37330 6960 37606
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 6380 35834 6408 37062
rect 6368 35828 6420 35834
rect 6368 35770 6420 35776
rect 6276 35624 6328 35630
rect 6276 35566 6328 35572
rect 6092 35488 6144 35494
rect 6092 35430 6144 35436
rect 6000 32904 6052 32910
rect 6000 32846 6052 32852
rect 6012 32026 6040 32846
rect 6000 32020 6052 32026
rect 6000 31962 6052 31968
rect 6104 29714 6132 35430
rect 6288 35154 6316 35566
rect 6276 35148 6328 35154
rect 6276 35090 6328 35096
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 6276 32292 6328 32298
rect 6276 32234 6328 32240
rect 6552 32292 6604 32298
rect 6552 32234 6604 32240
rect 6288 31346 6316 32234
rect 6564 31890 6592 32234
rect 7392 31890 7420 32710
rect 6552 31884 6604 31890
rect 6552 31826 6604 31832
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7668 31414 7696 44639
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 50300 44092 50596 44112
rect 50356 44090 50380 44092
rect 50436 44090 50460 44092
rect 50516 44090 50540 44092
rect 50378 44038 50380 44090
rect 50442 44038 50454 44090
rect 50516 44038 50518 44090
rect 50356 44036 50380 44038
rect 50436 44036 50460 44038
rect 50516 44036 50540 44038
rect 50300 44016 50596 44036
rect 40500 43920 40552 43926
rect 40500 43862 40552 43868
rect 19432 43852 19484 43858
rect 19432 43794 19484 43800
rect 24216 43852 24268 43858
rect 24216 43794 24268 43800
rect 25596 43852 25648 43858
rect 25596 43794 25648 43800
rect 39028 43852 39080 43858
rect 39028 43794 39080 43800
rect 17040 43716 17092 43722
rect 17040 43658 17092 43664
rect 10784 43240 10836 43246
rect 10784 43182 10836 43188
rect 9680 43172 9732 43178
rect 9680 43114 9732 43120
rect 8024 43104 8076 43110
rect 8024 43046 8076 43052
rect 8036 42090 8064 43046
rect 9692 42770 9720 43114
rect 9680 42764 9732 42770
rect 9680 42706 9732 42712
rect 10692 42696 10744 42702
rect 10692 42638 10744 42644
rect 9956 42288 10008 42294
rect 9956 42230 10008 42236
rect 8024 42084 8076 42090
rect 8024 42026 8076 42032
rect 9588 42084 9640 42090
rect 9588 42026 9640 42032
rect 8036 41682 8064 42026
rect 9496 42016 9548 42022
rect 9496 41958 9548 41964
rect 9508 41750 9536 41958
rect 9600 41834 9628 42026
rect 9600 41806 9812 41834
rect 9784 41750 9812 41806
rect 8116 41744 8168 41750
rect 8116 41686 8168 41692
rect 9496 41744 9548 41750
rect 9496 41686 9548 41692
rect 9772 41744 9824 41750
rect 9772 41686 9824 41692
rect 8024 41676 8076 41682
rect 8024 41618 8076 41624
rect 8024 40928 8076 40934
rect 8024 40870 8076 40876
rect 7840 39840 7892 39846
rect 7840 39782 7892 39788
rect 7748 32768 7800 32774
rect 7748 32710 7800 32716
rect 7472 31408 7524 31414
rect 7472 31350 7524 31356
rect 7656 31408 7708 31414
rect 7656 31350 7708 31356
rect 6276 31340 6328 31346
rect 6276 31282 6328 31288
rect 6092 29708 6144 29714
rect 6092 29650 6144 29656
rect 5908 28416 5960 28422
rect 5908 28358 5960 28364
rect 5908 26580 5960 26586
rect 5908 26522 5960 26528
rect 5448 25696 5500 25702
rect 5448 25638 5500 25644
rect 5460 25158 5488 25638
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5460 24614 5488 25094
rect 5724 24676 5776 24682
rect 5724 24618 5776 24624
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5460 24274 5488 24550
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 5460 23866 5488 24210
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5460 22710 5488 23802
rect 5736 23662 5764 24618
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 5828 23866 5856 24142
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 4816 19774 4936 19802
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4528 15496 4580 15502
rect 4580 15444 4660 15450
rect 4528 15438 4660 15444
rect 4540 15422 4660 15438
rect 3974 15328 4030 15337
rect 3974 15263 4030 15272
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4632 15094 4660 15422
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 3712 14878 3832 14906
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 6905 3372 8434
rect 3330 6896 3386 6905
rect 3330 6831 3386 6840
rect 3712 6361 3740 13126
rect 3698 6352 3754 6361
rect 3698 6287 3754 6296
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3252 4078 3280 5102
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3252 2990 3280 4014
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3804 1465 3832 14878
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 14113 4016 14758
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 3974 14104 4030 14113
rect 4220 14096 4516 14116
rect 3974 14039 4030 14048
rect 4632 14006 4660 15030
rect 4816 14074 4844 19774
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 4908 17134 4936 19178
rect 5644 18902 5672 19178
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4908 14657 4936 15098
rect 4894 14648 4950 14657
rect 4894 14583 4950 14592
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 3988 12889 4016 13670
rect 4080 13569 4108 13670
rect 4066 13560 4122 13569
rect 4066 13495 4122 13504
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 3974 12880 4030 12889
rect 3974 12815 4030 12824
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4066 12336 4122 12345
rect 4066 12271 4068 12280
rect 4120 12271 4122 12280
rect 4068 12242 4120 12248
rect 4172 12152 4200 12582
rect 4080 12124 4200 12152
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3988 11121 4016 11766
rect 4080 11665 4108 12124
rect 4632 12102 4660 12582
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 4632 11558 4660 12038
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 3974 11112 4030 11121
rect 3974 11047 4030 11056
rect 4172 10996 4200 11494
rect 4080 10968 4200 10996
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3988 9897 4016 10746
rect 4080 10577 4108 10968
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4632 10470 4660 11494
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4172 10010 4200 10406
rect 4080 9982 4200 10010
rect 3974 9888 4030 9897
rect 3974 9823 4030 9832
rect 4080 9353 4108 9982
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4632 9518 4660 10406
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4160 9376 4212 9382
rect 4066 9344 4122 9353
rect 4160 9318 4212 9324
rect 4066 9279 4122 9288
rect 4172 8922 4200 9318
rect 3988 8894 4200 8922
rect 3988 8129 4016 8894
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4080 8673 4108 8774
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4066 8664 4122 8673
rect 4220 8656 4516 8676
rect 4066 8599 4122 8608
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 3974 8120 4030 8129
rect 3974 8055 4030 8064
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4080 7449 4108 7890
rect 4172 7886 4200 8230
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4632 7546 4660 7822
rect 4816 7546 4844 8230
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4066 7440 4122 7449
rect 4816 7410 4844 7482
rect 4066 7375 4122 7384
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4724 6866 4752 7278
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4816 6458 4844 7346
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5681 4016 6054
rect 3974 5672 4030 5681
rect 3974 5607 4030 5616
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4816 5370 4844 6394
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4066 5128 4122 5137
rect 4066 5063 4122 5072
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4457 4016 4966
rect 4080 4826 4108 5063
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3974 4448 4030 4457
rect 3974 4383 4030 4392
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4816 4282 4844 5306
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4080 3913 4108 3946
rect 4160 3936 4212 3942
rect 4066 3904 4122 3913
rect 4160 3878 4212 3884
rect 4066 3839 4122 3848
rect 3976 3528 4028 3534
rect 4172 3482 4200 3878
rect 3976 3470 4028 3476
rect 3988 3369 4016 3470
rect 4080 3454 4200 3482
rect 3974 3360 4030 3369
rect 3974 3295 4030 3304
rect 4080 2145 4108 3454
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4816 2990 4844 4218
rect 5000 3194 5028 18566
rect 5092 18426 5120 18770
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5184 17814 5212 18158
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5092 16046 5120 17614
rect 5184 17066 5212 17750
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5276 16658 5304 18158
rect 5736 18034 5764 22578
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5828 18290 5856 19858
rect 5920 19310 5948 26522
rect 6288 26042 6316 31282
rect 7484 29073 7512 31350
rect 7656 31272 7708 31278
rect 7656 31214 7708 31220
rect 7668 30394 7696 31214
rect 7760 30802 7788 32710
rect 7748 30796 7800 30802
rect 7748 30738 7800 30744
rect 7656 30388 7708 30394
rect 7656 30330 7708 30336
rect 7470 29064 7526 29073
rect 7470 28999 7526 29008
rect 7562 28792 7618 28801
rect 7562 28727 7618 28736
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6840 26586 6868 28358
rect 7576 26790 7604 28727
rect 7656 27872 7708 27878
rect 7656 27814 7708 27820
rect 7564 26784 7616 26790
rect 7564 26726 7616 26732
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7024 25362 7052 25774
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23662 6960 24006
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 5460 18006 5764 18034
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5368 16794 5396 17546
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5460 12986 5488 18006
rect 6288 17746 6316 18158
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6012 16250 6040 17682
rect 6288 17338 6316 17682
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6380 15706 6408 18702
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5552 11558 5580 15642
rect 6748 15638 6776 15846
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5736 12782 5764 13330
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7546 6040 7686
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5092 3534 5120 4422
rect 6196 4146 6224 15370
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6840 12850 6868 13398
rect 6932 13326 6960 21830
rect 7024 16046 7052 25298
rect 7300 22030 7328 25842
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7484 23730 7512 24686
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7300 21894 7328 21966
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7116 15858 7144 21286
rect 7576 19242 7604 26726
rect 7668 26450 7696 27814
rect 7656 26444 7708 26450
rect 7656 26386 7708 26392
rect 7748 25696 7800 25702
rect 7748 25638 7800 25644
rect 7760 25362 7788 25638
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7852 24750 7880 39782
rect 8036 39642 8064 40870
rect 8024 39636 8076 39642
rect 8024 39578 8076 39584
rect 8036 38418 8064 39578
rect 8128 38554 8156 41686
rect 9968 41682 9996 42230
rect 10416 42152 10468 42158
rect 10416 42094 10468 42100
rect 10232 42016 10284 42022
rect 10232 41958 10284 41964
rect 8300 41676 8352 41682
rect 8300 41618 8352 41624
rect 8668 41676 8720 41682
rect 8668 41618 8720 41624
rect 9956 41676 10008 41682
rect 9956 41618 10008 41624
rect 8312 41070 8340 41618
rect 8680 41562 8708 41618
rect 8680 41546 8892 41562
rect 8680 41540 8904 41546
rect 8680 41534 8852 41540
rect 8852 41482 8904 41488
rect 9956 41540 10008 41546
rect 9956 41482 10008 41488
rect 9128 41472 9180 41478
rect 9128 41414 9180 41420
rect 9140 41070 9168 41414
rect 9968 41070 9996 41482
rect 10244 41274 10272 41958
rect 10428 41857 10456 42094
rect 10414 41848 10470 41857
rect 10704 41818 10732 42638
rect 10796 42294 10824 43182
rect 12624 43172 12676 43178
rect 12624 43114 12676 43120
rect 11704 43104 11756 43110
rect 11704 43046 11756 43052
rect 11716 42702 11744 43046
rect 11704 42696 11756 42702
rect 11704 42638 11756 42644
rect 12176 42622 12572 42650
rect 12176 42566 12204 42622
rect 12164 42560 12216 42566
rect 12164 42502 12216 42508
rect 12256 42560 12308 42566
rect 12256 42502 12308 42508
rect 10784 42288 10836 42294
rect 10784 42230 10836 42236
rect 11334 42120 11390 42129
rect 11334 42055 11390 42064
rect 10414 41783 10416 41792
rect 10468 41783 10470 41792
rect 10692 41812 10744 41818
rect 10416 41754 10468 41760
rect 10692 41754 10744 41760
rect 10968 41812 11020 41818
rect 10968 41754 11020 41760
rect 10428 41723 10456 41754
rect 10980 41682 11008 41754
rect 10416 41676 10468 41682
rect 10416 41618 10468 41624
rect 10968 41676 11020 41682
rect 10968 41618 11020 41624
rect 10428 41478 10456 41618
rect 10416 41472 10468 41478
rect 10416 41414 10468 41420
rect 10232 41268 10284 41274
rect 10232 41210 10284 41216
rect 10980 41206 11008 41618
rect 10968 41200 11020 41206
rect 10968 41142 11020 41148
rect 8300 41064 8352 41070
rect 8300 41006 8352 41012
rect 9128 41064 9180 41070
rect 9128 41006 9180 41012
rect 9956 41064 10008 41070
rect 9956 41006 10008 41012
rect 8852 40996 8904 41002
rect 8852 40938 8904 40944
rect 8760 39364 8812 39370
rect 8760 39306 8812 39312
rect 8116 38548 8168 38554
rect 8116 38490 8168 38496
rect 8772 38418 8800 39306
rect 8024 38412 8076 38418
rect 8024 38354 8076 38360
rect 8760 38412 8812 38418
rect 8760 38354 8812 38360
rect 8300 37392 8352 37398
rect 8300 37334 8352 37340
rect 8208 36236 8260 36242
rect 8208 36178 8260 36184
rect 8220 35086 8248 36178
rect 8312 35154 8340 37334
rect 8864 36718 8892 40938
rect 9968 40730 9996 41006
rect 10508 40928 10560 40934
rect 10508 40870 10560 40876
rect 10520 40730 10548 40870
rect 9956 40724 10008 40730
rect 9956 40666 10008 40672
rect 10508 40724 10560 40730
rect 10508 40666 10560 40672
rect 9772 40044 9824 40050
rect 9772 39986 9824 39992
rect 9784 39846 9812 39986
rect 9772 39840 9824 39846
rect 9772 39782 9824 39788
rect 9784 39438 9812 39782
rect 9772 39432 9824 39438
rect 9772 39374 9824 39380
rect 9784 39098 9812 39374
rect 9772 39092 9824 39098
rect 9772 39034 9824 39040
rect 9772 38820 9824 38826
rect 9772 38762 9824 38768
rect 8852 36712 8904 36718
rect 8852 36654 8904 36660
rect 9784 35222 9812 38762
rect 9968 38554 9996 40666
rect 11152 40520 11204 40526
rect 11152 40462 11204 40468
rect 11164 40186 11192 40462
rect 11152 40180 11204 40186
rect 11152 40122 11204 40128
rect 10692 40112 10744 40118
rect 10692 40054 10744 40060
rect 10704 39982 10732 40054
rect 10692 39976 10744 39982
rect 10692 39918 10744 39924
rect 10876 39976 10928 39982
rect 10876 39918 10928 39924
rect 10888 39370 10916 39918
rect 10600 39364 10652 39370
rect 10600 39306 10652 39312
rect 10876 39364 10928 39370
rect 10876 39306 10928 39312
rect 9956 38548 10008 38554
rect 9956 38490 10008 38496
rect 10416 38480 10468 38486
rect 10416 38422 10468 38428
rect 10048 38276 10100 38282
rect 10048 38218 10100 38224
rect 9864 38004 9916 38010
rect 9864 37946 9916 37952
rect 9876 37330 9904 37946
rect 10060 37874 10088 38218
rect 10048 37868 10100 37874
rect 10048 37810 10100 37816
rect 10060 37466 10088 37810
rect 10140 37732 10192 37738
rect 10140 37674 10192 37680
rect 10048 37460 10100 37466
rect 10048 37402 10100 37408
rect 9864 37324 9916 37330
rect 9864 37266 9916 37272
rect 9876 36310 9904 37266
rect 9864 36304 9916 36310
rect 9864 36246 9916 36252
rect 10152 35630 10180 37674
rect 10140 35624 10192 35630
rect 10140 35566 10192 35572
rect 10324 35556 10376 35562
rect 10324 35498 10376 35504
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 9772 35216 9824 35222
rect 9772 35158 9824 35164
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 8208 35080 8260 35086
rect 8208 35022 8260 35028
rect 8220 33454 8248 35022
rect 9128 35012 9180 35018
rect 9128 34954 9180 34960
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 9048 33522 9076 33934
rect 9036 33516 9088 33522
rect 9036 33458 9088 33464
rect 8208 33448 8260 33454
rect 8208 33390 8260 33396
rect 8300 33312 8352 33318
rect 8300 33254 8352 33260
rect 8208 32972 8260 32978
rect 8208 32914 8260 32920
rect 8220 32570 8248 32914
rect 7932 32564 7984 32570
rect 7932 32506 7984 32512
rect 8208 32564 8260 32570
rect 8208 32506 8260 32512
rect 7944 32298 7972 32506
rect 8116 32428 8168 32434
rect 8116 32370 8168 32376
rect 8024 32360 8076 32366
rect 8024 32302 8076 32308
rect 7932 32292 7984 32298
rect 7932 32234 7984 32240
rect 7944 29646 7972 32234
rect 8036 31482 8064 32302
rect 8128 32026 8156 32370
rect 8208 32224 8260 32230
rect 8208 32166 8260 32172
rect 8220 32026 8248 32166
rect 8116 32020 8168 32026
rect 8116 31962 8168 31968
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8024 31476 8076 31482
rect 8024 31418 8076 31424
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 8312 28948 8340 33254
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 8668 32768 8720 32774
rect 8668 32710 8720 32716
rect 8680 32230 8708 32710
rect 8760 32564 8812 32570
rect 8760 32506 8812 32512
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8576 31680 8628 31686
rect 8576 31622 8628 31628
rect 8588 29170 8616 31622
rect 8680 31482 8708 32166
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 8576 29164 8628 29170
rect 8576 29106 8628 29112
rect 8128 28920 8340 28948
rect 8128 25974 8156 28920
rect 8484 28416 8536 28422
rect 8484 28358 8536 28364
rect 8496 28218 8524 28358
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8772 28098 8800 32506
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 8864 31686 8892 31758
rect 8852 31680 8904 31686
rect 8852 31622 8904 31628
rect 8680 28070 8800 28098
rect 8484 28008 8536 28014
rect 8484 27950 8536 27956
rect 8496 27674 8524 27950
rect 8484 27668 8536 27674
rect 8484 27610 8536 27616
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8392 26852 8444 26858
rect 8392 26794 8444 26800
rect 8116 25968 8168 25974
rect 8116 25910 8168 25916
rect 8404 25838 8432 26794
rect 8588 26042 8616 26862
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 8680 25974 8708 28070
rect 8760 27940 8812 27946
rect 8760 27882 8812 27888
rect 8772 27606 8800 27882
rect 8760 27600 8812 27606
rect 8760 27542 8812 27548
rect 8668 25968 8720 25974
rect 8668 25910 8720 25916
rect 8392 25832 8444 25838
rect 8392 25774 8444 25780
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 7840 24744 7892 24750
rect 8024 24744 8076 24750
rect 7840 24686 7892 24692
rect 7944 24704 8024 24732
rect 7944 23662 7972 24704
rect 8024 24686 8076 24692
rect 8208 24676 8260 24682
rect 8208 24618 8260 24624
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7196 19236 7248 19242
rect 7196 19178 7248 19184
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7208 18766 7236 19178
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7208 18358 7236 18702
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7300 17066 7328 18294
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7300 15978 7328 17002
rect 7392 16726 7420 19110
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7024 15830 7144 15858
rect 7024 14278 7052 15830
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6564 4826 6592 12786
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6932 11694 6960 11834
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10810 6868 10950
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9518 6868 10066
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9586 6960 9998
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 7750 6868 9454
rect 7024 7954 7052 14214
rect 7208 13394 7236 14418
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9586 7420 9862
rect 7484 9602 7512 12854
rect 7576 12782 7604 13330
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 10266 7604 10474
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7380 9580 7432 9586
rect 7484 9574 7604 9602
rect 7380 9522 7432 9528
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7300 8022 7328 9454
rect 7484 8634 7512 9454
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6840 6254 6868 7686
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7116 6322 7144 6666
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 4826 6868 6190
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 7576 4010 7604 9574
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 7750 7696 8366
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 7410 7696 7686
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7760 5710 7788 23462
rect 7944 19378 7972 23598
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8128 21486 8156 22034
rect 8220 21554 8248 24618
rect 8312 24206 8340 25094
rect 8680 24750 8708 25774
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 8852 23656 8904 23662
rect 8852 23598 8904 23604
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8588 22234 8616 22510
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8864 21622 8892 23598
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18834 8616 19110
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8588 18222 8616 18770
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8864 18290 8892 18702
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 7944 17814 7972 18158
rect 8116 18080 8168 18086
rect 8114 18048 8116 18057
rect 8168 18048 8170 18057
rect 8114 17983 8170 17992
rect 8588 17882 8616 18158
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 8864 17270 8892 18226
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8956 16998 8984 32846
rect 9140 31668 9168 34954
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 9404 34536 9456 34542
rect 9404 34478 9456 34484
rect 9416 33046 9444 34478
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 9404 33040 9456 33046
rect 9404 32982 9456 32988
rect 9048 31640 9168 31668
rect 9048 28966 9076 31640
rect 9220 30592 9272 30598
rect 9220 30534 9272 30540
rect 9036 28960 9088 28966
rect 9036 28902 9088 28908
rect 9126 27568 9182 27577
rect 9126 27503 9128 27512
rect 9180 27503 9182 27512
rect 9128 27474 9180 27480
rect 9232 26926 9260 30534
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 9312 27668 9364 27674
rect 9312 27610 9364 27616
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 9324 26042 9352 27610
rect 9416 26994 9444 27950
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 9324 25838 9352 25978
rect 9312 25832 9364 25838
rect 9312 25774 9364 25780
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9048 21486 9076 21830
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9048 19378 9076 21422
rect 9508 19922 9536 33798
rect 9770 31512 9826 31521
rect 9770 31447 9772 31456
rect 9824 31447 9826 31456
rect 9772 31418 9824 31424
rect 9588 31204 9640 31210
rect 9588 31146 9640 31152
rect 9600 30870 9628 31146
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9588 30864 9640 30870
rect 9588 30806 9640 30812
rect 9692 30190 9720 31078
rect 9680 30184 9732 30190
rect 9732 30132 9812 30138
rect 9680 30126 9812 30132
rect 9692 30110 9812 30126
rect 9784 30054 9812 30110
rect 9772 30048 9824 30054
rect 9772 29990 9824 29996
rect 9680 28008 9732 28014
rect 9680 27950 9732 27956
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9600 26382 9628 27270
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9600 24206 9628 24550
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9600 23798 9628 24142
rect 9588 23792 9640 23798
rect 9588 23734 9640 23740
rect 9600 22710 9628 23734
rect 9692 22982 9720 27950
rect 9784 24410 9812 29990
rect 9876 28150 9904 34546
rect 10244 33998 10272 35430
rect 10336 35154 10364 35498
rect 10324 35148 10376 35154
rect 10324 35090 10376 35096
rect 10428 34678 10456 38422
rect 10612 37806 10640 39306
rect 10968 38888 11020 38894
rect 10968 38830 11020 38836
rect 11244 38888 11296 38894
rect 11244 38830 11296 38836
rect 10980 38486 11008 38830
rect 11256 38554 11284 38830
rect 11244 38548 11296 38554
rect 11244 38490 11296 38496
rect 10968 38480 11020 38486
rect 10968 38422 11020 38428
rect 10784 38412 10836 38418
rect 10784 38354 10836 38360
rect 10600 37800 10652 37806
rect 10600 37742 10652 37748
rect 10796 36718 10824 38354
rect 10876 38344 10928 38350
rect 10876 38286 10928 38292
rect 10888 37806 10916 38286
rect 10980 37874 11008 38422
rect 11256 38418 11284 38490
rect 11244 38412 11296 38418
rect 11244 38354 11296 38360
rect 10968 37868 11020 37874
rect 10968 37810 11020 37816
rect 10876 37800 10928 37806
rect 10876 37742 10928 37748
rect 10888 36922 10916 37742
rect 10980 37398 11008 37810
rect 10968 37392 11020 37398
rect 10968 37334 11020 37340
rect 10876 36916 10928 36922
rect 10876 36858 10928 36864
rect 10784 36712 10836 36718
rect 10784 36654 10836 36660
rect 10600 36304 10652 36310
rect 10600 36246 10652 36252
rect 10612 34678 10640 36246
rect 10796 35714 10824 36654
rect 11060 36168 11112 36174
rect 11060 36110 11112 36116
rect 10796 35686 11008 35714
rect 10980 35630 11008 35686
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10980 35018 11008 35566
rect 11072 35222 11100 36110
rect 11060 35216 11112 35222
rect 11060 35158 11112 35164
rect 10968 35012 11020 35018
rect 10968 34954 11020 34960
rect 10416 34672 10468 34678
rect 10416 34614 10468 34620
rect 10600 34672 10652 34678
rect 10600 34614 10652 34620
rect 10612 34066 10640 34614
rect 10980 34490 11008 34954
rect 11152 34536 11204 34542
rect 10980 34484 11152 34490
rect 10980 34478 11204 34484
rect 10980 34462 11192 34478
rect 10600 34060 10652 34066
rect 10600 34002 10652 34008
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 10980 33402 11008 34462
rect 10888 33386 11008 33402
rect 10876 33380 11008 33386
rect 10928 33374 11008 33380
rect 10876 33322 10928 33328
rect 10968 33312 11020 33318
rect 10968 33254 11020 33260
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 10060 32502 10088 32710
rect 10048 32496 10100 32502
rect 10048 32438 10100 32444
rect 10060 31278 10088 32438
rect 10048 31272 10100 31278
rect 10048 31214 10100 31220
rect 10600 30388 10652 30394
rect 10600 30330 10652 30336
rect 10612 30190 10640 30330
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 9864 28144 9916 28150
rect 9864 28086 9916 28092
rect 10600 27532 10652 27538
rect 10600 27474 10652 27480
rect 10612 25702 10640 27474
rect 10980 27402 11008 33254
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 11152 31204 11204 31210
rect 11152 31146 11204 31152
rect 11060 30796 11112 30802
rect 11060 30738 11112 30744
rect 11072 30326 11100 30738
rect 11060 30320 11112 30326
rect 11060 30262 11112 30268
rect 11164 29714 11192 31146
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 11256 27946 11284 31826
rect 11348 28150 11376 42055
rect 12268 41818 12296 42502
rect 12544 42362 12572 42622
rect 12532 42356 12584 42362
rect 12532 42298 12584 42304
rect 12636 42158 12664 43114
rect 17052 42838 17080 43658
rect 19444 43450 19472 43794
rect 23848 43784 23900 43790
rect 23848 43726 23900 43732
rect 23860 43654 23888 43726
rect 23848 43648 23900 43654
rect 23848 43590 23900 43596
rect 19432 43444 19484 43450
rect 19432 43386 19484 43392
rect 18236 43308 18288 43314
rect 18236 43250 18288 43256
rect 17684 43104 17736 43110
rect 17684 43046 17736 43052
rect 17040 42832 17092 42838
rect 17040 42774 17092 42780
rect 14096 42764 14148 42770
rect 14096 42706 14148 42712
rect 15660 42764 15712 42770
rect 15660 42706 15712 42712
rect 13636 42220 13688 42226
rect 13636 42162 13688 42168
rect 12624 42152 12676 42158
rect 12624 42094 12676 42100
rect 12532 42016 12584 42022
rect 12530 41984 12532 41993
rect 12584 41984 12586 41993
rect 12530 41919 12586 41928
rect 12256 41812 12308 41818
rect 12256 41754 12308 41760
rect 11520 41744 11572 41750
rect 11520 41686 11572 41692
rect 11532 41478 11560 41686
rect 11520 41472 11572 41478
rect 11520 41414 11572 41420
rect 13360 41472 13412 41478
rect 13360 41414 13412 41420
rect 13084 41268 13136 41274
rect 13084 41210 13136 41216
rect 12808 41132 12860 41138
rect 12808 41074 12860 41080
rect 12716 41064 12768 41070
rect 12716 41006 12768 41012
rect 12624 40384 12676 40390
rect 12624 40326 12676 40332
rect 11704 39840 11756 39846
rect 11704 39782 11756 39788
rect 11716 39574 11744 39782
rect 11704 39568 11756 39574
rect 11704 39510 11756 39516
rect 12636 39506 12664 40326
rect 12728 39574 12756 41006
rect 12820 40730 12848 41074
rect 12808 40724 12860 40730
rect 12808 40666 12860 40672
rect 12900 40520 12952 40526
rect 12900 40462 12952 40468
rect 12912 40186 12940 40462
rect 12900 40180 12952 40186
rect 12900 40122 12952 40128
rect 12716 39568 12768 39574
rect 12716 39510 12768 39516
rect 12912 39506 12940 40122
rect 12992 39976 13044 39982
rect 12992 39918 13044 39924
rect 13004 39574 13032 39918
rect 12992 39568 13044 39574
rect 12992 39510 13044 39516
rect 12624 39500 12676 39506
rect 12624 39442 12676 39448
rect 12900 39500 12952 39506
rect 12900 39442 12952 39448
rect 11520 39092 11572 39098
rect 11520 39034 11572 39040
rect 11532 38894 11560 39034
rect 11520 38888 11572 38894
rect 11520 38830 11572 38836
rect 11980 38412 12032 38418
rect 11980 38354 12032 38360
rect 12164 38412 12216 38418
rect 12164 38354 12216 38360
rect 11428 37936 11480 37942
rect 11428 37878 11480 37884
rect 11440 37330 11468 37878
rect 11992 37330 12020 38354
rect 12176 38010 12204 38354
rect 12164 38004 12216 38010
rect 12164 37946 12216 37952
rect 12636 37806 12664 39442
rect 13096 38554 13124 41210
rect 13372 39982 13400 41414
rect 13648 40934 13676 42162
rect 13740 41682 13860 41698
rect 13740 41676 13872 41682
rect 13740 41670 13820 41676
rect 13740 41478 13768 41670
rect 13820 41618 13872 41624
rect 13728 41472 13780 41478
rect 13728 41414 13780 41420
rect 13636 40928 13688 40934
rect 13636 40870 13688 40876
rect 14004 40928 14056 40934
rect 14004 40870 14056 40876
rect 14016 40730 14044 40870
rect 14004 40724 14056 40730
rect 14004 40666 14056 40672
rect 13360 39976 13412 39982
rect 13360 39918 13412 39924
rect 13372 39846 13400 39918
rect 13268 39840 13320 39846
rect 13268 39782 13320 39788
rect 13360 39840 13412 39846
rect 13360 39782 13412 39788
rect 13280 38894 13308 39782
rect 13268 38888 13320 38894
rect 13268 38830 13320 38836
rect 13084 38548 13136 38554
rect 13084 38490 13136 38496
rect 12624 37800 12676 37806
rect 12624 37742 12676 37748
rect 11428 37324 11480 37330
rect 11428 37266 11480 37272
rect 11980 37324 12032 37330
rect 11980 37266 12032 37272
rect 11520 35488 11572 35494
rect 11520 35430 11572 35436
rect 11532 35086 11560 35430
rect 12348 35284 12400 35290
rect 12348 35226 12400 35232
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 12360 32842 12388 35226
rect 13176 34060 13228 34066
rect 13176 34002 13228 34008
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12820 33862 12848 33934
rect 12808 33856 12860 33862
rect 12808 33798 12860 33804
rect 12820 33454 12848 33798
rect 12532 33448 12584 33454
rect 12532 33390 12584 33396
rect 12808 33448 12860 33454
rect 12808 33390 12860 33396
rect 12348 32836 12400 32842
rect 12348 32778 12400 32784
rect 12072 32224 12124 32230
rect 12072 32166 12124 32172
rect 12084 31890 12112 32166
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 12164 30864 12216 30870
rect 12164 30806 12216 30812
rect 12176 30598 12204 30806
rect 12164 30592 12216 30598
rect 12164 30534 12216 30540
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11532 29306 11560 30194
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 12084 29850 12112 30126
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11704 28484 11756 28490
rect 11704 28426 11756 28432
rect 11336 28144 11388 28150
rect 11336 28086 11388 28092
rect 11244 27940 11296 27946
rect 11244 27882 11296 27888
rect 11152 27872 11204 27878
rect 11152 27814 11204 27820
rect 11164 27674 11192 27814
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 11348 27130 11376 28086
rect 11716 27470 11744 28426
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 11704 27464 11756 27470
rect 11704 27406 11756 27412
rect 11336 27124 11388 27130
rect 11336 27066 11388 27072
rect 11716 26976 11744 27406
rect 11624 26948 11744 26976
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 9968 24750 9996 25638
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 11072 24682 11100 25434
rect 11060 24676 11112 24682
rect 11060 24618 11112 24624
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9968 24274 9996 24550
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10232 23588 10284 23594
rect 10232 23530 10284 23536
rect 10244 23322 10272 23530
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9588 22704 9640 22710
rect 9588 22646 9640 22652
rect 9692 21690 9720 22918
rect 9954 22808 10010 22817
rect 9954 22743 10010 22752
rect 9968 22506 9996 22743
rect 9956 22500 10008 22506
rect 9956 22442 10008 22448
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9784 21146 9812 21966
rect 9968 21146 9996 22442
rect 10244 22098 10272 23258
rect 10692 23248 10744 23254
rect 10692 23190 10744 23196
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9784 19922 9812 21082
rect 10704 21010 10732 23190
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10704 20398 10732 20946
rect 10888 20398 10916 21422
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 9496 19916 9548 19922
rect 9772 19916 9824 19922
rect 9548 19876 9720 19904
rect 9496 19858 9548 19864
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9692 19310 9720 19876
rect 9772 19858 9824 19864
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9680 19304 9732 19310
rect 9600 19264 9680 19292
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9232 18034 9260 18634
rect 9600 18057 9628 19264
rect 9680 19246 9732 19252
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9692 18086 9720 18838
rect 9680 18080 9732 18086
rect 9586 18048 9642 18057
rect 9232 18006 9352 18034
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 9048 17134 9076 17682
rect 9232 17134 9260 17818
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 9232 16726 9260 17070
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9324 16046 9352 18006
rect 9680 18022 9732 18028
rect 9586 17983 9642 17992
rect 9600 17338 9628 17983
rect 9692 17746 9720 18022
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9416 17134 9444 17206
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8772 15706 8800 15846
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7852 13530 7880 14894
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7944 13394 7972 15302
rect 8772 15094 8800 15642
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 9508 14618 9536 16662
rect 9692 16658 9720 17546
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9784 16046 9812 19722
rect 10060 19718 10088 19858
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10336 19514 10364 19654
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9876 15570 9904 17002
rect 10060 16658 10088 18090
rect 10152 16658 10180 19314
rect 10520 19310 10548 19858
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10428 18698 10456 18838
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10796 17882 10824 18634
rect 10888 18086 10916 20334
rect 10980 19310 11008 20742
rect 11072 19990 11100 20810
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10980 18902 11008 19246
rect 11072 18970 11100 19246
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 11164 18222 11192 24006
rect 11336 23588 11388 23594
rect 11336 23530 11388 23536
rect 11348 22098 11376 23530
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11244 21616 11296 21622
rect 11244 21558 11296 21564
rect 11256 19854 11284 21558
rect 11624 21146 11652 26948
rect 11796 26784 11848 26790
rect 11796 26726 11848 26732
rect 11704 24744 11756 24750
rect 11704 24686 11756 24692
rect 11716 24070 11744 24686
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11704 23180 11756 23186
rect 11808 23168 11836 26726
rect 11980 25968 12032 25974
rect 11980 25910 12032 25916
rect 11992 25498 12020 25910
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 12084 25378 12112 27610
rect 12360 26858 12388 32778
rect 12544 32774 12572 33390
rect 12900 33040 12952 33046
rect 12900 32982 12952 32988
rect 12532 32768 12584 32774
rect 12532 32710 12584 32716
rect 12808 32224 12860 32230
rect 12808 32166 12860 32172
rect 12714 32056 12770 32065
rect 12714 31991 12770 32000
rect 12728 31958 12756 31991
rect 12716 31952 12768 31958
rect 12716 31894 12768 31900
rect 12820 31890 12848 32166
rect 12808 31884 12860 31890
rect 12808 31826 12860 31832
rect 12716 31816 12768 31822
rect 12714 31784 12716 31793
rect 12768 31784 12770 31793
rect 12714 31719 12770 31728
rect 12912 31414 12940 32982
rect 12992 32292 13044 32298
rect 12992 32234 13044 32240
rect 13004 31958 13032 32234
rect 12992 31952 13044 31958
rect 12992 31894 13044 31900
rect 12992 31816 13044 31822
rect 12992 31758 13044 31764
rect 13004 31686 13032 31758
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 12900 31408 12952 31414
rect 12900 31350 12952 31356
rect 13004 31210 13032 31622
rect 13188 31414 13216 34002
rect 13372 33046 13400 39782
rect 14004 38820 14056 38826
rect 14004 38762 14056 38768
rect 14016 38418 14044 38762
rect 14004 38412 14056 38418
rect 14004 38354 14056 38360
rect 13544 37392 13596 37398
rect 13544 37334 13596 37340
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13464 34542 13492 35430
rect 13452 34536 13504 34542
rect 13452 34478 13504 34484
rect 13360 33040 13412 33046
rect 13360 32982 13412 32988
rect 13464 31906 13492 34478
rect 13556 34202 13584 37334
rect 13636 35624 13688 35630
rect 13636 35566 13688 35572
rect 13544 34196 13596 34202
rect 13544 34138 13596 34144
rect 13648 33658 13676 35566
rect 13912 34944 13964 34950
rect 13912 34886 13964 34892
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13924 33454 13952 34886
rect 13912 33448 13964 33454
rect 13912 33390 13964 33396
rect 14016 33114 14044 38354
rect 14004 33108 14056 33114
rect 14004 33050 14056 33056
rect 13912 32768 13964 32774
rect 13912 32710 13964 32716
rect 13924 32609 13952 32710
rect 13542 32600 13598 32609
rect 13542 32535 13598 32544
rect 13910 32600 13966 32609
rect 13910 32535 13966 32544
rect 13556 32366 13584 32535
rect 13544 32360 13596 32366
rect 13596 32320 13676 32348
rect 13544 32302 13596 32308
rect 13372 31878 13492 31906
rect 13176 31408 13228 31414
rect 13176 31350 13228 31356
rect 12992 31204 13044 31210
rect 12992 31146 13044 31152
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12912 30190 12940 30670
rect 12900 30184 12952 30190
rect 12900 30126 12952 30132
rect 13004 30054 13032 31146
rect 13188 30394 13216 31350
rect 13372 30802 13400 31878
rect 13648 31754 13676 32320
rect 13728 32292 13780 32298
rect 13728 32234 13780 32240
rect 13636 31748 13688 31754
rect 13636 31690 13688 31696
rect 13740 31686 13768 32234
rect 13820 31816 13872 31822
rect 13818 31784 13820 31793
rect 13872 31784 13874 31793
rect 13818 31719 13874 31728
rect 13728 31680 13780 31686
rect 13728 31622 13780 31628
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13740 30802 13768 31214
rect 13360 30796 13412 30802
rect 13360 30738 13412 30744
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13372 30598 13400 30738
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 13176 30388 13228 30394
rect 13176 30330 13228 30336
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 13372 29170 13400 30534
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13544 29096 13596 29102
rect 13544 29038 13596 29044
rect 13176 28688 13228 28694
rect 13176 28630 13228 28636
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 12624 28484 12676 28490
rect 12624 28426 12676 28432
rect 12636 27538 12664 28426
rect 13004 27878 13032 28494
rect 13084 28008 13136 28014
rect 13084 27950 13136 27956
rect 13096 27878 13124 27950
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 12624 27532 12676 27538
rect 12624 27474 12676 27480
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 11992 25362 12112 25378
rect 11980 25356 12112 25362
rect 12032 25350 12112 25356
rect 11980 25298 12032 25304
rect 11992 23254 12020 25298
rect 12360 24886 12388 26794
rect 12348 24880 12400 24886
rect 12348 24822 12400 24828
rect 12360 23866 12388 24822
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 11980 23248 12032 23254
rect 11980 23190 12032 23196
rect 11756 23140 11836 23168
rect 12164 23180 12216 23186
rect 11704 23122 11756 23128
rect 12164 23122 12216 23128
rect 12176 22982 12204 23122
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 11992 21894 12020 22034
rect 12176 21894 12204 22918
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11624 21010 11652 21082
rect 11900 21010 11928 21490
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19514 11284 19790
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 10876 18080 10928 18086
rect 11256 18034 11284 19450
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11348 18834 11376 18906
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 10876 18022 10928 18028
rect 11072 18006 11284 18034
rect 11072 17898 11100 18006
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10888 17870 11100 17898
rect 10888 17814 10916 17870
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10876 17808 10928 17814
rect 11060 17808 11112 17814
rect 10876 17750 10928 17756
rect 10980 17756 11060 17762
rect 10980 17750 11112 17756
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10428 17066 10456 17682
rect 10520 17542 10548 17750
rect 10980 17734 11100 17750
rect 11256 17746 11284 18006
rect 11348 17746 11376 18770
rect 11244 17740 11296 17746
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10888 17134 10916 17614
rect 10980 17134 11008 17734
rect 11244 17682 11296 17688
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10506 16688 10562 16697
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10140 16652 10192 16658
rect 10506 16623 10508 16632
rect 10140 16594 10192 16600
rect 10560 16623 10562 16632
rect 10692 16652 10744 16658
rect 10508 16594 10560 16600
rect 10692 16594 10744 16600
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 13938 8156 14282
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12238 8064 12582
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8220 11898 8248 14010
rect 9508 13938 9536 14554
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8864 12782 8892 13126
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8864 12646 8892 12718
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 12442 8892 12582
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 10612 11694 10640 15982
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 7944 11218 7972 11630
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7944 10810 7972 11154
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8036 9654 8064 11086
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 8128 4622 8156 11562
rect 10704 11354 10732 16594
rect 11348 15978 11376 16594
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11348 15434 11376 15914
rect 11440 15706 11468 16594
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 13870 11008 14758
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10980 13394 11008 13806
rect 11624 13530 11652 20946
rect 11900 20602 11928 20946
rect 11992 20806 12020 21830
rect 13004 21570 13032 27814
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13096 26926 13124 27270
rect 13188 27130 13216 28630
rect 13556 28098 13584 29038
rect 13740 28626 13768 30738
rect 13832 30394 13860 31719
rect 13820 30388 13872 30394
rect 13820 30330 13872 30336
rect 14108 29850 14136 42706
rect 15016 42696 15068 42702
rect 15016 42638 15068 42644
rect 14186 41848 14242 41857
rect 15028 41818 15056 42638
rect 15292 42084 15344 42090
rect 15292 42026 15344 42032
rect 15200 42016 15252 42022
rect 15200 41958 15252 41964
rect 14186 41783 14242 41792
rect 15016 41812 15068 41818
rect 14200 41478 14228 41783
rect 15016 41754 15068 41760
rect 14648 41744 14700 41750
rect 14700 41692 14964 41698
rect 14648 41686 14964 41692
rect 14660 41670 14964 41686
rect 14936 41614 14964 41670
rect 14924 41608 14976 41614
rect 14924 41550 14976 41556
rect 14188 41472 14240 41478
rect 14188 41414 14240 41420
rect 14188 40112 14240 40118
rect 14188 40054 14240 40060
rect 14200 38554 14228 40054
rect 14648 39840 14700 39846
rect 14648 39782 14700 39788
rect 14660 38962 14688 39782
rect 15028 39030 15056 41754
rect 15212 41274 15240 41958
rect 15200 41268 15252 41274
rect 15200 41210 15252 41216
rect 15016 39024 15068 39030
rect 15016 38966 15068 38972
rect 14648 38956 14700 38962
rect 14648 38898 14700 38904
rect 14832 38888 14884 38894
rect 14832 38830 14884 38836
rect 15016 38888 15068 38894
rect 15016 38830 15068 38836
rect 14188 38548 14240 38554
rect 14188 38490 14240 38496
rect 14200 38010 14228 38490
rect 14464 38480 14516 38486
rect 14464 38422 14516 38428
rect 14188 38004 14240 38010
rect 14188 37946 14240 37952
rect 14280 38004 14332 38010
rect 14280 37946 14332 37952
rect 14292 37806 14320 37946
rect 14476 37874 14504 38422
rect 14844 38418 14872 38830
rect 15028 38729 15056 38830
rect 15014 38720 15070 38729
rect 15014 38655 15070 38664
rect 14832 38412 14884 38418
rect 14832 38354 14884 38360
rect 14844 38214 14872 38354
rect 15200 38276 15252 38282
rect 15200 38218 15252 38224
rect 14832 38208 14884 38214
rect 14832 38150 14884 38156
rect 15212 37874 15240 38218
rect 14464 37868 14516 37874
rect 14464 37810 14516 37816
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 14280 37800 14332 37806
rect 14280 37742 14332 37748
rect 15304 37738 15332 42026
rect 15672 41478 15700 42706
rect 17052 42702 17080 42774
rect 17696 42702 17724 43046
rect 17040 42696 17092 42702
rect 17040 42638 17092 42644
rect 17684 42696 17736 42702
rect 17684 42638 17736 42644
rect 17960 42696 18012 42702
rect 17960 42638 18012 42644
rect 16394 42256 16450 42265
rect 17052 42242 17080 42638
rect 17592 42560 17644 42566
rect 17592 42502 17644 42508
rect 17604 42401 17632 42502
rect 17590 42392 17646 42401
rect 17590 42327 17646 42336
rect 17498 42256 17554 42265
rect 17052 42226 17264 42242
rect 16394 42191 16450 42200
rect 16856 42220 16908 42226
rect 16408 42158 16436 42191
rect 17052 42220 17276 42226
rect 17052 42214 17224 42220
rect 16856 42162 16908 42168
rect 17498 42191 17500 42200
rect 17224 42162 17276 42168
rect 17552 42191 17554 42200
rect 17500 42162 17552 42168
rect 16396 42152 16448 42158
rect 16396 42094 16448 42100
rect 16580 42152 16632 42158
rect 16580 42094 16632 42100
rect 16592 42022 16620 42094
rect 16580 42016 16632 42022
rect 16580 41958 16632 41964
rect 16868 41818 16896 42162
rect 17512 41834 17540 42162
rect 17684 42152 17736 42158
rect 17684 42094 17736 42100
rect 17592 42016 17644 42022
rect 17696 41970 17724 42094
rect 17644 41964 17724 41970
rect 17592 41958 17724 41964
rect 17776 42016 17828 42022
rect 17776 41958 17828 41964
rect 17866 41984 17922 41993
rect 17604 41942 17724 41958
rect 16856 41812 16908 41818
rect 17512 41806 17632 41834
rect 16856 41754 16908 41760
rect 15660 41472 15712 41478
rect 15660 41414 15712 41420
rect 16396 40928 16448 40934
rect 16396 40870 16448 40876
rect 16408 40526 16436 40870
rect 16488 40588 16540 40594
rect 16488 40530 16540 40536
rect 16396 40520 16448 40526
rect 16396 40462 16448 40468
rect 16408 39506 16436 40462
rect 16396 39500 16448 39506
rect 16396 39442 16448 39448
rect 15752 39432 15804 39438
rect 15752 39374 15804 39380
rect 15474 38720 15530 38729
rect 15474 38655 15530 38664
rect 15384 38344 15436 38350
rect 15384 38286 15436 38292
rect 15292 37732 15344 37738
rect 15292 37674 15344 37680
rect 15396 37398 15424 38286
rect 15384 37392 15436 37398
rect 15384 37334 15436 37340
rect 15488 37330 15516 38655
rect 15568 37664 15620 37670
rect 15568 37606 15620 37612
rect 15580 37466 15608 37606
rect 15568 37460 15620 37466
rect 15568 37402 15620 37408
rect 15476 37324 15528 37330
rect 15476 37266 15528 37272
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 14936 36582 14964 37062
rect 15488 36786 15516 37266
rect 15476 36780 15528 36786
rect 15476 36722 15528 36728
rect 14924 36576 14976 36582
rect 14924 36518 14976 36524
rect 14936 35698 14964 36518
rect 15488 36378 15516 36722
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 14556 35624 14608 35630
rect 14556 35566 14608 35572
rect 14280 34536 14332 34542
rect 14280 34478 14332 34484
rect 14292 34134 14320 34478
rect 14568 34406 14596 35566
rect 15016 35556 15068 35562
rect 15016 35498 15068 35504
rect 15028 35154 15056 35498
rect 15016 35148 15068 35154
rect 15016 35090 15068 35096
rect 15764 34678 15792 39374
rect 16500 38554 16528 40530
rect 16868 40118 16896 41754
rect 17604 41682 17632 41806
rect 17316 41676 17368 41682
rect 17316 41618 17368 41624
rect 17500 41676 17552 41682
rect 17500 41618 17552 41624
rect 17592 41676 17644 41682
rect 17592 41618 17644 41624
rect 17328 41478 17356 41618
rect 17316 41472 17368 41478
rect 17316 41414 17368 41420
rect 17512 41274 17540 41618
rect 17500 41268 17552 41274
rect 17500 41210 17552 41216
rect 16948 41064 17000 41070
rect 16948 41006 17000 41012
rect 16856 40112 16908 40118
rect 16856 40054 16908 40060
rect 16672 39432 16724 39438
rect 16672 39374 16724 39380
rect 16684 39098 16712 39374
rect 16672 39092 16724 39098
rect 16672 39034 16724 39040
rect 16960 38894 16988 41006
rect 17696 40050 17724 41942
rect 17788 41818 17816 41958
rect 17866 41919 17922 41928
rect 17776 41812 17828 41818
rect 17776 41754 17828 41760
rect 17880 41682 17908 41919
rect 17972 41818 18000 42638
rect 18050 42392 18106 42401
rect 18050 42327 18106 42336
rect 17960 41812 18012 41818
rect 17960 41754 18012 41760
rect 17868 41676 17920 41682
rect 17868 41618 17920 41624
rect 18064 41546 18092 42327
rect 18052 41540 18104 41546
rect 18052 41482 18104 41488
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 17972 41206 18000 41414
rect 18248 41274 18276 43250
rect 18328 43240 18380 43246
rect 18328 43182 18380 43188
rect 18340 42770 18368 43182
rect 19248 43104 19300 43110
rect 19248 43046 19300 43052
rect 23480 43104 23532 43110
rect 23480 43046 23532 43052
rect 18420 42900 18472 42906
rect 18420 42842 18472 42848
rect 18328 42764 18380 42770
rect 18328 42706 18380 42712
rect 18432 42362 18460 42842
rect 19260 42566 19288 43046
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19984 42900 20036 42906
rect 19984 42842 20036 42848
rect 19340 42696 19392 42702
rect 19340 42638 19392 42644
rect 19248 42560 19300 42566
rect 19248 42502 19300 42508
rect 18420 42356 18472 42362
rect 18420 42298 18472 42304
rect 18328 42220 18380 42226
rect 18328 42162 18380 42168
rect 18340 41818 18368 42162
rect 19352 42158 19380 42638
rect 19340 42152 19392 42158
rect 19340 42094 19392 42100
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 18328 41812 18380 41818
rect 18328 41754 18380 41760
rect 18512 41472 18564 41478
rect 18512 41414 18564 41420
rect 18524 41274 18552 41414
rect 18236 41268 18288 41274
rect 18236 41210 18288 41216
rect 18512 41268 18564 41274
rect 18512 41210 18564 41216
rect 17960 41200 18012 41206
rect 17960 41142 18012 41148
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 18236 40384 18288 40390
rect 18236 40326 18288 40332
rect 18420 40384 18472 40390
rect 18420 40326 18472 40332
rect 17684 40044 17736 40050
rect 17684 39986 17736 39992
rect 17408 39568 17460 39574
rect 17408 39510 17460 39516
rect 16672 38888 16724 38894
rect 16672 38830 16724 38836
rect 16948 38888 17000 38894
rect 16948 38830 17000 38836
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 16592 38554 16620 38694
rect 16488 38548 16540 38554
rect 16488 38490 16540 38496
rect 16580 38548 16632 38554
rect 16580 38490 16632 38496
rect 16592 38418 16620 38490
rect 15936 38412 15988 38418
rect 15936 38354 15988 38360
rect 16580 38412 16632 38418
rect 16580 38354 16632 38360
rect 15948 37806 15976 38354
rect 16396 38004 16448 38010
rect 16396 37946 16448 37952
rect 16488 38004 16540 38010
rect 16488 37946 16540 37952
rect 15936 37800 15988 37806
rect 15934 37768 15936 37777
rect 16304 37800 16356 37806
rect 15988 37768 15990 37777
rect 16304 37742 16356 37748
rect 15934 37703 15990 37712
rect 16316 37670 16344 37742
rect 16304 37664 16356 37670
rect 16304 37606 16356 37612
rect 16408 35154 16436 37946
rect 16500 37466 16528 37946
rect 16580 37800 16632 37806
rect 16578 37768 16580 37777
rect 16632 37768 16634 37777
rect 16578 37703 16634 37712
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16580 37460 16632 37466
rect 16580 37402 16632 37408
rect 16592 37346 16620 37402
rect 16500 37318 16620 37346
rect 16500 37194 16528 37318
rect 16488 37188 16540 37194
rect 16488 37130 16540 37136
rect 16500 36718 16528 37130
rect 16488 36712 16540 36718
rect 16488 36654 16540 36660
rect 16500 36242 16528 36654
rect 16488 36236 16540 36242
rect 16488 36178 16540 36184
rect 16488 36032 16540 36038
rect 16488 35974 16540 35980
rect 16396 35148 16448 35154
rect 16396 35090 16448 35096
rect 15752 34672 15804 34678
rect 15752 34614 15804 34620
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 14280 34128 14332 34134
rect 14280 34070 14332 34076
rect 14568 33658 14596 34342
rect 15764 34202 15792 34614
rect 15752 34196 15804 34202
rect 15752 34138 15804 34144
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14568 33454 14596 33594
rect 14556 33448 14608 33454
rect 14556 33390 14608 33396
rect 14740 33380 14792 33386
rect 14740 33322 14792 33328
rect 14752 32502 14780 33322
rect 14832 33312 14884 33318
rect 14832 33254 14884 33260
rect 14740 32496 14792 32502
rect 14740 32438 14792 32444
rect 14844 32230 14872 33254
rect 15200 32360 15252 32366
rect 15200 32302 15252 32308
rect 14832 32224 14884 32230
rect 14832 32166 14884 32172
rect 15212 31754 15240 32302
rect 15200 31748 15252 31754
rect 15200 31690 15252 31696
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 14462 30152 14518 30161
rect 14462 30087 14464 30096
rect 14516 30087 14518 30096
rect 14464 30058 14516 30064
rect 15028 30054 15056 30670
rect 15212 30598 15240 31690
rect 16212 31680 16264 31686
rect 16212 31622 16264 31628
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15292 30184 15344 30190
rect 15120 30144 15292 30172
rect 15016 30048 15068 30054
rect 15016 29990 15068 29996
rect 14096 29844 14148 29850
rect 14096 29786 14148 29792
rect 13912 29708 13964 29714
rect 13912 29650 13964 29656
rect 13924 28762 13952 29650
rect 15028 29102 15056 29990
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 14188 29028 14240 29034
rect 14188 28970 14240 28976
rect 13912 28756 13964 28762
rect 13912 28698 13964 28704
rect 13728 28620 13780 28626
rect 13728 28562 13780 28568
rect 13556 28082 13676 28098
rect 13556 28076 13688 28082
rect 13556 28070 13636 28076
rect 13636 28018 13688 28024
rect 13740 27674 13768 28562
rect 13924 28490 13952 28698
rect 13912 28484 13964 28490
rect 13912 28426 13964 28432
rect 13924 28014 13952 28426
rect 13912 28008 13964 28014
rect 13912 27950 13964 27956
rect 13728 27668 13780 27674
rect 13728 27610 13780 27616
rect 13176 27124 13228 27130
rect 13176 27066 13228 27072
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 13188 24954 13216 27066
rect 14200 26994 14228 28970
rect 15016 28960 15068 28966
rect 15120 28914 15148 30144
rect 15292 30126 15344 30132
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 15068 28908 15148 28914
rect 15016 28902 15148 28908
rect 15028 28886 15148 28902
rect 15028 27878 15056 28886
rect 15016 27872 15068 27878
rect 15016 27814 15068 27820
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 13176 24948 13228 24954
rect 13176 24890 13228 24896
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 13360 24880 13412 24886
rect 13358 24848 13360 24857
rect 13412 24848 13414 24857
rect 13358 24783 13414 24792
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 13096 23730 13124 24550
rect 13556 24410 13584 24754
rect 14200 24750 14228 24890
rect 14278 24848 14334 24857
rect 14278 24783 14334 24792
rect 14292 24750 14320 24783
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13740 22982 13768 24550
rect 14004 24336 14056 24342
rect 14004 24278 14056 24284
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 14016 22574 14044 24278
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14108 23662 14136 23802
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 13004 21542 13216 21570
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 21010 12480 21286
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 19922 12756 20334
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11808 18086 11836 19654
rect 12164 18896 12216 18902
rect 12164 18838 12216 18844
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 12176 17814 12204 18838
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11256 12918 11284 13262
rect 12268 13190 12296 16390
rect 12360 16114 12388 16526
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12452 15570 12480 18294
rect 12728 17882 12756 19858
rect 12912 18222 12940 20946
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 13004 18034 13032 21542
rect 13188 21486 13216 21542
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13096 21078 13124 21422
rect 13084 21072 13136 21078
rect 13084 21014 13136 21020
rect 13740 20058 13768 22510
rect 14108 21690 14136 23598
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13556 18222 13584 18294
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 12912 18006 13032 18034
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16114 12572 16934
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12636 14482 12664 17614
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12728 15706 12756 15982
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 12544 12782 12572 14214
rect 12728 14006 12756 14758
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 10888 12646 10916 12718
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 11992 12442 12020 12718
rect 12544 12646 12572 12718
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12636 12374 12664 13262
rect 12728 13190 12756 13942
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12624 12368 12676 12374
rect 12624 12310 12676 12316
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 11898 12572 12174
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8312 9450 8340 10066
rect 9140 9722 9168 11222
rect 11348 10266 11376 11494
rect 12636 11218 12664 12106
rect 12728 11898 12756 13126
rect 12912 12714 12940 18006
rect 13188 16250 13216 18090
rect 13464 18086 13492 18158
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13280 16454 13308 16594
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13648 15638 13676 18294
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14108 16590 14136 17070
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13832 15570 13860 16526
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13004 13530 13032 14894
rect 13556 14822 13584 15438
rect 13924 14958 13952 16050
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 13004 12306 13032 13466
rect 13556 12306 13584 14758
rect 13924 14482 13952 14894
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 12912 11898 12940 12038
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12728 11354 12756 11834
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 9048 8498 9076 9454
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9042 10548 9318
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 10520 8430 10548 8978
rect 10968 8560 11020 8566
rect 11072 8514 11100 9862
rect 11348 9722 11376 10202
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11020 8508 11100 8514
rect 10968 8502 11100 8508
rect 10980 8486 11100 8502
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 7478 9444 8230
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8404 6458 8432 7278
rect 9876 6866 9904 7414
rect 10888 6866 10916 7822
rect 10980 7546 11008 8366
rect 11440 7954 11468 8910
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 12268 7002 12296 8978
rect 12360 8498 12388 9046
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12452 8430 12480 9318
rect 12544 8634 12572 9998
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 12636 9178 12664 9386
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12636 8430 12664 8842
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 8022 12664 8366
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7002 12848 7686
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 9876 6254 9904 6802
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 10244 6322 10272 6734
rect 10980 6390 11008 6734
rect 11624 6458 11652 6734
rect 11716 6458 11744 6802
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 13188 6118 13216 9386
rect 13372 8906 13400 9590
rect 13464 9382 13492 12038
rect 13832 11354 13860 14350
rect 14108 11626 14136 15982
rect 14200 15366 14228 24550
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14292 18766 14320 22918
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 14384 19718 14412 22510
rect 14462 21448 14518 21457
rect 14462 21383 14464 21392
rect 14516 21383 14518 21392
rect 14464 21354 14516 21360
rect 14476 21146 14504 21354
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14476 21010 14504 21082
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14752 20806 14780 22918
rect 14844 22710 14872 23598
rect 14832 22704 14884 22710
rect 14832 22646 14884 22652
rect 15028 21010 15056 27814
rect 15396 25702 15424 29990
rect 15936 27532 15988 27538
rect 15936 27474 15988 27480
rect 15948 27130 15976 27474
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 15672 24818 15700 26726
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15212 20874 15240 23190
rect 15764 23118 15792 24142
rect 15856 24070 15884 24210
rect 15948 24070 15976 25638
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 16040 24614 16068 24686
rect 16028 24608 16080 24614
rect 16028 24550 16080 24556
rect 16040 24410 16068 24550
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15844 24064 15896 24070
rect 15844 24006 15896 24012
rect 15936 24064 15988 24070
rect 15936 24006 15988 24012
rect 15856 23594 15884 24006
rect 16040 23798 16068 24346
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 15844 23588 15896 23594
rect 15844 23530 15896 23536
rect 15856 23497 15884 23530
rect 15842 23488 15898 23497
rect 15842 23423 15898 23432
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 19990 14780 20742
rect 15304 20398 15332 20878
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14464 18624 14516 18630
rect 14462 18592 14464 18601
rect 14516 18592 14518 18601
rect 14462 18527 14518 18536
rect 14844 18426 14872 20198
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14384 16726 14412 17070
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 10674 13860 11086
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 9110 13492 9318
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 14200 8838 14228 14758
rect 14292 13326 14320 16526
rect 14384 15706 14412 16662
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 14618 14412 14894
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14384 12306 14412 14554
rect 14476 14482 14504 15438
rect 14936 14822 14964 19654
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15028 17202 15056 18158
rect 15212 18086 15240 18362
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15120 16794 15148 17478
rect 15488 17134 15516 22918
rect 15764 22574 15792 23054
rect 15752 22568 15804 22574
rect 15752 22510 15804 22516
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15580 19378 15608 19790
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 18154 15792 18566
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15120 16046 15148 16730
rect 15212 16726 15240 17002
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15212 16046 15240 16662
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15580 15570 15608 16934
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16040 15570 16068 16186
rect 16224 15570 16252 31622
rect 16408 31210 16436 35090
rect 16500 35086 16528 35974
rect 16488 35080 16540 35086
rect 16488 35022 16540 35028
rect 16500 31754 16528 35022
rect 16580 34944 16632 34950
rect 16684 34932 16712 38830
rect 16856 38752 16908 38758
rect 16856 38694 16908 38700
rect 16868 37806 16896 38694
rect 17420 38554 17448 39510
rect 18248 39506 18276 40326
rect 18236 39500 18288 39506
rect 18236 39442 18288 39448
rect 18432 39302 18460 40326
rect 19996 40118 20024 42842
rect 23112 42764 23164 42770
rect 23112 42706 23164 42712
rect 20260 42084 20312 42090
rect 20260 42026 20312 42032
rect 20272 41818 20300 42026
rect 23124 42022 23152 42706
rect 23388 42696 23440 42702
rect 23388 42638 23440 42644
rect 23296 42560 23348 42566
rect 23296 42502 23348 42508
rect 23308 42362 23336 42502
rect 23296 42356 23348 42362
rect 23296 42298 23348 42304
rect 23308 42158 23336 42298
rect 23296 42152 23348 42158
rect 23296 42094 23348 42100
rect 23400 42106 23428 42638
rect 23492 42294 23520 43046
rect 23860 42702 23888 43590
rect 24228 43178 24256 43794
rect 25608 43654 25636 43794
rect 29000 43784 29052 43790
rect 29000 43726 29052 43732
rect 25596 43648 25648 43654
rect 25596 43590 25648 43596
rect 24216 43172 24268 43178
rect 24216 43114 24268 43120
rect 25228 43104 25280 43110
rect 25228 43046 25280 43052
rect 25240 42906 25268 43046
rect 25228 42900 25280 42906
rect 25228 42842 25280 42848
rect 25240 42770 25268 42842
rect 25608 42838 25636 43590
rect 26976 43240 27028 43246
rect 26976 43182 27028 43188
rect 26516 43104 26568 43110
rect 26516 43046 26568 43052
rect 25596 42832 25648 42838
rect 25596 42774 25648 42780
rect 25228 42764 25280 42770
rect 25228 42706 25280 42712
rect 23848 42696 23900 42702
rect 23848 42638 23900 42644
rect 23572 42560 23624 42566
rect 23572 42502 23624 42508
rect 23480 42288 23532 42294
rect 23480 42230 23532 42236
rect 23584 42226 23612 42502
rect 23664 42356 23716 42362
rect 23664 42298 23716 42304
rect 23572 42220 23624 42226
rect 23572 42162 23624 42168
rect 23400 42078 23520 42106
rect 23112 42016 23164 42022
rect 23112 41958 23164 41964
rect 20260 41812 20312 41818
rect 20260 41754 20312 41760
rect 23492 41682 23520 42078
rect 23572 42016 23624 42022
rect 23572 41958 23624 41964
rect 23388 41676 23440 41682
rect 23388 41618 23440 41624
rect 23480 41676 23532 41682
rect 23480 41618 23532 41624
rect 23400 41274 23428 41618
rect 23584 41614 23612 41958
rect 23572 41608 23624 41614
rect 23572 41550 23624 41556
rect 23480 41472 23532 41478
rect 23676 41426 23704 42298
rect 23756 42084 23808 42090
rect 23756 42026 23808 42032
rect 23768 41818 23796 42026
rect 23756 41812 23808 41818
rect 23756 41754 23808 41760
rect 23480 41414 23532 41420
rect 23388 41268 23440 41274
rect 23388 41210 23440 41216
rect 20904 41064 20956 41070
rect 20904 41006 20956 41012
rect 19984 40112 20036 40118
rect 19984 40054 20036 40060
rect 19340 39976 19392 39982
rect 19340 39918 19392 39924
rect 19352 39438 19380 39918
rect 19996 39914 20024 40054
rect 19984 39908 20036 39914
rect 19984 39850 20036 39856
rect 20444 39840 20496 39846
rect 20444 39782 20496 39788
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19340 39432 19392 39438
rect 19340 39374 19392 39380
rect 18052 39296 18104 39302
rect 18052 39238 18104 39244
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18972 39296 19024 39302
rect 18972 39238 19024 39244
rect 18064 38894 18092 39238
rect 18984 38894 19012 39238
rect 20456 39030 20484 39782
rect 20444 39024 20496 39030
rect 20444 38966 20496 38972
rect 19340 38956 19392 38962
rect 19340 38898 19392 38904
rect 18052 38888 18104 38894
rect 18052 38830 18104 38836
rect 18972 38888 19024 38894
rect 18972 38830 19024 38836
rect 17408 38548 17460 38554
rect 17408 38490 17460 38496
rect 16948 38276 17000 38282
rect 16948 38218 17000 38224
rect 16856 37800 16908 37806
rect 16856 37742 16908 37748
rect 16960 37330 16988 38218
rect 18420 38208 18472 38214
rect 18420 38150 18472 38156
rect 18432 37942 18460 38150
rect 18420 37936 18472 37942
rect 18420 37878 18472 37884
rect 17684 37800 17736 37806
rect 17684 37742 17736 37748
rect 17696 37330 17724 37742
rect 17776 37392 17828 37398
rect 17776 37334 17828 37340
rect 16948 37324 17000 37330
rect 16948 37266 17000 37272
rect 17684 37324 17736 37330
rect 17684 37266 17736 37272
rect 17224 36712 17276 36718
rect 17224 36654 17276 36660
rect 17236 36378 17264 36654
rect 17224 36372 17276 36378
rect 17224 36314 17276 36320
rect 16764 36304 16816 36310
rect 16764 36246 16816 36252
rect 16776 36174 16804 36246
rect 16764 36168 16816 36174
rect 16764 36110 16816 36116
rect 16764 36032 16816 36038
rect 16764 35974 16816 35980
rect 16632 34904 16712 34932
rect 16580 34886 16632 34892
rect 16488 31748 16540 31754
rect 16488 31690 16540 31696
rect 16500 31278 16528 31690
rect 16488 31272 16540 31278
rect 16488 31214 16540 31220
rect 16396 31204 16448 31210
rect 16396 31146 16448 31152
rect 16304 30796 16356 30802
rect 16304 30738 16356 30744
rect 16316 30394 16344 30738
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16592 29782 16620 34886
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 16684 32026 16712 33050
rect 16672 32020 16724 32026
rect 16672 31962 16724 31968
rect 16776 30802 16804 35974
rect 17224 33040 17276 33046
rect 17224 32982 17276 32988
rect 17236 32570 17264 32982
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 17788 30870 17816 37334
rect 18432 37330 18460 37878
rect 18984 37806 19012 38830
rect 19248 38548 19300 38554
rect 19248 38490 19300 38496
rect 19260 38457 19288 38490
rect 19246 38448 19302 38457
rect 19246 38383 19302 38392
rect 18972 37800 19024 37806
rect 18972 37742 19024 37748
rect 19248 37800 19300 37806
rect 19248 37742 19300 37748
rect 19260 37398 19288 37742
rect 19248 37392 19300 37398
rect 19248 37334 19300 37340
rect 18420 37324 18472 37330
rect 18420 37266 18472 37272
rect 18236 36916 18288 36922
rect 18236 36858 18288 36864
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 18064 32774 18092 32846
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 18064 32065 18092 32710
rect 18050 32056 18106 32065
rect 18050 31991 18052 32000
rect 18104 31991 18106 32000
rect 18052 31962 18104 31968
rect 18064 31822 18092 31962
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 18064 30870 18092 31282
rect 17776 30864 17828 30870
rect 17776 30806 17828 30812
rect 18052 30864 18104 30870
rect 18052 30806 18104 30812
rect 16764 30796 16816 30802
rect 16764 30738 16816 30744
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 16684 30054 16712 30534
rect 17224 30320 17276 30326
rect 17224 30262 17276 30268
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16672 30048 16724 30054
rect 16672 29990 16724 29996
rect 16580 29776 16632 29782
rect 16580 29718 16632 29724
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16592 28558 16620 29446
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16396 28008 16448 28014
rect 16396 27950 16448 27956
rect 16408 27538 16436 27950
rect 16592 27946 16620 28494
rect 16684 28150 16712 29990
rect 16776 29170 16804 30194
rect 17236 30122 17264 30262
rect 18248 30258 18276 36858
rect 18432 36786 18460 37266
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 19352 36582 19380 38898
rect 20812 38752 20864 38758
rect 20812 38694 20864 38700
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 20536 38412 20588 38418
rect 20536 38354 20588 38360
rect 20548 38010 20576 38354
rect 20536 38004 20588 38010
rect 20536 37946 20588 37952
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 20824 37330 20852 38694
rect 20916 37330 20944 41006
rect 21732 40928 21784 40934
rect 21732 40870 21784 40876
rect 21180 38956 21232 38962
rect 21180 38898 21232 38904
rect 21192 38758 21220 38898
rect 21180 38752 21232 38758
rect 21180 38694 21232 38700
rect 21192 38593 21220 38694
rect 21178 38584 21234 38593
rect 21178 38519 21234 38528
rect 21192 37942 21220 38519
rect 21180 37936 21232 37942
rect 21180 37878 21232 37884
rect 21088 37460 21140 37466
rect 21088 37402 21140 37408
rect 20812 37324 20864 37330
rect 20812 37266 20864 37272
rect 20904 37324 20956 37330
rect 20904 37266 20956 37272
rect 21100 36718 21128 37402
rect 21364 37120 21416 37126
rect 21364 37062 21416 37068
rect 21376 36854 21404 37062
rect 21364 36848 21416 36854
rect 21364 36790 21416 36796
rect 21744 36718 21772 40870
rect 23400 40118 23428 41210
rect 23388 40112 23440 40118
rect 23388 40054 23440 40060
rect 23492 39982 23520 41414
rect 23584 41398 23704 41426
rect 23584 40050 23612 41398
rect 23664 41064 23716 41070
rect 23664 41006 23716 41012
rect 23676 40662 23704 41006
rect 23664 40656 23716 40662
rect 23664 40598 23716 40604
rect 23572 40044 23624 40050
rect 23572 39986 23624 39992
rect 23480 39976 23532 39982
rect 23480 39918 23532 39924
rect 23572 39908 23624 39914
rect 23572 39850 23624 39856
rect 23296 39840 23348 39846
rect 23296 39782 23348 39788
rect 23308 39506 23336 39782
rect 23584 39506 23612 39850
rect 23296 39500 23348 39506
rect 23296 39442 23348 39448
rect 23572 39500 23624 39506
rect 23572 39442 23624 39448
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 22284 38480 22336 38486
rect 22284 38422 22336 38428
rect 21824 37324 21876 37330
rect 21824 37266 21876 37272
rect 19892 36712 19944 36718
rect 20168 36712 20220 36718
rect 19944 36660 20024 36666
rect 19892 36654 20024 36660
rect 20168 36654 20220 36660
rect 21088 36712 21140 36718
rect 21088 36654 21140 36660
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 19904 36638 20024 36654
rect 19340 36576 19392 36582
rect 19340 36518 19392 36524
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19996 34542 20024 36638
rect 20180 36582 20208 36654
rect 20168 36576 20220 36582
rect 20168 36518 20220 36524
rect 20720 36576 20772 36582
rect 20720 36518 20772 36524
rect 21548 36576 21600 36582
rect 21548 36518 21600 36524
rect 20732 35698 20760 36518
rect 20996 36168 21048 36174
rect 20996 36110 21048 36116
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 21008 36038 21036 36110
rect 20996 36032 21048 36038
rect 20996 35974 21048 35980
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 21008 35630 21036 35974
rect 20996 35624 21048 35630
rect 20996 35566 21048 35572
rect 20720 35080 20772 35086
rect 20720 35022 20772 35028
rect 19984 34536 20036 34542
rect 19984 34478 20036 34484
rect 20628 34536 20680 34542
rect 20732 34490 20760 35022
rect 20680 34484 20760 34490
rect 20628 34478 20760 34484
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 18880 34060 18932 34066
rect 18880 34002 18932 34008
rect 18696 33992 18748 33998
rect 18696 33934 18748 33940
rect 18708 33658 18736 33934
rect 18696 33652 18748 33658
rect 18696 33594 18748 33600
rect 18708 32978 18736 33594
rect 18696 32972 18748 32978
rect 18696 32914 18748 32920
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18420 32496 18472 32502
rect 18420 32438 18472 32444
rect 18432 31872 18460 32438
rect 18616 32366 18644 32846
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18788 32224 18840 32230
rect 18892 32178 18920 34002
rect 19352 33658 19380 34342
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19708 34060 19760 34066
rect 19444 34020 19708 34048
rect 19340 33652 19392 33658
rect 19340 33594 19392 33600
rect 19352 33454 19380 33594
rect 19340 33448 19392 33454
rect 19340 33390 19392 33396
rect 19340 33312 19392 33318
rect 19340 33254 19392 33260
rect 19248 32972 19300 32978
rect 19248 32914 19300 32920
rect 19260 32774 19288 32914
rect 19248 32768 19300 32774
rect 19248 32710 19300 32716
rect 18970 32600 19026 32609
rect 18970 32535 19026 32544
rect 18984 32502 19012 32535
rect 18972 32496 19024 32502
rect 19260 32450 19288 32710
rect 18972 32438 19024 32444
rect 18840 32172 18920 32178
rect 18788 32166 18920 32172
rect 18800 32150 18920 32166
rect 18512 31884 18564 31890
rect 18432 31844 18512 31872
rect 18512 31826 18564 31832
rect 18892 30802 18920 32150
rect 18984 30870 19012 32438
rect 19076 32422 19288 32450
rect 18972 30864 19024 30870
rect 18972 30806 19024 30812
rect 18880 30796 18932 30802
rect 18880 30738 18932 30744
rect 19076 30666 19104 32422
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19168 30870 19196 31826
rect 19246 31512 19302 31521
rect 19246 31447 19248 31456
rect 19300 31447 19302 31456
rect 19248 31418 19300 31424
rect 19156 30864 19208 30870
rect 19156 30806 19208 30812
rect 19064 30660 19116 30666
rect 19064 30602 19116 30608
rect 19352 30326 19380 33254
rect 19444 32978 19472 34020
rect 19708 34002 19760 34008
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19432 32972 19484 32978
rect 19432 32914 19484 32920
rect 19444 32502 19472 32914
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19432 32360 19484 32366
rect 19708 32360 19760 32366
rect 19432 32302 19484 32308
rect 19522 32328 19578 32337
rect 19444 31346 19472 32302
rect 19760 32320 19932 32348
rect 19708 32302 19760 32308
rect 19522 32263 19524 32272
rect 19576 32263 19578 32272
rect 19524 32234 19576 32240
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19708 31952 19760 31958
rect 19706 31920 19708 31929
rect 19760 31920 19762 31929
rect 19706 31855 19762 31864
rect 19904 31754 19932 32320
rect 19892 31748 19944 31754
rect 19892 31690 19944 31696
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19432 31204 19484 31210
rect 19432 31146 19484 31152
rect 19444 30394 19472 31146
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18420 30252 18472 30258
rect 18420 30194 18472 30200
rect 17224 30116 17276 30122
rect 17224 30058 17276 30064
rect 17236 30025 17264 30058
rect 17512 30054 17540 30194
rect 18326 30152 18382 30161
rect 18052 30116 18104 30122
rect 18326 30087 18328 30096
rect 18052 30058 18104 30064
rect 18380 30087 18382 30096
rect 18328 30058 18380 30064
rect 17500 30048 17552 30054
rect 17222 30016 17278 30025
rect 17500 29990 17552 29996
rect 17222 29951 17278 29960
rect 17512 29850 17540 29990
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 18064 29782 18092 30058
rect 18052 29776 18104 29782
rect 18052 29718 18104 29724
rect 17316 29708 17368 29714
rect 17316 29650 17368 29656
rect 18144 29708 18196 29714
rect 18144 29650 18196 29656
rect 17328 29510 17356 29650
rect 17500 29572 17552 29578
rect 17500 29514 17552 29520
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 16764 29164 16816 29170
rect 16764 29106 16816 29112
rect 17132 28960 17184 28966
rect 17132 28902 17184 28908
rect 17144 28422 17172 28902
rect 17132 28416 17184 28422
rect 17132 28358 17184 28364
rect 16672 28144 16724 28150
rect 16672 28086 16724 28092
rect 16580 27940 16632 27946
rect 16580 27882 16632 27888
rect 16396 27532 16448 27538
rect 16396 27474 16448 27480
rect 16304 25832 16356 25838
rect 16304 25774 16356 25780
rect 16316 25362 16344 25774
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16408 24682 16436 27474
rect 17144 27470 17172 28358
rect 17328 27606 17356 29446
rect 17512 28626 17540 29514
rect 18156 29306 18184 29650
rect 18432 29594 18460 30194
rect 19340 30184 19392 30190
rect 19340 30126 19392 30132
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18878 30016 18934 30025
rect 18340 29566 18460 29594
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 17500 28620 17552 28626
rect 17500 28562 17552 28568
rect 18340 28218 18368 29566
rect 18420 29504 18472 29510
rect 18420 29446 18472 29452
rect 18432 28966 18460 29446
rect 18708 29238 18736 29990
rect 18878 29951 18934 29960
rect 18892 29782 18920 29951
rect 18880 29776 18932 29782
rect 18880 29718 18932 29724
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 19352 29102 19380 30126
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19708 29776 19760 29782
rect 19892 29776 19944 29782
rect 19760 29736 19892 29764
rect 19708 29718 19760 29724
rect 19892 29718 19944 29724
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 28422 18460 28902
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18328 28212 18380 28218
rect 18328 28154 18380 28160
rect 17316 27600 17368 27606
rect 17316 27542 17368 27548
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 16948 27328 17000 27334
rect 16948 27270 17000 27276
rect 16868 26994 16896 27270
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16856 26784 16908 26790
rect 16960 26772 16988 27270
rect 16908 26744 16988 26772
rect 16856 26726 16908 26732
rect 16868 26586 16896 26726
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 17144 26450 17172 27406
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17880 26518 17908 27270
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17868 26512 17920 26518
rect 17868 26454 17920 26460
rect 17132 26444 17184 26450
rect 17132 26386 17184 26392
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16684 25974 16712 26318
rect 16672 25968 16724 25974
rect 16672 25910 16724 25916
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16396 24676 16448 24682
rect 16396 24618 16448 24624
rect 16500 24410 16528 25230
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 16868 24274 16896 24550
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16684 21486 16712 22374
rect 16776 22098 16804 24142
rect 16960 23866 16988 24686
rect 16948 23860 17000 23866
rect 16948 23802 17000 23808
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17236 21690 17264 21966
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 21010 16712 21422
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16776 21010 16804 21354
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16776 20602 16804 20946
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16776 19854 16804 19994
rect 16960 19854 16988 20266
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16776 19514 16804 19790
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16408 18222 16436 18770
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 16726 16528 17614
rect 16684 17134 16712 18022
rect 16776 17270 16804 19450
rect 17052 18630 17080 19858
rect 17604 19310 17632 26454
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17788 24206 17816 26250
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17880 23526 17908 25298
rect 17972 24070 18000 25774
rect 18144 25696 18196 25702
rect 18144 25638 18196 25644
rect 18156 25430 18184 25638
rect 18144 25424 18196 25430
rect 18144 25366 18196 25372
rect 18156 24682 18184 25366
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18340 24818 18368 25094
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17880 23186 17908 23462
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17040 18624 17092 18630
rect 17132 18624 17184 18630
rect 17040 18566 17092 18572
rect 17130 18592 17132 18601
rect 17184 18592 17186 18601
rect 17052 17678 17080 18566
rect 17130 18527 17186 18536
rect 17880 18086 17908 19110
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16672 17128 16724 17134
rect 16724 17088 16804 17116
rect 16672 17070 16724 17076
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16776 16658 16804 17088
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16316 16182 16344 16458
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 15028 13938 15056 14758
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14476 10606 14504 11290
rect 14568 11218 14596 11562
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 15028 10266 15056 11834
rect 15212 10810 15240 15370
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15672 14618 15700 14894
rect 16224 14618 16252 15506
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16224 13938 16252 14554
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11354 15424 11630
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15304 10690 15332 11018
rect 15212 10662 15332 10690
rect 15212 10470 15240 10662
rect 16224 10606 16252 11086
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 15028 7546 15056 10202
rect 15212 9586 15240 10406
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15580 9586 15608 9998
rect 16224 9586 16252 10542
rect 16408 10266 16436 16594
rect 16868 15638 16896 17274
rect 17512 16794 17540 17546
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 16948 16584 17000 16590
rect 17000 16532 17816 16538
rect 16948 16526 17816 16532
rect 16960 16522 17816 16526
rect 16960 16516 17828 16522
rect 16960 16510 17776 16516
rect 17776 16458 17828 16464
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 17144 15706 17172 15914
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 13802 16712 14758
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16684 13462 16712 13738
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16672 12300 16724 12306
rect 16776 12288 16804 13738
rect 16724 12260 16804 12288
rect 16672 12242 16724 12248
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 15212 9042 15240 9522
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 16132 8498 16160 9522
rect 16224 9178 16252 9522
rect 16408 9518 16436 10202
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16500 8634 16528 10406
rect 16868 9450 16896 15302
rect 17880 14822 17908 18022
rect 17972 17746 18000 24006
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 18064 23662 18092 23802
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 19786 18184 20198
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 18156 18902 18184 19722
rect 18432 18970 18460 28358
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18616 22166 18644 22374
rect 18604 22160 18656 22166
rect 18602 22128 18604 22137
rect 18656 22128 18658 22137
rect 18602 22063 18658 22072
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18524 18290 18552 18702
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18708 17898 18736 22442
rect 19352 21690 19380 29038
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19892 28416 19944 28422
rect 19892 28358 19944 28364
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19444 27878 19472 28018
rect 19904 28014 19932 28358
rect 19892 28008 19944 28014
rect 19892 27950 19944 27956
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19444 25770 19472 27814
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19432 25764 19484 25770
rect 19432 25706 19484 25712
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19444 23866 19472 24754
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19996 22250 20024 34478
rect 20640 34462 20760 34478
rect 21284 34474 21312 36110
rect 21364 35556 21416 35562
rect 21364 35498 21416 35504
rect 21376 35290 21404 35498
rect 21364 35284 21416 35290
rect 21364 35226 21416 35232
rect 21376 34542 21404 35226
rect 21364 34536 21416 34542
rect 21560 34524 21588 36518
rect 21744 35766 21772 36654
rect 21732 35760 21784 35766
rect 21732 35702 21784 35708
rect 21836 35154 21864 37266
rect 22008 36032 22060 36038
rect 22008 35974 22060 35980
rect 22020 35494 22048 35974
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 21732 35148 21784 35154
rect 21732 35090 21784 35096
rect 21824 35148 21876 35154
rect 21824 35090 21876 35096
rect 21744 34542 21772 35090
rect 21364 34478 21416 34484
rect 21468 34496 21588 34524
rect 21732 34536 21784 34542
rect 21272 34468 21324 34474
rect 21272 34410 21324 34416
rect 20260 34400 20312 34406
rect 20260 34342 20312 34348
rect 20168 34060 20220 34066
rect 20168 34002 20220 34008
rect 20180 33862 20208 34002
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 20180 33658 20208 33798
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 20076 33448 20128 33454
rect 20076 33390 20128 33396
rect 20088 32570 20116 33390
rect 20168 32904 20220 32910
rect 20168 32846 20220 32852
rect 20076 32564 20128 32570
rect 20076 32506 20128 32512
rect 20180 31346 20208 32846
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20272 29306 20300 34342
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20640 33862 20668 33934
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20640 33386 20668 33798
rect 20628 33380 20680 33386
rect 20628 33322 20680 33328
rect 21364 32972 21416 32978
rect 21468 32960 21496 34496
rect 21732 34478 21784 34484
rect 21836 34406 21864 35090
rect 22008 35080 22060 35086
rect 22008 35022 22060 35028
rect 21824 34400 21876 34406
rect 21824 34342 21876 34348
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 21548 34060 21600 34066
rect 21548 34002 21600 34008
rect 21560 32978 21588 34002
rect 21416 32932 21496 32960
rect 21548 32972 21600 32978
rect 21364 32914 21416 32920
rect 21548 32914 21600 32920
rect 20352 32768 20404 32774
rect 20352 32710 20404 32716
rect 20364 31958 20392 32710
rect 21836 32450 21864 34138
rect 22020 32978 22048 35022
rect 22008 32972 22060 32978
rect 22008 32914 22060 32920
rect 21468 32422 21864 32450
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 20352 31952 20404 31958
rect 20352 31894 20404 31900
rect 21008 31890 21036 32166
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 20536 31816 20588 31822
rect 20536 31758 20588 31764
rect 20350 30968 20406 30977
rect 20350 30903 20352 30912
rect 20404 30903 20406 30912
rect 20444 30932 20496 30938
rect 20352 30874 20404 30880
rect 20444 30874 20496 30880
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20272 28762 20300 29242
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20456 24188 20484 30874
rect 20548 24818 20576 31758
rect 20628 31272 20680 31278
rect 20628 31214 20680 31220
rect 20640 29510 20668 31214
rect 20996 31204 21048 31210
rect 20996 31146 21048 31152
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20640 27470 20668 29446
rect 21008 28218 21036 31146
rect 21088 30320 21140 30326
rect 21088 30262 21140 30268
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20732 24698 20760 28154
rect 20996 27940 21048 27946
rect 20996 27882 21048 27888
rect 21008 27538 21036 27882
rect 20996 27532 21048 27538
rect 20996 27474 21048 27480
rect 21100 26926 21128 30262
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 20824 25498 20852 26862
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 19904 22222 20024 22250
rect 20088 24160 20484 24188
rect 20640 24670 20760 24698
rect 19904 22114 19932 22222
rect 19812 22086 19932 22114
rect 19812 21894 19840 22086
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18800 20534 18828 21422
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18800 20330 18828 20470
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 18800 18766 18828 20266
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18984 18154 19012 18770
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18708 17870 18828 17898
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17972 15570 18000 16730
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16960 14074 16988 14282
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17052 12306 17080 12582
rect 17144 12442 17172 13262
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17788 11014 17816 13806
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18156 12306 18184 12582
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 11218 18644 11494
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 17960 11144 18012 11150
rect 17880 11104 17960 11132
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16592 8430 16620 9046
rect 17880 8838 17908 11104
rect 17960 11086 18012 11092
rect 18708 9110 18736 17750
rect 18800 14006 18828 17870
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 19076 13870 19104 14214
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19168 13734 19196 20198
rect 19444 19310 19472 20266
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19444 17678 19472 18770
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19996 16726 20024 20266
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 20088 16182 20116 24160
rect 20640 20602 20668 24670
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20732 24206 20760 24550
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20732 23254 20760 24142
rect 20720 23248 20772 23254
rect 20720 23190 20772 23196
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20180 18902 20208 20334
rect 20640 19514 20668 20538
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20732 17746 20760 21966
rect 20824 21486 20852 22510
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20916 17746 20944 19450
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 16658 20944 17478
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19352 14074 19380 14962
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 20548 13462 20576 15914
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 20536 13456 20588 13462
rect 20536 13398 20588 13404
rect 19352 12986 19380 13398
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 20640 10198 20668 16390
rect 20824 16114 20852 16594
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 21008 16046 21036 24278
rect 21100 22982 21128 26862
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 21100 22506 21128 22918
rect 21192 22710 21220 23054
rect 21180 22704 21232 22710
rect 21180 22646 21232 22652
rect 21088 22500 21140 22506
rect 21088 22442 21140 22448
rect 21468 22114 21496 32422
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21548 31884 21600 31890
rect 21548 31826 21600 31832
rect 21560 31346 21588 31826
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 21548 31136 21600 31142
rect 21548 31078 21600 31084
rect 21560 30190 21588 31078
rect 21640 30864 21692 30870
rect 21640 30806 21692 30812
rect 21652 30258 21680 30806
rect 21640 30252 21692 30258
rect 21640 30194 21692 30200
rect 21548 30184 21600 30190
rect 21548 30126 21600 30132
rect 21560 26926 21588 30126
rect 21548 26920 21600 26926
rect 21548 26862 21600 26868
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21560 26450 21588 26726
rect 21548 26444 21600 26450
rect 21548 26386 21600 26392
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21376 22086 21496 22114
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 21100 21894 21128 21966
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21100 20942 21128 21830
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21100 20534 21128 20878
rect 21192 20602 21220 21898
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21284 21350 21312 21490
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 21192 20398 21220 20538
rect 21180 20392 21232 20398
rect 21180 20334 21232 20340
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21192 18358 21220 18770
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21192 18154 21220 18294
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 21192 17338 21220 18090
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 21100 16658 21128 17002
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21192 16250 21220 16594
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 14618 20760 14962
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20824 13530 20852 15846
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21100 14618 21128 15642
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20732 11694 20760 11834
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20824 9654 20852 13466
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21192 12374 21220 12786
rect 21180 12368 21232 12374
rect 21180 12310 21232 12316
rect 21284 12102 21312 21286
rect 21376 20058 21404 22086
rect 21652 22030 21680 22510
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21744 18630 21772 32302
rect 22296 31958 22324 38422
rect 22468 35760 22520 35766
rect 22468 35702 22520 35708
rect 22480 35222 22508 35702
rect 22940 35630 22968 39374
rect 23572 38820 23624 38826
rect 23572 38762 23624 38768
rect 22928 35624 22980 35630
rect 22928 35566 22980 35572
rect 22468 35216 22520 35222
rect 22468 35158 22520 35164
rect 23584 33402 23612 38762
rect 23676 36038 23704 40598
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35154 23704 35974
rect 23664 35148 23716 35154
rect 23664 35090 23716 35096
rect 23492 33374 23612 33402
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22284 31952 22336 31958
rect 22284 31894 22336 31900
rect 22652 30864 22704 30870
rect 22652 30806 22704 30812
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22204 26586 22232 26930
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 22574 21956 23462
rect 21916 22568 21968 22574
rect 21916 22510 21968 22516
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 22100 21480 22152 21486
rect 22100 21422 22152 21428
rect 22020 20806 22048 21422
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22020 20534 22048 20742
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 22112 20466 22140 21422
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 14414 21496 17614
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21376 13530 21404 13806
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21560 12986 21588 18022
rect 22296 17626 22324 27406
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 22388 26586 22416 26726
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22388 22166 22416 26522
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22480 23662 22508 24074
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22572 23526 22600 23557
rect 22560 23520 22612 23526
rect 22558 23488 22560 23497
rect 22612 23488 22614 23497
rect 22558 23423 22614 23432
rect 22572 23254 22600 23423
rect 22560 23248 22612 23254
rect 22560 23190 22612 23196
rect 22664 22982 22692 30806
rect 22756 30190 22784 32506
rect 23492 32026 23520 33374
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23480 32020 23532 32026
rect 23480 31962 23532 31968
rect 23480 30728 23532 30734
rect 23480 30670 23532 30676
rect 23492 30258 23520 30670
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 22744 30184 22796 30190
rect 22744 30126 22796 30132
rect 22756 30054 22784 30126
rect 22744 30048 22796 30054
rect 22744 29990 22796 29996
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22376 22160 22428 22166
rect 22376 22102 22428 22108
rect 22664 21622 22692 22918
rect 22652 21616 22704 21622
rect 22652 21558 22704 21564
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22664 21010 22692 21354
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22756 20602 22784 29990
rect 23584 27334 23612 33254
rect 23768 32434 23796 39238
rect 23860 39030 23888 42638
rect 24584 42356 24636 42362
rect 24584 42298 24636 42304
rect 25412 42356 25464 42362
rect 25412 42298 25464 42304
rect 23940 42288 23992 42294
rect 23940 42230 23992 42236
rect 23952 41750 23980 42230
rect 24596 42158 24624 42298
rect 24584 42152 24636 42158
rect 24584 42094 24636 42100
rect 23940 41744 23992 41750
rect 23940 41686 23992 41692
rect 24676 41744 24728 41750
rect 24676 41686 24728 41692
rect 24492 41676 24544 41682
rect 24492 41618 24544 41624
rect 23940 41540 23992 41546
rect 23940 41482 23992 41488
rect 23952 41274 23980 41482
rect 24504 41478 24532 41618
rect 24492 41472 24544 41478
rect 24492 41414 24544 41420
rect 23940 41268 23992 41274
rect 23940 41210 23992 41216
rect 24124 41064 24176 41070
rect 24124 41006 24176 41012
rect 24136 40934 24164 41006
rect 24124 40928 24176 40934
rect 24124 40870 24176 40876
rect 23940 40384 23992 40390
rect 23940 40326 23992 40332
rect 23952 39506 23980 40326
rect 24504 40066 24532 41414
rect 24688 41070 24716 41686
rect 25424 41682 25452 42298
rect 25412 41676 25464 41682
rect 25412 41618 25464 41624
rect 25608 41478 25636 42774
rect 26528 42566 26556 43046
rect 26988 42702 27016 43182
rect 29012 42770 29040 43726
rect 36820 43716 36872 43722
rect 36820 43658 36872 43664
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 36832 43450 36860 43658
rect 37648 43648 37700 43654
rect 37648 43590 37700 43596
rect 36820 43444 36872 43450
rect 36820 43386 36872 43392
rect 29092 43308 29144 43314
rect 29092 43250 29144 43256
rect 30472 43308 30524 43314
rect 30472 43250 30524 43256
rect 29104 42770 29132 43250
rect 29736 43172 29788 43178
rect 29736 43114 29788 43120
rect 29000 42764 29052 42770
rect 29000 42706 29052 42712
rect 29092 42764 29144 42770
rect 29092 42706 29144 42712
rect 26976 42696 27028 42702
rect 26976 42638 27028 42644
rect 26516 42560 26568 42566
rect 26516 42502 26568 42508
rect 25872 42220 25924 42226
rect 25872 42162 25924 42168
rect 25688 42152 25740 42158
rect 25688 42094 25740 42100
rect 25700 42022 25728 42094
rect 25884 42022 25912 42162
rect 25688 42016 25740 42022
rect 25688 41958 25740 41964
rect 25872 42016 25924 42022
rect 25872 41958 25924 41964
rect 25700 41750 25728 41958
rect 25688 41744 25740 41750
rect 25688 41686 25740 41692
rect 26240 41676 26292 41682
rect 26240 41618 26292 41624
rect 25504 41472 25556 41478
rect 25504 41414 25556 41420
rect 25596 41472 25648 41478
rect 25596 41414 25648 41420
rect 25516 41138 25544 41414
rect 26252 41206 26280 41618
rect 26528 41546 26556 42502
rect 27252 42084 27304 42090
rect 27252 42026 27304 42032
rect 26792 41608 26844 41614
rect 26792 41550 26844 41556
rect 26516 41540 26568 41546
rect 26516 41482 26568 41488
rect 26240 41200 26292 41206
rect 26240 41142 26292 41148
rect 25504 41132 25556 41138
rect 25504 41074 25556 41080
rect 24676 41064 24728 41070
rect 24676 41006 24728 41012
rect 24584 40928 24636 40934
rect 24584 40870 24636 40876
rect 25228 40928 25280 40934
rect 25228 40870 25280 40876
rect 24596 40594 24624 40870
rect 24766 40760 24822 40769
rect 24766 40695 24822 40704
rect 24584 40588 24636 40594
rect 24584 40530 24636 40536
rect 24504 40038 24624 40066
rect 24596 39982 24624 40038
rect 24584 39976 24636 39982
rect 24584 39918 24636 39924
rect 23940 39500 23992 39506
rect 23940 39442 23992 39448
rect 23952 39302 23980 39442
rect 23940 39296 23992 39302
rect 23940 39238 23992 39244
rect 23848 39024 23900 39030
rect 23848 38966 23900 38972
rect 23860 38894 23888 38925
rect 24780 38894 24808 40695
rect 25240 40594 25268 40870
rect 25228 40588 25280 40594
rect 25228 40530 25280 40536
rect 25044 40384 25096 40390
rect 25044 40326 25096 40332
rect 24860 40044 24912 40050
rect 24860 39986 24912 39992
rect 24872 39914 24900 39986
rect 24860 39908 24912 39914
rect 24860 39850 24912 39856
rect 24872 39506 24900 39850
rect 25056 39506 25084 40326
rect 25516 40118 25544 41074
rect 26252 41070 26280 41142
rect 26240 41064 26292 41070
rect 26240 41006 26292 41012
rect 25688 40928 25740 40934
rect 25688 40870 25740 40876
rect 25872 40928 25924 40934
rect 25872 40870 25924 40876
rect 25700 40662 25728 40870
rect 25688 40656 25740 40662
rect 25688 40598 25740 40604
rect 25700 40458 25728 40598
rect 25688 40452 25740 40458
rect 25688 40394 25740 40400
rect 25504 40112 25556 40118
rect 25504 40054 25556 40060
rect 25688 40112 25740 40118
rect 25688 40054 25740 40060
rect 24860 39500 24912 39506
rect 24860 39442 24912 39448
rect 25044 39500 25096 39506
rect 25044 39442 25096 39448
rect 23848 38888 23900 38894
rect 23846 38856 23848 38865
rect 24400 38888 24452 38894
rect 23900 38856 23902 38865
rect 24400 38830 24452 38836
rect 24768 38888 24820 38894
rect 25228 38888 25280 38894
rect 24768 38830 24820 38836
rect 25226 38856 25228 38865
rect 25280 38856 25282 38865
rect 23846 38791 23902 38800
rect 23860 38418 23888 38791
rect 24412 38758 24440 38830
rect 25226 38791 25282 38800
rect 24400 38752 24452 38758
rect 23938 38720 23994 38729
rect 24400 38694 24452 38700
rect 24582 38720 24638 38729
rect 23938 38655 23994 38664
rect 23952 38486 23980 38655
rect 23940 38480 23992 38486
rect 23940 38422 23992 38428
rect 24412 38418 24440 38694
rect 24582 38655 24638 38664
rect 24596 38418 24624 38655
rect 23848 38412 23900 38418
rect 23848 38354 23900 38360
rect 24400 38412 24452 38418
rect 24400 38354 24452 38360
rect 24584 38412 24636 38418
rect 24584 38354 24636 38360
rect 25240 38350 25268 38791
rect 25412 38752 25464 38758
rect 25412 38694 25464 38700
rect 25424 38554 25452 38694
rect 25412 38548 25464 38554
rect 25412 38490 25464 38496
rect 25228 38344 25280 38350
rect 25228 38286 25280 38292
rect 24124 38208 24176 38214
rect 24124 38150 24176 38156
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23768 27470 23796 31214
rect 23756 27464 23808 27470
rect 23756 27406 23808 27412
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23584 26042 23612 27270
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 23584 24274 23612 25298
rect 23572 24268 23624 24274
rect 23572 24210 23624 24216
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22756 20398 22784 20538
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23768 18970 23796 20198
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23768 17814 23796 18906
rect 23860 17882 23888 32846
rect 23940 32428 23992 32434
rect 23940 32370 23992 32376
rect 23952 31142 23980 32370
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23952 28014 23980 31078
rect 24044 30870 24072 31282
rect 24032 30864 24084 30870
rect 24032 30806 24084 30812
rect 23940 28008 23992 28014
rect 23940 27950 23992 27956
rect 24136 27538 24164 38150
rect 25504 37800 25556 37806
rect 25504 37742 25556 37748
rect 25412 37732 25464 37738
rect 25412 37674 25464 37680
rect 25424 37466 25452 37674
rect 25516 37670 25544 37742
rect 25504 37664 25556 37670
rect 25504 37606 25556 37612
rect 25412 37460 25464 37466
rect 25412 37402 25464 37408
rect 24768 37188 24820 37194
rect 24768 37130 24820 37136
rect 24676 34400 24728 34406
rect 24676 34342 24728 34348
rect 24400 33448 24452 33454
rect 24400 33390 24452 33396
rect 24412 32978 24440 33390
rect 24400 32972 24452 32978
rect 24400 32914 24452 32920
rect 24492 32972 24544 32978
rect 24492 32914 24544 32920
rect 24216 32904 24268 32910
rect 24216 32846 24268 32852
rect 24228 32774 24256 32846
rect 24216 32768 24268 32774
rect 24216 32710 24268 32716
rect 24504 32434 24532 32914
rect 24492 32428 24544 32434
rect 24492 32370 24544 32376
rect 24688 32230 24716 34342
rect 24780 32366 24808 37130
rect 25424 36854 25452 37402
rect 25412 36848 25464 36854
rect 25412 36790 25464 36796
rect 25424 36718 25452 36790
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 24860 36644 24912 36650
rect 24860 36586 24912 36592
rect 24872 36242 24900 36586
rect 25412 36576 25464 36582
rect 25412 36518 25464 36524
rect 24860 36236 24912 36242
rect 24860 36178 24912 36184
rect 24952 36236 25004 36242
rect 24952 36178 25004 36184
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24768 32360 24820 32366
rect 24766 32328 24768 32337
rect 24820 32328 24822 32337
rect 24766 32263 24822 32272
rect 24676 32224 24728 32230
rect 24676 32166 24728 32172
rect 24584 31680 24636 31686
rect 24584 31622 24636 31628
rect 24492 30320 24544 30326
rect 24492 30262 24544 30268
rect 24504 30190 24532 30262
rect 24596 30190 24624 31622
rect 24688 31278 24716 32166
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 24492 30184 24544 30190
rect 24492 30126 24544 30132
rect 24584 30184 24636 30190
rect 24584 30126 24636 30132
rect 24504 29306 24532 30126
rect 24872 29850 24900 32370
rect 24964 32026 24992 36178
rect 25320 36100 25372 36106
rect 25320 36042 25372 36048
rect 25136 35148 25188 35154
rect 25136 35090 25188 35096
rect 25148 34746 25176 35090
rect 25136 34740 25188 34746
rect 25136 34682 25188 34688
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 25056 33318 25084 33458
rect 25228 33448 25280 33454
rect 25228 33390 25280 33396
rect 25044 33312 25096 33318
rect 25044 33254 25096 33260
rect 25240 32366 25268 33390
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25332 32212 25360 36042
rect 25424 35630 25452 36518
rect 25516 36310 25544 37606
rect 25596 36712 25648 36718
rect 25596 36654 25648 36660
rect 25608 36582 25636 36654
rect 25596 36576 25648 36582
rect 25596 36518 25648 36524
rect 25504 36304 25556 36310
rect 25504 36246 25556 36252
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25240 32184 25360 32212
rect 24952 32020 25004 32026
rect 24952 31962 25004 31968
rect 24964 31906 24992 31962
rect 24964 31890 25084 31906
rect 24952 31884 25084 31890
rect 25004 31878 25084 31884
rect 24952 31826 25004 31832
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24676 29504 24728 29510
rect 24676 29446 24728 29452
rect 24492 29300 24544 29306
rect 24492 29242 24544 29248
rect 24688 29034 24716 29446
rect 24676 29028 24728 29034
rect 24676 28970 24728 28976
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24124 25832 24176 25838
rect 24124 25774 24176 25780
rect 24136 25362 24164 25774
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 24044 23798 24072 25094
rect 24492 24744 24544 24750
rect 24492 24686 24544 24692
rect 24504 24410 24532 24686
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 24136 23254 24164 24210
rect 24216 23520 24268 23526
rect 24216 23462 24268 23468
rect 24124 23248 24176 23254
rect 24124 23190 24176 23196
rect 24228 23100 24256 23462
rect 24136 23072 24256 23100
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23952 20806 23980 21286
rect 23940 20800 23992 20806
rect 23938 20768 23940 20777
rect 23992 20768 23994 20777
rect 23938 20703 23994 20712
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 24044 18630 24072 18770
rect 24136 18698 24164 23072
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 24044 18426 24072 18566
rect 24032 18420 24084 18426
rect 24032 18362 24084 18368
rect 24044 17882 24072 18362
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 23756 17808 23808 17814
rect 23756 17750 23808 17756
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22204 17610 22324 17626
rect 22192 17604 22324 17610
rect 22244 17598 22324 17604
rect 22192 17546 22244 17552
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21744 16658 21772 16934
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21652 16046 21680 16186
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21652 15638 21680 15982
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21744 15026 21772 16594
rect 21836 15570 21864 17274
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21928 16658 21956 16730
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 22112 16130 22140 17478
rect 22388 17134 22416 17682
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 22558 17368 22614 17377
rect 22558 17303 22614 17312
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22572 16998 22600 17303
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 16794 22600 16934
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 22020 16114 22140 16130
rect 22008 16108 22140 16114
rect 22060 16102 22140 16108
rect 22008 16050 22060 16056
rect 21916 16040 21968 16046
rect 21914 16008 21916 16017
rect 22560 16040 22612 16046
rect 21968 16008 21970 16017
rect 22560 15982 22612 15988
rect 21914 15943 21970 15952
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 22020 15706 22048 15914
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 22020 14414 22048 15642
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 22008 13796 22060 13802
rect 22008 13738 22060 13744
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 22020 12714 22048 13738
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 22112 12170 22140 15846
rect 22572 15570 22600 15982
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22940 14550 22968 15846
rect 23308 15502 23336 16390
rect 23676 16046 23704 17614
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 24136 15706 24164 18634
rect 24228 16658 24256 18702
rect 24688 17066 24716 28970
rect 24964 27656 24992 31214
rect 25056 30394 25084 31878
rect 25240 30802 25268 32184
rect 25424 32042 25452 35566
rect 25504 34740 25556 34746
rect 25504 34682 25556 34688
rect 25332 32014 25452 32042
rect 25228 30796 25280 30802
rect 25228 30738 25280 30744
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 25044 30048 25096 30054
rect 25044 29990 25096 29996
rect 25056 29714 25084 29990
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 25240 28014 25268 28358
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 24964 27628 25084 27656
rect 24860 27600 24912 27606
rect 25056 27588 25084 27628
rect 25136 27600 25188 27606
rect 25056 27560 25136 27588
rect 24860 27542 24912 27548
rect 25136 27542 25188 27548
rect 24872 19922 24900 27542
rect 25332 27010 25360 32014
rect 25412 29096 25464 29102
rect 25412 29038 25464 29044
rect 25424 28150 25452 29038
rect 25412 28144 25464 28150
rect 25412 28086 25464 28092
rect 25332 26982 25452 27010
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25148 26602 25176 26726
rect 25148 26574 25268 26602
rect 25240 25702 25268 26574
rect 25332 26042 25360 26862
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 25240 24614 25268 25638
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25044 24132 25096 24138
rect 25044 24074 25096 24080
rect 25056 23186 25084 24074
rect 25240 23526 25268 24550
rect 25332 24274 25360 24550
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 25424 23746 25452 26982
rect 25516 26330 25544 34682
rect 25596 32360 25648 32366
rect 25596 32302 25648 32308
rect 25608 30870 25636 32302
rect 25700 31929 25728 40054
rect 25780 39296 25832 39302
rect 25780 39238 25832 39244
rect 25792 38894 25820 39238
rect 25780 38888 25832 38894
rect 25780 38830 25832 38836
rect 25884 38593 25912 40870
rect 26608 40384 26660 40390
rect 26608 40326 26660 40332
rect 26516 40112 26568 40118
rect 26516 40054 26568 40060
rect 26528 39982 26556 40054
rect 26620 39982 26648 40326
rect 26516 39976 26568 39982
rect 26516 39918 26568 39924
rect 26608 39976 26660 39982
rect 26608 39918 26660 39924
rect 26148 39840 26200 39846
rect 26148 39782 26200 39788
rect 26516 39840 26568 39846
rect 26516 39782 26568 39788
rect 25964 39024 26016 39030
rect 25964 38966 26016 38972
rect 25870 38584 25926 38593
rect 25870 38519 25926 38528
rect 25884 38350 25912 38519
rect 25872 38344 25924 38350
rect 25872 38286 25924 38292
rect 25884 36106 25912 38286
rect 25872 36100 25924 36106
rect 25872 36042 25924 36048
rect 25872 34944 25924 34950
rect 25872 34886 25924 34892
rect 25884 34746 25912 34886
rect 25872 34740 25924 34746
rect 25872 34682 25924 34688
rect 25884 34542 25912 34682
rect 25872 34536 25924 34542
rect 25872 34478 25924 34484
rect 25976 33522 26004 38966
rect 26160 38894 26188 39782
rect 26528 39574 26556 39782
rect 26516 39568 26568 39574
rect 26516 39510 26568 39516
rect 26804 39302 26832 41550
rect 27264 40662 27292 42026
rect 29748 41682 29776 43114
rect 30380 42696 30432 42702
rect 30380 42638 30432 42644
rect 30392 41682 30420 42638
rect 30484 42022 30512 43250
rect 34796 43172 34848 43178
rect 34796 43114 34848 43120
rect 34152 43104 34204 43110
rect 34152 43046 34204 43052
rect 34164 42702 34192 43046
rect 34152 42696 34204 42702
rect 34152 42638 34204 42644
rect 34428 42696 34480 42702
rect 34428 42638 34480 42644
rect 31576 42560 31628 42566
rect 31576 42502 31628 42508
rect 31588 42226 31616 42502
rect 31576 42220 31628 42226
rect 31576 42162 31628 42168
rect 30472 42016 30524 42022
rect 30472 41958 30524 41964
rect 30564 42016 30616 42022
rect 30564 41958 30616 41964
rect 30576 41750 30604 41958
rect 30564 41744 30616 41750
rect 30564 41686 30616 41692
rect 29736 41676 29788 41682
rect 29736 41618 29788 41624
rect 30380 41676 30432 41682
rect 30380 41618 30432 41624
rect 30932 41676 30984 41682
rect 30932 41618 30984 41624
rect 29748 41562 29776 41618
rect 29748 41534 29960 41562
rect 29828 41268 29880 41274
rect 29828 41210 29880 41216
rect 29840 41177 29868 41210
rect 29826 41168 29882 41177
rect 27344 41132 27396 41138
rect 27620 41132 27672 41138
rect 27396 41092 27620 41120
rect 27344 41074 27396 41080
rect 29826 41103 29882 41112
rect 27620 41074 27672 41080
rect 28632 40724 28684 40730
rect 28632 40666 28684 40672
rect 27252 40656 27304 40662
rect 27252 40598 27304 40604
rect 27620 40588 27672 40594
rect 27540 40548 27620 40576
rect 27540 40118 27568 40548
rect 27620 40530 27672 40536
rect 28264 40384 28316 40390
rect 28264 40326 28316 40332
rect 28356 40384 28408 40390
rect 28356 40326 28408 40332
rect 27528 40112 27580 40118
rect 27528 40054 27580 40060
rect 28276 39817 28304 40326
rect 28368 40118 28396 40326
rect 28644 40118 28672 40666
rect 28724 40520 28776 40526
rect 28816 40520 28868 40526
rect 28776 40480 28816 40508
rect 28724 40462 28776 40468
rect 28816 40462 28868 40468
rect 29000 40520 29052 40526
rect 29000 40462 29052 40468
rect 28356 40112 28408 40118
rect 28356 40054 28408 40060
rect 28632 40112 28684 40118
rect 28632 40054 28684 40060
rect 28262 39808 28318 39817
rect 28262 39743 28318 39752
rect 26976 39500 27028 39506
rect 26976 39442 27028 39448
rect 26884 39432 26936 39438
rect 26884 39374 26936 39380
rect 26332 39296 26384 39302
rect 26332 39238 26384 39244
rect 26792 39296 26844 39302
rect 26792 39238 26844 39244
rect 26240 38956 26292 38962
rect 26240 38898 26292 38904
rect 26148 38888 26200 38894
rect 26148 38830 26200 38836
rect 26056 38820 26108 38826
rect 26056 38762 26108 38768
rect 26068 38706 26096 38762
rect 26252 38706 26280 38898
rect 26068 38678 26280 38706
rect 26148 37868 26200 37874
rect 26148 37810 26200 37816
rect 26056 37800 26108 37806
rect 26056 37742 26108 37748
rect 26068 37670 26096 37742
rect 26056 37664 26108 37670
rect 26056 37606 26108 37612
rect 26068 37466 26096 37606
rect 26160 37466 26188 37810
rect 26056 37460 26108 37466
rect 26056 37402 26108 37408
rect 26148 37460 26200 37466
rect 26148 37402 26200 37408
rect 26068 37262 26096 37402
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 26068 35714 26096 37198
rect 26148 36236 26200 36242
rect 26148 36178 26200 36184
rect 26160 35834 26188 36178
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26148 35828 26200 35834
rect 26148 35770 26200 35776
rect 26068 35686 26188 35714
rect 26056 33652 26108 33658
rect 26056 33594 26108 33600
rect 26068 33522 26096 33594
rect 25964 33516 26016 33522
rect 25964 33458 26016 33464
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 25872 33448 25924 33454
rect 25872 33390 25924 33396
rect 25780 33312 25832 33318
rect 25780 33254 25832 33260
rect 25792 33114 25820 33254
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 25686 31920 25742 31929
rect 25686 31855 25742 31864
rect 25596 30864 25648 30870
rect 25596 30806 25648 30812
rect 25884 29646 25912 33390
rect 26056 33380 26108 33386
rect 26056 33322 26108 33328
rect 25964 33108 26016 33114
rect 25964 33050 26016 33056
rect 25976 30938 26004 33050
rect 26068 32978 26096 33322
rect 26056 32972 26108 32978
rect 26056 32914 26108 32920
rect 25964 30932 26016 30938
rect 25964 30874 26016 30880
rect 25872 29640 25924 29646
rect 25872 29582 25924 29588
rect 25516 26302 25636 26330
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25516 25838 25544 26182
rect 25504 25832 25556 25838
rect 25504 25774 25556 25780
rect 25608 24154 25636 26302
rect 25332 23718 25452 23746
rect 25516 24126 25636 24154
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25240 22642 25268 23462
rect 25332 22778 25360 23718
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 25424 23254 25452 23598
rect 25412 23248 25464 23254
rect 25412 23190 25464 23196
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24780 18222 24808 19722
rect 24872 19242 24900 19858
rect 25042 19272 25098 19281
rect 24860 19236 24912 19242
rect 25042 19207 25098 19216
rect 24860 19178 24912 19184
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24780 18086 24808 18158
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24676 17060 24728 17066
rect 24676 17002 24728 17008
rect 24216 16652 24268 16658
rect 24216 16594 24268 16600
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 24780 15026 24808 18022
rect 24964 17202 24992 19110
rect 25056 18766 25084 19207
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25332 18426 25360 20470
rect 25412 20460 25464 20466
rect 25412 20402 25464 20408
rect 25424 20058 25452 20402
rect 25412 20052 25464 20058
rect 25412 19994 25464 20000
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25424 19281 25452 19858
rect 25410 19272 25466 19281
rect 25410 19207 25466 19216
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25332 18222 25360 18362
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25240 16998 25268 17138
rect 25332 17134 25360 18158
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24872 15337 24900 15370
rect 24858 15328 24914 15337
rect 24858 15263 24914 15272
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 22928 14544 22980 14550
rect 22928 14486 22980 14492
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 24044 13977 24072 14214
rect 24030 13968 24086 13977
rect 24030 13903 24032 13912
rect 24084 13903 24086 13912
rect 24032 13874 24084 13880
rect 22652 13796 22704 13802
rect 22652 13738 22704 13744
rect 22664 13394 22692 13738
rect 24044 13462 24072 13874
rect 24032 13456 24084 13462
rect 24032 13398 24084 13404
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22296 12442 22324 12718
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21100 11150 21128 11290
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21100 10606 21128 11086
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21376 10266 21404 10542
rect 21744 10266 21772 11834
rect 22388 11694 22416 13262
rect 23400 12782 23428 13262
rect 24872 12986 24900 15263
rect 25240 13530 25268 16934
rect 25516 15162 25544 24126
rect 26160 21146 26188 35686
rect 26252 35018 26280 35974
rect 26240 35012 26292 35018
rect 26240 34954 26292 34960
rect 26344 32910 26372 39238
rect 26792 38888 26844 38894
rect 26698 38856 26754 38865
rect 26608 38820 26660 38826
rect 26792 38830 26844 38836
rect 26698 38791 26700 38800
rect 26608 38762 26660 38768
rect 26752 38791 26754 38800
rect 26700 38762 26752 38768
rect 26620 38418 26648 38762
rect 26804 38729 26832 38830
rect 26790 38720 26846 38729
rect 26790 38655 26846 38664
rect 26896 38486 26924 39374
rect 26988 39030 27016 39442
rect 27252 39432 27304 39438
rect 27250 39400 27252 39409
rect 27304 39400 27306 39409
rect 27250 39335 27306 39344
rect 27436 39092 27488 39098
rect 27436 39034 27488 39040
rect 26976 39024 27028 39030
rect 26976 38966 27028 38972
rect 26884 38480 26936 38486
rect 26884 38422 26936 38428
rect 26608 38412 26660 38418
rect 26608 38354 26660 38360
rect 26884 38208 26936 38214
rect 26884 38150 26936 38156
rect 26896 37806 26924 38150
rect 26884 37800 26936 37806
rect 26884 37742 26936 37748
rect 27068 37732 27120 37738
rect 27068 37674 27120 37680
rect 26700 37664 26752 37670
rect 26700 37606 26752 37612
rect 26712 37330 26740 37606
rect 26700 37324 26752 37330
rect 26700 37266 26752 37272
rect 26608 36916 26660 36922
rect 26608 36858 26660 36864
rect 26620 36378 26648 36858
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 27080 36174 27108 37674
rect 27448 37330 27476 39034
rect 27526 38584 27582 38593
rect 27526 38519 27528 38528
rect 27580 38519 27582 38528
rect 27528 38490 27580 38496
rect 28356 38344 28408 38350
rect 28356 38286 28408 38292
rect 28368 37398 28396 38286
rect 29012 37398 29040 40462
rect 29828 39636 29880 39642
rect 29828 39578 29880 39584
rect 29840 39506 29868 39578
rect 29932 39506 29960 41534
rect 30654 41168 30710 41177
rect 30654 41103 30710 41112
rect 30668 41070 30696 41103
rect 30656 41064 30708 41070
rect 30656 41006 30708 41012
rect 30012 40996 30064 41002
rect 30012 40938 30064 40944
rect 30024 40594 30052 40938
rect 30012 40588 30064 40594
rect 30012 40530 30064 40536
rect 30944 39982 30972 41618
rect 31588 41614 31616 42162
rect 32588 42084 32640 42090
rect 32588 42026 32640 42032
rect 31668 41744 31720 41750
rect 31668 41686 31720 41692
rect 31576 41608 31628 41614
rect 31576 41550 31628 41556
rect 31680 41426 31708 41686
rect 31588 41398 31708 41426
rect 31588 41274 31616 41398
rect 31576 41268 31628 41274
rect 31576 41210 31628 41216
rect 31576 40928 31628 40934
rect 31576 40870 31628 40876
rect 31588 40186 31616 40870
rect 31576 40180 31628 40186
rect 31576 40122 31628 40128
rect 30564 39976 30616 39982
rect 30564 39918 30616 39924
rect 30748 39976 30800 39982
rect 30748 39918 30800 39924
rect 30932 39976 30984 39982
rect 30932 39918 30984 39924
rect 31116 39976 31168 39982
rect 31116 39918 31168 39924
rect 30576 39642 30604 39918
rect 30564 39636 30616 39642
rect 30564 39578 30616 39584
rect 29828 39500 29880 39506
rect 29828 39442 29880 39448
rect 29920 39500 29972 39506
rect 29920 39442 29972 39448
rect 29736 39432 29788 39438
rect 29736 39374 29788 39380
rect 29748 39098 29776 39374
rect 29736 39092 29788 39098
rect 29736 39034 29788 39040
rect 29828 39092 29880 39098
rect 29828 39034 29880 39040
rect 29840 38978 29868 39034
rect 29472 38950 29868 38978
rect 29472 38894 29500 38950
rect 29460 38888 29512 38894
rect 29460 38830 29512 38836
rect 29644 38888 29696 38894
rect 29644 38830 29696 38836
rect 29656 38554 29684 38830
rect 29644 38548 29696 38554
rect 29644 38490 29696 38496
rect 30654 38448 30710 38457
rect 30654 38383 30656 38392
rect 30708 38383 30710 38392
rect 30656 38354 30708 38360
rect 29092 38276 29144 38282
rect 29092 38218 29144 38224
rect 29104 37942 29132 38218
rect 30668 37942 30696 38354
rect 30760 38214 30788 39918
rect 31128 39846 31156 39918
rect 31116 39840 31168 39846
rect 31116 39782 31168 39788
rect 31024 39568 31076 39574
rect 31022 39536 31024 39545
rect 31076 39536 31078 39545
rect 31128 39506 31156 39782
rect 31392 39636 31444 39642
rect 31392 39578 31444 39584
rect 31022 39471 31078 39480
rect 31116 39500 31168 39506
rect 31116 39442 31168 39448
rect 30840 39296 30892 39302
rect 30840 39238 30892 39244
rect 30748 38208 30800 38214
rect 30748 38150 30800 38156
rect 29092 37936 29144 37942
rect 29092 37878 29144 37884
rect 30656 37936 30708 37942
rect 30656 37878 30708 37884
rect 30760 37806 30788 38150
rect 29092 37800 29144 37806
rect 29092 37742 29144 37748
rect 29276 37800 29328 37806
rect 29276 37742 29328 37748
rect 30748 37800 30800 37806
rect 30748 37742 30800 37748
rect 29104 37505 29132 37742
rect 29090 37496 29146 37505
rect 29090 37431 29146 37440
rect 28356 37392 28408 37398
rect 28356 37334 28408 37340
rect 29000 37392 29052 37398
rect 29000 37334 29052 37340
rect 27252 37324 27304 37330
rect 27252 37266 27304 37272
rect 27436 37324 27488 37330
rect 27436 37266 27488 37272
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 27172 36038 27200 36722
rect 27160 36032 27212 36038
rect 27160 35974 27212 35980
rect 27264 35630 27292 37266
rect 27448 36786 27476 37266
rect 27436 36780 27488 36786
rect 27436 36722 27488 36728
rect 27436 36168 27488 36174
rect 29288 36122 29316 37742
rect 30380 37732 30432 37738
rect 30380 37674 30432 37680
rect 30288 37664 30340 37670
rect 30288 37606 30340 37612
rect 30300 36174 30328 37606
rect 30392 37398 30420 37674
rect 30380 37392 30432 37398
rect 30380 37334 30432 37340
rect 30852 37330 30880 39238
rect 31404 39098 31432 39578
rect 31392 39092 31444 39098
rect 31392 39034 31444 39040
rect 31484 38412 31536 38418
rect 31484 38354 31536 38360
rect 30840 37324 30892 37330
rect 30840 37266 30892 37272
rect 30564 37188 30616 37194
rect 30564 37130 30616 37136
rect 30472 37120 30524 37126
rect 30472 37062 30524 37068
rect 30484 36922 30512 37062
rect 30472 36916 30524 36922
rect 30472 36858 30524 36864
rect 27436 36110 27488 36116
rect 27448 36038 27476 36110
rect 29196 36106 29316 36122
rect 30288 36168 30340 36174
rect 30288 36110 30340 36116
rect 27528 36100 27580 36106
rect 27528 36042 27580 36048
rect 29184 36100 29316 36106
rect 29236 36094 29316 36100
rect 29184 36042 29236 36048
rect 27436 36032 27488 36038
rect 27436 35974 27488 35980
rect 27540 35766 27568 36042
rect 27528 35760 27580 35766
rect 27528 35702 27580 35708
rect 27252 35624 27304 35630
rect 27252 35566 27304 35572
rect 28632 35624 28684 35630
rect 28632 35566 28684 35572
rect 28644 35494 28672 35566
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 28632 35488 28684 35494
rect 28632 35430 28684 35436
rect 26424 34672 26476 34678
rect 26424 34614 26476 34620
rect 26436 34542 26464 34614
rect 26424 34536 26476 34542
rect 26424 34478 26476 34484
rect 26528 33998 26556 35430
rect 27896 35216 27948 35222
rect 27896 35158 27948 35164
rect 26700 35148 26752 35154
rect 26700 35090 26752 35096
rect 26516 33992 26568 33998
rect 26516 33934 26568 33940
rect 26528 33674 26556 33934
rect 26712 33810 26740 35090
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27816 34785 27844 35022
rect 27802 34776 27858 34785
rect 27802 34711 27858 34720
rect 26976 34672 27028 34678
rect 26976 34614 27028 34620
rect 26792 34400 26844 34406
rect 26792 34342 26844 34348
rect 26804 34066 26832 34342
rect 26792 34060 26844 34066
rect 26792 34002 26844 34008
rect 26712 33782 26832 33810
rect 26528 33658 26740 33674
rect 26528 33652 26752 33658
rect 26528 33646 26700 33652
rect 26700 33594 26752 33600
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26804 31686 26832 33782
rect 26988 32570 27016 34614
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 26976 32564 27028 32570
rect 26976 32506 27028 32512
rect 27068 32564 27120 32570
rect 27068 32506 27120 32512
rect 26976 32360 27028 32366
rect 26976 32302 27028 32308
rect 26792 31680 26844 31686
rect 26792 31622 26844 31628
rect 26804 31278 26832 31622
rect 26792 31272 26844 31278
rect 26792 31214 26844 31220
rect 26792 31136 26844 31142
rect 26792 31078 26844 31084
rect 26804 30802 26832 31078
rect 26792 30796 26844 30802
rect 26792 30738 26844 30744
rect 26988 30682 27016 32302
rect 26896 30654 27016 30682
rect 26700 29300 26752 29306
rect 26700 29242 26752 29248
rect 26712 28626 26740 29242
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26608 27940 26660 27946
rect 26608 27882 26660 27888
rect 26620 27826 26648 27882
rect 26620 27798 26740 27826
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26252 27130 26280 27270
rect 26620 27130 26648 27610
rect 26712 27538 26740 27798
rect 26700 27532 26752 27538
rect 26700 27474 26752 27480
rect 26240 27124 26292 27130
rect 26240 27066 26292 27072
rect 26608 27124 26660 27130
rect 26608 27066 26660 27072
rect 26620 26450 26648 27066
rect 26608 26444 26660 26450
rect 26608 26386 26660 26392
rect 26516 25832 26568 25838
rect 26516 25774 26568 25780
rect 26528 25498 26556 25774
rect 26516 25492 26568 25498
rect 26516 25434 26568 25440
rect 26712 25378 26740 27474
rect 26792 26240 26844 26246
rect 26792 26182 26844 26188
rect 26528 25350 26740 25378
rect 26804 25362 26832 26182
rect 26792 25356 26844 25362
rect 26528 24274 26556 25350
rect 26792 25298 26844 25304
rect 26516 24268 26568 24274
rect 26516 24210 26568 24216
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 26252 23866 26280 24142
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 26528 23798 26556 24210
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 26712 23186 26740 24006
rect 26896 23730 26924 30654
rect 26976 30592 27028 30598
rect 26976 30534 27028 30540
rect 26988 29170 27016 30534
rect 27080 30122 27108 32506
rect 27068 30116 27120 30122
rect 27068 30058 27120 30064
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 26988 28966 27016 29106
rect 26976 28960 27028 28966
rect 26976 28902 27028 28908
rect 26988 28082 27016 28902
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 27172 26586 27200 32914
rect 27264 30598 27292 33594
rect 27356 31822 27384 34546
rect 27804 32768 27856 32774
rect 27804 32710 27856 32716
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 27540 31414 27568 31962
rect 27816 31958 27844 32710
rect 27804 31952 27856 31958
rect 27724 31912 27804 31940
rect 27620 31884 27672 31890
rect 27620 31826 27672 31832
rect 27632 31793 27660 31826
rect 27724 31822 27752 31912
rect 27804 31894 27856 31900
rect 27712 31816 27764 31822
rect 27618 31784 27674 31793
rect 27712 31758 27764 31764
rect 27618 31719 27674 31728
rect 27344 31408 27396 31414
rect 27344 31350 27396 31356
rect 27528 31408 27580 31414
rect 27528 31350 27580 31356
rect 27356 31142 27384 31350
rect 27344 31136 27396 31142
rect 27344 31078 27396 31084
rect 27526 30968 27582 30977
rect 27724 30938 27752 31758
rect 27526 30903 27582 30912
rect 27712 30932 27764 30938
rect 27540 30870 27568 30903
rect 27712 30874 27764 30880
rect 27528 30864 27580 30870
rect 27528 30806 27580 30812
rect 27252 30592 27304 30598
rect 27252 30534 27304 30540
rect 27436 28416 27488 28422
rect 27436 28358 27488 28364
rect 27448 27538 27476 28358
rect 27804 28008 27856 28014
rect 27804 27950 27856 27956
rect 27816 27606 27844 27950
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 27436 27532 27488 27538
rect 27436 27474 27488 27480
rect 27160 26580 27212 26586
rect 27160 26522 27212 26528
rect 27804 26444 27856 26450
rect 27804 26386 27856 26392
rect 27816 26042 27844 26386
rect 27804 26036 27856 26042
rect 27804 25978 27856 25984
rect 26884 23724 26936 23730
rect 26884 23666 26936 23672
rect 27160 23588 27212 23594
rect 27160 23530 27212 23536
rect 26700 23180 26752 23186
rect 26700 23122 26752 23128
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 26804 22642 26832 22918
rect 26792 22636 26844 22642
rect 26792 22578 26844 22584
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26252 20602 26280 20810
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26252 20398 26280 20538
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25792 19310 25820 19926
rect 25688 19304 25740 19310
rect 25688 19246 25740 19252
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25700 19174 25728 19246
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 17678 25728 19110
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25792 18358 25820 18634
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25780 18352 25832 18358
rect 25780 18294 25832 18300
rect 25792 18222 25820 18294
rect 25884 18222 25912 18362
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 26252 17882 26280 20334
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26712 19174 26740 19654
rect 26804 19242 26832 20878
rect 26792 19236 26844 19242
rect 26792 19178 26844 19184
rect 26700 19168 26752 19174
rect 26700 19110 26752 19116
rect 26424 18148 26476 18154
rect 26424 18090 26476 18096
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26252 17678 26280 17818
rect 26436 17746 26464 18090
rect 26332 17740 26384 17746
rect 26332 17682 26384 17688
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 26252 15706 26280 17614
rect 26344 17134 26372 17682
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26792 17060 26844 17066
rect 26792 17002 26844 17008
rect 26240 15700 26292 15706
rect 26240 15642 26292 15648
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25700 14958 25728 15302
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 25700 13394 25728 14894
rect 26252 14618 26280 15642
rect 26804 15570 26832 17002
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26792 14884 26844 14890
rect 26792 14826 26844 14832
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 24872 12442 24900 12922
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 25148 11762 25176 13330
rect 26252 13258 26280 14554
rect 26804 14482 26832 14826
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26252 12986 26280 13194
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26804 12850 26832 13126
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 24400 11688 24452 11694
rect 24400 11630 24452 11636
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22296 10810 22324 11086
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 23584 10674 23612 10950
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 21376 9586 21404 10202
rect 24412 9654 24440 11630
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26252 10674 26280 11494
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26528 10606 26556 12786
rect 26516 10600 26568 10606
rect 26516 10542 26568 10548
rect 26528 10130 26556 10542
rect 26792 10464 26844 10470
rect 26792 10406 26844 10412
rect 26804 10130 26832 10406
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26528 9722 26556 10066
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 7954 16252 8230
rect 16592 8106 16620 8366
rect 16592 8090 16712 8106
rect 16592 8084 16724 8090
rect 16592 8078 16672 8084
rect 16672 8026 16724 8032
rect 16776 7970 16804 8774
rect 17880 8634 17908 8774
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17144 8430 17172 8570
rect 18064 8498 18092 8910
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18708 8430 18736 9046
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22112 8634 22140 8774
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22296 8498 22324 9318
rect 23216 8974 23244 9454
rect 24412 9042 24440 9590
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 16948 8424 17000 8430
rect 17132 8424 17184 8430
rect 17000 8384 17080 8412
rect 16948 8366 17000 8372
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16592 7942 16804 7970
rect 16592 7886 16620 7942
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 6322 13860 7210
rect 15028 7002 15056 7482
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 16592 6866 16620 7822
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16960 6866 16988 7142
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17052 6798 17080 8384
rect 17132 8366 17184 8372
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 20548 8090 20576 8298
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 22296 7954 22324 8434
rect 22756 8362 22784 8774
rect 23124 8634 23152 8910
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 23584 7750 23612 8298
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 22848 7410 22876 7686
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 22848 6866 22876 7346
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 23584 6798 23612 7686
rect 23952 7002 23980 7822
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 23584 5642 23612 6734
rect 23572 5636 23624 5642
rect 23572 5578 23624 5584
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 27172 4146 27200 23530
rect 27712 23180 27764 23186
rect 27712 23122 27764 23128
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27632 22098 27660 22714
rect 27724 22098 27752 23122
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27908 20602 27936 35158
rect 28172 35148 28224 35154
rect 28172 35090 28224 35096
rect 28184 34134 28212 35090
rect 28172 34128 28224 34134
rect 28172 34070 28224 34076
rect 28356 34128 28408 34134
rect 28356 34070 28408 34076
rect 27988 34060 28040 34066
rect 27988 34002 28040 34008
rect 28000 21146 28028 34002
rect 28264 33856 28316 33862
rect 28264 33798 28316 33804
rect 28276 33658 28304 33798
rect 28264 33652 28316 33658
rect 28264 33594 28316 33600
rect 28264 32768 28316 32774
rect 28264 32710 28316 32716
rect 28080 28620 28132 28626
rect 28080 28562 28132 28568
rect 28092 28218 28120 28562
rect 28080 28212 28132 28218
rect 28080 28154 28132 28160
rect 28276 25430 28304 32710
rect 28368 31210 28396 34070
rect 28356 31204 28408 31210
rect 28356 31146 28408 31152
rect 28644 28558 28672 35430
rect 28906 35184 28962 35193
rect 28906 35119 28908 35128
rect 28960 35119 28962 35128
rect 28908 35090 28960 35096
rect 28722 34640 28778 34649
rect 28722 34575 28778 34584
rect 28632 28552 28684 28558
rect 28632 28494 28684 28500
rect 28264 25424 28316 25430
rect 28264 25366 28316 25372
rect 28736 24410 28764 34575
rect 28920 34474 28948 35090
rect 29196 34542 29224 36042
rect 29460 35624 29512 35630
rect 29460 35566 29512 35572
rect 30012 35624 30064 35630
rect 30012 35566 30064 35572
rect 29472 35494 29500 35566
rect 30024 35494 30052 35566
rect 29460 35488 29512 35494
rect 29460 35430 29512 35436
rect 30012 35488 30064 35494
rect 30012 35430 30064 35436
rect 29550 34776 29606 34785
rect 29550 34711 29606 34720
rect 29564 34542 29592 34711
rect 30300 34626 30328 36110
rect 30576 35698 30604 37130
rect 31496 37126 31524 38354
rect 31576 37936 31628 37942
rect 31576 37878 31628 37884
rect 31588 37670 31616 37878
rect 31576 37664 31628 37670
rect 31576 37606 31628 37612
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 31496 36242 31524 37062
rect 31484 36236 31536 36242
rect 31484 36178 31536 36184
rect 30840 35828 30892 35834
rect 30840 35770 30892 35776
rect 30932 35828 30984 35834
rect 30932 35770 30984 35776
rect 30564 35692 30616 35698
rect 30564 35634 30616 35640
rect 30380 35148 30432 35154
rect 30380 35090 30432 35096
rect 30392 34746 30420 35090
rect 30380 34740 30432 34746
rect 30380 34682 30432 34688
rect 30748 34740 30800 34746
rect 30748 34682 30800 34688
rect 30300 34598 30420 34626
rect 30760 34610 30788 34682
rect 30852 34610 30880 35770
rect 30944 35698 30972 35770
rect 31392 35760 31444 35766
rect 31588 35748 31616 37606
rect 31680 37330 31708 41398
rect 32220 40044 32272 40050
rect 32220 39986 32272 39992
rect 32232 39953 32260 39986
rect 32600 39982 32628 42026
rect 32680 40996 32732 41002
rect 32680 40938 32732 40944
rect 32692 40050 32720 40938
rect 32956 40520 33008 40526
rect 32956 40462 33008 40468
rect 32968 40050 32996 40462
rect 32680 40044 32732 40050
rect 32680 39986 32732 39992
rect 32956 40044 33008 40050
rect 32956 39986 33008 39992
rect 34060 40044 34112 40050
rect 34060 39986 34112 39992
rect 32588 39976 32640 39982
rect 32218 39944 32274 39953
rect 32128 39908 32180 39914
rect 32588 39918 32640 39924
rect 33416 39976 33468 39982
rect 33416 39918 33468 39924
rect 32218 39879 32274 39888
rect 32128 39850 32180 39856
rect 31760 39840 31812 39846
rect 31760 39782 31812 39788
rect 31772 39438 31800 39782
rect 31760 39432 31812 39438
rect 31760 39374 31812 39380
rect 32140 37874 32168 39850
rect 32232 39506 32260 39879
rect 32220 39500 32272 39506
rect 32220 39442 32272 39448
rect 32864 38344 32916 38350
rect 32916 38292 33272 38298
rect 32864 38286 33272 38292
rect 32876 38270 33272 38286
rect 33244 38214 33272 38270
rect 33140 38208 33192 38214
rect 33140 38150 33192 38156
rect 33232 38208 33284 38214
rect 33232 38150 33284 38156
rect 33152 38026 33180 38150
rect 33152 37998 33272 38026
rect 33244 37942 33272 37998
rect 32680 37936 32732 37942
rect 32680 37878 32732 37884
rect 33232 37936 33284 37942
rect 33232 37878 33284 37884
rect 32128 37868 32180 37874
rect 32128 37810 32180 37816
rect 31668 37324 31720 37330
rect 31668 37266 31720 37272
rect 32404 36644 32456 36650
rect 32404 36586 32456 36592
rect 32220 36304 32272 36310
rect 32272 36264 32352 36292
rect 32220 36246 32272 36252
rect 32324 35834 32352 36264
rect 32416 36242 32444 36586
rect 32404 36236 32456 36242
rect 32404 36178 32456 36184
rect 31668 35828 31720 35834
rect 31668 35770 31720 35776
rect 32220 35828 32272 35834
rect 32220 35770 32272 35776
rect 32312 35828 32364 35834
rect 32312 35770 32364 35776
rect 31392 35702 31444 35708
rect 31496 35720 31616 35748
rect 30932 35692 30984 35698
rect 30932 35634 30984 35640
rect 31024 35624 31076 35630
rect 31024 35566 31076 35572
rect 31036 35494 31064 35566
rect 31404 35494 31432 35702
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 31392 35488 31444 35494
rect 31392 35430 31444 35436
rect 29184 34536 29236 34542
rect 29184 34478 29236 34484
rect 29552 34536 29604 34542
rect 29552 34478 29604 34484
rect 28908 34468 28960 34474
rect 28908 34410 28960 34416
rect 29196 33862 29224 34478
rect 30288 34468 30340 34474
rect 30288 34410 30340 34416
rect 30300 34202 30328 34410
rect 30392 34406 30420 34598
rect 30748 34604 30800 34610
rect 30748 34546 30800 34552
rect 30840 34604 30892 34610
rect 30840 34546 30892 34552
rect 30380 34400 30432 34406
rect 30380 34342 30432 34348
rect 30288 34196 30340 34202
rect 30288 34138 30340 34144
rect 29184 33856 29236 33862
rect 29184 33798 29236 33804
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 28828 30326 28856 32846
rect 29642 30832 29698 30841
rect 29642 30767 29698 30776
rect 28816 30320 28868 30326
rect 28816 30262 28868 30268
rect 28998 30152 29054 30161
rect 28998 30087 29054 30096
rect 28906 29472 28962 29481
rect 28906 29407 28962 29416
rect 28920 28218 28948 29407
rect 29012 29306 29040 30087
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 28908 28212 28960 28218
rect 28908 28154 28960 28160
rect 28998 28112 29054 28121
rect 28998 28047 29054 28056
rect 29012 27674 29040 28047
rect 29000 27668 29052 27674
rect 29000 27610 29052 27616
rect 28906 26752 28962 26761
rect 28906 26687 28962 26696
rect 28920 26042 28948 26687
rect 28908 26036 28960 26042
rect 28908 25978 28960 25984
rect 28998 25528 29054 25537
rect 28998 25463 29054 25472
rect 29012 24886 29040 25463
rect 29000 24880 29052 24886
rect 29000 24822 29052 24828
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28736 23866 28764 24346
rect 29000 24200 29052 24206
rect 28998 24168 29000 24177
rect 29052 24168 29054 24177
rect 28998 24103 29054 24112
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 29090 22808 29146 22817
rect 29090 22743 29092 22752
rect 29144 22743 29146 22752
rect 29092 22714 29144 22720
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27896 20596 27948 20602
rect 27896 20538 27948 20544
rect 27540 20058 27568 20538
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 28000 19854 28028 21082
rect 29090 20088 29146 20097
rect 29090 20023 29146 20032
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 27710 18728 27766 18737
rect 27710 18663 27766 18672
rect 27724 18426 27752 18663
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27724 18222 27752 18362
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27724 17882 27752 18158
rect 27712 17876 27764 17882
rect 27712 17818 27764 17824
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27264 16250 27292 17070
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27540 15638 27568 15846
rect 27528 15632 27580 15638
rect 27528 15574 27580 15580
rect 29104 14958 29132 20023
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 28998 14784 29054 14793
rect 28998 14719 29054 14728
rect 29012 13870 29040 14719
rect 29104 14550 29132 14894
rect 29092 14544 29144 14550
rect 29092 14486 29144 14492
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27724 13394 27752 13670
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 28092 12986 28120 13806
rect 28080 12980 28132 12986
rect 28080 12922 28132 12928
rect 29656 11898 29684 30767
rect 31036 26994 31064 35430
rect 31496 29238 31524 35720
rect 31576 35624 31628 35630
rect 31680 35612 31708 35770
rect 32232 35630 32260 35770
rect 32692 35766 32720 37878
rect 33140 36848 33192 36854
rect 33140 36790 33192 36796
rect 32680 35760 32732 35766
rect 32680 35702 32732 35708
rect 31628 35584 31708 35612
rect 32220 35624 32272 35630
rect 31576 35566 31628 35572
rect 32220 35566 32272 35572
rect 33152 35306 33180 36790
rect 32784 35290 33180 35306
rect 32772 35284 33180 35290
rect 32824 35278 33180 35284
rect 32772 35226 32824 35232
rect 33244 35154 33272 37878
rect 33428 37738 33456 39918
rect 34072 38758 34100 39986
rect 34152 39432 34204 39438
rect 34152 39374 34204 39380
rect 34164 38758 34192 39374
rect 34060 38752 34112 38758
rect 34060 38694 34112 38700
rect 34152 38752 34204 38758
rect 34152 38694 34204 38700
rect 34440 37942 34468 42638
rect 34808 42158 34836 43114
rect 35440 42764 35492 42770
rect 35440 42706 35492 42712
rect 35348 42560 35400 42566
rect 35348 42502 35400 42508
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 34796 42152 34848 42158
rect 34796 42094 34848 42100
rect 34808 41138 34836 42094
rect 35360 41750 35388 42502
rect 35348 41744 35400 41750
rect 35348 41686 35400 41692
rect 35452 41682 35480 42706
rect 35532 42628 35584 42634
rect 35532 42570 35584 42576
rect 35440 41676 35492 41682
rect 35440 41618 35492 41624
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 34796 41132 34848 41138
rect 34796 41074 34848 41080
rect 34610 40760 34666 40769
rect 34610 40695 34666 40704
rect 34624 40662 34652 40695
rect 34612 40656 34664 40662
rect 34612 40598 34664 40604
rect 35348 40588 35400 40594
rect 35348 40530 35400 40536
rect 34796 40384 34848 40390
rect 34796 40326 34848 40332
rect 34808 40118 34836 40326
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34796 40112 34848 40118
rect 34796 40054 34848 40060
rect 34612 39364 34664 39370
rect 34612 39306 34664 39312
rect 34624 39098 34652 39306
rect 34704 39296 34756 39302
rect 34704 39238 34756 39244
rect 34612 39092 34664 39098
rect 34612 39034 34664 39040
rect 34716 39030 34744 39238
rect 34704 39024 34756 39030
rect 34704 38966 34756 38972
rect 34808 38962 34836 40054
rect 35360 40050 35388 40530
rect 35348 40044 35400 40050
rect 35348 39986 35400 39992
rect 35070 39536 35126 39545
rect 35360 39506 35388 39986
rect 35544 39930 35572 42570
rect 36728 42152 36780 42158
rect 37280 42152 37332 42158
rect 36780 42100 36952 42106
rect 36728 42094 36952 42100
rect 37280 42094 37332 42100
rect 35900 42084 35952 42090
rect 36740 42078 36952 42094
rect 35900 42026 35952 42032
rect 35624 40588 35676 40594
rect 35624 40530 35676 40536
rect 35716 40588 35768 40594
rect 35716 40530 35768 40536
rect 35636 40118 35664 40530
rect 35728 40390 35756 40530
rect 35716 40384 35768 40390
rect 35716 40326 35768 40332
rect 35624 40112 35676 40118
rect 35624 40054 35676 40060
rect 35728 39982 35756 40326
rect 35912 40186 35940 42026
rect 36924 42022 36952 42078
rect 36912 42016 36964 42022
rect 36912 41958 36964 41964
rect 35992 41676 36044 41682
rect 35992 41618 36044 41624
rect 36268 41676 36320 41682
rect 36268 41618 36320 41624
rect 36004 41138 36032 41618
rect 36280 41290 36308 41618
rect 36096 41262 36308 41290
rect 35992 41132 36044 41138
rect 35992 41074 36044 41080
rect 35900 40180 35952 40186
rect 35900 40122 35952 40128
rect 35716 39976 35768 39982
rect 35544 39902 35664 39930
rect 35716 39918 35768 39924
rect 35532 39840 35584 39846
rect 35532 39782 35584 39788
rect 35544 39574 35572 39782
rect 35532 39568 35584 39574
rect 35532 39510 35584 39516
rect 35070 39471 35126 39480
rect 35348 39500 35400 39506
rect 35084 39370 35112 39471
rect 35348 39442 35400 39448
rect 35072 39364 35124 39370
rect 35072 39306 35124 39312
rect 35360 39302 35388 39442
rect 35348 39296 35400 39302
rect 35348 39238 35400 39244
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34796 38956 34848 38962
rect 34796 38898 34848 38904
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34428 37936 34480 37942
rect 34428 37878 34480 37884
rect 33416 37732 33468 37738
rect 33416 37674 33468 37680
rect 34440 37330 34468 37878
rect 35636 37777 35664 39902
rect 35808 39840 35860 39846
rect 35808 39782 35860 39788
rect 35820 39506 35848 39782
rect 36096 39658 36124 41262
rect 36176 41200 36228 41206
rect 36176 41142 36228 41148
rect 36188 40730 36216 41142
rect 36268 41064 36320 41070
rect 36268 41006 36320 41012
rect 36452 41064 36504 41070
rect 36452 41006 36504 41012
rect 36636 41064 36688 41070
rect 36636 41006 36688 41012
rect 36280 40730 36308 41006
rect 36176 40724 36228 40730
rect 36176 40666 36228 40672
rect 36268 40724 36320 40730
rect 36268 40666 36320 40672
rect 35912 39630 36124 39658
rect 36176 39636 36228 39642
rect 35808 39500 35860 39506
rect 35808 39442 35860 39448
rect 35912 38026 35940 39630
rect 36176 39578 36228 39584
rect 36084 39500 36136 39506
rect 36188 39488 36216 39578
rect 36136 39460 36216 39488
rect 36084 39442 36136 39448
rect 36464 38350 36492 41006
rect 36648 40934 36676 41006
rect 36544 40928 36596 40934
rect 36544 40870 36596 40876
rect 36636 40928 36688 40934
rect 36636 40870 36688 40876
rect 36556 40662 36584 40870
rect 36544 40656 36596 40662
rect 36544 40598 36596 40604
rect 36636 40588 36688 40594
rect 36636 40530 36688 40536
rect 36648 39438 36676 40530
rect 36820 40384 36872 40390
rect 36820 40326 36872 40332
rect 36832 40118 36860 40326
rect 36820 40112 36872 40118
rect 36820 40054 36872 40060
rect 36832 39642 36860 40054
rect 36924 39982 36952 41958
rect 37292 41818 37320 42094
rect 37280 41812 37332 41818
rect 37280 41754 37332 41760
rect 37660 41750 37688 43590
rect 39040 43246 39068 43794
rect 39396 43716 39448 43722
rect 39396 43658 39448 43664
rect 39028 43240 39080 43246
rect 39028 43182 39080 43188
rect 38476 43172 38528 43178
rect 38476 43114 38528 43120
rect 38568 43172 38620 43178
rect 38568 43114 38620 43120
rect 37832 42560 37884 42566
rect 37832 42502 37884 42508
rect 37844 42090 37872 42502
rect 37740 42084 37792 42090
rect 37740 42026 37792 42032
rect 37832 42084 37884 42090
rect 37832 42026 37884 42032
rect 37096 41744 37148 41750
rect 37648 41744 37700 41750
rect 37096 41686 37148 41692
rect 37278 41712 37334 41721
rect 37108 40934 37136 41686
rect 37648 41686 37700 41692
rect 37278 41647 37334 41656
rect 37292 41614 37320 41647
rect 37280 41608 37332 41614
rect 37280 41550 37332 41556
rect 37648 41540 37700 41546
rect 37648 41482 37700 41488
rect 37464 41472 37516 41478
rect 37464 41414 37516 41420
rect 37096 40928 37148 40934
rect 37096 40870 37148 40876
rect 37476 40662 37504 41414
rect 37464 40656 37516 40662
rect 37464 40598 37516 40604
rect 37660 40390 37688 41482
rect 37752 41070 37780 42026
rect 38108 41744 38160 41750
rect 38108 41686 38160 41692
rect 38120 41478 38148 41686
rect 38292 41540 38344 41546
rect 38292 41482 38344 41488
rect 38108 41472 38160 41478
rect 38108 41414 38160 41420
rect 37740 41064 37792 41070
rect 37740 41006 37792 41012
rect 38304 40662 38332 41482
rect 38488 41138 38516 43114
rect 38580 42906 38608 43114
rect 39040 43110 39068 43182
rect 39028 43104 39080 43110
rect 39028 43046 39080 43052
rect 38568 42900 38620 42906
rect 38568 42842 38620 42848
rect 38936 42016 38988 42022
rect 38936 41958 38988 41964
rect 38660 41744 38712 41750
rect 38658 41712 38660 41721
rect 38712 41712 38714 41721
rect 38658 41647 38714 41656
rect 38568 41200 38620 41206
rect 38568 41142 38620 41148
rect 38476 41132 38528 41138
rect 38476 41074 38528 41080
rect 37924 40656 37976 40662
rect 37924 40598 37976 40604
rect 38292 40656 38344 40662
rect 38580 40610 38608 41142
rect 38660 41132 38712 41138
rect 38660 41074 38712 41080
rect 38672 41041 38700 41074
rect 38658 41032 38714 41041
rect 38658 40967 38714 40976
rect 38292 40598 38344 40604
rect 37648 40384 37700 40390
rect 37648 40326 37700 40332
rect 37936 40118 37964 40598
rect 38488 40582 38608 40610
rect 38488 40526 38516 40582
rect 38476 40520 38528 40526
rect 38476 40462 38528 40468
rect 38568 40384 38620 40390
rect 38568 40326 38620 40332
rect 38660 40384 38712 40390
rect 38660 40326 38712 40332
rect 37924 40112 37976 40118
rect 37924 40054 37976 40060
rect 36912 39976 36964 39982
rect 36912 39918 36964 39924
rect 38200 39976 38252 39982
rect 38200 39918 38252 39924
rect 38384 39976 38436 39982
rect 38384 39918 38436 39924
rect 38108 39908 38160 39914
rect 38108 39850 38160 39856
rect 38120 39681 38148 39850
rect 38212 39846 38240 39918
rect 38396 39846 38424 39918
rect 38200 39840 38252 39846
rect 38200 39782 38252 39788
rect 38384 39840 38436 39846
rect 38384 39782 38436 39788
rect 38106 39672 38162 39681
rect 36820 39636 36872 39642
rect 38106 39607 38162 39616
rect 38476 39636 38528 39642
rect 36820 39578 36872 39584
rect 38476 39578 38528 39584
rect 36636 39432 36688 39438
rect 36636 39374 36688 39380
rect 37740 39432 37792 39438
rect 37740 39374 37792 39380
rect 36648 39302 36676 39374
rect 36636 39296 36688 39302
rect 36636 39238 36688 39244
rect 36912 39296 36964 39302
rect 36912 39238 36964 39244
rect 36924 38758 36952 39238
rect 37648 39024 37700 39030
rect 37648 38966 37700 38972
rect 37096 38888 37148 38894
rect 37096 38830 37148 38836
rect 37660 38842 37688 38966
rect 37752 38962 37780 39374
rect 37924 39092 37976 39098
rect 37924 39034 37976 39040
rect 37740 38956 37792 38962
rect 37740 38898 37792 38904
rect 37936 38842 37964 39034
rect 38488 38894 38516 39578
rect 38580 39574 38608 40326
rect 38672 40186 38700 40326
rect 38660 40180 38712 40186
rect 38660 40122 38712 40128
rect 38948 39982 38976 41958
rect 39028 41132 39080 41138
rect 39028 41074 39080 41080
rect 39040 41041 39068 41074
rect 39026 41032 39082 41041
rect 39026 40967 39082 40976
rect 39028 40928 39080 40934
rect 39026 40896 39028 40905
rect 39120 40928 39172 40934
rect 39080 40896 39082 40905
rect 39120 40870 39172 40876
rect 39026 40831 39082 40840
rect 39132 40730 39160 40870
rect 39120 40724 39172 40730
rect 39120 40666 39172 40672
rect 39408 40526 39436 43658
rect 40512 43246 40540 43862
rect 48044 43852 48096 43858
rect 48044 43794 48096 43800
rect 49792 43852 49844 43858
rect 49792 43794 49844 43800
rect 47676 43784 47728 43790
rect 47676 43726 47728 43732
rect 46756 43648 46808 43654
rect 46756 43590 46808 43596
rect 45468 43444 45520 43450
rect 45468 43386 45520 43392
rect 40500 43240 40552 43246
rect 40500 43182 40552 43188
rect 43444 43240 43496 43246
rect 43444 43182 43496 43188
rect 40512 42906 40540 43182
rect 40500 42900 40552 42906
rect 40500 42842 40552 42848
rect 43456 42702 43484 43182
rect 43720 43104 43772 43110
rect 43720 43046 43772 43052
rect 43444 42696 43496 42702
rect 43444 42638 43496 42644
rect 39764 42152 39816 42158
rect 39764 42094 39816 42100
rect 39396 40520 39448 40526
rect 39396 40462 39448 40468
rect 38936 39976 38988 39982
rect 38936 39918 38988 39924
rect 38568 39568 38620 39574
rect 38568 39510 38620 39516
rect 39488 39092 39540 39098
rect 39488 39034 39540 39040
rect 36912 38752 36964 38758
rect 36912 38694 36964 38700
rect 37108 38593 37136 38830
rect 37660 38814 37964 38842
rect 38476 38888 38528 38894
rect 38476 38830 38528 38836
rect 36542 38584 36598 38593
rect 36542 38519 36598 38528
rect 37094 38584 37150 38593
rect 37094 38519 37150 38528
rect 36556 38418 36584 38519
rect 36544 38412 36596 38418
rect 36544 38354 36596 38360
rect 36452 38344 36504 38350
rect 36452 38286 36504 38292
rect 35912 37998 36216 38026
rect 35912 37856 35940 37998
rect 36188 37874 36216 37998
rect 35820 37828 35940 37856
rect 35992 37868 36044 37874
rect 35622 37768 35678 37777
rect 35622 37703 35678 37712
rect 34428 37324 34480 37330
rect 34428 37266 34480 37272
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 34612 37120 34664 37126
rect 34612 37062 34664 37068
rect 34624 36786 34652 37062
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34612 36780 34664 36786
rect 34612 36722 34664 36728
rect 33690 36408 33746 36417
rect 33690 36343 33692 36352
rect 33744 36343 33746 36352
rect 33692 36314 33744 36320
rect 34152 36236 34204 36242
rect 34152 36178 34204 36184
rect 33416 35556 33468 35562
rect 33416 35498 33468 35504
rect 33508 35556 33560 35562
rect 33508 35498 33560 35504
rect 33428 35154 33456 35498
rect 33232 35148 33284 35154
rect 33232 35090 33284 35096
rect 33416 35148 33468 35154
rect 33416 35090 33468 35096
rect 32772 32632 32824 32638
rect 32772 32574 32824 32580
rect 32036 31408 32088 31414
rect 32036 31350 32088 31356
rect 31484 29232 31536 29238
rect 31484 29174 31536 29180
rect 31024 26988 31076 26994
rect 31024 26930 31076 26936
rect 32048 23322 32076 31350
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32036 23316 32088 23322
rect 32036 23258 32088 23264
rect 32416 15638 32444 31282
rect 32680 31204 32732 31210
rect 32680 31146 32732 31152
rect 32496 31068 32548 31074
rect 32496 31010 32548 31016
rect 32508 16522 32536 31010
rect 32588 31000 32640 31006
rect 32588 30942 32640 30948
rect 32496 16516 32548 16522
rect 32496 16458 32548 16464
rect 32600 16182 32628 30942
rect 32692 16590 32720 31146
rect 32784 18290 32812 32574
rect 33520 31482 33548 35498
rect 34164 34542 34192 36178
rect 34624 36038 34652 36722
rect 35452 36378 35480 37198
rect 35820 36718 35848 37828
rect 35992 37810 36044 37816
rect 36176 37868 36228 37874
rect 36176 37810 36228 37816
rect 36004 36854 36032 37810
rect 35992 36848 36044 36854
rect 35992 36790 36044 36796
rect 35624 36712 35676 36718
rect 35624 36654 35676 36660
rect 35808 36712 35860 36718
rect 35808 36654 35860 36660
rect 35992 36712 36044 36718
rect 35992 36654 36044 36660
rect 35440 36372 35492 36378
rect 35440 36314 35492 36320
rect 35348 36236 35400 36242
rect 35348 36178 35400 36184
rect 35256 36100 35308 36106
rect 35256 36042 35308 36048
rect 34612 36032 34664 36038
rect 34612 35974 34664 35980
rect 34152 34536 34204 34542
rect 34152 34478 34204 34484
rect 34624 33114 34652 35974
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35268 35834 35296 36042
rect 35360 35834 35388 36178
rect 35256 35828 35308 35834
rect 35256 35770 35308 35776
rect 35348 35828 35400 35834
rect 35348 35770 35400 35776
rect 35268 35562 35296 35770
rect 35256 35556 35308 35562
rect 35256 35498 35308 35504
rect 35636 35018 35664 36654
rect 35716 35692 35768 35698
rect 35820 35680 35848 36654
rect 36004 36417 36032 36654
rect 35990 36408 36046 36417
rect 35990 36343 36046 36352
rect 35898 36272 35954 36281
rect 36464 36242 36492 38286
rect 36636 38004 36688 38010
rect 36636 37946 36688 37952
rect 36648 37806 36676 37946
rect 36636 37800 36688 37806
rect 36542 37768 36598 37777
rect 36636 37742 36688 37748
rect 36542 37703 36544 37712
rect 36596 37703 36598 37712
rect 36544 37674 36596 37680
rect 37108 37398 37136 38519
rect 37738 38448 37794 38457
rect 37936 38418 37964 38814
rect 38488 38758 38516 38830
rect 38476 38752 38528 38758
rect 38476 38694 38528 38700
rect 38488 38418 38516 38694
rect 37738 38383 37740 38392
rect 37792 38383 37794 38392
rect 37924 38412 37976 38418
rect 37740 38354 37792 38360
rect 37924 38354 37976 38360
rect 38016 38412 38068 38418
rect 38016 38354 38068 38360
rect 38476 38412 38528 38418
rect 38660 38412 38712 38418
rect 38528 38372 38608 38400
rect 38476 38354 38528 38360
rect 38028 37806 38056 38354
rect 38580 38196 38608 38372
rect 38660 38354 38712 38360
rect 38672 38196 38700 38354
rect 38842 38312 38898 38321
rect 38842 38247 38844 38256
rect 38896 38247 38898 38256
rect 38844 38218 38896 38224
rect 39500 38214 39528 39034
rect 39580 38752 39632 38758
rect 39580 38694 39632 38700
rect 38580 38168 38700 38196
rect 39488 38208 39540 38214
rect 39488 38150 39540 38156
rect 38016 37800 38068 37806
rect 38016 37742 38068 37748
rect 38200 37664 38252 37670
rect 38200 37606 38252 37612
rect 37096 37392 37148 37398
rect 37096 37334 37148 37340
rect 38212 37330 38240 37606
rect 38290 37496 38346 37505
rect 38290 37431 38346 37440
rect 38304 37330 38332 37431
rect 38200 37324 38252 37330
rect 38200 37266 38252 37272
rect 38292 37324 38344 37330
rect 38292 37266 38344 37272
rect 39488 36780 39540 36786
rect 39488 36722 39540 36728
rect 36544 36576 36596 36582
rect 36544 36518 36596 36524
rect 36636 36576 36688 36582
rect 36636 36518 36688 36524
rect 36556 36378 36584 36518
rect 36544 36372 36596 36378
rect 36544 36314 36596 36320
rect 36648 36310 36676 36518
rect 36636 36304 36688 36310
rect 36636 36246 36688 36252
rect 37554 36272 37610 36281
rect 35898 36207 35954 36216
rect 35992 36236 36044 36242
rect 35912 36174 35940 36207
rect 35992 36178 36044 36184
rect 36452 36236 36504 36242
rect 37554 36207 37610 36216
rect 39120 36236 39172 36242
rect 36452 36178 36504 36184
rect 35900 36168 35952 36174
rect 35900 36110 35952 36116
rect 36004 35698 36032 36178
rect 37568 36174 37596 36207
rect 39120 36178 39172 36184
rect 37556 36168 37608 36174
rect 37556 36110 37608 36116
rect 38752 36032 38804 36038
rect 38658 36000 38714 36009
rect 38752 35974 38804 35980
rect 38658 35935 38714 35944
rect 38384 35828 38436 35834
rect 38384 35770 38436 35776
rect 38476 35828 38528 35834
rect 38476 35770 38528 35776
rect 38396 35737 38424 35770
rect 38382 35728 38438 35737
rect 35768 35652 35848 35680
rect 35992 35692 36044 35698
rect 35716 35634 35768 35640
rect 38382 35663 38438 35672
rect 35992 35634 36044 35640
rect 38488 35630 38516 35770
rect 38568 35692 38620 35698
rect 38672 35680 38700 35935
rect 38620 35652 38700 35680
rect 38568 35634 38620 35640
rect 38476 35624 38528 35630
rect 38396 35572 38476 35578
rect 38396 35566 38528 35572
rect 38396 35550 38516 35566
rect 38396 35494 38424 35550
rect 37832 35488 37884 35494
rect 37832 35430 37884 35436
rect 38016 35488 38068 35494
rect 38016 35430 38068 35436
rect 38384 35488 38436 35494
rect 38384 35430 38436 35436
rect 38476 35488 38528 35494
rect 38476 35430 38528 35436
rect 35624 35012 35676 35018
rect 35624 34954 35676 34960
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 37844 34746 37872 35430
rect 37832 34740 37884 34746
rect 37832 34682 37884 34688
rect 37844 34406 37872 34682
rect 37832 34400 37884 34406
rect 37832 34342 37884 34348
rect 34612 33108 34664 33114
rect 34612 33050 34664 33056
rect 38028 32366 38056 35430
rect 38488 35086 38516 35430
rect 38108 35080 38160 35086
rect 38108 35022 38160 35028
rect 38476 35080 38528 35086
rect 38476 35022 38528 35028
rect 38120 34950 38148 35022
rect 38568 35012 38620 35018
rect 38568 34954 38620 34960
rect 38108 34944 38160 34950
rect 38108 34886 38160 34892
rect 38292 34944 38344 34950
rect 38292 34886 38344 34892
rect 38304 32978 38332 34886
rect 38580 34746 38608 34954
rect 38568 34740 38620 34746
rect 38568 34682 38620 34688
rect 38384 34672 38436 34678
rect 38764 34626 38792 35974
rect 39132 35222 39160 36178
rect 39500 35698 39528 36722
rect 39592 36038 39620 38694
rect 39776 37398 39804 42094
rect 43732 41818 43760 43046
rect 44916 42900 44968 42906
rect 44916 42842 44968 42848
rect 44088 42764 44140 42770
rect 44088 42706 44140 42712
rect 44364 42764 44416 42770
rect 44364 42706 44416 42712
rect 43904 42696 43956 42702
rect 43904 42638 43956 42644
rect 43812 42016 43864 42022
rect 43812 41958 43864 41964
rect 43720 41812 43772 41818
rect 43720 41754 43772 41760
rect 43536 41676 43588 41682
rect 43536 41618 43588 41624
rect 39948 40996 40000 41002
rect 39948 40938 40000 40944
rect 40040 40996 40092 41002
rect 40040 40938 40092 40944
rect 42892 40996 42944 41002
rect 42892 40938 42944 40944
rect 39960 38214 39988 40938
rect 40052 40662 40080 40938
rect 42800 40928 42852 40934
rect 42800 40870 42852 40876
rect 40040 40656 40092 40662
rect 40040 40598 40092 40604
rect 42616 40656 42668 40662
rect 42616 40598 42668 40604
rect 41236 40588 41288 40594
rect 41236 40530 41288 40536
rect 40960 40520 41012 40526
rect 40960 40462 41012 40468
rect 40040 39976 40092 39982
rect 40040 39918 40092 39924
rect 39948 38208 40000 38214
rect 39948 38150 40000 38156
rect 39764 37392 39816 37398
rect 39764 37334 39816 37340
rect 39764 36848 39816 36854
rect 39764 36790 39816 36796
rect 39580 36032 39632 36038
rect 39580 35974 39632 35980
rect 39488 35692 39540 35698
rect 39488 35634 39540 35640
rect 39120 35216 39172 35222
rect 39120 35158 39172 35164
rect 39396 35148 39448 35154
rect 39396 35090 39448 35096
rect 39408 34950 39436 35090
rect 39776 35086 39804 36790
rect 39948 36032 40000 36038
rect 39948 35974 40000 35980
rect 39960 35873 39988 35974
rect 39946 35864 40002 35873
rect 39946 35799 40002 35808
rect 39960 35562 39988 35799
rect 39948 35556 40000 35562
rect 39948 35498 40000 35504
rect 39764 35080 39816 35086
rect 39764 35022 39816 35028
rect 39396 34944 39448 34950
rect 39396 34886 39448 34892
rect 39304 34740 39356 34746
rect 39356 34700 39436 34728
rect 39304 34682 39356 34688
rect 38436 34620 38792 34626
rect 38384 34614 38792 34620
rect 38396 34598 38792 34614
rect 39408 34610 39436 34700
rect 39396 34604 39448 34610
rect 39396 34546 39448 34552
rect 39960 34542 39988 35498
rect 38568 34536 38620 34542
rect 38568 34478 38620 34484
rect 39948 34536 40000 34542
rect 39948 34478 40000 34484
rect 38580 34406 38608 34478
rect 38568 34400 38620 34406
rect 38568 34342 38620 34348
rect 38292 32972 38344 32978
rect 38292 32914 38344 32920
rect 38016 32360 38068 32366
rect 38016 32302 38068 32308
rect 40052 32298 40080 39918
rect 40868 39500 40920 39506
rect 40868 39442 40920 39448
rect 40880 39137 40908 39442
rect 40972 39438 41000 40462
rect 41052 39840 41104 39846
rect 41052 39782 41104 39788
rect 40960 39432 41012 39438
rect 40960 39374 41012 39380
rect 40960 39296 41012 39302
rect 41064 39273 41092 39782
rect 41142 39536 41198 39545
rect 41142 39471 41198 39480
rect 40960 39238 41012 39244
rect 41050 39264 41106 39273
rect 40866 39128 40922 39137
rect 40866 39063 40922 39072
rect 40972 39001 41000 39238
rect 41050 39199 41106 39208
rect 40958 38992 41014 39001
rect 41156 38962 41184 39471
rect 40958 38927 41014 38936
rect 41144 38956 41196 38962
rect 41144 38898 41196 38904
rect 40868 38412 40920 38418
rect 40868 38354 40920 38360
rect 40880 38282 40908 38354
rect 41248 38350 41276 40530
rect 42248 40112 42300 40118
rect 42248 40054 42300 40060
rect 42260 39982 42288 40054
rect 41512 39976 41564 39982
rect 41512 39918 41564 39924
rect 42248 39976 42300 39982
rect 42248 39918 42300 39924
rect 41524 39846 41552 39918
rect 41512 39840 41564 39846
rect 41512 39782 41564 39788
rect 42248 39840 42300 39846
rect 42248 39782 42300 39788
rect 42260 39545 42288 39782
rect 42246 39536 42302 39545
rect 41696 39500 41748 39506
rect 42246 39471 42302 39480
rect 42432 39500 42484 39506
rect 41696 39442 41748 39448
rect 42432 39442 42484 39448
rect 41604 39364 41656 39370
rect 41604 39306 41656 39312
rect 41616 38894 41644 39306
rect 41604 38888 41656 38894
rect 41604 38830 41656 38836
rect 41708 38758 41736 39442
rect 42248 39432 42300 39438
rect 42444 39386 42472 39442
rect 42248 39374 42300 39380
rect 41880 39296 41932 39302
rect 41880 39238 41932 39244
rect 41892 39030 41920 39238
rect 41880 39024 41932 39030
rect 41880 38966 41932 38972
rect 42260 38894 42288 39374
rect 42352 39358 42472 39386
rect 42352 39273 42380 39358
rect 42524 39296 42576 39302
rect 42338 39264 42394 39273
rect 42524 39238 42576 39244
rect 42338 39199 42394 39208
rect 42248 38888 42300 38894
rect 42248 38830 42300 38836
rect 42536 38758 42564 39238
rect 42628 38944 42656 40598
rect 42812 40390 42840 40870
rect 42904 40662 42932 40938
rect 42984 40928 43036 40934
rect 42984 40870 43036 40876
rect 42892 40656 42944 40662
rect 42892 40598 42944 40604
rect 42708 40384 42760 40390
rect 42708 40326 42760 40332
rect 42800 40384 42852 40390
rect 42800 40326 42852 40332
rect 42720 40050 42748 40326
rect 42708 40044 42760 40050
rect 42708 39986 42760 39992
rect 42892 39296 42944 39302
rect 42892 39238 42944 39244
rect 42708 38956 42760 38962
rect 42628 38916 42708 38944
rect 42708 38898 42760 38904
rect 42904 38758 42932 39238
rect 42996 39001 43024 40870
rect 43548 40662 43576 41618
rect 43732 41070 43760 41754
rect 43824 41070 43852 41958
rect 43916 41682 43944 42638
rect 44100 42294 44128 42706
rect 44088 42288 44140 42294
rect 44088 42230 44140 42236
rect 44376 42158 44404 42706
rect 44548 42560 44600 42566
rect 44548 42502 44600 42508
rect 44364 42152 44416 42158
rect 44364 42094 44416 42100
rect 44456 42152 44508 42158
rect 44456 42094 44508 42100
rect 43904 41676 43956 41682
rect 43904 41618 43956 41624
rect 43720 41064 43772 41070
rect 43720 41006 43772 41012
rect 43812 41064 43864 41070
rect 43812 41006 43864 41012
rect 43824 40934 43852 41006
rect 43812 40928 43864 40934
rect 43812 40870 43864 40876
rect 44468 40662 44496 42094
rect 44560 41818 44588 42502
rect 44824 42152 44876 42158
rect 44824 42094 44876 42100
rect 44548 41812 44600 41818
rect 44548 41754 44600 41760
rect 44560 41546 44588 41754
rect 44732 41744 44784 41750
rect 44732 41686 44784 41692
rect 44638 41576 44694 41585
rect 44548 41540 44600 41546
rect 44638 41511 44694 41520
rect 44548 41482 44600 41488
rect 44652 41274 44680 41511
rect 44744 41274 44772 41686
rect 44640 41268 44692 41274
rect 44640 41210 44692 41216
rect 44732 41268 44784 41274
rect 44732 41210 44784 41216
rect 44836 41070 44864 42094
rect 44928 42090 44956 42842
rect 45284 42764 45336 42770
rect 45284 42706 45336 42712
rect 45100 42288 45152 42294
rect 45100 42230 45152 42236
rect 44916 42084 44968 42090
rect 44916 42026 44968 42032
rect 44928 41698 44956 42026
rect 45112 41818 45140 42230
rect 45296 42106 45324 42706
rect 45480 42634 45508 43386
rect 46768 43314 46796 43590
rect 46756 43308 46808 43314
rect 46756 43250 46808 43256
rect 47688 43110 47716 43726
rect 47676 43104 47728 43110
rect 47676 43046 47728 43052
rect 47860 43104 47912 43110
rect 47860 43046 47912 43052
rect 47688 42770 47716 43046
rect 46756 42764 46808 42770
rect 46756 42706 46808 42712
rect 47676 42764 47728 42770
rect 47676 42706 47728 42712
rect 45836 42696 45888 42702
rect 45836 42638 45888 42644
rect 45468 42628 45520 42634
rect 45468 42570 45520 42576
rect 45468 42152 45520 42158
rect 45192 42084 45244 42090
rect 45296 42078 45416 42106
rect 45468 42094 45520 42100
rect 45192 42026 45244 42032
rect 45100 41812 45152 41818
rect 45100 41754 45152 41760
rect 44928 41670 45140 41698
rect 45008 41472 45060 41478
rect 45008 41414 45060 41420
rect 44824 41064 44876 41070
rect 44824 41006 44876 41012
rect 43536 40656 43588 40662
rect 43536 40598 43588 40604
rect 44456 40656 44508 40662
rect 44456 40598 44508 40604
rect 45020 40594 45048 41414
rect 45112 41002 45140 41670
rect 45100 40996 45152 41002
rect 45100 40938 45152 40944
rect 45204 40662 45232 42026
rect 45388 40662 45416 42078
rect 45480 41274 45508 42094
rect 45848 41682 45876 42638
rect 45836 41676 45888 41682
rect 45836 41618 45888 41624
rect 45928 41676 45980 41682
rect 45928 41618 45980 41624
rect 45940 41585 45968 41618
rect 45926 41576 45982 41585
rect 45926 41511 45982 41520
rect 46768 41478 46796 42706
rect 47872 41682 47900 43046
rect 48056 42226 48084 43794
rect 49148 43784 49200 43790
rect 49148 43726 49200 43732
rect 48688 43376 48740 43382
rect 48688 43318 48740 43324
rect 48700 42702 48728 43318
rect 48964 43240 49016 43246
rect 48964 43182 49016 43188
rect 48688 42696 48740 42702
rect 48688 42638 48740 42644
rect 48044 42220 48096 42226
rect 48044 42162 48096 42168
rect 48700 42158 48728 42638
rect 48976 42226 49004 43182
rect 49056 42764 49108 42770
rect 49056 42706 49108 42712
rect 48964 42220 49016 42226
rect 48964 42162 49016 42168
rect 48688 42152 48740 42158
rect 48688 42094 48740 42100
rect 47860 41676 47912 41682
rect 47860 41618 47912 41624
rect 46756 41472 46808 41478
rect 46756 41414 46808 41420
rect 45468 41268 45520 41274
rect 45468 41210 45520 41216
rect 46294 40896 46350 40905
rect 46294 40831 46350 40840
rect 46308 40730 46336 40831
rect 46296 40724 46348 40730
rect 46296 40666 46348 40672
rect 45192 40656 45244 40662
rect 45192 40598 45244 40604
rect 45376 40656 45428 40662
rect 45376 40598 45428 40604
rect 43352 40588 43404 40594
rect 43352 40530 43404 40536
rect 45008 40588 45060 40594
rect 45008 40530 45060 40536
rect 43076 39840 43128 39846
rect 43076 39782 43128 39788
rect 43088 39522 43116 39782
rect 43088 39494 43300 39522
rect 43088 39302 43116 39494
rect 43272 39438 43300 39494
rect 43260 39432 43312 39438
rect 43260 39374 43312 39380
rect 43168 39364 43220 39370
rect 43168 39306 43220 39312
rect 43076 39296 43128 39302
rect 43076 39238 43128 39244
rect 42982 38992 43038 39001
rect 42982 38927 43038 38936
rect 41696 38752 41748 38758
rect 41696 38694 41748 38700
rect 42524 38752 42576 38758
rect 42524 38694 42576 38700
rect 42892 38752 42944 38758
rect 42892 38694 42944 38700
rect 41236 38344 41288 38350
rect 41236 38286 41288 38292
rect 40868 38276 40920 38282
rect 40868 38218 40920 38224
rect 41512 38208 41564 38214
rect 41512 38150 41564 38156
rect 42064 38208 42116 38214
rect 42064 38150 42116 38156
rect 41420 37868 41472 37874
rect 41420 37810 41472 37816
rect 40592 37800 40644 37806
rect 40592 37742 40644 37748
rect 40604 37330 40632 37742
rect 41432 37670 41460 37810
rect 41420 37664 41472 37670
rect 41420 37606 41472 37612
rect 40592 37324 40644 37330
rect 40592 37266 40644 37272
rect 40868 37120 40920 37126
rect 40868 37062 40920 37068
rect 40880 36650 40908 37062
rect 41326 36952 41382 36961
rect 41524 36922 41552 38150
rect 42076 37942 42104 38150
rect 42064 37936 42116 37942
rect 42064 37878 42116 37884
rect 41880 37800 41932 37806
rect 41880 37742 41932 37748
rect 41604 37664 41656 37670
rect 41604 37606 41656 37612
rect 41326 36887 41328 36896
rect 41380 36887 41382 36896
rect 41512 36916 41564 36922
rect 41328 36858 41380 36864
rect 41512 36858 41564 36864
rect 41420 36848 41472 36854
rect 41420 36790 41472 36796
rect 41328 36712 41380 36718
rect 41432 36700 41460 36790
rect 41380 36672 41460 36700
rect 41328 36654 41380 36660
rect 40868 36644 40920 36650
rect 40868 36586 40920 36592
rect 41512 36576 41564 36582
rect 41512 36518 41564 36524
rect 41328 36372 41380 36378
rect 41524 36360 41552 36518
rect 41380 36332 41552 36360
rect 41328 36314 41380 36320
rect 40684 36236 40736 36242
rect 40684 36178 40736 36184
rect 40224 36168 40276 36174
rect 40224 36110 40276 36116
rect 40236 36038 40264 36110
rect 40224 36032 40276 36038
rect 40224 35974 40276 35980
rect 40236 35193 40264 35974
rect 40696 35193 40724 36178
rect 40776 35828 40828 35834
rect 40776 35770 40828 35776
rect 40868 35828 40920 35834
rect 40868 35770 40920 35776
rect 40788 35630 40816 35770
rect 40880 35737 40908 35770
rect 41328 35760 41380 35766
rect 40866 35728 40922 35737
rect 41328 35702 41380 35708
rect 40866 35663 40922 35672
rect 40776 35624 40828 35630
rect 41236 35624 41288 35630
rect 40776 35566 40828 35572
rect 40880 35584 41236 35612
rect 40222 35184 40278 35193
rect 40222 35119 40278 35128
rect 40682 35184 40738 35193
rect 40682 35119 40738 35128
rect 40236 35086 40264 35119
rect 40224 35080 40276 35086
rect 40224 35022 40276 35028
rect 40880 35018 40908 35584
rect 41236 35566 41288 35572
rect 41234 35320 41290 35329
rect 41340 35290 41368 35702
rect 41510 35320 41566 35329
rect 41234 35255 41236 35264
rect 41288 35255 41290 35264
rect 41328 35284 41380 35290
rect 41236 35226 41288 35232
rect 41510 35255 41566 35264
rect 41328 35226 41380 35232
rect 41524 35222 41552 35255
rect 41512 35216 41564 35222
rect 41418 35184 41474 35193
rect 40972 35154 41276 35170
rect 40972 35148 41288 35154
rect 40972 35142 41236 35148
rect 40972 35086 41000 35142
rect 41512 35158 41564 35164
rect 41418 35119 41420 35128
rect 41236 35090 41288 35096
rect 41472 35119 41474 35128
rect 41420 35090 41472 35096
rect 40960 35080 41012 35086
rect 40960 35022 41012 35028
rect 40868 35012 40920 35018
rect 40868 34954 40920 34960
rect 40408 34944 40460 34950
rect 40408 34886 40460 34892
rect 40420 34678 40448 34886
rect 40408 34672 40460 34678
rect 40408 34614 40460 34620
rect 40040 32292 40092 32298
rect 40040 32234 40092 32240
rect 33508 31476 33560 31482
rect 33508 31418 33560 31424
rect 41616 31278 41644 37606
rect 41892 37330 41920 37742
rect 41880 37324 41932 37330
rect 41880 37266 41932 37272
rect 41696 36780 41748 36786
rect 41696 36722 41748 36728
rect 41708 36378 41736 36722
rect 42536 36582 42564 38694
rect 42616 37800 42668 37806
rect 42616 37742 42668 37748
rect 42628 37641 42656 37742
rect 42614 37632 42670 37641
rect 42614 37567 42670 37576
rect 42628 37398 42656 37567
rect 42616 37392 42668 37398
rect 42616 37334 42668 37340
rect 42524 36576 42576 36582
rect 42524 36518 42576 36524
rect 41696 36372 41748 36378
rect 41696 36314 41748 36320
rect 41788 36372 41840 36378
rect 41788 36314 41840 36320
rect 41800 36242 41828 36314
rect 41788 36236 41840 36242
rect 41788 36178 41840 36184
rect 42248 36236 42300 36242
rect 42248 36178 42300 36184
rect 41972 35760 42024 35766
rect 41972 35702 42024 35708
rect 41984 35222 42012 35702
rect 41972 35216 42024 35222
rect 42260 35193 42288 36178
rect 42522 35864 42578 35873
rect 42522 35799 42578 35808
rect 41972 35158 42024 35164
rect 42246 35184 42302 35193
rect 42246 35119 42248 35128
rect 42300 35119 42302 35128
rect 42248 35090 42300 35096
rect 42260 35059 42288 35090
rect 42536 35086 42564 35799
rect 42708 35556 42760 35562
rect 42708 35498 42760 35504
rect 42524 35080 42576 35086
rect 42524 35022 42576 35028
rect 42720 34746 42748 35498
rect 42708 34740 42760 34746
rect 42708 34682 42760 34688
rect 42064 34536 42116 34542
rect 42064 34478 42116 34484
rect 42076 34134 42104 34478
rect 42064 34128 42116 34134
rect 42064 34070 42116 34076
rect 43088 31822 43116 39238
rect 43180 38962 43208 39306
rect 43272 39273 43300 39374
rect 43258 39264 43314 39273
rect 43258 39199 43314 39208
rect 43168 38956 43220 38962
rect 43168 38898 43220 38904
rect 43260 38752 43312 38758
rect 43258 38720 43260 38729
rect 43312 38720 43314 38729
rect 43258 38655 43314 38664
rect 43364 37330 43392 40530
rect 43628 40384 43680 40390
rect 43628 40326 43680 40332
rect 43536 39976 43588 39982
rect 43536 39918 43588 39924
rect 43548 39506 43576 39918
rect 43536 39500 43588 39506
rect 43536 39442 43588 39448
rect 43534 39400 43590 39409
rect 43534 39335 43590 39344
rect 43548 39030 43576 39335
rect 43640 39030 43668 40326
rect 44640 40112 44692 40118
rect 44640 40054 44692 40060
rect 43996 39976 44048 39982
rect 43916 39936 43996 39964
rect 43720 39908 43772 39914
rect 43720 39850 43772 39856
rect 43732 39574 43760 39850
rect 43720 39568 43772 39574
rect 43720 39510 43772 39516
rect 43812 39568 43864 39574
rect 43812 39510 43864 39516
rect 43720 39432 43772 39438
rect 43824 39420 43852 39510
rect 43772 39392 43852 39420
rect 43720 39374 43772 39380
rect 43536 39024 43588 39030
rect 43536 38966 43588 38972
rect 43628 39024 43680 39030
rect 43628 38966 43680 38972
rect 43548 38894 43576 38966
rect 43536 38888 43588 38894
rect 43536 38830 43588 38836
rect 43916 38418 43944 39936
rect 43996 39918 44048 39924
rect 44272 39840 44324 39846
rect 44272 39782 44324 39788
rect 44548 39840 44600 39846
rect 44548 39782 44600 39788
rect 44088 39500 44140 39506
rect 44088 39442 44140 39448
rect 44180 39500 44232 39506
rect 44180 39442 44232 39448
rect 43994 39400 44050 39409
rect 44100 39370 44128 39442
rect 43994 39335 43996 39344
rect 44048 39335 44050 39344
rect 44088 39364 44140 39370
rect 43996 39306 44048 39312
rect 44088 39306 44140 39312
rect 44192 39273 44220 39442
rect 44178 39264 44234 39273
rect 44178 39199 44234 39208
rect 43996 39024 44048 39030
rect 43996 38966 44048 38972
rect 43904 38412 43956 38418
rect 43904 38354 43956 38360
rect 43444 37664 43496 37670
rect 43442 37632 43444 37641
rect 43496 37632 43498 37641
rect 43442 37567 43498 37576
rect 43352 37324 43404 37330
rect 43352 37266 43404 37272
rect 44008 36922 44036 38966
rect 44284 38962 44312 39782
rect 44456 39296 44508 39302
rect 44456 39238 44508 39244
rect 44468 39137 44496 39238
rect 44454 39128 44510 39137
rect 44454 39063 44510 39072
rect 44560 39030 44588 39782
rect 44652 39574 44680 40054
rect 44640 39568 44692 39574
rect 44640 39510 44692 39516
rect 44824 39500 44876 39506
rect 44824 39442 44876 39448
rect 44640 39432 44692 39438
rect 44638 39400 44640 39409
rect 44692 39400 44694 39409
rect 44836 39370 44864 39442
rect 44638 39335 44694 39344
rect 44824 39364 44876 39370
rect 44824 39306 44876 39312
rect 44548 39024 44600 39030
rect 44548 38966 44600 38972
rect 44272 38956 44324 38962
rect 44272 38898 44324 38904
rect 46020 38548 46072 38554
rect 46020 38490 46072 38496
rect 46112 38548 46164 38554
rect 46112 38490 46164 38496
rect 46032 37942 46060 38490
rect 46124 38321 46152 38490
rect 46110 38312 46166 38321
rect 46110 38247 46166 38256
rect 46296 38208 46348 38214
rect 46296 38150 46348 38156
rect 46020 37936 46072 37942
rect 46020 37878 46072 37884
rect 46308 37738 46336 38150
rect 44180 37732 44232 37738
rect 44180 37674 44232 37680
rect 46112 37732 46164 37738
rect 46112 37674 46164 37680
rect 46296 37732 46348 37738
rect 46296 37674 46348 37680
rect 43996 36916 44048 36922
rect 43996 36858 44048 36864
rect 44192 36718 44220 37674
rect 46124 37126 46152 37674
rect 46112 37120 46164 37126
rect 46112 37062 46164 37068
rect 46124 36718 46152 37062
rect 43996 36712 44048 36718
rect 43996 36654 44048 36660
rect 44180 36712 44232 36718
rect 44180 36654 44232 36660
rect 44548 36712 44600 36718
rect 44548 36654 44600 36660
rect 46112 36712 46164 36718
rect 46112 36654 46164 36660
rect 44008 36242 44036 36654
rect 44560 36378 44588 36654
rect 44548 36372 44600 36378
rect 44548 36314 44600 36320
rect 46018 36272 46074 36281
rect 43536 36236 43588 36242
rect 43536 36178 43588 36184
rect 43720 36236 43772 36242
rect 43720 36178 43772 36184
rect 43996 36236 44048 36242
rect 46018 36207 46020 36216
rect 43996 36178 44048 36184
rect 46072 36207 46074 36216
rect 46020 36178 46072 36184
rect 43548 36145 43576 36178
rect 43534 36136 43590 36145
rect 43534 36071 43590 36080
rect 43628 35692 43680 35698
rect 43628 35634 43680 35640
rect 43352 35488 43404 35494
rect 43352 35430 43404 35436
rect 43364 35018 43392 35430
rect 43352 35012 43404 35018
rect 43352 34954 43404 34960
rect 43640 34746 43668 35634
rect 43732 35222 43760 36178
rect 44916 36168 44968 36174
rect 44914 36136 44916 36145
rect 45836 36168 45888 36174
rect 44968 36136 44970 36145
rect 45836 36110 45888 36116
rect 44914 36071 44970 36080
rect 45848 36009 45876 36110
rect 45834 36000 45890 36009
rect 45834 35935 45890 35944
rect 43720 35216 43772 35222
rect 43720 35158 43772 35164
rect 43628 34740 43680 34746
rect 43628 34682 43680 34688
rect 46124 32502 46152 36654
rect 46768 34746 46796 41414
rect 48872 40044 48924 40050
rect 48872 39986 48924 39992
rect 47676 39976 47728 39982
rect 48136 39976 48188 39982
rect 47676 39918 47728 39924
rect 48056 39936 48136 39964
rect 47398 38992 47454 39001
rect 47398 38927 47400 38936
rect 47452 38927 47454 38936
rect 47400 38898 47452 38904
rect 47584 38888 47636 38894
rect 47584 38830 47636 38836
rect 47596 38758 47624 38830
rect 47584 38752 47636 38758
rect 47584 38694 47636 38700
rect 47688 38418 47716 39918
rect 48056 38894 48084 39936
rect 48136 39918 48188 39924
rect 48596 39840 48648 39846
rect 48594 39808 48596 39817
rect 48688 39840 48740 39846
rect 48648 39808 48650 39817
rect 48688 39782 48740 39788
rect 48594 39743 48650 39752
rect 48134 39672 48190 39681
rect 48134 39607 48190 39616
rect 48044 38888 48096 38894
rect 47858 38856 47914 38865
rect 48044 38830 48096 38836
rect 47858 38791 47860 38800
rect 47912 38791 47914 38800
rect 47860 38762 47912 38768
rect 48056 38729 48084 38830
rect 48148 38758 48176 39607
rect 48700 39574 48728 39782
rect 48688 39568 48740 39574
rect 48688 39510 48740 39516
rect 48780 39500 48832 39506
rect 48780 39442 48832 39448
rect 48688 39432 48740 39438
rect 48792 39409 48820 39442
rect 48688 39374 48740 39380
rect 48778 39400 48834 39409
rect 48700 39273 48728 39374
rect 48778 39335 48834 39344
rect 48686 39264 48742 39273
rect 48686 39199 48742 39208
rect 48884 39030 48912 39986
rect 48976 39506 49004 42162
rect 49068 42158 49096 42706
rect 49160 42634 49188 43726
rect 49240 43648 49292 43654
rect 49240 43590 49292 43596
rect 49252 43246 49280 43590
rect 49804 43246 49832 43794
rect 49240 43240 49292 43246
rect 49240 43182 49292 43188
rect 49792 43240 49844 43246
rect 49792 43182 49844 43188
rect 50804 43240 50856 43246
rect 50804 43182 50856 43188
rect 55772 43240 55824 43246
rect 55772 43182 55824 43188
rect 49332 43172 49384 43178
rect 49332 43114 49384 43120
rect 49344 42838 49372 43114
rect 49976 43104 50028 43110
rect 49976 43046 50028 43052
rect 49332 42832 49384 42838
rect 49332 42774 49384 42780
rect 49332 42696 49384 42702
rect 49332 42638 49384 42644
rect 49148 42628 49200 42634
rect 49148 42570 49200 42576
rect 49148 42288 49200 42294
rect 49148 42230 49200 42236
rect 49056 42152 49108 42158
rect 49056 42094 49108 42100
rect 49068 41818 49096 42094
rect 49160 42022 49188 42230
rect 49344 42158 49372 42638
rect 49988 42566 50016 43046
rect 50300 43004 50596 43024
rect 50356 43002 50380 43004
rect 50436 43002 50460 43004
rect 50516 43002 50540 43004
rect 50378 42950 50380 43002
rect 50442 42950 50454 43002
rect 50516 42950 50518 43002
rect 50356 42948 50380 42950
rect 50436 42948 50460 42950
rect 50516 42948 50540 42950
rect 50300 42928 50596 42948
rect 50816 42906 50844 43182
rect 55220 43172 55272 43178
rect 55220 43114 55272 43120
rect 50804 42900 50856 42906
rect 50804 42842 50856 42848
rect 50620 42764 50672 42770
rect 50620 42706 50672 42712
rect 49976 42560 50028 42566
rect 49976 42502 50028 42508
rect 49332 42152 49384 42158
rect 49332 42094 49384 42100
rect 49424 42084 49476 42090
rect 49424 42026 49476 42032
rect 49148 42016 49200 42022
rect 49148 41958 49200 41964
rect 49056 41812 49108 41818
rect 49056 41754 49108 41760
rect 49436 41002 49464 42026
rect 49424 40996 49476 41002
rect 49424 40938 49476 40944
rect 49148 39976 49200 39982
rect 49148 39918 49200 39924
rect 48964 39500 49016 39506
rect 48964 39442 49016 39448
rect 49160 39030 49188 39918
rect 49988 39574 50016 42502
rect 50632 42158 50660 42706
rect 55232 42702 55260 43114
rect 55784 42906 55812 43182
rect 55772 42900 55824 42906
rect 55772 42842 55824 42848
rect 53748 42696 53800 42702
rect 53748 42638 53800 42644
rect 55220 42696 55272 42702
rect 55220 42638 55272 42644
rect 51080 42560 51132 42566
rect 51080 42502 51132 42508
rect 51092 42362 51120 42502
rect 51080 42356 51132 42362
rect 51080 42298 51132 42304
rect 53760 42226 53788 42638
rect 55956 42560 56008 42566
rect 55956 42502 56008 42508
rect 53748 42220 53800 42226
rect 53748 42162 53800 42168
rect 50620 42152 50672 42158
rect 50620 42094 50672 42100
rect 52000 42152 52052 42158
rect 52000 42094 52052 42100
rect 50300 41916 50596 41936
rect 50356 41914 50380 41916
rect 50436 41914 50460 41916
rect 50516 41914 50540 41916
rect 50378 41862 50380 41914
rect 50442 41862 50454 41914
rect 50516 41862 50518 41914
rect 50356 41860 50380 41862
rect 50436 41860 50460 41862
rect 50516 41860 50540 41862
rect 50300 41840 50596 41860
rect 50632 41546 50660 42094
rect 51446 41984 51502 41993
rect 51446 41919 51502 41928
rect 51460 41750 51488 41919
rect 52012 41818 52040 42094
rect 52276 42016 52328 42022
rect 52276 41958 52328 41964
rect 51632 41812 51684 41818
rect 52000 41812 52052 41818
rect 51684 41772 51856 41800
rect 51632 41754 51684 41760
rect 51448 41744 51500 41750
rect 51448 41686 51500 41692
rect 51552 41682 51764 41698
rect 51552 41676 51776 41682
rect 51552 41670 51724 41676
rect 51552 41614 51580 41670
rect 51724 41618 51776 41624
rect 51540 41608 51592 41614
rect 51540 41550 51592 41556
rect 50620 41540 50672 41546
rect 50620 41482 50672 41488
rect 51828 41274 51856 41772
rect 52000 41754 52052 41760
rect 52184 41608 52236 41614
rect 52184 41550 52236 41556
rect 52196 41478 52224 41550
rect 52184 41472 52236 41478
rect 52184 41414 52236 41420
rect 51816 41268 51868 41274
rect 51816 41210 51868 41216
rect 50300 40828 50596 40848
rect 50356 40826 50380 40828
rect 50436 40826 50460 40828
rect 50516 40826 50540 40828
rect 50378 40774 50380 40826
rect 50442 40774 50454 40826
rect 50516 40774 50518 40826
rect 50356 40772 50380 40774
rect 50436 40772 50460 40774
rect 50516 40772 50540 40774
rect 50300 40752 50596 40772
rect 52288 40594 52316 41958
rect 53288 41676 53340 41682
rect 53288 41618 53340 41624
rect 52552 41472 52604 41478
rect 52552 41414 52604 41420
rect 52460 41064 52512 41070
rect 52564 41052 52592 41414
rect 53104 41268 53156 41274
rect 53104 41210 53156 41216
rect 53116 41070 53144 41210
rect 52512 41024 52592 41052
rect 52920 41064 52972 41070
rect 52460 41006 52512 41012
rect 52920 41006 52972 41012
rect 53104 41064 53156 41070
rect 53104 41006 53156 41012
rect 52276 40588 52328 40594
rect 52276 40530 52328 40536
rect 52184 39908 52236 39914
rect 52184 39850 52236 39856
rect 50300 39740 50596 39760
rect 50356 39738 50380 39740
rect 50436 39738 50460 39740
rect 50516 39738 50540 39740
rect 50378 39686 50380 39738
rect 50442 39686 50454 39738
rect 50516 39686 50518 39738
rect 50356 39684 50380 39686
rect 50436 39684 50460 39686
rect 50516 39684 50540 39686
rect 50300 39664 50596 39684
rect 52196 39658 52224 39850
rect 52288 39846 52316 40530
rect 52472 39982 52500 41006
rect 52932 40526 52960 41006
rect 53116 40594 53144 41006
rect 53104 40588 53156 40594
rect 53104 40530 53156 40536
rect 52920 40520 52972 40526
rect 52920 40462 52972 40468
rect 53300 40390 53328 41618
rect 53472 40996 53524 41002
rect 53472 40938 53524 40944
rect 53380 40928 53432 40934
rect 53378 40896 53380 40905
rect 53432 40896 53434 40905
rect 53378 40831 53434 40840
rect 53288 40384 53340 40390
rect 53288 40326 53340 40332
rect 52460 39976 52512 39982
rect 52460 39918 52512 39924
rect 52552 39976 52604 39982
rect 52552 39918 52604 39924
rect 52564 39846 52592 39918
rect 52276 39840 52328 39846
rect 52276 39782 52328 39788
rect 52552 39840 52604 39846
rect 52552 39782 52604 39788
rect 52196 39630 52316 39658
rect 49976 39568 50028 39574
rect 52000 39568 52052 39574
rect 49976 39510 50028 39516
rect 51998 39536 52000 39545
rect 52052 39536 52054 39545
rect 50988 39500 51040 39506
rect 50988 39442 51040 39448
rect 51724 39500 51776 39506
rect 51998 39471 52054 39480
rect 51724 39442 51776 39448
rect 49240 39432 49292 39438
rect 49240 39374 49292 39380
rect 49332 39432 49384 39438
rect 49332 39374 49384 39380
rect 48872 39024 48924 39030
rect 48686 38992 48742 39001
rect 48872 38966 48924 38972
rect 49148 39024 49200 39030
rect 49148 38966 49200 38972
rect 48686 38927 48742 38936
rect 48136 38752 48188 38758
rect 48042 38720 48098 38729
rect 48136 38694 48188 38700
rect 48412 38752 48464 38758
rect 48504 38752 48556 38758
rect 48464 38700 48504 38706
rect 48412 38694 48556 38700
rect 48424 38678 48544 38694
rect 48042 38655 48098 38664
rect 47676 38412 47728 38418
rect 47676 38354 47728 38360
rect 47676 38208 47728 38214
rect 47676 38150 47728 38156
rect 47768 38208 47820 38214
rect 47768 38150 47820 38156
rect 47688 37806 47716 38150
rect 47780 38010 47808 38150
rect 47768 38004 47820 38010
rect 47768 37946 47820 37952
rect 48700 37806 48728 38927
rect 49252 37942 49280 39374
rect 49344 39098 49372 39374
rect 50160 39296 50212 39302
rect 50160 39238 50212 39244
rect 49332 39092 49384 39098
rect 49332 39034 49384 39040
rect 50172 38418 50200 39238
rect 50300 38652 50596 38672
rect 50356 38650 50380 38652
rect 50436 38650 50460 38652
rect 50516 38650 50540 38652
rect 50378 38598 50380 38650
rect 50442 38598 50454 38650
rect 50516 38598 50518 38650
rect 50356 38596 50380 38598
rect 50436 38596 50460 38598
rect 50516 38596 50540 38598
rect 50300 38576 50596 38596
rect 50160 38412 50212 38418
rect 50160 38354 50212 38360
rect 50172 38282 50200 38354
rect 49700 38276 49752 38282
rect 49700 38218 49752 38224
rect 50160 38276 50212 38282
rect 50160 38218 50212 38224
rect 49240 37936 49292 37942
rect 49240 37878 49292 37884
rect 47676 37800 47728 37806
rect 47676 37742 47728 37748
rect 48688 37800 48740 37806
rect 48688 37742 48740 37748
rect 47032 37664 47084 37670
rect 47032 37606 47084 37612
rect 46848 36916 46900 36922
rect 46848 36858 46900 36864
rect 46860 36718 46888 36858
rect 46940 36848 46992 36854
rect 46940 36790 46992 36796
rect 46848 36712 46900 36718
rect 46848 36654 46900 36660
rect 46952 36310 46980 36790
rect 47044 36718 47072 37606
rect 47216 37324 47268 37330
rect 47216 37266 47268 37272
rect 47228 36854 47256 37266
rect 47306 36952 47362 36961
rect 47306 36887 47362 36896
rect 47320 36854 47348 36887
rect 47216 36848 47268 36854
rect 47216 36790 47268 36796
rect 47308 36848 47360 36854
rect 47308 36790 47360 36796
rect 47032 36712 47084 36718
rect 47032 36654 47084 36660
rect 46940 36304 46992 36310
rect 46940 36246 46992 36252
rect 46940 36168 46992 36174
rect 47044 36156 47072 36654
rect 47688 36242 47716 37742
rect 48700 37398 48728 37742
rect 49712 37398 49740 38218
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 48688 37392 48740 37398
rect 48688 37334 48740 37340
rect 49700 37392 49752 37398
rect 49700 37334 49752 37340
rect 51000 37330 51028 39442
rect 51736 38418 51764 39442
rect 51816 38480 51868 38486
rect 51868 38428 52224 38434
rect 51816 38422 52224 38428
rect 51724 38412 51776 38418
rect 51828 38406 52224 38422
rect 51724 38354 51776 38360
rect 51540 38344 51592 38350
rect 51540 38286 51592 38292
rect 51816 38344 51868 38350
rect 51816 38286 51868 38292
rect 50988 37324 51040 37330
rect 50988 37266 51040 37272
rect 50344 37256 50396 37262
rect 49988 37216 50344 37244
rect 49240 36780 49292 36786
rect 49240 36722 49292 36728
rect 48412 36712 48464 36718
rect 48412 36654 48464 36660
rect 47676 36236 47728 36242
rect 47676 36178 47728 36184
rect 46992 36128 47072 36156
rect 46940 36110 46992 36116
rect 48424 34746 48452 36654
rect 49056 36236 49108 36242
rect 49056 36178 49108 36184
rect 48964 35828 49016 35834
rect 48964 35770 49016 35776
rect 48976 35562 49004 35770
rect 49068 35698 49096 36178
rect 49148 36032 49200 36038
rect 49148 35974 49200 35980
rect 49056 35692 49108 35698
rect 49056 35634 49108 35640
rect 48964 35556 49016 35562
rect 48964 35498 49016 35504
rect 49068 35494 49096 35634
rect 49056 35488 49108 35494
rect 49056 35430 49108 35436
rect 48962 35048 49018 35057
rect 48962 34983 49018 34992
rect 48872 34944 48924 34950
rect 48872 34886 48924 34892
rect 48884 34746 48912 34886
rect 46756 34740 46808 34746
rect 46756 34682 46808 34688
rect 48412 34740 48464 34746
rect 48412 34682 48464 34688
rect 48872 34740 48924 34746
rect 48872 34682 48924 34688
rect 46662 34640 46718 34649
rect 46662 34575 46664 34584
rect 46716 34575 46718 34584
rect 48424 34626 48452 34682
rect 48424 34598 48636 34626
rect 46664 34546 46716 34552
rect 48320 34400 48372 34406
rect 48424 34388 48452 34598
rect 48608 34406 48636 34598
rect 48884 34542 48912 34682
rect 48976 34610 49004 34983
rect 48964 34604 49016 34610
rect 48964 34546 49016 34552
rect 48872 34536 48924 34542
rect 48872 34478 48924 34484
rect 48372 34360 48452 34388
rect 48504 34400 48556 34406
rect 48320 34342 48372 34348
rect 48504 34342 48556 34348
rect 48596 34400 48648 34406
rect 48596 34342 48648 34348
rect 46112 32496 46164 32502
rect 46112 32438 46164 32444
rect 48516 32026 48544 34342
rect 49068 32638 49096 35430
rect 49160 35193 49188 35974
rect 49252 35612 49280 36722
rect 49700 36712 49752 36718
rect 49700 36654 49752 36660
rect 49516 36032 49568 36038
rect 49516 35974 49568 35980
rect 49424 35624 49476 35630
rect 49252 35584 49424 35612
rect 49252 35494 49280 35584
rect 49424 35566 49476 35572
rect 49528 35494 49556 35974
rect 49712 35834 49740 36654
rect 49988 36378 50016 37216
rect 50344 37198 50396 37204
rect 50986 37224 51042 37233
rect 50986 37159 51042 37168
rect 51000 37126 51028 37159
rect 50988 37120 51040 37126
rect 50988 37062 51040 37068
rect 50712 36848 50764 36854
rect 50712 36790 50764 36796
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 49976 36372 50028 36378
rect 49976 36314 50028 36320
rect 49790 36272 49846 36281
rect 50724 36242 50752 36790
rect 50804 36712 50856 36718
rect 50802 36680 50804 36689
rect 50856 36680 50858 36689
rect 50802 36615 50858 36624
rect 49790 36207 49846 36216
rect 50160 36236 50212 36242
rect 49804 36174 49832 36207
rect 50160 36178 50212 36184
rect 50712 36236 50764 36242
rect 50712 36178 50764 36184
rect 49792 36168 49844 36174
rect 49792 36110 49844 36116
rect 49700 35828 49752 35834
rect 49700 35770 49752 35776
rect 49712 35630 49740 35770
rect 49700 35624 49752 35630
rect 49700 35566 49752 35572
rect 50172 35494 50200 36178
rect 50816 35834 50844 36615
rect 51552 36310 51580 38286
rect 51632 38004 51684 38010
rect 51632 37946 51684 37952
rect 51644 36922 51672 37946
rect 51828 37874 51856 38286
rect 51816 37868 51868 37874
rect 51816 37810 51868 37816
rect 51724 37392 51776 37398
rect 51724 37334 51776 37340
rect 51632 36916 51684 36922
rect 51632 36858 51684 36864
rect 51736 36718 51764 37334
rect 51828 36922 51856 37810
rect 52000 37800 52052 37806
rect 52000 37742 52052 37748
rect 51908 37732 51960 37738
rect 51908 37674 51960 37680
rect 51920 37641 51948 37674
rect 51906 37632 51962 37641
rect 51906 37567 51962 37576
rect 52012 37330 52040 37742
rect 52196 37670 52224 38406
rect 52288 37788 52316 39630
rect 52564 39506 52592 39782
rect 53300 39658 53328 40326
rect 53208 39630 53328 39658
rect 53208 39574 53236 39630
rect 53196 39568 53248 39574
rect 53196 39510 53248 39516
rect 53484 39506 53512 40938
rect 53760 39982 53788 42162
rect 55968 42158 55996 42502
rect 56152 42226 56180 45440
rect 67272 44192 67324 44198
rect 67272 44134 67324 44140
rect 61936 43852 61988 43858
rect 61936 43794 61988 43800
rect 63040 43852 63092 43858
rect 63040 43794 63092 43800
rect 61108 43308 61160 43314
rect 61108 43250 61160 43256
rect 56232 43240 56284 43246
rect 56232 43182 56284 43188
rect 59544 43240 59596 43246
rect 59544 43182 59596 43188
rect 56244 42770 56272 43182
rect 56600 43172 56652 43178
rect 56600 43114 56652 43120
rect 57888 43172 57940 43178
rect 57888 43114 57940 43120
rect 56232 42764 56284 42770
rect 56232 42706 56284 42712
rect 56140 42220 56192 42226
rect 56140 42162 56192 42168
rect 55956 42152 56008 42158
rect 55034 42120 55090 42129
rect 55956 42094 56008 42100
rect 55034 42055 55036 42064
rect 55088 42055 55090 42064
rect 55036 42026 55088 42032
rect 55404 42016 55456 42022
rect 55968 41993 55996 42094
rect 56244 42022 56272 42706
rect 56232 42016 56284 42022
rect 55404 41958 55456 41964
rect 55954 41984 56010 41993
rect 54576 41676 54628 41682
rect 54576 41618 54628 41624
rect 54588 41274 54616 41618
rect 55416 41478 55444 41958
rect 56232 41958 56284 41964
rect 55954 41919 56010 41928
rect 54668 41472 54720 41478
rect 54668 41414 54720 41420
rect 55404 41472 55456 41478
rect 55404 41414 55456 41420
rect 55496 41472 55548 41478
rect 55496 41414 55548 41420
rect 54576 41268 54628 41274
rect 54576 41210 54628 41216
rect 54484 41064 54536 41070
rect 54484 41006 54536 41012
rect 54496 40746 54524 41006
rect 54680 40746 54708 41414
rect 55508 41070 55536 41414
rect 55496 41064 55548 41070
rect 55496 41006 55548 41012
rect 56612 41002 56640 43114
rect 57900 42770 57928 43114
rect 57888 42764 57940 42770
rect 57888 42706 57940 42712
rect 58532 42696 58584 42702
rect 58532 42638 58584 42644
rect 58544 42566 58572 42638
rect 59452 42628 59504 42634
rect 59452 42570 59504 42576
rect 58532 42560 58584 42566
rect 58532 42502 58584 42508
rect 58544 42158 58572 42502
rect 59464 42294 59492 42570
rect 59176 42288 59228 42294
rect 59176 42230 59228 42236
rect 59452 42288 59504 42294
rect 59452 42230 59504 42236
rect 58532 42152 58584 42158
rect 58532 42094 58584 42100
rect 59188 41818 59216 42230
rect 58808 41812 58860 41818
rect 58808 41754 58860 41760
rect 59176 41812 59228 41818
rect 59176 41754 59228 41760
rect 57152 41676 57204 41682
rect 57152 41618 57204 41624
rect 57164 41002 57192 41618
rect 55128 40996 55180 41002
rect 55128 40938 55180 40944
rect 56600 40996 56652 41002
rect 56600 40938 56652 40944
rect 57060 40996 57112 41002
rect 57060 40938 57112 40944
rect 57152 40996 57204 41002
rect 57152 40938 57204 40944
rect 54496 40718 54708 40746
rect 55140 40594 55168 40938
rect 55956 40928 56008 40934
rect 55876 40888 55956 40916
rect 55772 40656 55824 40662
rect 55772 40598 55824 40604
rect 54760 40588 54812 40594
rect 54760 40530 54812 40536
rect 55128 40588 55180 40594
rect 55128 40530 55180 40536
rect 53748 39976 53800 39982
rect 53748 39918 53800 39924
rect 54024 39976 54076 39982
rect 54024 39918 54076 39924
rect 54116 39976 54168 39982
rect 54116 39918 54168 39924
rect 52552 39500 52604 39506
rect 52552 39442 52604 39448
rect 52828 39500 52880 39506
rect 52828 39442 52880 39448
rect 53472 39500 53524 39506
rect 53472 39442 53524 39448
rect 52840 38894 52868 39442
rect 53380 39092 53432 39098
rect 53380 39034 53432 39040
rect 53286 38992 53342 39001
rect 53286 38927 53342 38936
rect 53300 38894 53328 38927
rect 53392 38894 53420 39034
rect 52828 38888 52880 38894
rect 52828 38830 52880 38836
rect 53288 38888 53340 38894
rect 53288 38830 53340 38836
rect 53380 38888 53432 38894
rect 53380 38830 53432 38836
rect 52552 38820 52604 38826
rect 52552 38762 52604 38768
rect 52564 38554 52592 38762
rect 53392 38554 53420 38830
rect 52552 38548 52604 38554
rect 52552 38490 52604 38496
rect 53380 38548 53432 38554
rect 53380 38490 53432 38496
rect 52828 38208 52880 38214
rect 52828 38150 52880 38156
rect 53104 38208 53156 38214
rect 53104 38150 53156 38156
rect 53380 38208 53432 38214
rect 53380 38150 53432 38156
rect 52644 37800 52696 37806
rect 52288 37760 52644 37788
rect 52644 37742 52696 37748
rect 52092 37664 52144 37670
rect 52092 37606 52144 37612
rect 52184 37664 52236 37670
rect 52184 37606 52236 37612
rect 52104 37466 52132 37606
rect 52840 37466 52868 38150
rect 52092 37460 52144 37466
rect 52092 37402 52144 37408
rect 52828 37460 52880 37466
rect 52828 37402 52880 37408
rect 53116 37330 53144 38150
rect 53392 37874 53420 38150
rect 53380 37868 53432 37874
rect 53380 37810 53432 37816
rect 53484 37330 53512 39442
rect 53760 39080 53788 39918
rect 54036 39574 54064 39918
rect 54024 39568 54076 39574
rect 54024 39510 54076 39516
rect 54128 39080 54156 39918
rect 54574 39536 54630 39545
rect 54772 39506 54800 40530
rect 55784 40186 55812 40598
rect 55876 40594 55904 40888
rect 55956 40870 56008 40876
rect 57072 40662 57100 40938
rect 58820 40905 58848 41754
rect 59556 41750 59584 43182
rect 61120 43110 61148 43250
rect 60832 43104 60884 43110
rect 60832 43046 60884 43052
rect 61108 43104 61160 43110
rect 61108 43046 61160 43052
rect 60844 42770 60872 43046
rect 60832 42764 60884 42770
rect 60832 42706 60884 42712
rect 61120 42702 61148 43046
rect 61108 42696 61160 42702
rect 61108 42638 61160 42644
rect 60372 42560 60424 42566
rect 60372 42502 60424 42508
rect 60832 42560 60884 42566
rect 60832 42502 60884 42508
rect 59636 42016 59688 42022
rect 59636 41958 59688 41964
rect 59544 41744 59596 41750
rect 59544 41686 59596 41692
rect 59648 41682 59676 41958
rect 59636 41676 59688 41682
rect 59636 41618 59688 41624
rect 60384 41614 60412 42502
rect 60372 41608 60424 41614
rect 60372 41550 60424 41556
rect 60648 41200 60700 41206
rect 60646 41168 60648 41177
rect 60700 41168 60702 41177
rect 60646 41103 60702 41112
rect 60844 41070 60872 42502
rect 61948 42226 61976 43794
rect 62212 43648 62264 43654
rect 62212 43590 62264 43596
rect 62224 42770 62252 43590
rect 62212 42764 62264 42770
rect 62212 42706 62264 42712
rect 63052 42362 63080 43794
rect 63500 43716 63552 43722
rect 63500 43658 63552 43664
rect 63512 42770 63540 43658
rect 65660 43548 65956 43568
rect 65716 43546 65740 43548
rect 65796 43546 65820 43548
rect 65876 43546 65900 43548
rect 65738 43494 65740 43546
rect 65802 43494 65814 43546
rect 65876 43494 65878 43546
rect 65716 43492 65740 43494
rect 65796 43492 65820 43494
rect 65876 43492 65900 43494
rect 65660 43472 65956 43492
rect 66260 43376 66312 43382
rect 66260 43318 66312 43324
rect 66168 43104 66220 43110
rect 66168 43046 66220 43052
rect 63500 42764 63552 42770
rect 63500 42706 63552 42712
rect 64604 42764 64656 42770
rect 64604 42706 64656 42712
rect 63040 42356 63092 42362
rect 63040 42298 63092 42304
rect 61016 42220 61068 42226
rect 61016 42162 61068 42168
rect 61936 42220 61988 42226
rect 61936 42162 61988 42168
rect 63868 42220 63920 42226
rect 63868 42162 63920 42168
rect 61028 41682 61056 42162
rect 61568 42152 61620 42158
rect 61752 42152 61804 42158
rect 61620 42112 61752 42140
rect 61568 42094 61620 42100
rect 61752 42094 61804 42100
rect 62028 42084 62080 42090
rect 62028 42026 62080 42032
rect 61016 41676 61068 41682
rect 61016 41618 61068 41624
rect 62040 41546 62068 42026
rect 63880 41818 63908 42162
rect 63868 41812 63920 41818
rect 63868 41754 63920 41760
rect 63592 41676 63644 41682
rect 63592 41618 63644 41624
rect 62580 41608 62632 41614
rect 62580 41550 62632 41556
rect 62028 41540 62080 41546
rect 62028 41482 62080 41488
rect 62040 41206 62068 41482
rect 62028 41200 62080 41206
rect 62028 41142 62080 41148
rect 60832 41064 60884 41070
rect 60832 41006 60884 41012
rect 61568 41064 61620 41070
rect 61568 41006 61620 41012
rect 57242 40896 57298 40905
rect 57242 40831 57298 40840
rect 58806 40896 58862 40905
rect 58806 40831 58862 40840
rect 57060 40656 57112 40662
rect 57060 40598 57112 40604
rect 55864 40588 55916 40594
rect 55864 40530 55916 40536
rect 54852 40180 54904 40186
rect 54852 40122 54904 40128
rect 55772 40180 55824 40186
rect 55772 40122 55824 40128
rect 54864 39506 54892 40122
rect 55876 40066 55904 40530
rect 57256 40526 57284 40831
rect 57244 40520 57296 40526
rect 57244 40462 57296 40468
rect 56876 40384 56928 40390
rect 56876 40326 56928 40332
rect 57336 40384 57388 40390
rect 57336 40326 57388 40332
rect 57796 40384 57848 40390
rect 57796 40326 57848 40332
rect 56888 40118 56916 40326
rect 55784 40038 55904 40066
rect 56876 40112 56928 40118
rect 56876 40054 56928 40060
rect 56048 40044 56100 40050
rect 55496 39976 55548 39982
rect 55496 39918 55548 39924
rect 55404 39568 55456 39574
rect 55404 39510 55456 39516
rect 54574 39471 54630 39480
rect 54760 39500 54812 39506
rect 54588 39302 54616 39471
rect 54760 39442 54812 39448
rect 54852 39500 54904 39506
rect 54852 39442 54904 39448
rect 55416 39302 55444 39510
rect 55508 39302 55536 39918
rect 54576 39296 54628 39302
rect 54576 39238 54628 39244
rect 55404 39296 55456 39302
rect 55404 39238 55456 39244
rect 55496 39296 55548 39302
rect 55496 39238 55548 39244
rect 53760 39052 54156 39080
rect 53564 38820 53616 38826
rect 53564 38762 53616 38768
rect 53576 38010 53604 38762
rect 53748 38752 53800 38758
rect 53748 38694 53800 38700
rect 53564 38004 53616 38010
rect 53564 37946 53616 37952
rect 53656 37800 53708 37806
rect 53656 37742 53708 37748
rect 53668 37330 53696 37742
rect 52000 37324 52052 37330
rect 52000 37266 52052 37272
rect 53012 37324 53064 37330
rect 53012 37266 53064 37272
rect 53104 37324 53156 37330
rect 53104 37266 53156 37272
rect 53472 37324 53524 37330
rect 53472 37266 53524 37272
rect 53656 37324 53708 37330
rect 53656 37266 53708 37272
rect 52460 37120 52512 37126
rect 52460 37062 52512 37068
rect 51816 36916 51868 36922
rect 51816 36858 51868 36864
rect 51724 36712 51776 36718
rect 51724 36654 51776 36660
rect 51632 36576 51684 36582
rect 51632 36518 51684 36524
rect 51172 36304 51224 36310
rect 51172 36246 51224 36252
rect 51540 36304 51592 36310
rect 51644 36281 51672 36518
rect 52472 36310 52500 37062
rect 52460 36304 52512 36310
rect 51540 36246 51592 36252
rect 51630 36272 51686 36281
rect 51184 36174 51212 36246
rect 52460 36246 52512 36252
rect 51630 36207 51686 36216
rect 51172 36168 51224 36174
rect 51172 36110 51224 36116
rect 50804 35828 50856 35834
rect 50804 35770 50856 35776
rect 50988 35556 51040 35562
rect 50988 35498 51040 35504
rect 49240 35488 49292 35494
rect 49240 35430 49292 35436
rect 49516 35488 49568 35494
rect 49516 35430 49568 35436
rect 50160 35488 50212 35494
rect 50160 35430 50212 35436
rect 49146 35184 49202 35193
rect 49146 35119 49202 35128
rect 49252 32774 49280 35430
rect 49424 35080 49476 35086
rect 49424 35022 49476 35028
rect 49332 34944 49384 34950
rect 49332 34886 49384 34892
rect 49344 32910 49372 34886
rect 49436 34785 49464 35022
rect 49528 34950 49556 35430
rect 50300 35388 50596 35408
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 51000 35272 51028 35498
rect 50724 35244 51028 35272
rect 50434 35184 50490 35193
rect 49884 35148 49936 35154
rect 50434 35119 50436 35128
rect 49884 35090 49936 35096
rect 50488 35119 50490 35128
rect 50436 35090 50488 35096
rect 49700 35080 49752 35086
rect 49700 35022 49752 35028
rect 49712 34950 49740 35022
rect 49896 34950 49924 35090
rect 49516 34944 49568 34950
rect 49516 34886 49568 34892
rect 49700 34944 49752 34950
rect 49700 34886 49752 34892
rect 49884 34944 49936 34950
rect 49884 34886 49936 34892
rect 49422 34776 49478 34785
rect 49422 34711 49478 34720
rect 50250 34776 50306 34785
rect 50250 34711 50252 34720
rect 49436 34542 49464 34711
rect 50304 34711 50306 34720
rect 50252 34682 50304 34688
rect 49792 34672 49844 34678
rect 49790 34640 49792 34649
rect 49844 34640 49846 34649
rect 50724 34626 50752 35244
rect 51184 35154 51212 36110
rect 51264 36100 51316 36106
rect 51264 36042 51316 36048
rect 51276 35193 51304 36042
rect 52000 35760 52052 35766
rect 52000 35702 52052 35708
rect 51448 35624 51500 35630
rect 51448 35566 51500 35572
rect 51262 35184 51318 35193
rect 51172 35148 51224 35154
rect 51262 35119 51318 35128
rect 51172 35090 51224 35096
rect 51184 34950 51212 35090
rect 51276 34950 51304 35119
rect 51460 35018 51488 35566
rect 52012 35222 52040 35702
rect 53024 35630 53052 37266
rect 53484 36854 53512 37266
rect 53472 36848 53524 36854
rect 53472 36790 53524 36796
rect 53760 36786 53788 38694
rect 54036 37874 54064 39052
rect 55784 38894 55812 40038
rect 56048 39986 56100 39992
rect 56060 39574 56088 39986
rect 56048 39568 56100 39574
rect 56048 39510 56100 39516
rect 57348 39506 57376 40326
rect 57808 40118 57836 40326
rect 57796 40112 57848 40118
rect 57796 40054 57848 40060
rect 57336 39500 57388 39506
rect 57336 39442 57388 39448
rect 56138 39400 56194 39409
rect 55864 39364 55916 39370
rect 56138 39335 56194 39344
rect 55864 39306 55916 39312
rect 55680 38888 55732 38894
rect 55772 38888 55824 38894
rect 55680 38830 55732 38836
rect 55770 38856 55772 38865
rect 55824 38856 55826 38865
rect 55692 38706 55720 38830
rect 55876 38826 55904 39306
rect 56048 39296 56100 39302
rect 56048 39238 56100 39244
rect 56060 38894 56088 39238
rect 56152 38962 56180 39335
rect 56230 39264 56286 39273
rect 56230 39199 56286 39208
rect 56244 39030 56272 39199
rect 56232 39024 56284 39030
rect 56232 38966 56284 38972
rect 56140 38956 56192 38962
rect 56140 38898 56192 38904
rect 56048 38888 56100 38894
rect 56048 38830 56100 38836
rect 55770 38791 55826 38800
rect 55864 38820 55916 38826
rect 55864 38762 55916 38768
rect 56060 38706 56088 38830
rect 55692 38678 56088 38706
rect 54024 37868 54076 37874
rect 54024 37810 54076 37816
rect 53932 37800 53984 37806
rect 53932 37742 53984 37748
rect 53748 36780 53800 36786
rect 53748 36722 53800 36728
rect 53944 36718 53972 37742
rect 53656 36712 53708 36718
rect 53656 36654 53708 36660
rect 53932 36712 53984 36718
rect 53932 36654 53984 36660
rect 53288 36032 53340 36038
rect 53288 35974 53340 35980
rect 53196 35692 53248 35698
rect 53196 35634 53248 35640
rect 53012 35624 53064 35630
rect 53012 35566 53064 35572
rect 53208 35222 53236 35634
rect 53300 35630 53328 35974
rect 53668 35834 53696 36654
rect 53656 35828 53708 35834
rect 53656 35770 53708 35776
rect 53288 35624 53340 35630
rect 53288 35566 53340 35572
rect 53840 35488 53892 35494
rect 53840 35430 53892 35436
rect 52000 35216 52052 35222
rect 52000 35158 52052 35164
rect 53196 35216 53248 35222
rect 53196 35158 53248 35164
rect 51816 35148 51868 35154
rect 51816 35090 51868 35096
rect 52092 35148 52144 35154
rect 52092 35090 52144 35096
rect 52644 35148 52696 35154
rect 52644 35090 52696 35096
rect 51724 35080 51776 35086
rect 51724 35022 51776 35028
rect 51448 35012 51500 35018
rect 51448 34954 51500 34960
rect 51736 34950 51764 35022
rect 51828 34950 51856 35090
rect 51172 34944 51224 34950
rect 51172 34886 51224 34892
rect 51264 34944 51316 34950
rect 51264 34886 51316 34892
rect 51540 34944 51592 34950
rect 51540 34886 51592 34892
rect 51724 34944 51776 34950
rect 51724 34886 51776 34892
rect 51816 34944 51868 34950
rect 51816 34886 51868 34892
rect 49790 34575 49846 34584
rect 50632 34598 50752 34626
rect 50632 34542 50660 34598
rect 49424 34536 49476 34542
rect 49424 34478 49476 34484
rect 50620 34536 50672 34542
rect 50620 34478 50672 34484
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 51552 34202 51580 34886
rect 52104 34746 52132 35090
rect 52656 35057 52684 35090
rect 52642 35048 52698 35057
rect 52642 34983 52698 34992
rect 53472 35012 53524 35018
rect 53472 34954 53524 34960
rect 53484 34898 53512 34954
rect 53208 34870 53512 34898
rect 53208 34746 53236 34870
rect 52092 34740 52144 34746
rect 52092 34682 52144 34688
rect 53196 34740 53248 34746
rect 53196 34682 53248 34688
rect 53852 34610 53880 35430
rect 53840 34604 53892 34610
rect 53840 34546 53892 34552
rect 53932 34400 53984 34406
rect 54036 34388 54064 37810
rect 55312 37324 55364 37330
rect 55312 37266 55364 37272
rect 54392 37120 54444 37126
rect 54392 37062 54444 37068
rect 54852 37120 54904 37126
rect 54852 37062 54904 37068
rect 54404 36922 54432 37062
rect 54392 36916 54444 36922
rect 54392 36858 54444 36864
rect 54484 36916 54536 36922
rect 54484 36858 54536 36864
rect 54300 36780 54352 36786
rect 54300 36722 54352 36728
rect 54208 36712 54260 36718
rect 54206 36680 54208 36689
rect 54260 36680 54262 36689
rect 54206 36615 54262 36624
rect 54312 36242 54340 36722
rect 54496 36378 54524 36858
rect 54864 36650 54892 37062
rect 54852 36644 54904 36650
rect 54852 36586 54904 36592
rect 55036 36576 55088 36582
rect 55036 36518 55088 36524
rect 54484 36372 54536 36378
rect 54484 36314 54536 36320
rect 54300 36236 54352 36242
rect 54300 36178 54352 36184
rect 54852 36100 54904 36106
rect 54852 36042 54904 36048
rect 54864 35834 54892 36042
rect 55048 36038 55076 36518
rect 55036 36032 55088 36038
rect 55036 35974 55088 35980
rect 55048 35834 55076 35974
rect 54852 35828 54904 35834
rect 54852 35770 54904 35776
rect 55036 35828 55088 35834
rect 55036 35770 55088 35776
rect 55048 35630 55076 35770
rect 55036 35624 55088 35630
rect 55036 35566 55088 35572
rect 55220 35556 55272 35562
rect 55220 35498 55272 35504
rect 53984 34360 54064 34388
rect 55128 34400 55180 34406
rect 53932 34342 53984 34348
rect 55128 34342 55180 34348
rect 51540 34196 51592 34202
rect 51540 34138 51592 34144
rect 55140 33046 55168 34342
rect 55128 33040 55180 33046
rect 55128 32982 55180 32988
rect 49332 32904 49384 32910
rect 49332 32846 49384 32852
rect 49240 32768 49292 32774
rect 49240 32710 49292 32716
rect 49056 32632 49108 32638
rect 49056 32574 49108 32580
rect 55140 32502 55168 32982
rect 55232 32570 55260 35498
rect 55324 34542 55352 37266
rect 55692 37233 55720 38678
rect 57808 38554 57836 40054
rect 57796 38548 57848 38554
rect 57796 38490 57848 38496
rect 58716 38004 58768 38010
rect 58716 37946 58768 37952
rect 57704 37868 57756 37874
rect 57704 37810 57756 37816
rect 57152 37664 57204 37670
rect 57152 37606 57204 37612
rect 57242 37632 57298 37641
rect 57058 37496 57114 37505
rect 57058 37431 57060 37440
rect 57112 37431 57114 37440
rect 57060 37402 57112 37408
rect 57164 37369 57192 37606
rect 57242 37567 57298 37576
rect 57256 37466 57284 37567
rect 57716 37466 57744 37810
rect 58624 37800 58676 37806
rect 58624 37742 58676 37748
rect 57794 37496 57850 37505
rect 57244 37460 57296 37466
rect 57244 37402 57296 37408
rect 57704 37460 57756 37466
rect 57794 37431 57796 37440
rect 57704 37402 57756 37408
rect 57848 37431 57850 37440
rect 57796 37402 57848 37408
rect 57150 37360 57206 37369
rect 57150 37295 57206 37304
rect 57716 37262 57744 37402
rect 57704 37256 57756 37262
rect 55678 37224 55734 37233
rect 57704 37198 57756 37204
rect 55678 37159 55734 37168
rect 56600 36576 56652 36582
rect 56600 36518 56652 36524
rect 56612 36174 56640 36518
rect 58636 36310 58664 37742
rect 58728 37330 58756 37946
rect 58716 37324 58768 37330
rect 58716 37266 58768 37272
rect 58624 36304 58676 36310
rect 58624 36246 58676 36252
rect 58728 36242 58756 37266
rect 58716 36236 58768 36242
rect 58716 36178 58768 36184
rect 56600 36168 56652 36174
rect 56600 36110 56652 36116
rect 56876 36168 56928 36174
rect 58820 36122 58848 40831
rect 60740 40656 60792 40662
rect 60740 40598 60792 40604
rect 60752 39982 60780 40598
rect 60740 39976 60792 39982
rect 60740 39918 60792 39924
rect 60844 38758 60872 41006
rect 61580 40934 61608 41006
rect 62592 40934 62620 41550
rect 63040 41472 63092 41478
rect 63040 41414 63092 41420
rect 63052 41206 63080 41414
rect 63500 41268 63552 41274
rect 63500 41210 63552 41216
rect 63040 41200 63092 41206
rect 63132 41200 63184 41206
rect 63040 41142 63092 41148
rect 63130 41168 63132 41177
rect 63184 41168 63186 41177
rect 63130 41103 63186 41112
rect 63040 41064 63092 41070
rect 63040 41006 63092 41012
rect 61568 40928 61620 40934
rect 61568 40870 61620 40876
rect 61844 40928 61896 40934
rect 61844 40870 61896 40876
rect 62580 40928 62632 40934
rect 62580 40870 62632 40876
rect 61580 40186 61608 40870
rect 61568 40180 61620 40186
rect 61568 40122 61620 40128
rect 61660 39568 61712 39574
rect 61660 39510 61712 39516
rect 61672 39302 61700 39510
rect 61856 39506 61884 40870
rect 62592 40594 62620 40870
rect 62948 40656 63000 40662
rect 62948 40598 63000 40604
rect 62304 40588 62356 40594
rect 62304 40530 62356 40536
rect 62580 40588 62632 40594
rect 62580 40530 62632 40536
rect 61936 40044 61988 40050
rect 61936 39986 61988 39992
rect 61844 39500 61896 39506
rect 61844 39442 61896 39448
rect 61948 39409 61976 39986
rect 62210 39536 62266 39545
rect 62210 39471 62212 39480
rect 62264 39471 62266 39480
rect 62212 39442 62264 39448
rect 61934 39400 61990 39409
rect 61934 39335 61990 39344
rect 61660 39296 61712 39302
rect 61660 39238 61712 39244
rect 62120 39092 62172 39098
rect 62120 39034 62172 39040
rect 62132 38826 62160 39034
rect 62316 38894 62344 40530
rect 62764 40520 62816 40526
rect 62764 40462 62816 40468
rect 62672 40452 62724 40458
rect 62672 40394 62724 40400
rect 62684 40186 62712 40394
rect 62672 40180 62724 40186
rect 62672 40122 62724 40128
rect 62776 39302 62804 40462
rect 62960 40390 62988 40598
rect 62948 40384 63000 40390
rect 62948 40326 63000 40332
rect 63052 39506 63080 41006
rect 63316 40928 63368 40934
rect 63512 40882 63540 41210
rect 63368 40876 63540 40882
rect 63316 40870 63540 40876
rect 63328 40854 63540 40870
rect 63604 39545 63632 41618
rect 63880 40662 63908 41754
rect 64512 41540 64564 41546
rect 64512 41482 64564 41488
rect 64236 41064 64288 41070
rect 64288 41012 64460 41018
rect 64236 41006 64460 41012
rect 64248 41002 64460 41006
rect 64248 40996 64472 41002
rect 64248 40990 64420 40996
rect 64420 40938 64472 40944
rect 64328 40928 64380 40934
rect 64326 40896 64328 40905
rect 64380 40896 64382 40905
rect 64326 40831 64382 40840
rect 63868 40656 63920 40662
rect 63868 40598 63920 40604
rect 63776 40588 63828 40594
rect 63776 40530 63828 40536
rect 64420 40588 64472 40594
rect 64420 40530 64472 40536
rect 63590 39536 63646 39545
rect 63040 39500 63092 39506
rect 63040 39442 63092 39448
rect 63500 39500 63552 39506
rect 63590 39471 63646 39480
rect 63500 39442 63552 39448
rect 63224 39364 63276 39370
rect 63224 39306 63276 39312
rect 62764 39296 62816 39302
rect 62764 39238 62816 39244
rect 63236 38894 63264 39306
rect 63512 39302 63540 39442
rect 63500 39296 63552 39302
rect 63500 39238 63552 39244
rect 63788 38962 63816 40530
rect 64432 40050 64460 40530
rect 64420 40044 64472 40050
rect 64420 39986 64472 39992
rect 64524 38962 64552 41482
rect 64616 40662 64644 42706
rect 66076 42696 66128 42702
rect 66076 42638 66128 42644
rect 65660 42460 65956 42480
rect 65716 42458 65740 42460
rect 65796 42458 65820 42460
rect 65876 42458 65900 42460
rect 65738 42406 65740 42458
rect 65802 42406 65814 42458
rect 65876 42406 65878 42458
rect 65716 42404 65740 42406
rect 65796 42404 65820 42406
rect 65876 42404 65900 42406
rect 65660 42384 65956 42404
rect 65708 42288 65760 42294
rect 65708 42230 65760 42236
rect 65720 41682 65748 42230
rect 66088 42226 66116 42638
rect 66076 42220 66128 42226
rect 66076 42162 66128 42168
rect 65984 42084 66036 42090
rect 65984 42026 66036 42032
rect 65708 41676 65760 41682
rect 65708 41618 65760 41624
rect 65996 41478 66024 42026
rect 66180 42022 66208 43046
rect 66272 42226 66300 43318
rect 66536 43240 66588 43246
rect 66536 43182 66588 43188
rect 66904 43240 66956 43246
rect 66904 43182 66956 43188
rect 66260 42220 66312 42226
rect 66260 42162 66312 42168
rect 66548 42090 66576 43182
rect 66812 42628 66864 42634
rect 66812 42570 66864 42576
rect 66536 42084 66588 42090
rect 66536 42026 66588 42032
rect 66168 42016 66220 42022
rect 66168 41958 66220 41964
rect 65984 41472 66036 41478
rect 65984 41414 66036 41420
rect 65660 41372 65956 41392
rect 65716 41370 65740 41372
rect 65796 41370 65820 41372
rect 65876 41370 65900 41372
rect 65738 41318 65740 41370
rect 65802 41318 65814 41370
rect 65876 41318 65878 41370
rect 65716 41316 65740 41318
rect 65796 41316 65820 41318
rect 65876 41316 65900 41318
rect 65660 41296 65956 41316
rect 64696 41268 64748 41274
rect 64696 41210 64748 41216
rect 64708 40662 64736 41210
rect 64604 40656 64656 40662
rect 64604 40598 64656 40604
rect 64696 40656 64748 40662
rect 64696 40598 64748 40604
rect 64602 39536 64658 39545
rect 64602 39471 64604 39480
rect 64656 39471 64658 39480
rect 64604 39442 64656 39448
rect 64708 39302 64736 40598
rect 65660 40284 65956 40304
rect 65716 40282 65740 40284
rect 65796 40282 65820 40284
rect 65876 40282 65900 40284
rect 65738 40230 65740 40282
rect 65802 40230 65814 40282
rect 65876 40230 65878 40282
rect 65716 40228 65740 40230
rect 65796 40228 65820 40230
rect 65876 40228 65900 40230
rect 65660 40208 65956 40228
rect 64788 39840 64840 39846
rect 64788 39782 64840 39788
rect 64696 39296 64748 39302
rect 64696 39238 64748 39244
rect 63776 38956 63828 38962
rect 63776 38898 63828 38904
rect 64052 38956 64104 38962
rect 64052 38898 64104 38904
rect 64512 38956 64564 38962
rect 64512 38898 64564 38904
rect 62304 38888 62356 38894
rect 62304 38830 62356 38836
rect 63224 38888 63276 38894
rect 63224 38830 63276 38836
rect 63684 38888 63736 38894
rect 63684 38830 63736 38836
rect 62120 38820 62172 38826
rect 62120 38762 62172 38768
rect 60832 38752 60884 38758
rect 60832 38694 60884 38700
rect 59820 38412 59872 38418
rect 59820 38354 59872 38360
rect 59832 37262 59860 38354
rect 60280 38344 60332 38350
rect 60280 38286 60332 38292
rect 60292 37806 60320 38286
rect 61844 38276 61896 38282
rect 61844 38218 61896 38224
rect 61752 38004 61804 38010
rect 61752 37946 61804 37952
rect 60280 37800 60332 37806
rect 60280 37742 60332 37748
rect 59820 37256 59872 37262
rect 59820 37198 59872 37204
rect 56876 36110 56928 36116
rect 55956 36100 56008 36106
rect 55956 36042 56008 36048
rect 55680 35828 55732 35834
rect 55680 35770 55732 35776
rect 55692 35630 55720 35770
rect 55968 35630 55996 36042
rect 55680 35624 55732 35630
rect 55680 35566 55732 35572
rect 55956 35624 56008 35630
rect 55956 35566 56008 35572
rect 56600 35624 56652 35630
rect 56600 35566 56652 35572
rect 56140 35216 56192 35222
rect 56192 35176 56456 35204
rect 56140 35158 56192 35164
rect 56428 35086 56456 35176
rect 55956 35080 56008 35086
rect 55954 35048 55956 35057
rect 56048 35080 56100 35086
rect 56008 35048 56010 35057
rect 56048 35022 56100 35028
rect 56324 35080 56376 35086
rect 56324 35022 56376 35028
rect 56416 35080 56468 35086
rect 56416 35022 56468 35028
rect 55954 34983 56010 34992
rect 55588 34944 55640 34950
rect 55588 34886 55640 34892
rect 55312 34536 55364 34542
rect 55312 34478 55364 34484
rect 55600 34474 55628 34886
rect 56060 34626 56088 35022
rect 56336 34746 56364 35022
rect 56324 34740 56376 34746
rect 56324 34682 56376 34688
rect 56060 34598 56180 34626
rect 56152 34542 56180 34598
rect 56612 34542 56640 35566
rect 56782 34640 56838 34649
rect 56782 34575 56784 34584
rect 56836 34575 56838 34584
rect 56784 34546 56836 34552
rect 56140 34536 56192 34542
rect 56140 34478 56192 34484
rect 56600 34536 56652 34542
rect 56600 34478 56652 34484
rect 55588 34468 55640 34474
rect 55588 34410 55640 34416
rect 56612 32842 56640 34478
rect 56600 32836 56652 32842
rect 56600 32778 56652 32784
rect 55220 32564 55272 32570
rect 55220 32506 55272 32512
rect 55128 32496 55180 32502
rect 55128 32438 55180 32444
rect 48504 32020 48556 32026
rect 48504 31962 48556 31968
rect 43076 31816 43128 31822
rect 43076 31758 43128 31764
rect 41604 31272 41656 31278
rect 56600 31272 56652 31278
rect 41604 31214 41656 31220
rect 56598 31240 56600 31249
rect 56888 31249 56916 36110
rect 58728 36094 58848 36122
rect 58256 35828 58308 35834
rect 58256 35770 58308 35776
rect 57060 35216 57112 35222
rect 57060 35158 57112 35164
rect 57072 34785 57100 35158
rect 57428 34944 57480 34950
rect 57428 34886 57480 34892
rect 57058 34776 57114 34785
rect 57440 34746 57468 34886
rect 57058 34711 57114 34720
rect 57428 34740 57480 34746
rect 57428 34682 57480 34688
rect 56652 31240 56654 31249
rect 56598 31175 56654 31184
rect 56874 31240 56930 31249
rect 56874 31175 56930 31184
rect 56322 30832 56378 30841
rect 56322 30767 56378 30776
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32680 16584 32732 16590
rect 32680 16526 32732 16532
rect 32588 16176 32640 16182
rect 32588 16118 32640 16124
rect 32404 15632 32456 15638
rect 32404 15574 32456 15580
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 27908 9586 27936 9862
rect 27896 9580 27948 9586
rect 27896 9522 27948 9528
rect 27712 9376 27764 9382
rect 27712 9318 27764 9324
rect 27724 9178 27752 9318
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 29920 5568 29972 5574
rect 29920 5510 29972 5516
rect 29932 4865 29960 5510
rect 29918 4856 29974 4865
rect 29918 4791 29974 4800
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 28080 4140 28132 4146
rect 28080 4082 28132 4088
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4066 2136 4122 2145
rect 4220 2128 4516 2148
rect 4066 2071 4122 2080
rect 3790 1456 3846 1465
rect 3790 1391 3846 1400
rect 28092 800 28120 4082
rect 56336 3466 56364 30767
rect 57440 27169 57468 34682
rect 58268 34542 58296 35770
rect 58348 35556 58400 35562
rect 58348 35498 58400 35504
rect 58360 35222 58388 35498
rect 58348 35216 58400 35222
rect 58348 35158 58400 35164
rect 58728 35154 58756 36094
rect 60292 35766 60320 37742
rect 60556 37460 60608 37466
rect 60556 37402 60608 37408
rect 60568 36106 60596 37402
rect 61764 37330 61792 37946
rect 61856 37806 61884 38218
rect 61844 37800 61896 37806
rect 61844 37742 61896 37748
rect 61856 37466 61884 37742
rect 62120 37732 62172 37738
rect 62120 37674 62172 37680
rect 61844 37460 61896 37466
rect 61844 37402 61896 37408
rect 61752 37324 61804 37330
rect 61752 37266 61804 37272
rect 60660 36922 60780 36938
rect 60648 36916 60792 36922
rect 60700 36910 60740 36916
rect 60648 36858 60700 36864
rect 60740 36858 60792 36864
rect 61108 36712 61160 36718
rect 61108 36654 61160 36660
rect 61120 36378 61148 36654
rect 62132 36650 62160 37674
rect 63696 37330 63724 38830
rect 64064 37398 64092 38898
rect 64800 38894 64828 39782
rect 65524 39432 65576 39438
rect 65524 39374 65576 39380
rect 65536 38962 65564 39374
rect 65660 39196 65956 39216
rect 65716 39194 65740 39196
rect 65796 39194 65820 39196
rect 65876 39194 65900 39196
rect 65738 39142 65740 39194
rect 65802 39142 65814 39194
rect 65876 39142 65878 39194
rect 65716 39140 65740 39142
rect 65796 39140 65820 39142
rect 65876 39140 65900 39142
rect 65660 39120 65956 39140
rect 65524 38956 65576 38962
rect 65524 38898 65576 38904
rect 64788 38888 64840 38894
rect 64788 38830 64840 38836
rect 65996 38758 66024 41414
rect 66180 40118 66208 41958
rect 66720 40928 66772 40934
rect 66720 40870 66772 40876
rect 66732 40594 66760 40870
rect 66720 40588 66772 40594
rect 66720 40530 66772 40536
rect 66168 40112 66220 40118
rect 66168 40054 66220 40060
rect 66536 39568 66588 39574
rect 66536 39510 66588 39516
rect 66548 39409 66576 39510
rect 66732 39506 66760 40530
rect 66824 40458 66852 42570
rect 66916 42226 66944 43182
rect 66996 42560 67048 42566
rect 66996 42502 67048 42508
rect 66904 42220 66956 42226
rect 66904 42162 66956 42168
rect 67008 41682 67036 42502
rect 66996 41676 67048 41682
rect 66996 41618 67048 41624
rect 66812 40452 66864 40458
rect 66812 40394 66864 40400
rect 66824 40050 66852 40394
rect 67284 40050 67312 44134
rect 81020 44092 81316 44112
rect 81076 44090 81100 44092
rect 81156 44090 81180 44092
rect 81236 44090 81260 44092
rect 81098 44038 81100 44090
rect 81162 44038 81174 44090
rect 81236 44038 81238 44090
rect 81076 44036 81100 44038
rect 81156 44036 81180 44038
rect 81236 44036 81260 44038
rect 81020 44016 81316 44036
rect 69112 43852 69164 43858
rect 69112 43794 69164 43800
rect 70308 43852 70360 43858
rect 70308 43794 70360 43800
rect 68652 41676 68704 41682
rect 68652 41618 68704 41624
rect 68100 41608 68152 41614
rect 68100 41550 68152 41556
rect 68112 41274 68140 41550
rect 68664 41274 68692 41618
rect 69020 41472 69072 41478
rect 69020 41414 69072 41420
rect 69032 41274 69060 41414
rect 68100 41268 68152 41274
rect 68100 41210 68152 41216
rect 68652 41268 68704 41274
rect 68652 41210 68704 41216
rect 69020 41268 69072 41274
rect 69020 41210 69072 41216
rect 68112 41070 68140 41210
rect 68100 41064 68152 41070
rect 68100 41006 68152 41012
rect 68376 40928 68428 40934
rect 68376 40870 68428 40876
rect 69020 40928 69072 40934
rect 69020 40870 69072 40876
rect 68388 40050 68416 40870
rect 68468 40588 68520 40594
rect 68468 40530 68520 40536
rect 68480 40089 68508 40530
rect 68652 40384 68704 40390
rect 68652 40326 68704 40332
rect 68466 40080 68522 40089
rect 66812 40044 66864 40050
rect 66812 39986 66864 39992
rect 67272 40044 67324 40050
rect 67272 39986 67324 39992
rect 67732 40044 67784 40050
rect 67732 39986 67784 39992
rect 68376 40044 68428 40050
rect 68466 40015 68522 40024
rect 68376 39986 68428 39992
rect 67180 39840 67232 39846
rect 67180 39782 67232 39788
rect 66720 39500 66772 39506
rect 66720 39442 66772 39448
rect 66534 39400 66590 39409
rect 66534 39335 66536 39344
rect 66588 39335 66590 39344
rect 66536 39306 66588 39312
rect 65984 38752 66036 38758
rect 65984 38694 66036 38700
rect 65524 38548 65576 38554
rect 65524 38490 65576 38496
rect 64420 38344 64472 38350
rect 64420 38286 64472 38292
rect 65156 38344 65208 38350
rect 65156 38286 65208 38292
rect 64432 38010 64460 38286
rect 64512 38208 64564 38214
rect 64512 38150 64564 38156
rect 64880 38208 64932 38214
rect 64880 38150 64932 38156
rect 64420 38004 64472 38010
rect 64420 37946 64472 37952
rect 64524 37874 64552 38150
rect 64512 37868 64564 37874
rect 64512 37810 64564 37816
rect 64892 37738 64920 38150
rect 65168 38010 65196 38286
rect 65156 38004 65208 38010
rect 65156 37946 65208 37952
rect 65168 37806 65196 37946
rect 65156 37800 65208 37806
rect 65156 37742 65208 37748
rect 64880 37732 64932 37738
rect 64880 37674 64932 37680
rect 64788 37460 64840 37466
rect 64788 37402 64840 37408
rect 64052 37392 64104 37398
rect 64052 37334 64104 37340
rect 62580 37324 62632 37330
rect 62580 37266 62632 37272
rect 63592 37324 63644 37330
rect 63592 37266 63644 37272
rect 63684 37324 63736 37330
rect 63684 37266 63736 37272
rect 64328 37324 64380 37330
rect 64328 37266 64380 37272
rect 62120 36644 62172 36650
rect 62120 36586 62172 36592
rect 61108 36372 61160 36378
rect 61108 36314 61160 36320
rect 62212 36236 62264 36242
rect 62212 36178 62264 36184
rect 62120 36168 62172 36174
rect 62120 36110 62172 36116
rect 60556 36100 60608 36106
rect 60556 36042 60608 36048
rect 62132 35766 62160 36110
rect 62224 36038 62252 36178
rect 62212 36032 62264 36038
rect 62212 35974 62264 35980
rect 59544 35760 59596 35766
rect 59544 35702 59596 35708
rect 60280 35760 60332 35766
rect 60280 35702 60332 35708
rect 62120 35760 62172 35766
rect 62120 35702 62172 35708
rect 58808 35216 58860 35222
rect 58808 35158 58860 35164
rect 58716 35148 58768 35154
rect 58716 35090 58768 35096
rect 58440 35080 58492 35086
rect 58820 35034 58848 35158
rect 58492 35028 58848 35034
rect 58440 35022 58848 35028
rect 58452 35006 58848 35022
rect 58808 34944 58860 34950
rect 58808 34886 58860 34892
rect 58900 34944 58952 34950
rect 58900 34886 58952 34892
rect 59084 34944 59136 34950
rect 59084 34886 59136 34892
rect 58622 34640 58678 34649
rect 58622 34575 58624 34584
rect 58676 34575 58678 34584
rect 58624 34546 58676 34552
rect 58256 34536 58308 34542
rect 58256 34478 58308 34484
rect 58440 30184 58492 30190
rect 58438 30152 58440 30161
rect 58492 30152 58494 30161
rect 58438 30087 58494 30096
rect 58440 29844 58492 29850
rect 58440 29786 58492 29792
rect 58452 29481 58480 29786
rect 58438 29472 58494 29481
rect 58438 29407 58494 29416
rect 58440 28076 58492 28082
rect 58438 28044 58440 28053
rect 58492 28044 58494 28053
rect 58438 27979 58494 27988
rect 56414 27160 56470 27169
rect 56414 27095 56470 27104
rect 57426 27160 57482 27169
rect 57426 27095 57482 27104
rect 56428 4865 56456 27095
rect 58440 26852 58492 26858
rect 58438 26820 58440 26829
rect 58492 26820 58494 26829
rect 58438 26755 58494 26764
rect 58440 26648 58492 26654
rect 58440 26590 58492 26596
rect 58452 25605 58480 26590
rect 58438 25596 58494 25605
rect 58360 25554 58438 25582
rect 58070 24168 58126 24177
rect 58070 24103 58126 24112
rect 58084 23361 58112 24103
rect 58360 23497 58388 25554
rect 58438 25531 58494 25540
rect 58438 24168 58494 24177
rect 58820 24154 58848 34886
rect 58912 30190 58940 34886
rect 58992 34536 59044 34542
rect 58992 34478 59044 34484
rect 58900 30184 58952 30190
rect 58900 30126 58952 30132
rect 58494 24126 58848 24154
rect 58438 24103 58494 24112
rect 59004 23662 59032 34478
rect 59096 29850 59124 34886
rect 59452 34604 59504 34610
rect 59452 34546 59504 34552
rect 59176 34536 59228 34542
rect 59176 34478 59228 34484
rect 59360 34536 59412 34542
rect 59360 34478 59412 34484
rect 59084 29844 59136 29850
rect 59084 29786 59136 29792
rect 58440 23656 58492 23662
rect 58440 23598 58492 23604
rect 58992 23656 59044 23662
rect 58992 23598 59044 23604
rect 58346 23488 58402 23497
rect 58346 23423 58402 23432
rect 58070 23352 58126 23361
rect 58070 23287 58126 23296
rect 58452 22817 58480 23598
rect 58438 22808 58494 22817
rect 58438 22743 58494 22752
rect 59188 20330 59216 34478
rect 59372 31550 59400 34478
rect 59360 31544 59412 31550
rect 59360 31486 59412 31492
rect 59360 27668 59412 27674
rect 59360 27610 59412 27616
rect 59372 26858 59400 27610
rect 59360 26852 59412 26858
rect 59360 26794 59412 26800
rect 59464 26654 59492 34546
rect 59556 34406 59584 35702
rect 61292 35284 61344 35290
rect 61292 35226 61344 35232
rect 59636 35080 59688 35086
rect 59636 35022 59688 35028
rect 59648 34542 59676 35022
rect 61304 34950 61332 35226
rect 62132 35170 62160 35702
rect 62040 35154 62160 35170
rect 62028 35148 62160 35154
rect 62080 35142 62160 35148
rect 62028 35090 62080 35096
rect 62028 35012 62080 35018
rect 62028 34954 62080 34960
rect 59728 34944 59780 34950
rect 59728 34886 59780 34892
rect 61292 34944 61344 34950
rect 61292 34886 61344 34892
rect 61750 34912 61806 34921
rect 59636 34536 59688 34542
rect 59636 34478 59688 34484
rect 59544 34400 59596 34406
rect 59544 34342 59596 34348
rect 59636 34400 59688 34406
rect 59636 34342 59688 34348
rect 59648 28098 59676 34342
rect 59740 31618 59768 34886
rect 61750 34847 61806 34856
rect 61764 34542 61792 34847
rect 62040 34746 62068 34954
rect 62028 34740 62080 34746
rect 62028 34682 62080 34688
rect 61936 34672 61988 34678
rect 61936 34614 61988 34620
rect 61752 34536 61804 34542
rect 61752 34478 61804 34484
rect 61948 33658 61976 34614
rect 61936 33652 61988 33658
rect 61936 33594 61988 33600
rect 62224 33590 62252 35974
rect 62304 35080 62356 35086
rect 62304 35022 62356 35028
rect 62316 34649 62344 35022
rect 62592 34678 62620 37266
rect 63604 36718 63632 37266
rect 63696 36802 63724 37266
rect 63696 36774 63816 36802
rect 63788 36718 63816 36774
rect 63592 36712 63644 36718
rect 63592 36654 63644 36660
rect 63776 36712 63828 36718
rect 63776 36654 63828 36660
rect 62948 35760 63000 35766
rect 62948 35702 63000 35708
rect 63776 35760 63828 35766
rect 63776 35702 63828 35708
rect 62960 35630 62988 35702
rect 62948 35624 63000 35630
rect 62948 35566 63000 35572
rect 62580 34672 62632 34678
rect 62302 34640 62358 34649
rect 62580 34614 62632 34620
rect 62302 34575 62358 34584
rect 62960 34542 62988 35566
rect 63788 35494 63816 35702
rect 63776 35488 63828 35494
rect 63776 35430 63828 35436
rect 63040 35216 63092 35222
rect 63040 35158 63092 35164
rect 63052 35057 63080 35158
rect 63038 35048 63094 35057
rect 63038 34983 63094 34992
rect 64340 34678 64368 37266
rect 64512 36712 64564 36718
rect 64512 36654 64564 36660
rect 64524 36038 64552 36654
rect 64604 36576 64656 36582
rect 64604 36518 64656 36524
rect 64512 36032 64564 36038
rect 64512 35974 64564 35980
rect 64524 35154 64552 35974
rect 64512 35148 64564 35154
rect 64512 35090 64564 35096
rect 64616 34950 64644 36518
rect 64800 36310 64828 37402
rect 65432 36712 65484 36718
rect 65432 36654 65484 36660
rect 64788 36304 64840 36310
rect 64788 36246 64840 36252
rect 65444 35494 65472 36654
rect 65536 36174 65564 38490
rect 65660 38108 65956 38128
rect 65716 38106 65740 38108
rect 65796 38106 65820 38108
rect 65876 38106 65900 38108
rect 65738 38054 65740 38106
rect 65802 38054 65814 38106
rect 65876 38054 65878 38106
rect 65716 38052 65740 38054
rect 65796 38052 65820 38054
rect 65876 38052 65900 38054
rect 65660 38032 65956 38052
rect 67192 37466 67220 39782
rect 67284 38758 67312 39986
rect 67640 39500 67692 39506
rect 67640 39442 67692 39448
rect 67652 39098 67680 39442
rect 67744 39302 67772 39986
rect 68480 39982 68508 40015
rect 68468 39976 68520 39982
rect 68468 39918 68520 39924
rect 68560 39908 68612 39914
rect 68560 39850 68612 39856
rect 67732 39296 67784 39302
rect 67732 39238 67784 39244
rect 67640 39092 67692 39098
rect 67640 39034 67692 39040
rect 67272 38752 67324 38758
rect 67272 38694 67324 38700
rect 67640 38480 67692 38486
rect 67640 38422 67692 38428
rect 67652 38214 67680 38422
rect 67640 38208 67692 38214
rect 67640 38150 67692 38156
rect 67456 37664 67508 37670
rect 67456 37606 67508 37612
rect 67180 37460 67232 37466
rect 67180 37402 67232 37408
rect 67468 37330 67496 37606
rect 66260 37324 66312 37330
rect 66260 37266 66312 37272
rect 66444 37324 66496 37330
rect 66444 37266 66496 37272
rect 66628 37324 66680 37330
rect 66628 37266 66680 37272
rect 67456 37324 67508 37330
rect 67456 37266 67508 37272
rect 66168 37256 66220 37262
rect 66168 37198 66220 37204
rect 66180 37126 66208 37198
rect 65984 37120 66036 37126
rect 65984 37062 66036 37068
rect 66168 37120 66220 37126
rect 66168 37062 66220 37068
rect 65660 37020 65956 37040
rect 65716 37018 65740 37020
rect 65796 37018 65820 37020
rect 65876 37018 65900 37020
rect 65738 36966 65740 37018
rect 65802 36966 65814 37018
rect 65876 36966 65878 37018
rect 65716 36964 65740 36966
rect 65796 36964 65820 36966
rect 65876 36964 65900 36966
rect 65660 36944 65956 36964
rect 65996 36242 66024 37062
rect 66168 36712 66220 36718
rect 66168 36654 66220 36660
rect 65984 36236 66036 36242
rect 65984 36178 66036 36184
rect 65524 36168 65576 36174
rect 65524 36110 65576 36116
rect 65660 35932 65956 35952
rect 65716 35930 65740 35932
rect 65796 35930 65820 35932
rect 65876 35930 65900 35932
rect 65738 35878 65740 35930
rect 65802 35878 65814 35930
rect 65876 35878 65878 35930
rect 65716 35876 65740 35878
rect 65796 35876 65820 35878
rect 65876 35876 65900 35878
rect 65660 35856 65956 35876
rect 66180 35630 66208 36654
rect 66168 35624 66220 35630
rect 66168 35566 66220 35572
rect 65432 35488 65484 35494
rect 65432 35430 65484 35436
rect 66272 34950 66300 37266
rect 66456 36718 66484 37266
rect 66640 36786 66668 37266
rect 66720 37256 66772 37262
rect 66720 37198 66772 37204
rect 66628 36780 66680 36786
rect 66628 36722 66680 36728
rect 66444 36712 66496 36718
rect 66444 36654 66496 36660
rect 66732 35154 66760 37198
rect 67744 37126 67772 39238
rect 68572 39001 68600 39850
rect 68558 38992 68614 39001
rect 68558 38927 68614 38936
rect 68572 38894 68600 38927
rect 68560 38888 68612 38894
rect 68466 38856 68522 38865
rect 68560 38830 68612 38836
rect 68466 38791 68522 38800
rect 68480 38758 68508 38791
rect 68468 38752 68520 38758
rect 68468 38694 68520 38700
rect 68664 38554 68692 40326
rect 69032 39930 69060 40870
rect 69124 40186 69152 43794
rect 69756 43648 69808 43654
rect 69756 43590 69808 43596
rect 69388 43240 69440 43246
rect 69388 43182 69440 43188
rect 69204 42764 69256 42770
rect 69204 42706 69256 42712
rect 69296 42764 69348 42770
rect 69296 42706 69348 42712
rect 69216 42226 69244 42706
rect 69308 42362 69336 42706
rect 69400 42566 69428 43182
rect 69664 43104 69716 43110
rect 69664 43046 69716 43052
rect 69676 42634 69704 43046
rect 69664 42628 69716 42634
rect 69664 42570 69716 42576
rect 69388 42560 69440 42566
rect 69388 42502 69440 42508
rect 69296 42356 69348 42362
rect 69296 42298 69348 42304
rect 69676 42226 69704 42570
rect 69204 42220 69256 42226
rect 69204 42162 69256 42168
rect 69664 42220 69716 42226
rect 69664 42162 69716 42168
rect 69216 41682 69244 42162
rect 69768 42158 69796 43590
rect 70320 43450 70348 43794
rect 96380 43548 96676 43568
rect 96436 43546 96460 43548
rect 96516 43546 96540 43548
rect 96596 43546 96620 43548
rect 96458 43494 96460 43546
rect 96522 43494 96534 43546
rect 96596 43494 96598 43546
rect 96436 43492 96460 43494
rect 96516 43492 96540 43494
rect 96596 43492 96620 43494
rect 96380 43472 96676 43492
rect 70308 43444 70360 43450
rect 70308 43386 70360 43392
rect 81020 43004 81316 43024
rect 81076 43002 81100 43004
rect 81156 43002 81180 43004
rect 81236 43002 81260 43004
rect 81098 42950 81100 43002
rect 81162 42950 81174 43002
rect 81236 42950 81238 43002
rect 81076 42948 81100 42950
rect 81156 42948 81180 42950
rect 81236 42948 81260 42950
rect 81020 42928 81316 42948
rect 71412 42764 71464 42770
rect 71412 42706 71464 42712
rect 70400 42696 70452 42702
rect 70400 42638 70452 42644
rect 70032 42560 70084 42566
rect 70032 42502 70084 42508
rect 69756 42152 69808 42158
rect 69756 42094 69808 42100
rect 69768 41750 69796 42094
rect 69756 41744 69808 41750
rect 69756 41686 69808 41692
rect 70044 41682 70072 42502
rect 70308 42084 70360 42090
rect 70308 42026 70360 42032
rect 69204 41676 69256 41682
rect 69204 41618 69256 41624
rect 69848 41676 69900 41682
rect 69848 41618 69900 41624
rect 70032 41676 70084 41682
rect 70032 41618 70084 41624
rect 69388 41132 69440 41138
rect 69388 41074 69440 41080
rect 69400 40594 69428 41074
rect 69860 40594 69888 41618
rect 70044 41478 70072 41618
rect 70320 41614 70348 42026
rect 70308 41608 70360 41614
rect 70308 41550 70360 41556
rect 70032 41472 70084 41478
rect 70032 41414 70084 41420
rect 70320 41002 70348 41550
rect 70412 41138 70440 42638
rect 71136 42152 71188 42158
rect 71136 42094 71188 42100
rect 71148 41138 71176 42094
rect 71424 42022 71452 42706
rect 96380 42460 96676 42480
rect 96436 42458 96460 42460
rect 96516 42458 96540 42460
rect 96596 42458 96620 42460
rect 96458 42406 96460 42458
rect 96522 42406 96534 42458
rect 96596 42406 96598 42458
rect 96436 42404 96460 42406
rect 96516 42404 96540 42406
rect 96596 42404 96620 42406
rect 96380 42384 96676 42404
rect 72516 42220 72568 42226
rect 72516 42162 72568 42168
rect 71412 42016 71464 42022
rect 71412 41958 71464 41964
rect 71424 41682 71452 41958
rect 71412 41676 71464 41682
rect 71412 41618 71464 41624
rect 72528 41478 72556 42162
rect 81020 41916 81316 41936
rect 81076 41914 81100 41916
rect 81156 41914 81180 41916
rect 81236 41914 81260 41916
rect 81098 41862 81100 41914
rect 81162 41862 81174 41914
rect 81236 41862 81238 41914
rect 81076 41860 81100 41862
rect 81156 41860 81180 41862
rect 81236 41860 81260 41862
rect 81020 41840 81316 41860
rect 78220 41608 78272 41614
rect 78220 41550 78272 41556
rect 71596 41472 71648 41478
rect 71596 41414 71648 41420
rect 72516 41472 72568 41478
rect 72516 41414 72568 41420
rect 77944 41472 77996 41478
rect 77944 41414 77996 41420
rect 70400 41132 70452 41138
rect 70400 41074 70452 41080
rect 71136 41132 71188 41138
rect 71136 41074 71188 41080
rect 70492 41064 70544 41070
rect 70492 41006 70544 41012
rect 70308 40996 70360 41002
rect 70308 40938 70360 40944
rect 70124 40656 70176 40662
rect 70124 40598 70176 40604
rect 69388 40588 69440 40594
rect 69388 40530 69440 40536
rect 69848 40588 69900 40594
rect 69848 40530 69900 40536
rect 69400 40390 69428 40530
rect 69860 40390 69888 40530
rect 69388 40384 69440 40390
rect 69388 40326 69440 40332
rect 69848 40384 69900 40390
rect 69848 40326 69900 40332
rect 70032 40384 70084 40390
rect 70032 40326 70084 40332
rect 69112 40180 69164 40186
rect 69112 40122 69164 40128
rect 69400 40050 69428 40326
rect 69388 40044 69440 40050
rect 69388 39986 69440 39992
rect 69940 40044 69992 40050
rect 69940 39986 69992 39992
rect 68940 39902 69060 39930
rect 69388 39908 69440 39914
rect 68744 39024 68796 39030
rect 68940 39012 68968 39902
rect 69388 39850 69440 39856
rect 69400 39506 69428 39850
rect 69664 39840 69716 39846
rect 69664 39782 69716 39788
rect 69676 39642 69704 39782
rect 69664 39636 69716 39642
rect 69664 39578 69716 39584
rect 69020 39500 69072 39506
rect 69020 39442 69072 39448
rect 69388 39500 69440 39506
rect 69388 39442 69440 39448
rect 68796 38984 68968 39012
rect 68744 38966 68796 38972
rect 68744 38752 68796 38758
rect 68742 38720 68744 38729
rect 68796 38720 68798 38729
rect 68742 38655 68798 38664
rect 68652 38548 68704 38554
rect 68652 38490 68704 38496
rect 68928 38208 68980 38214
rect 68928 38150 68980 38156
rect 67732 37120 67784 37126
rect 67732 37062 67784 37068
rect 68652 37120 68704 37126
rect 68652 37062 68704 37068
rect 68664 36718 68692 37062
rect 68652 36712 68704 36718
rect 68652 36654 68704 36660
rect 68664 36378 68692 36654
rect 68652 36372 68704 36378
rect 68652 36314 68704 36320
rect 68940 35766 68968 38150
rect 69032 38010 69060 39442
rect 69952 39370 69980 39986
rect 70044 39982 70072 40326
rect 70136 40186 70164 40598
rect 70400 40520 70452 40526
rect 70400 40462 70452 40468
rect 70124 40180 70176 40186
rect 70124 40122 70176 40128
rect 70308 40180 70360 40186
rect 70308 40122 70360 40128
rect 70320 40050 70348 40122
rect 70308 40044 70360 40050
rect 70308 39986 70360 39992
rect 70412 39982 70440 40462
rect 70504 40186 70532 41006
rect 71608 40934 71636 41414
rect 71688 41200 71740 41206
rect 71688 41142 71740 41148
rect 71596 40928 71648 40934
rect 71596 40870 71648 40876
rect 70492 40180 70544 40186
rect 70492 40122 70544 40128
rect 71410 40080 71466 40089
rect 71410 40015 71466 40024
rect 71424 39982 71452 40015
rect 70032 39976 70084 39982
rect 70032 39918 70084 39924
rect 70400 39976 70452 39982
rect 70400 39918 70452 39924
rect 71412 39976 71464 39982
rect 71412 39918 71464 39924
rect 70952 39840 71004 39846
rect 70952 39782 71004 39788
rect 70964 39370 70992 39782
rect 69940 39364 69992 39370
rect 69940 39306 69992 39312
rect 70952 39364 71004 39370
rect 70952 39306 71004 39312
rect 70964 39098 70992 39306
rect 69112 39092 69164 39098
rect 69112 39034 69164 39040
rect 70952 39092 71004 39098
rect 70952 39034 71004 39040
rect 69124 39001 69152 39034
rect 69110 38992 69166 39001
rect 69110 38927 69166 38936
rect 71424 38894 71452 39918
rect 71700 39846 71728 41142
rect 71964 40996 72016 41002
rect 71964 40938 72016 40944
rect 71976 40390 72004 40938
rect 72528 40730 72556 41414
rect 77852 41064 77904 41070
rect 77852 41006 77904 41012
rect 74264 40928 74316 40934
rect 74264 40870 74316 40876
rect 76840 40928 76892 40934
rect 76840 40870 76892 40876
rect 77576 40928 77628 40934
rect 77576 40870 77628 40876
rect 72516 40724 72568 40730
rect 72516 40666 72568 40672
rect 71964 40384 72016 40390
rect 71964 40326 72016 40332
rect 73988 40384 74040 40390
rect 73988 40326 74040 40332
rect 71872 39976 71924 39982
rect 71872 39918 71924 39924
rect 72606 39944 72662 39953
rect 71688 39840 71740 39846
rect 71688 39782 71740 39788
rect 71412 38888 71464 38894
rect 69478 38856 69534 38865
rect 71412 38830 71464 38836
rect 69478 38791 69480 38800
rect 69532 38791 69534 38800
rect 69480 38762 69532 38768
rect 69756 38752 69808 38758
rect 69756 38694 69808 38700
rect 70308 38752 70360 38758
rect 70308 38694 70360 38700
rect 69020 38004 69072 38010
rect 69020 37946 69072 37952
rect 69032 37806 69060 37946
rect 69020 37800 69072 37806
rect 69020 37742 69072 37748
rect 69572 37800 69624 37806
rect 69572 37742 69624 37748
rect 69032 36038 69060 37742
rect 69584 37398 69612 37742
rect 69572 37392 69624 37398
rect 69572 37334 69624 37340
rect 69112 37324 69164 37330
rect 69112 37266 69164 37272
rect 69020 36032 69072 36038
rect 69020 35974 69072 35980
rect 68928 35760 68980 35766
rect 68928 35702 68980 35708
rect 68940 35630 68968 35702
rect 68928 35624 68980 35630
rect 68928 35566 68980 35572
rect 69020 35624 69072 35630
rect 69020 35566 69072 35572
rect 66720 35148 66772 35154
rect 66720 35090 66772 35096
rect 64604 34944 64656 34950
rect 64696 34944 64748 34950
rect 64604 34886 64656 34892
rect 64694 34912 64696 34921
rect 66260 34944 66312 34950
rect 64748 34912 64750 34921
rect 64328 34672 64380 34678
rect 64328 34614 64380 34620
rect 64340 34542 64368 34614
rect 62948 34536 63000 34542
rect 62948 34478 63000 34484
rect 64328 34536 64380 34542
rect 64328 34478 64380 34484
rect 62672 34468 62724 34474
rect 62672 34410 62724 34416
rect 62684 34202 62712 34410
rect 62672 34196 62724 34202
rect 62672 34138 62724 34144
rect 62212 33584 62264 33590
rect 62212 33526 62264 33532
rect 64616 33522 64644 34886
rect 66260 34886 66312 34892
rect 64694 34847 64750 34856
rect 65660 34844 65956 34864
rect 65716 34842 65740 34844
rect 65796 34842 65820 34844
rect 65876 34842 65900 34844
rect 65738 34790 65740 34842
rect 65802 34790 65814 34842
rect 65876 34790 65878 34842
rect 65716 34788 65740 34790
rect 65796 34788 65820 34790
rect 65876 34788 65900 34790
rect 65660 34768 65956 34788
rect 64604 33516 64656 33522
rect 64604 33458 64656 33464
rect 69032 32434 69060 35566
rect 69124 35018 69152 37266
rect 69768 36718 69796 38694
rect 70320 38434 70348 38694
rect 70320 38418 70440 38434
rect 71884 38418 71912 39918
rect 72606 39879 72662 39888
rect 72620 39098 72648 39879
rect 74000 39098 74028 40326
rect 74276 40118 74304 40870
rect 75828 40588 75880 40594
rect 75828 40530 75880 40536
rect 74448 40520 74500 40526
rect 74448 40462 74500 40468
rect 74264 40112 74316 40118
rect 74264 40054 74316 40060
rect 74460 40032 74488 40462
rect 75840 40390 75868 40530
rect 75828 40384 75880 40390
rect 75828 40326 75880 40332
rect 74540 40044 74592 40050
rect 74460 40004 74540 40032
rect 74540 39986 74592 39992
rect 75840 39982 75868 40326
rect 75184 39976 75236 39982
rect 75184 39918 75236 39924
rect 75828 39976 75880 39982
rect 75828 39918 75880 39924
rect 75196 39098 75224 39918
rect 76196 39908 76248 39914
rect 76196 39850 76248 39856
rect 75828 39840 75880 39846
rect 75828 39782 75880 39788
rect 75840 39506 75868 39782
rect 76208 39642 76236 39850
rect 76656 39840 76708 39846
rect 76656 39782 76708 39788
rect 76196 39636 76248 39642
rect 76196 39578 76248 39584
rect 76472 39568 76524 39574
rect 76472 39510 76524 39516
rect 75828 39500 75880 39506
rect 75828 39442 75880 39448
rect 76484 39370 76512 39510
rect 76472 39364 76524 39370
rect 76472 39306 76524 39312
rect 76380 39296 76432 39302
rect 76380 39238 76432 39244
rect 72608 39092 72660 39098
rect 72608 39034 72660 39040
rect 73988 39092 74040 39098
rect 73988 39034 74040 39040
rect 75184 39092 75236 39098
rect 75184 39034 75236 39040
rect 72620 38894 72648 39034
rect 75734 38992 75790 39001
rect 75734 38927 75736 38936
rect 75788 38927 75790 38936
rect 75736 38898 75788 38904
rect 76392 38894 76420 39238
rect 72608 38888 72660 38894
rect 72608 38830 72660 38836
rect 76380 38888 76432 38894
rect 76380 38830 76432 38836
rect 76104 38820 76156 38826
rect 76104 38762 76156 38768
rect 70124 38412 70176 38418
rect 70320 38412 70452 38418
rect 70320 38406 70400 38412
rect 70124 38354 70176 38360
rect 70400 38354 70452 38360
rect 71872 38412 71924 38418
rect 71872 38354 71924 38360
rect 75736 38412 75788 38418
rect 75736 38354 75788 38360
rect 70032 38276 70084 38282
rect 70032 38218 70084 38224
rect 70044 37330 70072 38218
rect 70136 37330 70164 38354
rect 70308 38344 70360 38350
rect 70308 38286 70360 38292
rect 70320 38010 70348 38286
rect 70308 38004 70360 38010
rect 70308 37946 70360 37952
rect 70320 37330 70348 37946
rect 71688 37732 71740 37738
rect 71688 37674 71740 37680
rect 70676 37664 70728 37670
rect 70676 37606 70728 37612
rect 71136 37664 71188 37670
rect 71136 37606 71188 37612
rect 70032 37324 70084 37330
rect 70032 37266 70084 37272
rect 70124 37324 70176 37330
rect 70124 37266 70176 37272
rect 70308 37324 70360 37330
rect 70308 37266 70360 37272
rect 69940 37188 69992 37194
rect 69940 37130 69992 37136
rect 69952 36718 69980 37130
rect 69756 36712 69808 36718
rect 69756 36654 69808 36660
rect 69940 36712 69992 36718
rect 69940 36654 69992 36660
rect 70136 36582 70164 37266
rect 70320 36650 70348 37266
rect 70688 37126 70716 37606
rect 71148 37398 71176 37606
rect 71136 37392 71188 37398
rect 71136 37334 71188 37340
rect 70676 37120 70728 37126
rect 70676 37062 70728 37068
rect 71148 36922 71176 37334
rect 71700 37330 71728 37674
rect 71688 37324 71740 37330
rect 71688 37266 71740 37272
rect 71884 37312 71912 38354
rect 75644 38276 75696 38282
rect 75644 38218 75696 38224
rect 75656 37806 75684 38218
rect 75748 37874 75776 38354
rect 76116 38350 76144 38762
rect 76300 38758 76328 38789
rect 76288 38752 76340 38758
rect 76286 38720 76288 38729
rect 76340 38720 76342 38729
rect 76286 38655 76342 38664
rect 76104 38344 76156 38350
rect 76104 38286 76156 38292
rect 76116 38010 76144 38286
rect 76300 38214 76328 38655
rect 76392 38282 76420 38830
rect 76668 38758 76696 39782
rect 76656 38752 76708 38758
rect 76656 38694 76708 38700
rect 76380 38276 76432 38282
rect 76380 38218 76432 38224
rect 76288 38208 76340 38214
rect 76288 38150 76340 38156
rect 76104 38004 76156 38010
rect 76104 37946 76156 37952
rect 75736 37868 75788 37874
rect 75736 37810 75788 37816
rect 75644 37800 75696 37806
rect 75644 37742 75696 37748
rect 72056 37324 72108 37330
rect 71884 37284 72056 37312
rect 70952 36916 71004 36922
rect 70952 36858 71004 36864
rect 71136 36916 71188 36922
rect 71136 36858 71188 36864
rect 70964 36825 70992 36858
rect 70950 36816 71006 36825
rect 71148 36786 71176 36858
rect 71504 36848 71556 36854
rect 71504 36790 71556 36796
rect 70950 36751 71006 36760
rect 71136 36780 71188 36786
rect 71136 36722 71188 36728
rect 70308 36644 70360 36650
rect 70308 36586 70360 36592
rect 70584 36644 70636 36650
rect 70584 36586 70636 36592
rect 70124 36576 70176 36582
rect 70124 36518 70176 36524
rect 69572 36236 69624 36242
rect 69572 36178 69624 36184
rect 69584 35562 69612 36178
rect 70124 36032 70176 36038
rect 70124 35974 70176 35980
rect 70136 35766 70164 35974
rect 70124 35760 70176 35766
rect 69952 35720 70124 35748
rect 69572 35556 69624 35562
rect 69572 35498 69624 35504
rect 69848 35488 69900 35494
rect 69848 35430 69900 35436
rect 69294 35184 69350 35193
rect 69860 35154 69888 35430
rect 69294 35119 69296 35128
rect 69348 35119 69350 35128
rect 69848 35148 69900 35154
rect 69296 35090 69348 35096
rect 69848 35090 69900 35096
rect 69112 35012 69164 35018
rect 69112 34954 69164 34960
rect 69308 33386 69336 35090
rect 69952 34678 69980 35720
rect 70176 35720 70256 35748
rect 70124 35702 70176 35708
rect 70228 35630 70256 35720
rect 70596 35630 70624 36586
rect 71516 36310 71544 36790
rect 71596 36780 71648 36786
rect 71596 36722 71648 36728
rect 71504 36304 71556 36310
rect 71504 36246 71556 36252
rect 71608 36174 71636 36722
rect 71700 36242 71728 37266
rect 71688 36236 71740 36242
rect 71688 36178 71740 36184
rect 71596 36168 71648 36174
rect 71596 36110 71648 36116
rect 71320 35760 71372 35766
rect 71320 35702 71372 35708
rect 70124 35624 70176 35630
rect 70124 35566 70176 35572
rect 70216 35624 70268 35630
rect 70216 35566 70268 35572
rect 70584 35624 70636 35630
rect 70584 35566 70636 35572
rect 70676 35624 70728 35630
rect 70676 35566 70728 35572
rect 70032 35148 70084 35154
rect 70032 35090 70084 35096
rect 69940 34672 69992 34678
rect 69940 34614 69992 34620
rect 69952 34542 69980 34614
rect 69940 34536 69992 34542
rect 69940 34478 69992 34484
rect 70044 34066 70072 35090
rect 70136 34542 70164 35566
rect 70688 35306 70716 35566
rect 70860 35488 70912 35494
rect 70860 35430 70912 35436
rect 70596 35290 70716 35306
rect 70872 35290 70900 35430
rect 70584 35284 70716 35290
rect 70636 35278 70716 35284
rect 70860 35284 70912 35290
rect 70584 35226 70636 35232
rect 70860 35226 70912 35232
rect 71332 35193 71360 35702
rect 71318 35184 71374 35193
rect 71700 35154 71728 36178
rect 71318 35119 71374 35128
rect 71412 35148 71464 35154
rect 71412 35090 71464 35096
rect 71688 35148 71740 35154
rect 71688 35090 71740 35096
rect 71424 34746 71452 35090
rect 71596 35080 71648 35086
rect 71596 35022 71648 35028
rect 71608 34950 71636 35022
rect 71884 34950 71912 37284
rect 72056 37266 72108 37272
rect 75184 37256 75236 37262
rect 75184 37198 75236 37204
rect 75196 36854 75224 37198
rect 75184 36848 75236 36854
rect 71962 36816 72018 36825
rect 75184 36790 75236 36796
rect 71962 36751 71964 36760
rect 72016 36751 72018 36760
rect 71964 36722 72016 36728
rect 76852 36718 76880 40870
rect 77588 40594 77616 40870
rect 77864 40594 77892 41006
rect 77956 40730 77984 41414
rect 78128 41132 78180 41138
rect 78128 41074 78180 41080
rect 77944 40724 77996 40730
rect 77944 40666 77996 40672
rect 78140 40594 78168 41074
rect 78232 40662 78260 41550
rect 79784 41472 79836 41478
rect 79784 41414 79836 41420
rect 79796 41070 79824 41414
rect 96380 41372 96676 41392
rect 96436 41370 96460 41372
rect 96516 41370 96540 41372
rect 96596 41370 96620 41372
rect 96458 41318 96460 41370
rect 96522 41318 96534 41370
rect 96596 41318 96598 41370
rect 96436 41316 96460 41318
rect 96516 41316 96540 41318
rect 96596 41316 96620 41318
rect 96380 41296 96676 41316
rect 79784 41064 79836 41070
rect 79784 41006 79836 41012
rect 79876 40928 79928 40934
rect 79876 40870 79928 40876
rect 78220 40656 78272 40662
rect 78220 40598 78272 40604
rect 77576 40588 77628 40594
rect 77576 40530 77628 40536
rect 77668 40588 77720 40594
rect 77668 40530 77720 40536
rect 77852 40588 77904 40594
rect 77852 40530 77904 40536
rect 78128 40588 78180 40594
rect 78128 40530 78180 40536
rect 77680 40050 77708 40530
rect 78036 40384 78088 40390
rect 78036 40326 78088 40332
rect 78048 40118 78076 40326
rect 78140 40186 78168 40530
rect 78128 40180 78180 40186
rect 78128 40122 78180 40128
rect 78036 40112 78088 40118
rect 78036 40054 78088 40060
rect 77668 40044 77720 40050
rect 77668 39986 77720 39992
rect 77392 39908 77444 39914
rect 77392 39850 77444 39856
rect 77024 39840 77076 39846
rect 77024 39782 77076 39788
rect 77036 38826 77064 39782
rect 77300 39296 77352 39302
rect 77300 39238 77352 39244
rect 77024 38820 77076 38826
rect 77024 38762 77076 38768
rect 77036 38486 77064 38762
rect 76932 38480 76984 38486
rect 76932 38422 76984 38428
rect 77024 38480 77076 38486
rect 77024 38422 77076 38428
rect 77208 38480 77260 38486
rect 77208 38422 77260 38428
rect 76944 38332 76972 38422
rect 77220 38332 77248 38422
rect 77312 38418 77340 39238
rect 77404 38486 77432 39850
rect 77574 38992 77630 39001
rect 77574 38927 77576 38936
rect 77628 38927 77630 38936
rect 77576 38898 77628 38904
rect 77576 38752 77628 38758
rect 77574 38720 77576 38729
rect 77628 38720 77630 38729
rect 77574 38655 77630 38664
rect 77392 38480 77444 38486
rect 77392 38422 77444 38428
rect 77300 38412 77352 38418
rect 77300 38354 77352 38360
rect 77680 38350 77708 39986
rect 79888 39982 79916 40870
rect 81020 40828 81316 40848
rect 81076 40826 81100 40828
rect 81156 40826 81180 40828
rect 81236 40826 81260 40828
rect 81098 40774 81100 40826
rect 81162 40774 81174 40826
rect 81236 40774 81238 40826
rect 81076 40772 81100 40774
rect 81156 40772 81180 40774
rect 81236 40772 81260 40774
rect 81020 40752 81316 40772
rect 80796 40520 80848 40526
rect 80796 40462 80848 40468
rect 83648 40520 83700 40526
rect 83648 40462 83700 40468
rect 80244 40384 80296 40390
rect 80244 40326 80296 40332
rect 80256 39982 80284 40326
rect 79876 39976 79928 39982
rect 79876 39918 79928 39924
rect 80244 39976 80296 39982
rect 80244 39918 80296 39924
rect 79600 39840 79652 39846
rect 79600 39782 79652 39788
rect 78036 39500 78088 39506
rect 78036 39442 78088 39448
rect 79140 39500 79192 39506
rect 79140 39442 79192 39448
rect 79416 39500 79468 39506
rect 79416 39442 79468 39448
rect 78048 39409 78076 39442
rect 78034 39400 78090 39409
rect 78034 39335 78090 39344
rect 78954 39264 79010 39273
rect 78954 39199 79010 39208
rect 78968 39098 78996 39199
rect 79152 39137 79180 39442
rect 79138 39128 79194 39137
rect 78956 39092 79008 39098
rect 79138 39063 79194 39072
rect 78956 39034 79008 39040
rect 77760 38888 77812 38894
rect 79428 38865 79456 39442
rect 79612 39001 79640 39782
rect 79784 39024 79836 39030
rect 79598 38992 79654 39001
rect 79598 38927 79600 38936
rect 79652 38927 79654 38936
rect 79782 38992 79784 39001
rect 79836 38992 79838 39001
rect 79782 38927 79838 38936
rect 79600 38898 79652 38904
rect 77760 38830 77812 38836
rect 79414 38856 79470 38865
rect 77772 38554 77800 38830
rect 79888 38842 79916 39918
rect 80808 39642 80836 40462
rect 83660 40186 83688 40462
rect 84752 40384 84804 40390
rect 84752 40326 84804 40332
rect 83648 40180 83700 40186
rect 83648 40122 83700 40128
rect 84764 40118 84792 40326
rect 96380 40284 96676 40304
rect 96436 40282 96460 40284
rect 96516 40282 96540 40284
rect 96596 40282 96620 40284
rect 96458 40230 96460 40282
rect 96522 40230 96534 40282
rect 96596 40230 96598 40282
rect 96436 40228 96460 40230
rect 96516 40228 96540 40230
rect 96596 40228 96620 40230
rect 96380 40208 96676 40228
rect 84752 40112 84804 40118
rect 84752 40054 84804 40060
rect 83740 39976 83792 39982
rect 83740 39918 83792 39924
rect 85212 39976 85264 39982
rect 85212 39918 85264 39924
rect 81020 39740 81316 39760
rect 81076 39738 81100 39740
rect 81156 39738 81180 39740
rect 81236 39738 81260 39740
rect 81098 39686 81100 39738
rect 81162 39686 81174 39738
rect 81236 39686 81238 39738
rect 81076 39684 81100 39686
rect 81156 39684 81180 39686
rect 81236 39684 81260 39686
rect 81020 39664 81316 39684
rect 80796 39636 80848 39642
rect 80796 39578 80848 39584
rect 83752 39574 83780 39918
rect 83464 39568 83516 39574
rect 83464 39510 83516 39516
rect 83740 39568 83792 39574
rect 83740 39510 83792 39516
rect 80704 39500 80756 39506
rect 80704 39442 80756 39448
rect 80716 39273 80744 39442
rect 82912 39296 82964 39302
rect 80702 39264 80758 39273
rect 82912 39238 82964 39244
rect 80702 39199 80758 39208
rect 80426 39128 80482 39137
rect 80426 39063 80482 39072
rect 82728 39092 82780 39098
rect 80244 39024 80296 39030
rect 79796 38826 79916 38842
rect 79414 38791 79470 38800
rect 79784 38820 79916 38826
rect 79836 38814 79916 38820
rect 80164 38972 80244 38978
rect 80164 38966 80296 38972
rect 80164 38950 80284 38966
rect 80336 38956 80388 38962
rect 79784 38762 79836 38768
rect 78220 38752 78272 38758
rect 78218 38720 78220 38729
rect 78272 38720 78274 38729
rect 78218 38655 78274 38664
rect 77760 38548 77812 38554
rect 77760 38490 77812 38496
rect 78404 38412 78456 38418
rect 78404 38354 78456 38360
rect 76944 38304 77248 38332
rect 77668 38344 77720 38350
rect 77668 38286 77720 38292
rect 77484 38276 77536 38282
rect 77484 38218 77536 38224
rect 77116 38004 77168 38010
rect 77116 37946 77168 37952
rect 76932 37800 76984 37806
rect 76932 37742 76984 37748
rect 76944 37398 76972 37742
rect 76932 37392 76984 37398
rect 76932 37334 76984 37340
rect 77128 37312 77156 37946
rect 77496 37330 77524 38218
rect 78416 38214 78444 38354
rect 78404 38208 78456 38214
rect 78404 38150 78456 38156
rect 78416 37874 78444 38150
rect 78404 37868 78456 37874
rect 78404 37810 78456 37816
rect 80164 37670 80192 38950
rect 80336 38898 80388 38904
rect 80244 38820 80296 38826
rect 80348 38808 80376 38898
rect 80296 38780 80376 38808
rect 80244 38762 80296 38768
rect 80336 37868 80388 37874
rect 80336 37810 80388 37816
rect 77944 37664 77996 37670
rect 77944 37606 77996 37612
rect 80152 37664 80204 37670
rect 80152 37606 80204 37612
rect 77208 37324 77260 37330
rect 77128 37284 77208 37312
rect 77208 37266 77260 37272
rect 77484 37324 77536 37330
rect 77484 37266 77536 37272
rect 77956 37262 77984 37606
rect 80164 37482 80192 37606
rect 80072 37454 80192 37482
rect 78680 37324 78732 37330
rect 78680 37266 78732 37272
rect 77944 37256 77996 37262
rect 77944 37198 77996 37204
rect 77024 37120 77076 37126
rect 77024 37062 77076 37068
rect 77036 36922 77064 37062
rect 77024 36916 77076 36922
rect 77024 36858 77076 36864
rect 72608 36712 72660 36718
rect 72608 36654 72660 36660
rect 72792 36712 72844 36718
rect 72792 36654 72844 36660
rect 76840 36712 76892 36718
rect 76840 36654 76892 36660
rect 72516 36168 72568 36174
rect 72516 36110 72568 36116
rect 72528 35222 72556 36110
rect 72516 35216 72568 35222
rect 72516 35158 72568 35164
rect 72240 35148 72292 35154
rect 72240 35090 72292 35096
rect 72148 35080 72200 35086
rect 72148 35022 72200 35028
rect 71596 34944 71648 34950
rect 71596 34886 71648 34892
rect 71872 34944 71924 34950
rect 71872 34886 71924 34892
rect 71412 34740 71464 34746
rect 71412 34682 71464 34688
rect 72160 34610 72188 35022
rect 72252 34678 72280 35090
rect 72620 34746 72648 36654
rect 72804 36378 72832 36654
rect 74448 36644 74500 36650
rect 74448 36586 74500 36592
rect 72792 36372 72844 36378
rect 72792 36314 72844 36320
rect 72804 35630 72832 36314
rect 74460 35834 74488 36586
rect 74448 35828 74500 35834
rect 74448 35770 74500 35776
rect 72792 35624 72844 35630
rect 72792 35566 72844 35572
rect 77036 35494 77064 36858
rect 77208 36576 77260 36582
rect 77208 36518 77260 36524
rect 77852 36576 77904 36582
rect 77852 36518 77904 36524
rect 77220 35766 77248 36518
rect 77300 36236 77352 36242
rect 77300 36178 77352 36184
rect 77208 35760 77260 35766
rect 77208 35702 77260 35708
rect 77024 35488 77076 35494
rect 77024 35430 77076 35436
rect 77036 35154 77064 35430
rect 77024 35148 77076 35154
rect 77024 35090 77076 35096
rect 77220 34950 77248 35702
rect 76012 34944 76064 34950
rect 76012 34886 76064 34892
rect 77208 34944 77260 34950
rect 77208 34886 77260 34892
rect 72608 34740 72660 34746
rect 72608 34682 72660 34688
rect 72240 34672 72292 34678
rect 72240 34614 72292 34620
rect 72148 34604 72200 34610
rect 72148 34546 72200 34552
rect 70124 34536 70176 34542
rect 70124 34478 70176 34484
rect 70032 34060 70084 34066
rect 70032 34002 70084 34008
rect 69296 33380 69348 33386
rect 69296 33322 69348 33328
rect 76024 33318 76052 34886
rect 77312 34746 77340 36178
rect 77576 36168 77628 36174
rect 77576 36110 77628 36116
rect 77588 35698 77616 36110
rect 77864 35698 77892 36518
rect 77956 36378 77984 37198
rect 78220 36712 78272 36718
rect 78220 36654 78272 36660
rect 77944 36372 77996 36378
rect 77944 36314 77996 36320
rect 78232 36038 78260 36654
rect 78692 36378 78720 37266
rect 78680 36372 78732 36378
rect 78680 36314 78732 36320
rect 79968 36236 80020 36242
rect 79968 36178 80020 36184
rect 79692 36100 79744 36106
rect 79692 36042 79744 36048
rect 78220 36032 78272 36038
rect 78220 35974 78272 35980
rect 77576 35692 77628 35698
rect 77576 35634 77628 35640
rect 77852 35692 77904 35698
rect 77852 35634 77904 35640
rect 78128 35624 78180 35630
rect 78232 35612 78260 35974
rect 78180 35584 78260 35612
rect 78128 35566 78180 35572
rect 79704 35562 79732 36042
rect 79980 35698 80008 36178
rect 79968 35692 80020 35698
rect 79968 35634 80020 35640
rect 79692 35556 79744 35562
rect 79692 35498 79744 35504
rect 78588 35148 78640 35154
rect 78956 35148 79008 35154
rect 78588 35090 78640 35096
rect 78692 35108 78956 35136
rect 77760 35080 77812 35086
rect 77760 35022 77812 35028
rect 77772 34746 77800 35022
rect 77300 34740 77352 34746
rect 77300 34682 77352 34688
rect 77760 34740 77812 34746
rect 77760 34682 77812 34688
rect 78600 34406 78628 35090
rect 78692 35018 78720 35108
rect 78956 35090 79008 35096
rect 78680 35012 78732 35018
rect 78680 34954 78732 34960
rect 78968 34542 78996 35090
rect 79980 34746 80008 35634
rect 80072 35222 80100 37454
rect 80348 37398 80376 37810
rect 80336 37392 80388 37398
rect 80336 37334 80388 37340
rect 80152 36848 80204 36854
rect 80152 36790 80204 36796
rect 80164 35698 80192 36790
rect 80244 36032 80296 36038
rect 80244 35974 80296 35980
rect 80152 35692 80204 35698
rect 80152 35634 80204 35640
rect 80164 35494 80192 35634
rect 80152 35488 80204 35494
rect 80152 35430 80204 35436
rect 80256 35222 80284 35974
rect 80060 35216 80112 35222
rect 80060 35158 80112 35164
rect 80244 35216 80296 35222
rect 80244 35158 80296 35164
rect 80152 35148 80204 35154
rect 80152 35090 80204 35096
rect 80164 35034 80192 35090
rect 80348 35034 80376 37334
rect 80440 37126 80468 39063
rect 82728 39034 82780 39040
rect 80518 38856 80574 38865
rect 80518 38791 80574 38800
rect 80532 38758 80560 38791
rect 80520 38752 80572 38758
rect 80520 38694 80572 38700
rect 81020 38652 81316 38672
rect 81076 38650 81100 38652
rect 81156 38650 81180 38652
rect 81236 38650 81260 38652
rect 81098 38598 81100 38650
rect 81162 38598 81174 38650
rect 81236 38598 81238 38650
rect 81076 38596 81100 38598
rect 81156 38596 81180 38598
rect 81236 38596 81260 38598
rect 81020 38576 81316 38596
rect 82740 38486 82768 39034
rect 82924 39001 82952 39238
rect 83476 39098 83504 39510
rect 84384 39500 84436 39506
rect 84384 39442 84436 39448
rect 83738 39400 83794 39409
rect 83738 39335 83794 39344
rect 84016 39364 84068 39370
rect 83464 39092 83516 39098
rect 83464 39034 83516 39040
rect 82910 38992 82966 39001
rect 82910 38927 82966 38936
rect 82728 38480 82780 38486
rect 82728 38422 82780 38428
rect 82820 38208 82872 38214
rect 82820 38150 82872 38156
rect 82728 37800 82780 37806
rect 82728 37742 82780 37748
rect 82636 37732 82688 37738
rect 82636 37674 82688 37680
rect 81020 37564 81316 37584
rect 81076 37562 81100 37564
rect 81156 37562 81180 37564
rect 81236 37562 81260 37564
rect 81098 37510 81100 37562
rect 81162 37510 81174 37562
rect 81236 37510 81238 37562
rect 81076 37508 81100 37510
rect 81156 37508 81180 37510
rect 81236 37508 81260 37510
rect 81020 37488 81316 37508
rect 82648 37466 82676 37674
rect 82740 37466 82768 37742
rect 82832 37670 82860 38150
rect 82820 37664 82872 37670
rect 82820 37606 82872 37612
rect 82636 37460 82688 37466
rect 82636 37402 82688 37408
rect 82728 37460 82780 37466
rect 82728 37402 82780 37408
rect 80428 37120 80480 37126
rect 80428 37062 80480 37068
rect 80440 35834 80468 37062
rect 82176 36712 82228 36718
rect 82176 36654 82228 36660
rect 81020 36476 81316 36496
rect 81076 36474 81100 36476
rect 81156 36474 81180 36476
rect 81236 36474 81260 36476
rect 81098 36422 81100 36474
rect 81162 36422 81174 36474
rect 81236 36422 81238 36474
rect 81076 36420 81100 36422
rect 81156 36420 81180 36422
rect 81236 36420 81260 36422
rect 81020 36400 81316 36420
rect 82188 36378 82216 36654
rect 82176 36372 82228 36378
rect 82176 36314 82228 36320
rect 81348 36304 81400 36310
rect 81348 36246 81400 36252
rect 80428 35828 80480 35834
rect 80428 35770 80480 35776
rect 81020 35388 81316 35408
rect 81076 35386 81100 35388
rect 81156 35386 81180 35388
rect 81236 35386 81260 35388
rect 81098 35334 81100 35386
rect 81162 35334 81174 35386
rect 81236 35334 81238 35386
rect 81076 35332 81100 35334
rect 81156 35332 81180 35334
rect 81236 35332 81260 35334
rect 81020 35312 81316 35332
rect 80164 35006 80376 35034
rect 80520 34944 80572 34950
rect 80520 34886 80572 34892
rect 79968 34740 80020 34746
rect 79968 34682 80020 34688
rect 80532 34610 80560 34886
rect 80520 34604 80572 34610
rect 80520 34546 80572 34552
rect 81360 34542 81388 36246
rect 82832 36242 82860 37606
rect 82924 36922 82952 38927
rect 83476 38826 83504 39034
rect 83752 38962 83780 39335
rect 84016 39306 84068 39312
rect 83740 38956 83792 38962
rect 83740 38898 83792 38904
rect 83648 38888 83700 38894
rect 83648 38830 83700 38836
rect 83464 38820 83516 38826
rect 83464 38762 83516 38768
rect 83660 38554 83688 38830
rect 83648 38548 83700 38554
rect 83648 38490 83700 38496
rect 83556 38412 83608 38418
rect 83556 38354 83608 38360
rect 83188 37392 83240 37398
rect 83188 37334 83240 37340
rect 83200 36922 83228 37334
rect 83568 37126 83596 38354
rect 83752 38010 83780 38898
rect 84028 38554 84056 39306
rect 84396 39098 84424 39442
rect 84384 39092 84436 39098
rect 84384 39034 84436 39040
rect 85224 38894 85252 39918
rect 85396 39908 85448 39914
rect 85396 39850 85448 39856
rect 85948 39908 86000 39914
rect 85948 39850 86000 39856
rect 85408 39642 85436 39850
rect 85396 39636 85448 39642
rect 85396 39578 85448 39584
rect 85304 39092 85356 39098
rect 85304 39034 85356 39040
rect 85212 38888 85264 38894
rect 85212 38830 85264 38836
rect 84016 38548 84068 38554
rect 84016 38490 84068 38496
rect 84752 38208 84804 38214
rect 84752 38150 84804 38156
rect 83740 38004 83792 38010
rect 83740 37946 83792 37952
rect 84764 37874 84792 38150
rect 84752 37868 84804 37874
rect 84752 37810 84804 37816
rect 84764 37330 84792 37810
rect 85316 37806 85344 39034
rect 85408 38894 85436 39578
rect 85396 38888 85448 38894
rect 85396 38830 85448 38836
rect 85960 38418 85988 39850
rect 96380 39196 96676 39216
rect 96436 39194 96460 39196
rect 96516 39194 96540 39196
rect 96596 39194 96620 39196
rect 96458 39142 96460 39194
rect 96522 39142 96534 39194
rect 96596 39142 96598 39194
rect 96436 39140 96460 39142
rect 96516 39140 96540 39142
rect 96596 39140 96620 39142
rect 96380 39120 96676 39140
rect 86776 38888 86828 38894
rect 86776 38830 86828 38836
rect 86408 38752 86460 38758
rect 86408 38694 86460 38700
rect 86316 38480 86368 38486
rect 86316 38422 86368 38428
rect 85856 38412 85908 38418
rect 85856 38354 85908 38360
rect 85948 38412 86000 38418
rect 85948 38354 86000 38360
rect 85868 37874 85896 38354
rect 86328 38010 86356 38422
rect 86316 38004 86368 38010
rect 86316 37946 86368 37952
rect 85856 37868 85908 37874
rect 85856 37810 85908 37816
rect 85304 37800 85356 37806
rect 85304 37742 85356 37748
rect 84752 37324 84804 37330
rect 84752 37266 84804 37272
rect 85948 37324 86000 37330
rect 85948 37266 86000 37272
rect 86224 37324 86276 37330
rect 86224 37266 86276 37272
rect 83556 37120 83608 37126
rect 83556 37062 83608 37068
rect 82912 36916 82964 36922
rect 82912 36858 82964 36864
rect 83188 36916 83240 36922
rect 83188 36858 83240 36864
rect 82820 36236 82872 36242
rect 82820 36178 82872 36184
rect 82820 35828 82872 35834
rect 82820 35770 82872 35776
rect 82728 35624 82780 35630
rect 82728 35566 82780 35572
rect 82740 35494 82768 35566
rect 82728 35488 82780 35494
rect 82726 35456 82728 35465
rect 82780 35456 82782 35465
rect 82726 35391 82782 35400
rect 82832 35290 82860 35770
rect 82924 35698 82952 36858
rect 83568 36786 83596 37062
rect 83924 36916 83976 36922
rect 83924 36858 83976 36864
rect 83556 36780 83608 36786
rect 83556 36722 83608 36728
rect 83004 36576 83056 36582
rect 83004 36518 83056 36524
rect 83016 36106 83044 36518
rect 83568 36310 83596 36722
rect 83936 36718 83964 36858
rect 83924 36712 83976 36718
rect 83924 36654 83976 36660
rect 84200 36712 84252 36718
rect 84200 36654 84252 36660
rect 83556 36304 83608 36310
rect 83556 36246 83608 36252
rect 84212 36242 84240 36654
rect 84200 36236 84252 36242
rect 84200 36178 84252 36184
rect 83004 36100 83056 36106
rect 83004 36042 83056 36048
rect 83096 35760 83148 35766
rect 83096 35702 83148 35708
rect 82912 35692 82964 35698
rect 82912 35634 82964 35640
rect 83004 35556 83056 35562
rect 83004 35498 83056 35504
rect 83016 35290 83044 35498
rect 83108 35290 83136 35702
rect 84200 35692 84252 35698
rect 84200 35634 84252 35640
rect 83924 35624 83976 35630
rect 83924 35566 83976 35572
rect 83936 35494 83964 35566
rect 83924 35488 83976 35494
rect 83278 35456 83334 35465
rect 83924 35430 83976 35436
rect 83278 35391 83334 35400
rect 83292 35290 83320 35391
rect 82820 35284 82872 35290
rect 82820 35226 82872 35232
rect 83004 35284 83056 35290
rect 83004 35226 83056 35232
rect 83096 35284 83148 35290
rect 83096 35226 83148 35232
rect 83280 35284 83332 35290
rect 83280 35226 83332 35232
rect 83108 35154 83136 35226
rect 83096 35148 83148 35154
rect 83096 35090 83148 35096
rect 82176 35080 82228 35086
rect 82176 35022 82228 35028
rect 82188 34542 82216 35022
rect 83280 34944 83332 34950
rect 83280 34886 83332 34892
rect 83292 34542 83320 34886
rect 83936 34746 83964 35430
rect 84212 35018 84240 35634
rect 84384 35624 84436 35630
rect 84384 35566 84436 35572
rect 84396 35222 84424 35566
rect 84384 35216 84436 35222
rect 84384 35158 84436 35164
rect 84764 35154 84792 37266
rect 85960 36786 85988 37266
rect 85948 36780 86000 36786
rect 85948 36722 86000 36728
rect 86236 36310 86264 37266
rect 86224 36304 86276 36310
rect 86224 36246 86276 36252
rect 86328 36242 86356 37946
rect 86420 37398 86448 38694
rect 86788 38486 86816 38830
rect 87880 38752 87932 38758
rect 87880 38694 87932 38700
rect 86776 38480 86828 38486
rect 86776 38422 86828 38428
rect 87892 37874 87920 38694
rect 96380 38108 96676 38128
rect 96436 38106 96460 38108
rect 96516 38106 96540 38108
rect 96596 38106 96620 38108
rect 96458 38054 96460 38106
rect 96522 38054 96534 38106
rect 96596 38054 96598 38106
rect 96436 38052 96460 38054
rect 96516 38052 96540 38054
rect 96596 38052 96620 38054
rect 96380 38032 96676 38052
rect 87880 37868 87932 37874
rect 87880 37810 87932 37816
rect 86776 37800 86828 37806
rect 86776 37742 86828 37748
rect 86408 37392 86460 37398
rect 86408 37334 86460 37340
rect 86788 36650 86816 37742
rect 86868 37392 86920 37398
rect 86868 37334 86920 37340
rect 86880 36938 86908 37334
rect 87420 37324 87472 37330
rect 87420 37266 87472 37272
rect 86880 36922 87000 36938
rect 86880 36916 87012 36922
rect 86880 36910 86960 36916
rect 86776 36644 86828 36650
rect 86776 36586 86828 36592
rect 86788 36242 86816 36586
rect 86316 36236 86368 36242
rect 86316 36178 86368 36184
rect 86776 36236 86828 36242
rect 86776 36178 86828 36184
rect 86880 35834 86908 36910
rect 86960 36858 87012 36864
rect 87432 36786 87460 37266
rect 96380 37020 96676 37040
rect 96436 37018 96460 37020
rect 96516 37018 96540 37020
rect 96596 37018 96620 37020
rect 96458 36966 96460 37018
rect 96522 36966 96534 37018
rect 96596 36966 96598 37018
rect 96436 36964 96460 36966
rect 96516 36964 96540 36966
rect 96596 36964 96620 36966
rect 96380 36944 96676 36964
rect 87420 36780 87472 36786
rect 87420 36722 87472 36728
rect 86960 36712 87012 36718
rect 86960 36654 87012 36660
rect 86972 36378 87000 36654
rect 86960 36372 87012 36378
rect 86960 36314 87012 36320
rect 96380 35932 96676 35952
rect 96436 35930 96460 35932
rect 96516 35930 96540 35932
rect 96596 35930 96620 35932
rect 96458 35878 96460 35930
rect 96522 35878 96534 35930
rect 96596 35878 96598 35930
rect 96436 35876 96460 35878
rect 96516 35876 96540 35878
rect 96596 35876 96620 35878
rect 96380 35856 96676 35876
rect 86500 35828 86552 35834
rect 86500 35770 86552 35776
rect 86868 35828 86920 35834
rect 86868 35770 86920 35776
rect 85028 35488 85080 35494
rect 85028 35430 85080 35436
rect 84936 35216 84988 35222
rect 84936 35158 84988 35164
rect 84752 35148 84804 35154
rect 84752 35090 84804 35096
rect 84200 35012 84252 35018
rect 84200 34954 84252 34960
rect 83924 34740 83976 34746
rect 83924 34682 83976 34688
rect 78956 34536 79008 34542
rect 78956 34478 79008 34484
rect 81348 34536 81400 34542
rect 81348 34478 81400 34484
rect 82176 34536 82228 34542
rect 82176 34478 82228 34484
rect 83280 34536 83332 34542
rect 83280 34478 83332 34484
rect 84948 34406 84976 35158
rect 85040 35154 85068 35430
rect 86512 35290 86540 35770
rect 86880 35630 86908 35770
rect 86868 35624 86920 35630
rect 86868 35566 86920 35572
rect 88340 35624 88392 35630
rect 88340 35566 88392 35572
rect 86880 35306 86908 35566
rect 88248 35488 88300 35494
rect 88248 35430 88300 35436
rect 86500 35284 86552 35290
rect 86500 35226 86552 35232
rect 86788 35278 86908 35306
rect 85028 35148 85080 35154
rect 85028 35090 85080 35096
rect 85488 35080 85540 35086
rect 85488 35022 85540 35028
rect 85500 34610 85528 35022
rect 85948 34944 86000 34950
rect 85948 34886 86000 34892
rect 86132 34944 86184 34950
rect 86132 34886 86184 34892
rect 86684 34944 86736 34950
rect 86684 34886 86736 34892
rect 85764 34740 85816 34746
rect 85764 34682 85816 34688
rect 85488 34604 85540 34610
rect 85488 34546 85540 34552
rect 85776 34542 85804 34682
rect 85764 34536 85816 34542
rect 85764 34478 85816 34484
rect 78588 34400 78640 34406
rect 78588 34342 78640 34348
rect 84936 34400 84988 34406
rect 84936 34342 84988 34348
rect 81020 34300 81316 34320
rect 81076 34298 81100 34300
rect 81156 34298 81180 34300
rect 81236 34298 81260 34300
rect 81098 34246 81100 34298
rect 81162 34246 81174 34298
rect 81236 34246 81238 34298
rect 81076 34244 81100 34246
rect 81156 34244 81180 34246
rect 81236 34244 81260 34246
rect 81020 34224 81316 34244
rect 76012 33312 76064 33318
rect 76012 33254 76064 33260
rect 84016 32972 84068 32978
rect 84016 32914 84068 32920
rect 69020 32428 69072 32434
rect 69020 32370 69072 32376
rect 84028 32162 84056 32914
rect 84016 32156 84068 32162
rect 84016 32098 84068 32104
rect 59728 31612 59780 31618
rect 59728 31554 59780 31560
rect 59556 28082 59676 28098
rect 59544 28076 59676 28082
rect 59596 28070 59676 28076
rect 59544 28018 59596 28024
rect 59544 27940 59596 27946
rect 59544 27882 59596 27888
rect 59452 26648 59504 26654
rect 59452 26590 59504 26596
rect 59556 22098 59584 27882
rect 59360 22092 59412 22098
rect 59360 22034 59412 22040
rect 59544 22092 59596 22098
rect 59544 22034 59596 22040
rect 58440 20324 58492 20330
rect 58440 20266 58492 20272
rect 59176 20324 59228 20330
rect 59176 20266 59228 20272
rect 58452 20097 58480 20266
rect 58438 20088 58494 20097
rect 58438 20023 58494 20032
rect 59372 15230 59400 22034
rect 58440 15224 58492 15230
rect 58440 15166 58492 15172
rect 59360 15224 59412 15230
rect 59360 15166 59412 15172
rect 58452 14861 58480 15166
rect 58438 14852 58494 14861
rect 58438 14787 58494 14796
rect 84028 4865 84056 32098
rect 85960 20165 85988 34886
rect 86144 31226 86172 34886
rect 86696 32978 86724 34886
rect 86788 34746 86816 35278
rect 88260 35154 88288 35430
rect 86868 35148 86920 35154
rect 86868 35090 86920 35096
rect 87328 35148 87380 35154
rect 87328 35090 87380 35096
rect 88248 35148 88300 35154
rect 88248 35090 88300 35096
rect 86880 34746 86908 35090
rect 87236 35080 87288 35086
rect 87236 35022 87288 35028
rect 86776 34740 86828 34746
rect 86776 34682 86828 34688
rect 86868 34740 86920 34746
rect 86868 34682 86920 34688
rect 87052 34672 87104 34678
rect 87052 34614 87104 34620
rect 86960 34536 87012 34542
rect 86960 34478 87012 34484
rect 86684 32972 86736 32978
rect 86684 32914 86736 32920
rect 86052 31198 86172 31226
rect 86052 22885 86080 31198
rect 86868 31136 86920 31142
rect 86868 31078 86920 31084
rect 86132 31068 86184 31074
rect 86132 31010 86184 31016
rect 86144 30229 86172 31010
rect 86880 30954 86908 31078
rect 86972 31074 87000 34478
rect 86960 31068 87012 31074
rect 86960 31010 87012 31016
rect 86880 30926 87000 30954
rect 87064 30938 87092 34614
rect 87144 31612 87196 31618
rect 87144 31554 87196 31560
rect 86224 30864 86276 30870
rect 86222 30832 86224 30841
rect 86276 30832 86278 30841
rect 86222 30767 86278 30776
rect 86130 30220 86186 30229
rect 86130 30155 86186 30164
rect 86224 29572 86276 29578
rect 86222 29540 86224 29549
rect 86276 29540 86278 29549
rect 86222 29475 86278 29484
rect 86224 28212 86276 28218
rect 86222 28180 86224 28189
rect 86276 28180 86278 28189
rect 86222 28115 86278 28124
rect 86224 26784 86276 26790
rect 86222 26752 86224 26761
rect 86276 26752 86278 26761
rect 86222 26687 86278 26696
rect 86224 25628 86276 25634
rect 86222 25596 86224 25605
rect 86276 25596 86278 25605
rect 86222 25531 86278 25540
rect 86972 24274 87000 30926
rect 87052 30932 87104 30938
rect 87052 30874 87104 30880
rect 87064 28218 87092 30874
rect 87052 28212 87104 28218
rect 87052 28154 87104 28160
rect 87052 26988 87104 26994
rect 87052 26930 87104 26936
rect 87064 25514 87092 26930
rect 87156 25634 87184 31554
rect 87248 31210 87276 35022
rect 87236 31204 87288 31210
rect 87236 31146 87288 31152
rect 87248 29578 87276 31146
rect 87236 29572 87288 29578
rect 87236 29514 87288 29520
rect 87340 26994 87368 35090
rect 88248 35012 88300 35018
rect 88248 34954 88300 34960
rect 87512 34944 87564 34950
rect 87512 34886 87564 34892
rect 87420 34604 87472 34610
rect 87420 34546 87472 34552
rect 87432 31142 87460 34546
rect 87420 31136 87472 31142
rect 87420 31078 87472 31084
rect 87328 26988 87380 26994
rect 87328 26930 87380 26936
rect 87524 26874 87552 34886
rect 88260 34542 88288 34954
rect 88352 34746 88380 35566
rect 96380 34844 96676 34864
rect 96436 34842 96460 34844
rect 96516 34842 96540 34844
rect 96596 34842 96620 34844
rect 96458 34790 96460 34842
rect 96522 34790 96534 34842
rect 96596 34790 96598 34842
rect 96436 34788 96460 34790
rect 96516 34788 96540 34790
rect 96596 34788 96620 34790
rect 96380 34768 96676 34788
rect 88340 34740 88392 34746
rect 88340 34682 88392 34688
rect 87880 34536 87932 34542
rect 87880 34478 87932 34484
rect 88248 34536 88300 34542
rect 88248 34478 88300 34484
rect 87892 31618 87920 34478
rect 87880 31612 87932 31618
rect 87880 31554 87932 31560
rect 108304 31068 108356 31074
rect 108304 31010 108356 31016
rect 87248 26846 87552 26874
rect 87248 26790 87276 26846
rect 87236 26784 87288 26790
rect 87236 26726 87288 26732
rect 87144 25628 87196 25634
rect 87144 25570 87196 25576
rect 87064 25486 87184 25514
rect 86224 24268 86276 24274
rect 86222 24236 86224 24245
rect 86960 24268 87012 24274
rect 86276 24236 86278 24245
rect 86960 24210 87012 24216
rect 86222 24171 86278 24180
rect 86038 22876 86094 22885
rect 86038 22811 86094 22820
rect 85946 20156 86002 20165
rect 85946 20091 86002 20100
rect 87156 14890 87184 25486
rect 108316 23225 108344 31010
rect 108302 23216 108358 23225
rect 108302 23151 108358 23160
rect 86224 14884 86276 14890
rect 86222 14852 86224 14861
rect 87144 14884 87196 14890
rect 86276 14852 86278 14861
rect 87144 14826 87196 14832
rect 86222 14787 86278 14796
rect 56414 4856 56470 4865
rect 56414 4791 56470 4800
rect 84014 4856 84070 4865
rect 84014 4791 84070 4800
rect 56324 3460 56376 3466
rect 56324 3402 56376 3408
rect 84200 3460 84252 3466
rect 84200 3402 84252 3408
rect 84212 800 84240 3402
rect 3054 368 3110 377
rect 3054 303 3110 312
rect 28078 0 28134 800
rect 84198 0 84254 800
<< via2 >>
rect 4066 45872 4122 45928
rect 2410 45328 2466 45384
rect 7654 44648 7710 44704
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 3974 41656 4030 41712
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 3422 40432 3478 40488
rect 3330 36080 3386 36136
rect 3238 32680 3294 32736
rect 2870 20032 2926 20088
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4066 39908 4122 39944
rect 4066 39888 4068 39908
rect 4068 39888 4120 39908
rect 4120 39888 4122 39908
rect 3974 39344 4030 39400
rect 3514 36216 3570 36272
rect 3698 37440 3754 37496
rect 3606 30232 3662 30288
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4066 38664 4122 38720
rect 4066 38120 4122 38176
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 3790 31456 3846 31512
rect 3514 27920 3570 27976
rect 3514 26696 3570 26752
rect 3514 26016 3570 26072
rect 3330 22480 3386 22536
rect 3698 19488 3754 19544
rect 3422 18264 3478 18320
rect 3330 17720 3386 17776
rect 2686 2624 2742 2680
rect 2778 856 2834 912
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4066 36896 4122 36952
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4066 35672 4122 35728
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4066 34448 4122 34504
rect 4066 33904 4122 33960
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 3974 33224 4030 33280
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4066 32136 4122 32192
rect 6918 41112 6974 41168
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 3974 30912 4030 30968
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4066 29688 4122 29744
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 3974 29008 4030 29064
rect 4066 28464 4122 28520
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4066 27240 4122 27296
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 3974 25472 4030 25528
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 3974 24928 4030 24984
rect 3974 24248 4030 24304
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4066 23704 4122 23760
rect 4066 23024 4122 23080
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4066 21800 4122 21856
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 3974 21256 4030 21312
rect 4066 20712 4122 20768
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 3974 18808 4030 18864
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4066 17040 4122 17096
rect 4066 16496 4122 16552
rect 3882 15816 3938 15872
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 5630 35128 5686 35184
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 50300 44090 50356 44092
rect 50380 44090 50436 44092
rect 50460 44090 50516 44092
rect 50540 44090 50596 44092
rect 50300 44038 50326 44090
rect 50326 44038 50356 44090
rect 50380 44038 50390 44090
rect 50390 44038 50436 44090
rect 50460 44038 50506 44090
rect 50506 44038 50516 44090
rect 50540 44038 50570 44090
rect 50570 44038 50596 44090
rect 50300 44036 50356 44038
rect 50380 44036 50436 44038
rect 50460 44036 50516 44038
rect 50540 44036 50596 44038
rect 3974 15272 4030 15328
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 3330 6840 3386 6896
rect 3698 6296 3754 6352
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 3974 14048 4030 14104
rect 4894 14592 4950 14648
rect 4066 13504 4122 13560
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 3974 12824 4030 12880
rect 4066 12300 4122 12336
rect 4066 12280 4068 12300
rect 4068 12280 4120 12300
rect 4120 12280 4122 12300
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4066 11600 4122 11656
rect 3974 11056 4030 11112
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4066 10512 4122 10568
rect 3974 9832 4030 9888
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4066 9288 4122 9344
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4066 8608 4122 8664
rect 3974 8064 4030 8120
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4066 7384 4122 7440
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 3974 5616 4030 5672
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4066 5072 4122 5128
rect 3974 4392 4030 4448
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4066 3848 4122 3904
rect 3974 3304 4030 3360
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 7470 29008 7526 29064
rect 7562 28736 7618 28792
rect 10414 41812 10470 41848
rect 11334 42064 11390 42120
rect 10414 41792 10416 41812
rect 10416 41792 10468 41812
rect 10468 41792 10470 41812
rect 8114 18028 8116 18048
rect 8116 18028 8168 18048
rect 8168 18028 8170 18048
rect 8114 17992 8170 18028
rect 9126 27532 9182 27568
rect 9126 27512 9128 27532
rect 9128 27512 9180 27532
rect 9180 27512 9182 27532
rect 9770 31476 9826 31512
rect 9770 31456 9772 31476
rect 9772 31456 9824 31476
rect 9824 31456 9826 31476
rect 12530 41964 12532 41984
rect 12532 41964 12584 41984
rect 12584 41964 12586 41984
rect 12530 41928 12586 41964
rect 9954 22752 10010 22808
rect 9586 17992 9642 18048
rect 12714 32000 12770 32056
rect 12714 31764 12716 31784
rect 12716 31764 12768 31784
rect 12768 31764 12770 31784
rect 12714 31728 12770 31764
rect 13542 32544 13598 32600
rect 13910 32544 13966 32600
rect 13818 31764 13820 31784
rect 13820 31764 13872 31784
rect 13872 31764 13874 31784
rect 13818 31728 13874 31764
rect 10506 16652 10562 16688
rect 10506 16632 10508 16652
rect 10508 16632 10560 16652
rect 10560 16632 10562 16652
rect 14186 41792 14242 41848
rect 15014 38664 15070 38720
rect 16394 42200 16450 42256
rect 17590 42336 17646 42392
rect 17498 42220 17554 42256
rect 17498 42200 17500 42220
rect 17500 42200 17552 42220
rect 17552 42200 17554 42220
rect 15474 38664 15530 38720
rect 17866 41928 17922 41984
rect 18050 42336 18106 42392
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 15934 37748 15936 37768
rect 15936 37748 15988 37768
rect 15988 37748 15990 37768
rect 15934 37712 15990 37748
rect 16578 37748 16580 37768
rect 16580 37748 16632 37768
rect 16632 37748 16634 37768
rect 16578 37712 16634 37748
rect 14462 30116 14518 30152
rect 14462 30096 14464 30116
rect 14464 30096 14516 30116
rect 14516 30096 14518 30116
rect 13358 24828 13360 24848
rect 13360 24828 13412 24848
rect 13412 24828 13414 24848
rect 13358 24792 13414 24828
rect 14278 24792 14334 24848
rect 14462 21412 14518 21448
rect 14462 21392 14464 21412
rect 14464 21392 14516 21412
rect 14516 21392 14518 21412
rect 15842 23432 15898 23488
rect 14462 18572 14464 18592
rect 14464 18572 14516 18592
rect 14516 18572 14518 18592
rect 14462 18536 14518 18572
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19246 38392 19302 38448
rect 18050 32020 18106 32056
rect 18050 32000 18052 32020
rect 18052 32000 18104 32020
rect 18104 32000 18106 32020
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 21178 38528 21234 38584
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 18970 32544 19026 32600
rect 19246 31476 19302 31512
rect 19246 31456 19248 31476
rect 19248 31456 19300 31476
rect 19300 31456 19302 31476
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19522 32292 19578 32328
rect 19522 32272 19524 32292
rect 19524 32272 19576 32292
rect 19576 32272 19578 32292
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19706 31900 19708 31920
rect 19708 31900 19760 31920
rect 19760 31900 19762 31920
rect 19706 31864 19762 31900
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 18326 30116 18382 30152
rect 18326 30096 18328 30116
rect 18328 30096 18380 30116
rect 18380 30096 18382 30116
rect 17222 29960 17278 30016
rect 18878 29960 18934 30016
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 17130 18572 17132 18592
rect 17132 18572 17184 18592
rect 17184 18572 17186 18592
rect 17130 18536 17186 18572
rect 18602 22108 18604 22128
rect 18604 22108 18656 22128
rect 18656 22108 18658 22128
rect 18602 22072 18658 22108
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 20350 30932 20406 30968
rect 20350 30912 20352 30932
rect 20352 30912 20404 30932
rect 20404 30912 20406 30932
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 22558 23468 22560 23488
rect 22560 23468 22612 23488
rect 22612 23468 22614 23488
rect 22558 23432 22614 23468
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 24766 40704 24822 40760
rect 23846 38836 23848 38856
rect 23848 38836 23900 38856
rect 23900 38836 23902 38856
rect 23846 38800 23902 38836
rect 25226 38836 25228 38856
rect 25228 38836 25280 38856
rect 25280 38836 25282 38856
rect 25226 38800 25282 38836
rect 23938 38664 23994 38720
rect 24582 38664 24638 38720
rect 24766 32308 24768 32328
rect 24768 32308 24820 32328
rect 24820 32308 24822 32328
rect 24766 32272 24822 32308
rect 23938 20748 23940 20768
rect 23940 20748 23992 20768
rect 23992 20748 23994 20768
rect 23938 20712 23994 20748
rect 22558 17312 22614 17368
rect 21914 15988 21916 16008
rect 21916 15988 21968 16008
rect 21968 15988 21970 16008
rect 21914 15952 21970 15988
rect 25870 38528 25926 38584
rect 29826 41112 29882 41168
rect 28262 39752 28318 39808
rect 25686 31864 25742 31920
rect 25042 19216 25098 19272
rect 25410 19216 25466 19272
rect 24858 15272 24914 15328
rect 24030 13932 24086 13968
rect 24030 13912 24032 13932
rect 24032 13912 24084 13932
rect 24084 13912 24086 13932
rect 26698 38820 26754 38856
rect 26698 38800 26700 38820
rect 26700 38800 26752 38820
rect 26752 38800 26754 38820
rect 26790 38664 26846 38720
rect 27250 39380 27252 39400
rect 27252 39380 27304 39400
rect 27304 39380 27306 39400
rect 27250 39344 27306 39380
rect 27526 38548 27582 38584
rect 27526 38528 27528 38548
rect 27528 38528 27580 38548
rect 27580 38528 27582 38548
rect 30654 41112 30710 41168
rect 30654 38412 30710 38448
rect 30654 38392 30656 38412
rect 30656 38392 30708 38412
rect 30708 38392 30710 38412
rect 31022 39516 31024 39536
rect 31024 39516 31076 39536
rect 31076 39516 31078 39536
rect 31022 39480 31078 39516
rect 29090 37440 29146 37496
rect 27802 34720 27858 34776
rect 27618 31728 27674 31784
rect 27526 30912 27582 30968
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 28906 35148 28962 35184
rect 28906 35128 28908 35148
rect 28908 35128 28960 35148
rect 28960 35128 28962 35148
rect 28722 34584 28778 34640
rect 29550 34720 29606 34776
rect 32218 39888 32274 39944
rect 29642 30776 29698 30832
rect 28998 30096 29054 30152
rect 28906 29416 28962 29472
rect 28998 28056 29054 28112
rect 28906 26696 28962 26752
rect 28998 25472 29054 25528
rect 28998 24148 29000 24168
rect 29000 24148 29052 24168
rect 29052 24148 29054 24168
rect 28998 24112 29054 24148
rect 29090 22772 29146 22808
rect 29090 22752 29092 22772
rect 29092 22752 29144 22772
rect 29144 22752 29146 22772
rect 29090 20032 29146 20088
rect 27710 18672 27766 18728
rect 28998 14728 29054 14784
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34610 40704 34666 40760
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 35070 39480 35126 39536
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 37278 41656 37334 41712
rect 38658 41692 38660 41712
rect 38660 41692 38712 41712
rect 38712 41692 38714 41712
rect 38658 41656 38714 41692
rect 38658 40976 38714 41032
rect 38106 39616 38162 39672
rect 39026 40976 39082 41032
rect 39026 40876 39028 40896
rect 39028 40876 39080 40896
rect 39080 40876 39082 40896
rect 39026 40840 39082 40876
rect 36542 38528 36598 38584
rect 37094 38528 37150 38584
rect 35622 37712 35678 37768
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 33690 36372 33746 36408
rect 33690 36352 33692 36372
rect 33692 36352 33744 36372
rect 33744 36352 33746 36372
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 35990 36352 36046 36408
rect 35898 36216 35954 36272
rect 36542 37732 36598 37768
rect 36542 37712 36544 37732
rect 36544 37712 36596 37732
rect 36596 37712 36598 37732
rect 37738 38412 37794 38448
rect 37738 38392 37740 38412
rect 37740 38392 37792 38412
rect 37792 38392 37794 38412
rect 38842 38276 38898 38312
rect 38842 38256 38844 38276
rect 38844 38256 38896 38276
rect 38896 38256 38898 38276
rect 38290 37440 38346 37496
rect 37554 36216 37610 36272
rect 38658 35944 38714 36000
rect 38382 35672 38438 35728
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 39946 35808 40002 35864
rect 41142 39480 41198 39536
rect 40866 39072 40922 39128
rect 41050 39208 41106 39264
rect 40958 38936 41014 38992
rect 42246 39480 42302 39536
rect 42338 39208 42394 39264
rect 44638 41520 44694 41576
rect 45926 41520 45982 41576
rect 46294 40840 46350 40896
rect 42982 38936 43038 38992
rect 41326 36916 41382 36952
rect 41326 36896 41328 36916
rect 41328 36896 41380 36916
rect 41380 36896 41382 36916
rect 40866 35672 40922 35728
rect 40222 35128 40278 35184
rect 40682 35128 40738 35184
rect 41234 35284 41290 35320
rect 41234 35264 41236 35284
rect 41236 35264 41288 35284
rect 41288 35264 41290 35284
rect 41510 35264 41566 35320
rect 41418 35148 41474 35184
rect 41418 35128 41420 35148
rect 41420 35128 41472 35148
rect 41472 35128 41474 35148
rect 42614 37576 42670 37632
rect 42522 35808 42578 35864
rect 42246 35148 42302 35184
rect 42246 35128 42248 35148
rect 42248 35128 42300 35148
rect 42300 35128 42302 35148
rect 43258 39208 43314 39264
rect 43258 38700 43260 38720
rect 43260 38700 43312 38720
rect 43312 38700 43314 38720
rect 43258 38664 43314 38700
rect 43534 39344 43590 39400
rect 43994 39364 44050 39400
rect 43994 39344 43996 39364
rect 43996 39344 44048 39364
rect 44048 39344 44050 39364
rect 44178 39208 44234 39264
rect 43442 37612 43444 37632
rect 43444 37612 43496 37632
rect 43496 37612 43498 37632
rect 43442 37576 43498 37612
rect 44454 39072 44510 39128
rect 44638 39380 44640 39400
rect 44640 39380 44692 39400
rect 44692 39380 44694 39400
rect 44638 39344 44694 39380
rect 46110 38256 46166 38312
rect 46018 36236 46074 36272
rect 46018 36216 46020 36236
rect 46020 36216 46072 36236
rect 46072 36216 46074 36236
rect 43534 36080 43590 36136
rect 44914 36116 44916 36136
rect 44916 36116 44968 36136
rect 44968 36116 44970 36136
rect 44914 36080 44970 36116
rect 45834 35944 45890 36000
rect 47398 38956 47454 38992
rect 47398 38936 47400 38956
rect 47400 38936 47452 38956
rect 47452 38936 47454 38956
rect 48594 39788 48596 39808
rect 48596 39788 48648 39808
rect 48648 39788 48650 39808
rect 48594 39752 48650 39788
rect 48134 39616 48190 39672
rect 47858 38820 47914 38856
rect 47858 38800 47860 38820
rect 47860 38800 47912 38820
rect 47912 38800 47914 38820
rect 48778 39344 48834 39400
rect 48686 39208 48742 39264
rect 50300 43002 50356 43004
rect 50380 43002 50436 43004
rect 50460 43002 50516 43004
rect 50540 43002 50596 43004
rect 50300 42950 50326 43002
rect 50326 42950 50356 43002
rect 50380 42950 50390 43002
rect 50390 42950 50436 43002
rect 50460 42950 50506 43002
rect 50506 42950 50516 43002
rect 50540 42950 50570 43002
rect 50570 42950 50596 43002
rect 50300 42948 50356 42950
rect 50380 42948 50436 42950
rect 50460 42948 50516 42950
rect 50540 42948 50596 42950
rect 50300 41914 50356 41916
rect 50380 41914 50436 41916
rect 50460 41914 50516 41916
rect 50540 41914 50596 41916
rect 50300 41862 50326 41914
rect 50326 41862 50356 41914
rect 50380 41862 50390 41914
rect 50390 41862 50436 41914
rect 50460 41862 50506 41914
rect 50506 41862 50516 41914
rect 50540 41862 50570 41914
rect 50570 41862 50596 41914
rect 50300 41860 50356 41862
rect 50380 41860 50436 41862
rect 50460 41860 50516 41862
rect 50540 41860 50596 41862
rect 51446 41928 51502 41984
rect 50300 40826 50356 40828
rect 50380 40826 50436 40828
rect 50460 40826 50516 40828
rect 50540 40826 50596 40828
rect 50300 40774 50326 40826
rect 50326 40774 50356 40826
rect 50380 40774 50390 40826
rect 50390 40774 50436 40826
rect 50460 40774 50506 40826
rect 50506 40774 50516 40826
rect 50540 40774 50570 40826
rect 50570 40774 50596 40826
rect 50300 40772 50356 40774
rect 50380 40772 50436 40774
rect 50460 40772 50516 40774
rect 50540 40772 50596 40774
rect 50300 39738 50356 39740
rect 50380 39738 50436 39740
rect 50460 39738 50516 39740
rect 50540 39738 50596 39740
rect 50300 39686 50326 39738
rect 50326 39686 50356 39738
rect 50380 39686 50390 39738
rect 50390 39686 50436 39738
rect 50460 39686 50506 39738
rect 50506 39686 50516 39738
rect 50540 39686 50570 39738
rect 50570 39686 50596 39738
rect 50300 39684 50356 39686
rect 50380 39684 50436 39686
rect 50460 39684 50516 39686
rect 50540 39684 50596 39686
rect 53378 40876 53380 40896
rect 53380 40876 53432 40896
rect 53432 40876 53434 40896
rect 53378 40840 53434 40876
rect 51998 39516 52000 39536
rect 52000 39516 52052 39536
rect 52052 39516 52054 39536
rect 51998 39480 52054 39516
rect 48686 38936 48742 38992
rect 48042 38664 48098 38720
rect 50300 38650 50356 38652
rect 50380 38650 50436 38652
rect 50460 38650 50516 38652
rect 50540 38650 50596 38652
rect 50300 38598 50326 38650
rect 50326 38598 50356 38650
rect 50380 38598 50390 38650
rect 50390 38598 50436 38650
rect 50460 38598 50506 38650
rect 50506 38598 50516 38650
rect 50540 38598 50570 38650
rect 50570 38598 50596 38650
rect 50300 38596 50356 38598
rect 50380 38596 50436 38598
rect 50460 38596 50516 38598
rect 50540 38596 50596 38598
rect 47306 36896 47362 36952
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 48962 34992 49018 35048
rect 46662 34604 46718 34640
rect 46662 34584 46664 34604
rect 46664 34584 46716 34604
rect 46716 34584 46718 34604
rect 50986 37168 51042 37224
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 49790 36216 49846 36272
rect 50802 36660 50804 36680
rect 50804 36660 50856 36680
rect 50856 36660 50858 36680
rect 50802 36624 50858 36660
rect 51906 37576 51962 37632
rect 55034 42084 55090 42120
rect 55034 42064 55036 42084
rect 55036 42064 55088 42084
rect 55088 42064 55090 42084
rect 55954 41928 56010 41984
rect 53286 38936 53342 38992
rect 54574 39480 54630 39536
rect 60646 41148 60648 41168
rect 60648 41148 60700 41168
rect 60700 41148 60702 41168
rect 60646 41112 60702 41148
rect 65660 43546 65716 43548
rect 65740 43546 65796 43548
rect 65820 43546 65876 43548
rect 65900 43546 65956 43548
rect 65660 43494 65686 43546
rect 65686 43494 65716 43546
rect 65740 43494 65750 43546
rect 65750 43494 65796 43546
rect 65820 43494 65866 43546
rect 65866 43494 65876 43546
rect 65900 43494 65930 43546
rect 65930 43494 65956 43546
rect 65660 43492 65716 43494
rect 65740 43492 65796 43494
rect 65820 43492 65876 43494
rect 65900 43492 65956 43494
rect 57242 40840 57298 40896
rect 58806 40840 58862 40896
rect 51630 36216 51686 36272
rect 49146 35128 49202 35184
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 50434 35148 50490 35184
rect 50434 35128 50436 35148
rect 50436 35128 50488 35148
rect 50488 35128 50490 35148
rect 49422 34720 49478 34776
rect 50250 34740 50306 34776
rect 50250 34720 50252 34740
rect 50252 34720 50304 34740
rect 50304 34720 50306 34740
rect 49790 34620 49792 34640
rect 49792 34620 49844 34640
rect 49844 34620 49846 34640
rect 51262 35128 51318 35184
rect 56138 39344 56194 39400
rect 55770 38836 55772 38856
rect 55772 38836 55824 38856
rect 55824 38836 55826 38856
rect 55770 38800 55826 38836
rect 56230 39208 56286 39264
rect 49790 34584 49846 34620
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 52642 34992 52698 35048
rect 54206 36660 54208 36680
rect 54208 36660 54260 36680
rect 54260 36660 54262 36680
rect 54206 36624 54262 36660
rect 57058 37460 57114 37496
rect 57058 37440 57060 37460
rect 57060 37440 57112 37460
rect 57112 37440 57114 37460
rect 57242 37576 57298 37632
rect 57794 37460 57850 37496
rect 57794 37440 57796 37460
rect 57796 37440 57848 37460
rect 57848 37440 57850 37460
rect 57150 37304 57206 37360
rect 55678 37168 55734 37224
rect 63130 41148 63132 41168
rect 63132 41148 63184 41168
rect 63184 41148 63186 41168
rect 63130 41112 63186 41148
rect 62210 39500 62266 39536
rect 62210 39480 62212 39500
rect 62212 39480 62264 39500
rect 62264 39480 62266 39500
rect 61934 39344 61990 39400
rect 64326 40876 64328 40896
rect 64328 40876 64380 40896
rect 64380 40876 64382 40896
rect 64326 40840 64382 40876
rect 63590 39480 63646 39536
rect 65660 42458 65716 42460
rect 65740 42458 65796 42460
rect 65820 42458 65876 42460
rect 65900 42458 65956 42460
rect 65660 42406 65686 42458
rect 65686 42406 65716 42458
rect 65740 42406 65750 42458
rect 65750 42406 65796 42458
rect 65820 42406 65866 42458
rect 65866 42406 65876 42458
rect 65900 42406 65930 42458
rect 65930 42406 65956 42458
rect 65660 42404 65716 42406
rect 65740 42404 65796 42406
rect 65820 42404 65876 42406
rect 65900 42404 65956 42406
rect 65660 41370 65716 41372
rect 65740 41370 65796 41372
rect 65820 41370 65876 41372
rect 65900 41370 65956 41372
rect 65660 41318 65686 41370
rect 65686 41318 65716 41370
rect 65740 41318 65750 41370
rect 65750 41318 65796 41370
rect 65820 41318 65866 41370
rect 65866 41318 65876 41370
rect 65900 41318 65930 41370
rect 65930 41318 65956 41370
rect 65660 41316 65716 41318
rect 65740 41316 65796 41318
rect 65820 41316 65876 41318
rect 65900 41316 65956 41318
rect 64602 39500 64658 39536
rect 64602 39480 64604 39500
rect 64604 39480 64656 39500
rect 64656 39480 64658 39500
rect 65660 40282 65716 40284
rect 65740 40282 65796 40284
rect 65820 40282 65876 40284
rect 65900 40282 65956 40284
rect 65660 40230 65686 40282
rect 65686 40230 65716 40282
rect 65740 40230 65750 40282
rect 65750 40230 65796 40282
rect 65820 40230 65866 40282
rect 65866 40230 65876 40282
rect 65900 40230 65930 40282
rect 65930 40230 65956 40282
rect 65660 40228 65716 40230
rect 65740 40228 65796 40230
rect 65820 40228 65876 40230
rect 65900 40228 65956 40230
rect 55954 35028 55956 35048
rect 55956 35028 56008 35048
rect 56008 35028 56010 35048
rect 55954 34992 56010 35028
rect 56782 34604 56838 34640
rect 56782 34584 56784 34604
rect 56784 34584 56836 34604
rect 56836 34584 56838 34604
rect 57058 34720 57114 34776
rect 56598 31220 56600 31240
rect 56600 31220 56652 31240
rect 56652 31220 56654 31240
rect 56598 31184 56654 31220
rect 56874 31184 56930 31240
rect 56322 30776 56378 30832
rect 29918 4800 29974 4856
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 4066 2080 4122 2136
rect 3790 1400 3846 1456
rect 65660 39194 65716 39196
rect 65740 39194 65796 39196
rect 65820 39194 65876 39196
rect 65900 39194 65956 39196
rect 65660 39142 65686 39194
rect 65686 39142 65716 39194
rect 65740 39142 65750 39194
rect 65750 39142 65796 39194
rect 65820 39142 65866 39194
rect 65866 39142 65876 39194
rect 65900 39142 65930 39194
rect 65930 39142 65956 39194
rect 65660 39140 65716 39142
rect 65740 39140 65796 39142
rect 65820 39140 65876 39142
rect 65900 39140 65956 39142
rect 81020 44090 81076 44092
rect 81100 44090 81156 44092
rect 81180 44090 81236 44092
rect 81260 44090 81316 44092
rect 81020 44038 81046 44090
rect 81046 44038 81076 44090
rect 81100 44038 81110 44090
rect 81110 44038 81156 44090
rect 81180 44038 81226 44090
rect 81226 44038 81236 44090
rect 81260 44038 81290 44090
rect 81290 44038 81316 44090
rect 81020 44036 81076 44038
rect 81100 44036 81156 44038
rect 81180 44036 81236 44038
rect 81260 44036 81316 44038
rect 68466 40024 68522 40080
rect 66534 39364 66590 39400
rect 66534 39344 66536 39364
rect 66536 39344 66588 39364
rect 66588 39344 66590 39364
rect 58622 34604 58678 34640
rect 58622 34584 58624 34604
rect 58624 34584 58676 34604
rect 58676 34584 58678 34604
rect 58438 30132 58440 30152
rect 58440 30132 58492 30152
rect 58492 30132 58494 30152
rect 58438 30096 58494 30132
rect 58438 29416 58494 29472
rect 58438 28024 58440 28044
rect 58440 28024 58492 28044
rect 58492 28024 58494 28044
rect 58438 27988 58494 28024
rect 56414 27104 56470 27160
rect 57426 27104 57482 27160
rect 58438 26800 58440 26820
rect 58440 26800 58492 26820
rect 58492 26800 58494 26820
rect 58438 26764 58494 26800
rect 58070 24112 58126 24168
rect 58438 25540 58494 25596
rect 58438 24112 58494 24168
rect 58346 23432 58402 23488
rect 58070 23296 58126 23352
rect 58438 22752 58494 22808
rect 61750 34856 61806 34912
rect 62302 34584 62358 34640
rect 63038 34992 63094 35048
rect 65660 38106 65716 38108
rect 65740 38106 65796 38108
rect 65820 38106 65876 38108
rect 65900 38106 65956 38108
rect 65660 38054 65686 38106
rect 65686 38054 65716 38106
rect 65740 38054 65750 38106
rect 65750 38054 65796 38106
rect 65820 38054 65866 38106
rect 65866 38054 65876 38106
rect 65900 38054 65930 38106
rect 65930 38054 65956 38106
rect 65660 38052 65716 38054
rect 65740 38052 65796 38054
rect 65820 38052 65876 38054
rect 65900 38052 65956 38054
rect 65660 37018 65716 37020
rect 65740 37018 65796 37020
rect 65820 37018 65876 37020
rect 65900 37018 65956 37020
rect 65660 36966 65686 37018
rect 65686 36966 65716 37018
rect 65740 36966 65750 37018
rect 65750 36966 65796 37018
rect 65820 36966 65866 37018
rect 65866 36966 65876 37018
rect 65900 36966 65930 37018
rect 65930 36966 65956 37018
rect 65660 36964 65716 36966
rect 65740 36964 65796 36966
rect 65820 36964 65876 36966
rect 65900 36964 65956 36966
rect 65660 35930 65716 35932
rect 65740 35930 65796 35932
rect 65820 35930 65876 35932
rect 65900 35930 65956 35932
rect 65660 35878 65686 35930
rect 65686 35878 65716 35930
rect 65740 35878 65750 35930
rect 65750 35878 65796 35930
rect 65820 35878 65866 35930
rect 65866 35878 65876 35930
rect 65900 35878 65930 35930
rect 65930 35878 65956 35930
rect 65660 35876 65716 35878
rect 65740 35876 65796 35878
rect 65820 35876 65876 35878
rect 65900 35876 65956 35878
rect 68558 38936 68614 38992
rect 68466 38800 68522 38856
rect 96380 43546 96436 43548
rect 96460 43546 96516 43548
rect 96540 43546 96596 43548
rect 96620 43546 96676 43548
rect 96380 43494 96406 43546
rect 96406 43494 96436 43546
rect 96460 43494 96470 43546
rect 96470 43494 96516 43546
rect 96540 43494 96586 43546
rect 96586 43494 96596 43546
rect 96620 43494 96650 43546
rect 96650 43494 96676 43546
rect 96380 43492 96436 43494
rect 96460 43492 96516 43494
rect 96540 43492 96596 43494
rect 96620 43492 96676 43494
rect 81020 43002 81076 43004
rect 81100 43002 81156 43004
rect 81180 43002 81236 43004
rect 81260 43002 81316 43004
rect 81020 42950 81046 43002
rect 81046 42950 81076 43002
rect 81100 42950 81110 43002
rect 81110 42950 81156 43002
rect 81180 42950 81226 43002
rect 81226 42950 81236 43002
rect 81260 42950 81290 43002
rect 81290 42950 81316 43002
rect 81020 42948 81076 42950
rect 81100 42948 81156 42950
rect 81180 42948 81236 42950
rect 81260 42948 81316 42950
rect 96380 42458 96436 42460
rect 96460 42458 96516 42460
rect 96540 42458 96596 42460
rect 96620 42458 96676 42460
rect 96380 42406 96406 42458
rect 96406 42406 96436 42458
rect 96460 42406 96470 42458
rect 96470 42406 96516 42458
rect 96540 42406 96586 42458
rect 96586 42406 96596 42458
rect 96620 42406 96650 42458
rect 96650 42406 96676 42458
rect 96380 42404 96436 42406
rect 96460 42404 96516 42406
rect 96540 42404 96596 42406
rect 96620 42404 96676 42406
rect 81020 41914 81076 41916
rect 81100 41914 81156 41916
rect 81180 41914 81236 41916
rect 81260 41914 81316 41916
rect 81020 41862 81046 41914
rect 81046 41862 81076 41914
rect 81100 41862 81110 41914
rect 81110 41862 81156 41914
rect 81180 41862 81226 41914
rect 81226 41862 81236 41914
rect 81260 41862 81290 41914
rect 81290 41862 81316 41914
rect 81020 41860 81076 41862
rect 81100 41860 81156 41862
rect 81180 41860 81236 41862
rect 81260 41860 81316 41862
rect 68742 38700 68744 38720
rect 68744 38700 68796 38720
rect 68796 38700 68798 38720
rect 68742 38664 68798 38700
rect 71410 40024 71466 40080
rect 69110 38936 69166 38992
rect 69478 38820 69534 38856
rect 69478 38800 69480 38820
rect 69480 38800 69532 38820
rect 69532 38800 69534 38820
rect 64694 34892 64696 34912
rect 64696 34892 64748 34912
rect 64748 34892 64750 34912
rect 64694 34856 64750 34892
rect 65660 34842 65716 34844
rect 65740 34842 65796 34844
rect 65820 34842 65876 34844
rect 65900 34842 65956 34844
rect 65660 34790 65686 34842
rect 65686 34790 65716 34842
rect 65740 34790 65750 34842
rect 65750 34790 65796 34842
rect 65820 34790 65866 34842
rect 65866 34790 65876 34842
rect 65900 34790 65930 34842
rect 65930 34790 65956 34842
rect 65660 34788 65716 34790
rect 65740 34788 65796 34790
rect 65820 34788 65876 34790
rect 65900 34788 65956 34790
rect 72606 39888 72662 39944
rect 75734 38956 75790 38992
rect 75734 38936 75736 38956
rect 75736 38936 75788 38956
rect 75788 38936 75790 38956
rect 76286 38700 76288 38720
rect 76288 38700 76340 38720
rect 76340 38700 76342 38720
rect 76286 38664 76342 38700
rect 70950 36760 71006 36816
rect 69294 35148 69350 35184
rect 69294 35128 69296 35148
rect 69296 35128 69348 35148
rect 69348 35128 69350 35148
rect 71318 35128 71374 35184
rect 71962 36780 72018 36816
rect 71962 36760 71964 36780
rect 71964 36760 72016 36780
rect 72016 36760 72018 36780
rect 96380 41370 96436 41372
rect 96460 41370 96516 41372
rect 96540 41370 96596 41372
rect 96620 41370 96676 41372
rect 96380 41318 96406 41370
rect 96406 41318 96436 41370
rect 96460 41318 96470 41370
rect 96470 41318 96516 41370
rect 96540 41318 96586 41370
rect 96586 41318 96596 41370
rect 96620 41318 96650 41370
rect 96650 41318 96676 41370
rect 96380 41316 96436 41318
rect 96460 41316 96516 41318
rect 96540 41316 96596 41318
rect 96620 41316 96676 41318
rect 77574 38956 77630 38992
rect 77574 38936 77576 38956
rect 77576 38936 77628 38956
rect 77628 38936 77630 38956
rect 77574 38700 77576 38720
rect 77576 38700 77628 38720
rect 77628 38700 77630 38720
rect 77574 38664 77630 38700
rect 81020 40826 81076 40828
rect 81100 40826 81156 40828
rect 81180 40826 81236 40828
rect 81260 40826 81316 40828
rect 81020 40774 81046 40826
rect 81046 40774 81076 40826
rect 81100 40774 81110 40826
rect 81110 40774 81156 40826
rect 81180 40774 81226 40826
rect 81226 40774 81236 40826
rect 81260 40774 81290 40826
rect 81290 40774 81316 40826
rect 81020 40772 81076 40774
rect 81100 40772 81156 40774
rect 81180 40772 81236 40774
rect 81260 40772 81316 40774
rect 78034 39344 78090 39400
rect 78954 39208 79010 39264
rect 79138 39072 79194 39128
rect 79598 38956 79654 38992
rect 79598 38936 79600 38956
rect 79600 38936 79652 38956
rect 79652 38936 79654 38956
rect 79782 38972 79784 38992
rect 79784 38972 79836 38992
rect 79836 38972 79838 38992
rect 79782 38936 79838 38972
rect 79414 38800 79470 38856
rect 96380 40282 96436 40284
rect 96460 40282 96516 40284
rect 96540 40282 96596 40284
rect 96620 40282 96676 40284
rect 96380 40230 96406 40282
rect 96406 40230 96436 40282
rect 96460 40230 96470 40282
rect 96470 40230 96516 40282
rect 96540 40230 96586 40282
rect 96586 40230 96596 40282
rect 96620 40230 96650 40282
rect 96650 40230 96676 40282
rect 96380 40228 96436 40230
rect 96460 40228 96516 40230
rect 96540 40228 96596 40230
rect 96620 40228 96676 40230
rect 81020 39738 81076 39740
rect 81100 39738 81156 39740
rect 81180 39738 81236 39740
rect 81260 39738 81316 39740
rect 81020 39686 81046 39738
rect 81046 39686 81076 39738
rect 81100 39686 81110 39738
rect 81110 39686 81156 39738
rect 81180 39686 81226 39738
rect 81226 39686 81236 39738
rect 81260 39686 81290 39738
rect 81290 39686 81316 39738
rect 81020 39684 81076 39686
rect 81100 39684 81156 39686
rect 81180 39684 81236 39686
rect 81260 39684 81316 39686
rect 80702 39208 80758 39264
rect 80426 39072 80482 39128
rect 78218 38700 78220 38720
rect 78220 38700 78272 38720
rect 78272 38700 78274 38720
rect 78218 38664 78274 38700
rect 80518 38800 80574 38856
rect 81020 38650 81076 38652
rect 81100 38650 81156 38652
rect 81180 38650 81236 38652
rect 81260 38650 81316 38652
rect 81020 38598 81046 38650
rect 81046 38598 81076 38650
rect 81100 38598 81110 38650
rect 81110 38598 81156 38650
rect 81180 38598 81226 38650
rect 81226 38598 81236 38650
rect 81260 38598 81290 38650
rect 81290 38598 81316 38650
rect 81020 38596 81076 38598
rect 81100 38596 81156 38598
rect 81180 38596 81236 38598
rect 81260 38596 81316 38598
rect 83738 39344 83794 39400
rect 82910 38936 82966 38992
rect 81020 37562 81076 37564
rect 81100 37562 81156 37564
rect 81180 37562 81236 37564
rect 81260 37562 81316 37564
rect 81020 37510 81046 37562
rect 81046 37510 81076 37562
rect 81100 37510 81110 37562
rect 81110 37510 81156 37562
rect 81180 37510 81226 37562
rect 81226 37510 81236 37562
rect 81260 37510 81290 37562
rect 81290 37510 81316 37562
rect 81020 37508 81076 37510
rect 81100 37508 81156 37510
rect 81180 37508 81236 37510
rect 81260 37508 81316 37510
rect 81020 36474 81076 36476
rect 81100 36474 81156 36476
rect 81180 36474 81236 36476
rect 81260 36474 81316 36476
rect 81020 36422 81046 36474
rect 81046 36422 81076 36474
rect 81100 36422 81110 36474
rect 81110 36422 81156 36474
rect 81180 36422 81226 36474
rect 81226 36422 81236 36474
rect 81260 36422 81290 36474
rect 81290 36422 81316 36474
rect 81020 36420 81076 36422
rect 81100 36420 81156 36422
rect 81180 36420 81236 36422
rect 81260 36420 81316 36422
rect 81020 35386 81076 35388
rect 81100 35386 81156 35388
rect 81180 35386 81236 35388
rect 81260 35386 81316 35388
rect 81020 35334 81046 35386
rect 81046 35334 81076 35386
rect 81100 35334 81110 35386
rect 81110 35334 81156 35386
rect 81180 35334 81226 35386
rect 81226 35334 81236 35386
rect 81260 35334 81290 35386
rect 81290 35334 81316 35386
rect 81020 35332 81076 35334
rect 81100 35332 81156 35334
rect 81180 35332 81236 35334
rect 81260 35332 81316 35334
rect 96380 39194 96436 39196
rect 96460 39194 96516 39196
rect 96540 39194 96596 39196
rect 96620 39194 96676 39196
rect 96380 39142 96406 39194
rect 96406 39142 96436 39194
rect 96460 39142 96470 39194
rect 96470 39142 96516 39194
rect 96540 39142 96586 39194
rect 96586 39142 96596 39194
rect 96620 39142 96650 39194
rect 96650 39142 96676 39194
rect 96380 39140 96436 39142
rect 96460 39140 96516 39142
rect 96540 39140 96596 39142
rect 96620 39140 96676 39142
rect 82726 35436 82728 35456
rect 82728 35436 82780 35456
rect 82780 35436 82782 35456
rect 82726 35400 82782 35436
rect 83278 35400 83334 35456
rect 96380 38106 96436 38108
rect 96460 38106 96516 38108
rect 96540 38106 96596 38108
rect 96620 38106 96676 38108
rect 96380 38054 96406 38106
rect 96406 38054 96436 38106
rect 96460 38054 96470 38106
rect 96470 38054 96516 38106
rect 96540 38054 96586 38106
rect 96586 38054 96596 38106
rect 96620 38054 96650 38106
rect 96650 38054 96676 38106
rect 96380 38052 96436 38054
rect 96460 38052 96516 38054
rect 96540 38052 96596 38054
rect 96620 38052 96676 38054
rect 96380 37018 96436 37020
rect 96460 37018 96516 37020
rect 96540 37018 96596 37020
rect 96620 37018 96676 37020
rect 96380 36966 96406 37018
rect 96406 36966 96436 37018
rect 96460 36966 96470 37018
rect 96470 36966 96516 37018
rect 96540 36966 96586 37018
rect 96586 36966 96596 37018
rect 96620 36966 96650 37018
rect 96650 36966 96676 37018
rect 96380 36964 96436 36966
rect 96460 36964 96516 36966
rect 96540 36964 96596 36966
rect 96620 36964 96676 36966
rect 96380 35930 96436 35932
rect 96460 35930 96516 35932
rect 96540 35930 96596 35932
rect 96620 35930 96676 35932
rect 96380 35878 96406 35930
rect 96406 35878 96436 35930
rect 96460 35878 96470 35930
rect 96470 35878 96516 35930
rect 96540 35878 96586 35930
rect 96586 35878 96596 35930
rect 96620 35878 96650 35930
rect 96650 35878 96676 35930
rect 96380 35876 96436 35878
rect 96460 35876 96516 35878
rect 96540 35876 96596 35878
rect 96620 35876 96676 35878
rect 81020 34298 81076 34300
rect 81100 34298 81156 34300
rect 81180 34298 81236 34300
rect 81260 34298 81316 34300
rect 81020 34246 81046 34298
rect 81046 34246 81076 34298
rect 81100 34246 81110 34298
rect 81110 34246 81156 34298
rect 81180 34246 81226 34298
rect 81226 34246 81236 34298
rect 81260 34246 81290 34298
rect 81290 34246 81316 34298
rect 81020 34244 81076 34246
rect 81100 34244 81156 34246
rect 81180 34244 81236 34246
rect 81260 34244 81316 34246
rect 58438 20032 58494 20088
rect 58438 14796 58494 14852
rect 86222 30812 86224 30832
rect 86224 30812 86276 30832
rect 86276 30812 86278 30832
rect 86222 30776 86278 30812
rect 86130 30164 86186 30220
rect 86222 29520 86224 29540
rect 86224 29520 86276 29540
rect 86276 29520 86278 29540
rect 86222 29484 86278 29520
rect 86222 28160 86224 28180
rect 86224 28160 86276 28180
rect 86276 28160 86278 28180
rect 86222 28124 86278 28160
rect 86222 26732 86224 26752
rect 86224 26732 86276 26752
rect 86276 26732 86278 26752
rect 86222 26696 86278 26732
rect 86222 25576 86224 25596
rect 86224 25576 86276 25596
rect 86276 25576 86278 25596
rect 86222 25540 86278 25576
rect 96380 34842 96436 34844
rect 96460 34842 96516 34844
rect 96540 34842 96596 34844
rect 96620 34842 96676 34844
rect 96380 34790 96406 34842
rect 96406 34790 96436 34842
rect 96460 34790 96470 34842
rect 96470 34790 96516 34842
rect 96540 34790 96586 34842
rect 96586 34790 96596 34842
rect 96620 34790 96650 34842
rect 96650 34790 96676 34842
rect 96380 34788 96436 34790
rect 96460 34788 96516 34790
rect 96540 34788 96596 34790
rect 96620 34788 96676 34790
rect 86222 24216 86224 24236
rect 86224 24216 86276 24236
rect 86276 24216 86278 24236
rect 86222 24180 86278 24216
rect 86038 22820 86094 22876
rect 85946 20100 86002 20156
rect 108302 23160 108358 23216
rect 86222 14832 86224 14852
rect 86224 14832 86276 14852
rect 86276 14832 86278 14852
rect 86222 14796 86278 14832
rect 56414 4800 56470 4856
rect 84014 4800 84070 4856
rect 3054 312 3110 368
<< metal3 >>
rect 0 45930 800 45960
rect 4061 45930 4127 45933
rect 0 45928 4127 45930
rect 0 45872 4066 45928
rect 4122 45872 4127 45928
rect 0 45870 4127 45872
rect 0 45840 800 45870
rect 4061 45867 4127 45870
rect 0 45386 800 45416
rect 2405 45386 2471 45389
rect 0 45384 2471 45386
rect 0 45328 2410 45384
rect 2466 45328 2471 45384
rect 0 45326 2471 45328
rect 0 45296 800 45326
rect 2405 45323 2471 45326
rect 0 44706 800 44736
rect 7649 44706 7715 44709
rect 0 44704 7715 44706
rect 0 44648 7654 44704
rect 7710 44648 7715 44704
rect 0 44646 7715 44648
rect 0 44616 800 44646
rect 7649 44643 7715 44646
rect 0 44072 800 44192
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 50288 44096 50608 44097
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 44031 50608 44032
rect 81008 44096 81328 44097
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 44031 81328 44032
rect 4208 43552 4528 43553
rect 0 43392 800 43512
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 65648 43552 65968 43553
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43487 65968 43488
rect 96368 43552 96688 43553
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43487 96688 43488
rect 19568 43008 19888 43009
rect 0 42848 800 42968
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 50288 43008 50608 43009
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 42943 50608 42944
rect 81008 43008 81328 43009
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 42943 81328 42944
rect 4208 42464 4528 42465
rect 0 42304 800 42424
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 65648 42464 65968 42465
rect 65648 42400 65656 42464
rect 65720 42400 65736 42464
rect 65800 42400 65816 42464
rect 65880 42400 65896 42464
rect 65960 42400 65968 42464
rect 65648 42399 65968 42400
rect 96368 42464 96688 42465
rect 96368 42400 96376 42464
rect 96440 42400 96456 42464
rect 96520 42400 96536 42464
rect 96600 42400 96616 42464
rect 96680 42400 96688 42464
rect 96368 42399 96688 42400
rect 17585 42394 17651 42397
rect 18045 42394 18111 42397
rect 17585 42392 18111 42394
rect 17585 42336 17590 42392
rect 17646 42336 18050 42392
rect 18106 42336 18111 42392
rect 17585 42334 18111 42336
rect 17585 42331 17651 42334
rect 18045 42331 18111 42334
rect 16389 42258 16455 42261
rect 17493 42258 17559 42261
rect 16389 42256 17559 42258
rect 16389 42200 16394 42256
rect 16450 42200 17498 42256
rect 17554 42200 17559 42256
rect 16389 42198 17559 42200
rect 16389 42195 16455 42198
rect 17493 42195 17559 42198
rect 11329 42122 11395 42125
rect 55029 42122 55095 42125
rect 11329 42120 55095 42122
rect 11329 42064 11334 42120
rect 11390 42064 55034 42120
rect 55090 42064 55095 42120
rect 11329 42062 55095 42064
rect 11329 42059 11395 42062
rect 55029 42059 55095 42062
rect 12525 41986 12591 41989
rect 17861 41986 17927 41989
rect 12525 41984 17927 41986
rect 12525 41928 12530 41984
rect 12586 41928 17866 41984
rect 17922 41928 17927 41984
rect 12525 41926 17927 41928
rect 12525 41923 12591 41926
rect 17861 41923 17927 41926
rect 51441 41986 51507 41989
rect 55949 41986 56015 41989
rect 51441 41984 56015 41986
rect 51441 41928 51446 41984
rect 51502 41928 55954 41984
rect 56010 41928 56015 41984
rect 51441 41926 56015 41928
rect 51441 41923 51507 41926
rect 55949 41923 56015 41926
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 50288 41920 50608 41921
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 41855 50608 41856
rect 81008 41920 81328 41921
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 41855 81328 41856
rect 10409 41850 10475 41853
rect 14181 41850 14247 41853
rect 10409 41848 14247 41850
rect 10409 41792 10414 41848
rect 10470 41792 14186 41848
rect 14242 41792 14247 41848
rect 10409 41790 14247 41792
rect 10409 41787 10475 41790
rect 14181 41787 14247 41790
rect 0 41714 800 41744
rect 3969 41714 4035 41717
rect 0 41712 4035 41714
rect 0 41656 3974 41712
rect 4030 41656 4035 41712
rect 0 41654 4035 41656
rect 0 41624 800 41654
rect 3969 41651 4035 41654
rect 37273 41714 37339 41717
rect 38653 41714 38719 41717
rect 37273 41712 38719 41714
rect 37273 41656 37278 41712
rect 37334 41656 38658 41712
rect 38714 41656 38719 41712
rect 37273 41654 38719 41656
rect 37273 41651 37339 41654
rect 38653 41651 38719 41654
rect 44633 41578 44699 41581
rect 45921 41578 45987 41581
rect 44633 41576 45987 41578
rect 44633 41520 44638 41576
rect 44694 41520 45926 41576
rect 45982 41520 45987 41576
rect 44633 41518 45987 41520
rect 44633 41515 44699 41518
rect 45921 41515 45987 41518
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 65648 41376 65968 41377
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 41311 65968 41312
rect 96368 41376 96688 41377
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 41311 96688 41312
rect 0 41170 800 41200
rect 6913 41170 6979 41173
rect 0 41168 6979 41170
rect 0 41112 6918 41168
rect 6974 41112 6979 41168
rect 0 41110 6979 41112
rect 0 41080 800 41110
rect 6913 41107 6979 41110
rect 29821 41170 29887 41173
rect 30649 41170 30715 41173
rect 29821 41168 30715 41170
rect 29821 41112 29826 41168
rect 29882 41112 30654 41168
rect 30710 41112 30715 41168
rect 29821 41110 30715 41112
rect 29821 41107 29887 41110
rect 30649 41107 30715 41110
rect 60641 41170 60707 41173
rect 63125 41170 63191 41173
rect 60641 41168 63191 41170
rect 60641 41112 60646 41168
rect 60702 41112 63130 41168
rect 63186 41112 63191 41168
rect 60641 41110 63191 41112
rect 60641 41107 60707 41110
rect 63125 41107 63191 41110
rect 38653 41034 38719 41037
rect 39021 41034 39087 41037
rect 38653 41032 39087 41034
rect 38653 40976 38658 41032
rect 38714 40976 39026 41032
rect 39082 40976 39087 41032
rect 38653 40974 39087 40976
rect 38653 40971 38719 40974
rect 39021 40971 39087 40974
rect 39021 40898 39087 40901
rect 46289 40898 46355 40901
rect 39021 40896 46355 40898
rect 39021 40840 39026 40896
rect 39082 40840 46294 40896
rect 46350 40840 46355 40896
rect 39021 40838 46355 40840
rect 39021 40835 39087 40838
rect 46289 40835 46355 40838
rect 53373 40898 53439 40901
rect 57237 40898 57303 40901
rect 53373 40896 57303 40898
rect 53373 40840 53378 40896
rect 53434 40840 57242 40896
rect 57298 40840 57303 40896
rect 53373 40838 57303 40840
rect 53373 40835 53439 40838
rect 57237 40835 57303 40838
rect 58801 40898 58867 40901
rect 64321 40898 64387 40901
rect 58801 40896 64387 40898
rect 58801 40840 58806 40896
rect 58862 40840 64326 40896
rect 64382 40840 64387 40896
rect 58801 40838 64387 40840
rect 58801 40835 58867 40838
rect 64321 40835 64387 40838
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 50288 40832 50608 40833
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 40767 50608 40768
rect 81008 40832 81328 40833
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 40767 81328 40768
rect 24761 40762 24827 40765
rect 34605 40762 34671 40765
rect 24761 40760 34671 40762
rect 24761 40704 24766 40760
rect 24822 40704 34610 40760
rect 34666 40704 34671 40760
rect 24761 40702 34671 40704
rect 24761 40699 24827 40702
rect 34605 40699 34671 40702
rect 0 40490 800 40520
rect 3417 40490 3483 40493
rect 0 40488 3483 40490
rect 0 40432 3422 40488
rect 3478 40432 3483 40488
rect 0 40430 3483 40432
rect 0 40400 800 40430
rect 3417 40427 3483 40430
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 65648 40288 65968 40289
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 40223 65968 40224
rect 96368 40288 96688 40289
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 40223 96688 40224
rect 68461 40082 68527 40085
rect 71405 40082 71471 40085
rect 68461 40080 71471 40082
rect 68461 40024 68466 40080
rect 68522 40024 71410 40080
rect 71466 40024 71471 40080
rect 68461 40022 71471 40024
rect 68461 40019 68527 40022
rect 71405 40019 71471 40022
rect 0 39946 800 39976
rect 4061 39946 4127 39949
rect 0 39944 4127 39946
rect 0 39888 4066 39944
rect 4122 39888 4127 39944
rect 0 39886 4127 39888
rect 0 39856 800 39886
rect 4061 39883 4127 39886
rect 32213 39946 32279 39949
rect 72601 39946 72667 39949
rect 32213 39944 72667 39946
rect 32213 39888 32218 39944
rect 32274 39888 72606 39944
rect 72662 39888 72667 39944
rect 32213 39886 72667 39888
rect 32213 39883 32279 39886
rect 72601 39883 72667 39886
rect 28257 39810 28323 39813
rect 48589 39810 48655 39813
rect 28257 39808 48655 39810
rect 28257 39752 28262 39808
rect 28318 39752 48594 39808
rect 48650 39752 48655 39808
rect 28257 39750 48655 39752
rect 28257 39747 28323 39750
rect 48589 39747 48655 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 50288 39744 50608 39745
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 39679 50608 39680
rect 81008 39744 81328 39745
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 39679 81328 39680
rect 38101 39674 38167 39677
rect 48129 39674 48195 39677
rect 38101 39672 48195 39674
rect 38101 39616 38106 39672
rect 38162 39616 48134 39672
rect 48190 39616 48195 39672
rect 38101 39614 48195 39616
rect 38101 39611 38167 39614
rect 48129 39611 48195 39614
rect 31017 39538 31083 39541
rect 35065 39538 35131 39541
rect 31017 39536 35131 39538
rect 31017 39480 31022 39536
rect 31078 39480 35070 39536
rect 35126 39480 35131 39536
rect 31017 39478 35131 39480
rect 31017 39475 31083 39478
rect 35065 39475 35131 39478
rect 41137 39538 41203 39541
rect 42241 39538 42307 39541
rect 41137 39536 42307 39538
rect 41137 39480 41142 39536
rect 41198 39480 42246 39536
rect 42302 39480 42307 39536
rect 41137 39478 42307 39480
rect 41137 39475 41203 39478
rect 42241 39475 42307 39478
rect 51993 39538 52059 39541
rect 54569 39538 54635 39541
rect 51993 39536 54635 39538
rect 51993 39480 51998 39536
rect 52054 39480 54574 39536
rect 54630 39480 54635 39536
rect 51993 39478 54635 39480
rect 51993 39475 52059 39478
rect 54569 39475 54635 39478
rect 62205 39538 62271 39541
rect 63585 39538 63651 39541
rect 64597 39538 64663 39541
rect 62205 39536 64663 39538
rect 62205 39480 62210 39536
rect 62266 39480 63590 39536
rect 63646 39480 64602 39536
rect 64658 39480 64663 39536
rect 62205 39478 64663 39480
rect 62205 39475 62271 39478
rect 63585 39475 63651 39478
rect 64597 39475 64663 39478
rect 0 39402 800 39432
rect 3969 39402 4035 39405
rect 0 39400 4035 39402
rect 0 39344 3974 39400
rect 4030 39344 4035 39400
rect 0 39342 4035 39344
rect 0 39312 800 39342
rect 3969 39339 4035 39342
rect 27245 39402 27311 39405
rect 43529 39402 43595 39405
rect 27245 39400 43595 39402
rect 27245 39344 27250 39400
rect 27306 39344 43534 39400
rect 43590 39344 43595 39400
rect 27245 39342 43595 39344
rect 27245 39339 27311 39342
rect 43529 39339 43595 39342
rect 43989 39402 44055 39405
rect 44633 39402 44699 39405
rect 43989 39400 44699 39402
rect 43989 39344 43994 39400
rect 44050 39344 44638 39400
rect 44694 39344 44699 39400
rect 43989 39342 44699 39344
rect 43989 39339 44055 39342
rect 44633 39339 44699 39342
rect 48773 39402 48839 39405
rect 56133 39402 56199 39405
rect 48773 39400 56199 39402
rect 48773 39344 48778 39400
rect 48834 39344 56138 39400
rect 56194 39344 56199 39400
rect 48773 39342 56199 39344
rect 48773 39339 48839 39342
rect 56133 39339 56199 39342
rect 61929 39402 61995 39405
rect 66529 39402 66595 39405
rect 61929 39400 66595 39402
rect 61929 39344 61934 39400
rect 61990 39344 66534 39400
rect 66590 39344 66595 39400
rect 61929 39342 66595 39344
rect 61929 39339 61995 39342
rect 66529 39339 66595 39342
rect 78029 39402 78095 39405
rect 83733 39402 83799 39405
rect 78029 39400 83799 39402
rect 78029 39344 78034 39400
rect 78090 39344 83738 39400
rect 83794 39344 83799 39400
rect 78029 39342 83799 39344
rect 78029 39339 78095 39342
rect 83733 39339 83799 39342
rect 41045 39266 41111 39269
rect 42333 39266 42399 39269
rect 41045 39264 42399 39266
rect 41045 39208 41050 39264
rect 41106 39208 42338 39264
rect 42394 39208 42399 39264
rect 41045 39206 42399 39208
rect 41045 39203 41111 39206
rect 42333 39203 42399 39206
rect 43253 39266 43319 39269
rect 44173 39266 44239 39269
rect 43253 39264 44239 39266
rect 43253 39208 43258 39264
rect 43314 39208 44178 39264
rect 44234 39208 44239 39264
rect 43253 39206 44239 39208
rect 43253 39203 43319 39206
rect 44173 39203 44239 39206
rect 48681 39266 48747 39269
rect 56225 39266 56291 39269
rect 48681 39264 56291 39266
rect 48681 39208 48686 39264
rect 48742 39208 56230 39264
rect 56286 39208 56291 39264
rect 48681 39206 56291 39208
rect 48681 39203 48747 39206
rect 56225 39203 56291 39206
rect 78949 39266 79015 39269
rect 80697 39266 80763 39269
rect 78949 39264 80763 39266
rect 78949 39208 78954 39264
rect 79010 39208 80702 39264
rect 80758 39208 80763 39264
rect 78949 39206 80763 39208
rect 78949 39203 79015 39206
rect 80697 39203 80763 39206
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 65648 39200 65968 39201
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 39135 65968 39136
rect 96368 39200 96688 39201
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 39135 96688 39136
rect 40861 39130 40927 39133
rect 44449 39130 44515 39133
rect 40861 39128 44515 39130
rect 40861 39072 40866 39128
rect 40922 39072 44454 39128
rect 44510 39072 44515 39128
rect 40861 39070 44515 39072
rect 40861 39067 40927 39070
rect 44449 39067 44515 39070
rect 79133 39130 79199 39133
rect 80421 39130 80487 39133
rect 79133 39128 80487 39130
rect 79133 39072 79138 39128
rect 79194 39072 80426 39128
rect 80482 39072 80487 39128
rect 79133 39070 80487 39072
rect 79133 39067 79199 39070
rect 80421 39067 80487 39070
rect 40953 38994 41019 38997
rect 42977 38994 43043 38997
rect 40953 38992 43043 38994
rect 40953 38936 40958 38992
rect 41014 38936 42982 38992
rect 43038 38936 43043 38992
rect 40953 38934 43043 38936
rect 40953 38931 41019 38934
rect 42977 38931 43043 38934
rect 47393 38994 47459 38997
rect 48681 38994 48747 38997
rect 53281 38994 53347 38997
rect 47393 38992 53347 38994
rect 47393 38936 47398 38992
rect 47454 38936 48686 38992
rect 48742 38936 53286 38992
rect 53342 38936 53347 38992
rect 47393 38934 53347 38936
rect 47393 38931 47459 38934
rect 48681 38931 48747 38934
rect 53281 38931 53347 38934
rect 68553 38994 68619 38997
rect 69105 38994 69171 38997
rect 75729 38994 75795 38997
rect 68553 38992 75795 38994
rect 68553 38936 68558 38992
rect 68614 38936 69110 38992
rect 69166 38936 75734 38992
rect 75790 38936 75795 38992
rect 68553 38934 75795 38936
rect 68553 38931 68619 38934
rect 69105 38931 69171 38934
rect 75729 38931 75795 38934
rect 77569 38994 77635 38997
rect 79593 38994 79659 38997
rect 77569 38992 79659 38994
rect 77569 38936 77574 38992
rect 77630 38936 79598 38992
rect 79654 38936 79659 38992
rect 77569 38934 79659 38936
rect 77569 38931 77635 38934
rect 79593 38931 79659 38934
rect 79777 38994 79843 38997
rect 82905 38994 82971 38997
rect 79777 38992 82971 38994
rect 79777 38936 79782 38992
rect 79838 38936 82910 38992
rect 82966 38936 82971 38992
rect 79777 38934 82971 38936
rect 79777 38931 79843 38934
rect 82905 38931 82971 38934
rect 23841 38858 23907 38861
rect 25221 38858 25287 38861
rect 26693 38858 26759 38861
rect 23841 38856 26759 38858
rect 23841 38800 23846 38856
rect 23902 38800 25226 38856
rect 25282 38800 26698 38856
rect 26754 38800 26759 38856
rect 23841 38798 26759 38800
rect 23841 38795 23907 38798
rect 25221 38795 25287 38798
rect 26693 38795 26759 38798
rect 47853 38858 47919 38861
rect 55765 38858 55831 38861
rect 47853 38856 55831 38858
rect 47853 38800 47858 38856
rect 47914 38800 55770 38856
rect 55826 38800 55831 38856
rect 47853 38798 55831 38800
rect 47853 38795 47919 38798
rect 55765 38795 55831 38798
rect 68461 38858 68527 38861
rect 69473 38858 69539 38861
rect 68461 38856 69539 38858
rect 68461 38800 68466 38856
rect 68522 38800 69478 38856
rect 69534 38800 69539 38856
rect 68461 38798 69539 38800
rect 68461 38795 68527 38798
rect 69473 38795 69539 38798
rect 79409 38858 79475 38861
rect 80513 38858 80579 38861
rect 79409 38856 80579 38858
rect 79409 38800 79414 38856
rect 79470 38800 80518 38856
rect 80574 38800 80579 38856
rect 79409 38798 80579 38800
rect 79409 38795 79475 38798
rect 80513 38795 80579 38798
rect 0 38722 800 38752
rect 4061 38722 4127 38725
rect 0 38720 4127 38722
rect 0 38664 4066 38720
rect 4122 38664 4127 38720
rect 0 38662 4127 38664
rect 0 38632 800 38662
rect 4061 38659 4127 38662
rect 15009 38722 15075 38725
rect 15469 38722 15535 38725
rect 15009 38720 15535 38722
rect 15009 38664 15014 38720
rect 15070 38664 15474 38720
rect 15530 38664 15535 38720
rect 15009 38662 15535 38664
rect 15009 38659 15075 38662
rect 15469 38659 15535 38662
rect 23933 38722 23999 38725
rect 24577 38722 24643 38725
rect 26785 38722 26851 38725
rect 23933 38720 26851 38722
rect 23933 38664 23938 38720
rect 23994 38664 24582 38720
rect 24638 38664 26790 38720
rect 26846 38664 26851 38720
rect 23933 38662 26851 38664
rect 23933 38659 23999 38662
rect 24577 38659 24643 38662
rect 26785 38659 26851 38662
rect 43253 38722 43319 38725
rect 48037 38722 48103 38725
rect 43253 38720 48103 38722
rect 43253 38664 43258 38720
rect 43314 38664 48042 38720
rect 48098 38664 48103 38720
rect 43253 38662 48103 38664
rect 43253 38659 43319 38662
rect 48037 38659 48103 38662
rect 68737 38722 68803 38725
rect 76281 38722 76347 38725
rect 68737 38720 76347 38722
rect 68737 38664 68742 38720
rect 68798 38664 76286 38720
rect 76342 38664 76347 38720
rect 68737 38662 76347 38664
rect 68737 38659 68803 38662
rect 76281 38659 76347 38662
rect 77569 38722 77635 38725
rect 78213 38722 78279 38725
rect 77569 38720 78279 38722
rect 77569 38664 77574 38720
rect 77630 38664 78218 38720
rect 78274 38664 78279 38720
rect 77569 38662 78279 38664
rect 77569 38659 77635 38662
rect 78213 38659 78279 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 50288 38656 50608 38657
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 38591 50608 38592
rect 81008 38656 81328 38657
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 38591 81328 38592
rect 21173 38586 21239 38589
rect 25865 38586 25931 38589
rect 27521 38586 27587 38589
rect 21173 38584 25931 38586
rect 21173 38528 21178 38584
rect 21234 38528 25870 38584
rect 25926 38528 25931 38584
rect 21173 38526 25931 38528
rect 21173 38523 21239 38526
rect 25865 38523 25931 38526
rect 26006 38584 27587 38586
rect 26006 38528 27526 38584
rect 27582 38528 27587 38584
rect 26006 38526 27587 38528
rect 19241 38450 19307 38453
rect 26006 38450 26066 38526
rect 27521 38523 27587 38526
rect 36537 38586 36603 38589
rect 37089 38586 37155 38589
rect 36537 38584 37155 38586
rect 36537 38528 36542 38584
rect 36598 38528 37094 38584
rect 37150 38528 37155 38584
rect 36537 38526 37155 38528
rect 36537 38523 36603 38526
rect 37089 38523 37155 38526
rect 19241 38448 26066 38450
rect 19241 38392 19246 38448
rect 19302 38392 26066 38448
rect 19241 38390 26066 38392
rect 30649 38450 30715 38453
rect 37733 38450 37799 38453
rect 30649 38448 37799 38450
rect 30649 38392 30654 38448
rect 30710 38392 37738 38448
rect 37794 38392 37799 38448
rect 30649 38390 37799 38392
rect 19241 38387 19307 38390
rect 30649 38387 30715 38390
rect 37733 38387 37799 38390
rect 38837 38314 38903 38317
rect 46105 38314 46171 38317
rect 38837 38312 46171 38314
rect 38837 38256 38842 38312
rect 38898 38256 46110 38312
rect 46166 38256 46171 38312
rect 38837 38254 46171 38256
rect 38837 38251 38903 38254
rect 46105 38251 46171 38254
rect 0 38178 800 38208
rect 4061 38178 4127 38181
rect 0 38176 4127 38178
rect 0 38120 4066 38176
rect 4122 38120 4127 38176
rect 0 38118 4127 38120
rect 0 38088 800 38118
rect 4061 38115 4127 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 65648 38112 65968 38113
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 38047 65968 38048
rect 96368 38112 96688 38113
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 38047 96688 38048
rect 15929 37770 15995 37773
rect 16573 37770 16639 37773
rect 15929 37768 16639 37770
rect 15929 37712 15934 37768
rect 15990 37712 16578 37768
rect 16634 37712 16639 37768
rect 15929 37710 16639 37712
rect 15929 37707 15995 37710
rect 16573 37707 16639 37710
rect 35617 37770 35683 37773
rect 36537 37770 36603 37773
rect 35617 37768 36603 37770
rect 35617 37712 35622 37768
rect 35678 37712 36542 37768
rect 36598 37712 36603 37768
rect 35617 37710 36603 37712
rect 35617 37707 35683 37710
rect 36537 37707 36603 37710
rect 42609 37634 42675 37637
rect 43437 37634 43503 37637
rect 51901 37634 51967 37637
rect 57237 37634 57303 37637
rect 42609 37632 50170 37634
rect 42609 37576 42614 37632
rect 42670 37576 43442 37632
rect 43498 37576 50170 37632
rect 42609 37574 50170 37576
rect 42609 37571 42675 37574
rect 43437 37571 43503 37574
rect 19568 37568 19888 37569
rect 0 37498 800 37528
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 3693 37498 3759 37501
rect 0 37496 3759 37498
rect 0 37440 3698 37496
rect 3754 37440 3759 37496
rect 0 37438 3759 37440
rect 0 37408 800 37438
rect 3693 37435 3759 37438
rect 29085 37498 29151 37501
rect 38285 37498 38351 37501
rect 29085 37496 38351 37498
rect 29085 37440 29090 37496
rect 29146 37440 38290 37496
rect 38346 37440 38351 37496
rect 29085 37438 38351 37440
rect 29085 37435 29151 37438
rect 38285 37435 38351 37438
rect 50110 37362 50170 37574
rect 51901 37632 57303 37634
rect 51901 37576 51906 37632
rect 51962 37576 57242 37632
rect 57298 37576 57303 37632
rect 51901 37574 57303 37576
rect 51901 37571 51967 37574
rect 57237 37571 57303 37574
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 81008 37568 81328 37569
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 37503 81328 37504
rect 57053 37498 57119 37501
rect 57789 37498 57855 37501
rect 57053 37496 57855 37498
rect 57053 37440 57058 37496
rect 57114 37440 57794 37496
rect 57850 37440 57855 37496
rect 57053 37438 57855 37440
rect 57053 37435 57119 37438
rect 57789 37435 57855 37438
rect 57145 37362 57211 37365
rect 50110 37360 57211 37362
rect 50110 37304 57150 37360
rect 57206 37304 57211 37360
rect 50110 37302 57211 37304
rect 57145 37299 57211 37302
rect 50981 37226 51047 37229
rect 55673 37226 55739 37229
rect 50981 37224 55739 37226
rect 50981 37168 50986 37224
rect 51042 37168 55678 37224
rect 55734 37168 55739 37224
rect 50981 37166 55739 37168
rect 50981 37163 51047 37166
rect 55673 37163 55739 37166
rect 4208 37024 4528 37025
rect 0 36954 800 36984
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 65648 37024 65968 37025
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 36959 65968 36960
rect 96368 37024 96688 37025
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 36959 96688 36960
rect 4061 36954 4127 36957
rect 0 36952 4127 36954
rect 0 36896 4066 36952
rect 4122 36896 4127 36952
rect 0 36894 4127 36896
rect 0 36864 800 36894
rect 4061 36891 4127 36894
rect 41321 36954 41387 36957
rect 47301 36954 47367 36957
rect 41321 36952 47367 36954
rect 41321 36896 41326 36952
rect 41382 36896 47306 36952
rect 47362 36896 47367 36952
rect 41321 36894 47367 36896
rect 41321 36891 41387 36894
rect 47301 36891 47367 36894
rect 70945 36818 71011 36821
rect 71957 36818 72023 36821
rect 70945 36816 72023 36818
rect 70945 36760 70950 36816
rect 71006 36760 71962 36816
rect 72018 36760 72023 36816
rect 70945 36758 72023 36760
rect 70945 36755 71011 36758
rect 71957 36755 72023 36758
rect 17902 36620 17908 36684
rect 17972 36682 17978 36684
rect 50797 36682 50863 36685
rect 54201 36682 54267 36685
rect 17972 36622 20178 36682
rect 17972 36620 17978 36622
rect 20118 36546 20178 36622
rect 50797 36680 54267 36682
rect 50797 36624 50802 36680
rect 50858 36624 54206 36680
rect 54262 36624 54267 36680
rect 50797 36622 54267 36624
rect 50797 36619 50863 36622
rect 54201 36619 54267 36622
rect 26182 36546 26188 36548
rect 20118 36486 26188 36546
rect 26182 36484 26188 36486
rect 26252 36484 26258 36548
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 81008 36480 81328 36481
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 36415 81328 36416
rect 33685 36410 33751 36413
rect 35985 36410 36051 36413
rect 33685 36408 36051 36410
rect 33685 36352 33690 36408
rect 33746 36352 35990 36408
rect 36046 36352 36051 36408
rect 33685 36350 36051 36352
rect 33685 36347 33751 36350
rect 35985 36347 36051 36350
rect 0 36274 800 36304
rect 3509 36274 3575 36277
rect 17902 36274 17908 36276
rect 0 36272 3575 36274
rect 0 36216 3514 36272
rect 3570 36216 3575 36272
rect 0 36214 3575 36216
rect 0 36184 800 36214
rect 3509 36211 3575 36214
rect 9814 36214 17908 36274
rect 9814 36172 9874 36214
rect 17902 36212 17908 36214
rect 17972 36212 17978 36276
rect 26182 36212 26188 36276
rect 26252 36274 26258 36276
rect 35893 36274 35959 36277
rect 26252 36272 35959 36274
rect 26252 36216 35898 36272
rect 35954 36216 35959 36272
rect 26252 36214 35959 36216
rect 26252 36212 26258 36214
rect 35893 36211 35959 36214
rect 37549 36274 37615 36277
rect 46013 36274 46079 36277
rect 37549 36272 46079 36274
rect 37549 36216 37554 36272
rect 37610 36216 46018 36272
rect 46074 36216 46079 36272
rect 37549 36214 46079 36216
rect 37549 36211 37615 36214
rect 46013 36211 46079 36214
rect 49785 36274 49851 36277
rect 51625 36274 51691 36277
rect 49785 36272 51691 36274
rect 49785 36216 49790 36272
rect 49846 36216 51630 36272
rect 51686 36216 51691 36272
rect 49785 36214 51691 36216
rect 49785 36211 49851 36214
rect 51625 36211 51691 36214
rect 3325 36138 3391 36141
rect 9630 36138 9874 36172
rect 3325 36136 9874 36138
rect 3325 36080 3330 36136
rect 3386 36112 9874 36136
rect 43529 36138 43595 36141
rect 44909 36138 44975 36141
rect 43529 36136 44975 36138
rect 3386 36080 9690 36112
rect 3325 36078 9690 36080
rect 43529 36080 43534 36136
rect 43590 36080 44914 36136
rect 44970 36080 44975 36136
rect 43529 36078 44975 36080
rect 3325 36075 3391 36078
rect 43529 36075 43595 36078
rect 44909 36075 44975 36078
rect 38653 36002 38719 36005
rect 45829 36002 45895 36005
rect 38653 36000 45895 36002
rect 38653 35944 38658 36000
rect 38714 35944 45834 36000
rect 45890 35944 45895 36000
rect 38653 35942 45895 35944
rect 38653 35939 38719 35942
rect 45829 35939 45895 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 65648 35936 65968 35937
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 35871 65968 35872
rect 96368 35936 96688 35937
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 35871 96688 35872
rect 39941 35866 40007 35869
rect 42517 35866 42583 35869
rect 39941 35864 42583 35866
rect 39941 35808 39946 35864
rect 40002 35808 42522 35864
rect 42578 35808 42583 35864
rect 39941 35806 42583 35808
rect 39941 35803 40007 35806
rect 42517 35803 42583 35806
rect 0 35730 800 35760
rect 4061 35730 4127 35733
rect 0 35728 4127 35730
rect 0 35672 4066 35728
rect 4122 35672 4127 35728
rect 0 35670 4127 35672
rect 0 35640 800 35670
rect 4061 35667 4127 35670
rect 38377 35730 38443 35733
rect 40861 35730 40927 35733
rect 38377 35728 40927 35730
rect 38377 35672 38382 35728
rect 38438 35672 40866 35728
rect 40922 35672 40927 35728
rect 38377 35670 40927 35672
rect 38377 35667 38443 35670
rect 40861 35667 40927 35670
rect 82721 35458 82787 35461
rect 83273 35458 83339 35461
rect 82721 35456 83339 35458
rect 82721 35400 82726 35456
rect 82782 35400 83278 35456
rect 83334 35400 83339 35456
rect 82721 35398 83339 35400
rect 82721 35395 82787 35398
rect 83273 35395 83339 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 81008 35392 81328 35393
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 35327 81328 35328
rect 41229 35322 41295 35325
rect 41505 35322 41571 35325
rect 41229 35320 41571 35322
rect 41229 35264 41234 35320
rect 41290 35264 41510 35320
rect 41566 35264 41571 35320
rect 41229 35262 41571 35264
rect 41229 35259 41295 35262
rect 41505 35259 41571 35262
rect 0 35186 800 35216
rect 5625 35186 5691 35189
rect 0 35184 5691 35186
rect 0 35128 5630 35184
rect 5686 35128 5691 35184
rect 0 35126 5691 35128
rect 0 35096 800 35126
rect 5625 35123 5691 35126
rect 28901 35186 28967 35189
rect 40217 35186 40283 35189
rect 28901 35184 40283 35186
rect 28901 35128 28906 35184
rect 28962 35128 40222 35184
rect 40278 35128 40283 35184
rect 28901 35126 40283 35128
rect 28901 35123 28967 35126
rect 40217 35123 40283 35126
rect 40677 35186 40743 35189
rect 41413 35186 41479 35189
rect 42241 35186 42307 35189
rect 40677 35184 42307 35186
rect 40677 35128 40682 35184
rect 40738 35128 41418 35184
rect 41474 35128 42246 35184
rect 42302 35128 42307 35184
rect 40677 35126 42307 35128
rect 40677 35123 40743 35126
rect 41413 35123 41479 35126
rect 42241 35123 42307 35126
rect 49141 35186 49207 35189
rect 50429 35186 50495 35189
rect 51257 35186 51323 35189
rect 49141 35184 51323 35186
rect 49141 35128 49146 35184
rect 49202 35128 50434 35184
rect 50490 35128 51262 35184
rect 51318 35128 51323 35184
rect 49141 35126 51323 35128
rect 49141 35123 49207 35126
rect 50429 35123 50495 35126
rect 51257 35123 51323 35126
rect 69289 35186 69355 35189
rect 71313 35186 71379 35189
rect 69289 35184 71379 35186
rect 69289 35128 69294 35184
rect 69350 35128 71318 35184
rect 71374 35128 71379 35184
rect 69289 35126 71379 35128
rect 69289 35123 69355 35126
rect 71313 35123 71379 35126
rect 48957 35050 49023 35053
rect 52637 35050 52703 35053
rect 48957 35048 52703 35050
rect 48957 34992 48962 35048
rect 49018 34992 52642 35048
rect 52698 34992 52703 35048
rect 48957 34990 52703 34992
rect 48957 34987 49023 34990
rect 52637 34987 52703 34990
rect 55949 35050 56015 35053
rect 63033 35050 63099 35053
rect 55949 35048 63099 35050
rect 55949 34992 55954 35048
rect 56010 34992 63038 35048
rect 63094 34992 63099 35048
rect 55949 34990 63099 34992
rect 55949 34987 56015 34990
rect 63033 34987 63099 34990
rect 61745 34914 61811 34917
rect 64689 34914 64755 34917
rect 61745 34912 64755 34914
rect 61745 34856 61750 34912
rect 61806 34856 64694 34912
rect 64750 34856 64755 34912
rect 61745 34854 64755 34856
rect 61745 34851 61811 34854
rect 64689 34851 64755 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 65648 34848 65968 34849
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 34783 65968 34784
rect 96368 34848 96688 34849
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 34783 96688 34784
rect 27797 34778 27863 34781
rect 29545 34778 29611 34781
rect 27797 34776 29611 34778
rect 27797 34720 27802 34776
rect 27858 34720 29550 34776
rect 29606 34720 29611 34776
rect 27797 34718 29611 34720
rect 27797 34715 27863 34718
rect 29545 34715 29611 34718
rect 49417 34778 49483 34781
rect 50245 34778 50311 34781
rect 57053 34778 57119 34781
rect 49417 34776 57119 34778
rect 49417 34720 49422 34776
rect 49478 34720 50250 34776
rect 50306 34720 57058 34776
rect 57114 34720 57119 34776
rect 49417 34718 57119 34720
rect 49417 34715 49483 34718
rect 50245 34715 50311 34718
rect 57053 34715 57119 34718
rect 28717 34642 28783 34645
rect 46657 34642 46723 34645
rect 28717 34640 46723 34642
rect 28717 34584 28722 34640
rect 28778 34584 46662 34640
rect 46718 34584 46723 34640
rect 28717 34582 46723 34584
rect 28717 34579 28783 34582
rect 46657 34579 46723 34582
rect 49785 34642 49851 34645
rect 56777 34642 56843 34645
rect 49785 34640 56843 34642
rect 49785 34584 49790 34640
rect 49846 34584 56782 34640
rect 56838 34584 56843 34640
rect 49785 34582 56843 34584
rect 49785 34579 49851 34582
rect 56777 34579 56843 34582
rect 58617 34642 58683 34645
rect 62297 34642 62363 34645
rect 58617 34640 62363 34642
rect 58617 34584 58622 34640
rect 58678 34584 62302 34640
rect 62358 34584 62363 34640
rect 58617 34582 62363 34584
rect 58617 34579 58683 34582
rect 62297 34579 62363 34582
rect 0 34506 800 34536
rect 4061 34506 4127 34509
rect 0 34504 4127 34506
rect 0 34448 4066 34504
rect 4122 34448 4127 34504
rect 0 34446 4127 34448
rect 0 34416 800 34446
rect 4061 34443 4127 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 81008 34304 81328 34305
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 34239 81328 34240
rect 0 33962 800 33992
rect 4061 33962 4127 33965
rect 0 33960 4127 33962
rect 0 33904 4066 33960
rect 4122 33904 4127 33960
rect 0 33902 4127 33904
rect 0 33872 800 33902
rect 4061 33899 4127 33902
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 0 33282 800 33312
rect 3969 33282 4035 33285
rect 0 33280 4035 33282
rect 0 33224 3974 33280
rect 4030 33224 4035 33280
rect 0 33222 4035 33224
rect 0 33192 800 33222
rect 3969 33219 4035 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 0 32738 800 32768
rect 3233 32738 3299 32741
rect 0 32736 3299 32738
rect 0 32680 3238 32736
rect 3294 32680 3299 32736
rect 0 32678 3299 32680
rect 0 32648 800 32678
rect 3233 32675 3299 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 13537 32602 13603 32605
rect 13905 32602 13971 32605
rect 18965 32602 19031 32605
rect 13537 32600 19031 32602
rect 13537 32544 13542 32600
rect 13598 32544 13910 32600
rect 13966 32544 18970 32600
rect 19026 32544 19031 32600
rect 13537 32542 19031 32544
rect 13537 32539 13603 32542
rect 13905 32539 13971 32542
rect 18965 32539 19031 32542
rect 19517 32330 19583 32333
rect 24761 32330 24827 32333
rect 19517 32328 24827 32330
rect 19517 32272 19522 32328
rect 19578 32272 24766 32328
rect 24822 32272 24827 32328
rect 19517 32270 24827 32272
rect 19517 32267 19583 32270
rect 24761 32267 24827 32270
rect 0 32194 800 32224
rect 4061 32194 4127 32197
rect 0 32192 4127 32194
rect 0 32136 4066 32192
rect 4122 32136 4127 32192
rect 0 32134 4127 32136
rect 0 32104 800 32134
rect 4061 32131 4127 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 12709 32058 12775 32061
rect 18045 32058 18111 32061
rect 12709 32056 18111 32058
rect 12709 32000 12714 32056
rect 12770 32000 18050 32056
rect 18106 32000 18111 32056
rect 12709 31998 18111 32000
rect 12709 31995 12775 31998
rect 18045 31995 18111 31998
rect 19701 31922 19767 31925
rect 25681 31922 25747 31925
rect 19701 31920 25747 31922
rect 19701 31864 19706 31920
rect 19762 31864 25686 31920
rect 25742 31864 25747 31920
rect 19701 31862 25747 31864
rect 19701 31859 19767 31862
rect 25681 31859 25747 31862
rect 12709 31786 12775 31789
rect 13813 31786 13879 31789
rect 27613 31786 27679 31789
rect 12709 31784 27679 31786
rect 12709 31728 12714 31784
rect 12770 31728 13818 31784
rect 13874 31728 27618 31784
rect 27674 31728 27679 31784
rect 12709 31726 27679 31728
rect 12709 31723 12775 31726
rect 13813 31723 13879 31726
rect 27613 31723 27679 31726
rect 4208 31584 4528 31585
rect 0 31514 800 31544
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 3785 31514 3851 31517
rect 0 31512 3851 31514
rect 0 31456 3790 31512
rect 3846 31456 3851 31512
rect 0 31454 3851 31456
rect 0 31424 800 31454
rect 3785 31451 3851 31454
rect 9765 31514 9831 31517
rect 19241 31514 19307 31517
rect 9765 31512 19307 31514
rect 9765 31456 9770 31512
rect 9826 31456 19246 31512
rect 19302 31456 19307 31512
rect 9765 31454 19307 31456
rect 9765 31451 9831 31454
rect 19241 31451 19307 31454
rect 56593 31242 56659 31245
rect 56869 31242 56935 31245
rect 56593 31240 56935 31242
rect 56593 31184 56598 31240
rect 56654 31184 56874 31240
rect 56930 31184 56935 31240
rect 56593 31182 56935 31184
rect 56593 31179 56659 31182
rect 56869 31179 56935 31182
rect 19568 31040 19888 31041
rect 0 30970 800 31000
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 3969 30970 4035 30973
rect 0 30968 4035 30970
rect 0 30912 3974 30968
rect 4030 30912 4035 30968
rect 0 30910 4035 30912
rect 0 30880 800 30910
rect 3969 30907 4035 30910
rect 20345 30970 20411 30973
rect 27521 30970 27587 30973
rect 20345 30968 27587 30970
rect 20345 30912 20350 30968
rect 20406 30912 27526 30968
rect 27582 30912 27587 30968
rect 20345 30910 27587 30912
rect 20345 30907 20411 30910
rect 27521 30907 27587 30910
rect 29637 30834 29703 30837
rect 56317 30834 56383 30837
rect 86217 30834 86283 30837
rect 29637 30832 32108 30834
rect 29637 30776 29642 30832
rect 29698 30776 32108 30832
rect 29637 30774 32108 30776
rect 56317 30832 58604 30834
rect 56317 30776 56322 30832
rect 56378 30776 58604 30832
rect 56317 30774 58604 30776
rect 86217 30832 86388 30834
rect 86217 30776 86222 30832
rect 86278 30776 86388 30832
rect 86217 30774 86388 30776
rect 29637 30771 29703 30774
rect 56317 30771 56383 30774
rect 86217 30771 86283 30774
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 0 30290 800 30320
rect 3601 30290 3667 30293
rect 0 30288 3667 30290
rect 0 30232 3606 30288
rect 3662 30232 3667 30288
rect 0 30230 3667 30232
rect 0 30200 800 30230
rect 3601 30227 3667 30230
rect 86125 30222 86191 30225
rect 86125 30220 86388 30222
rect 86125 30164 86130 30220
rect 86186 30164 86388 30220
rect 86125 30162 86388 30164
rect 86125 30159 86191 30162
rect 14457 30154 14523 30157
rect 18321 30154 18387 30157
rect 14457 30152 18387 30154
rect 14457 30096 14462 30152
rect 14518 30096 18326 30152
rect 18382 30096 18387 30152
rect 14457 30094 18387 30096
rect 14457 30091 14523 30094
rect 18321 30091 18387 30094
rect 28993 30154 29059 30157
rect 28993 30152 32108 30154
rect 28993 30096 28998 30152
rect 29054 30096 32108 30152
rect 28993 30094 32108 30096
rect 28993 30091 29059 30094
rect 55622 30092 55628 30156
rect 55692 30154 55698 30156
rect 58433 30154 58499 30157
rect 55692 30152 58604 30154
rect 55692 30096 58438 30152
rect 58494 30096 58604 30152
rect 55692 30094 58604 30096
rect 55692 30092 55698 30094
rect 58433 30091 58499 30094
rect 17217 30018 17283 30021
rect 18873 30018 18939 30021
rect 17217 30016 18939 30018
rect 17217 29960 17222 30016
rect 17278 29960 18878 30016
rect 18934 29960 18939 30016
rect 17217 29958 18939 29960
rect 17217 29955 17283 29958
rect 18873 29955 18939 29958
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 0 29746 800 29776
rect 4061 29746 4127 29749
rect 0 29744 4127 29746
rect 0 29688 4066 29744
rect 4122 29688 4127 29744
rect 0 29686 4127 29688
rect 0 29656 800 29686
rect 4061 29683 4127 29686
rect 86217 29542 86283 29545
rect 86217 29540 86388 29542
rect 86217 29484 86222 29540
rect 86278 29484 86388 29540
rect 86217 29482 86388 29484
rect 86217 29479 86283 29482
rect 28901 29474 28967 29477
rect 28901 29472 32108 29474
rect 28901 29416 28906 29472
rect 28962 29416 32108 29472
rect 28901 29414 32108 29416
rect 28901 29411 28967 29414
rect 55806 29412 55812 29476
rect 55876 29474 55882 29476
rect 58433 29474 58499 29477
rect 55876 29472 58604 29474
rect 55876 29416 58438 29472
rect 58494 29416 58604 29472
rect 55876 29414 58604 29416
rect 55876 29412 55882 29414
rect 58433 29411 58499 29414
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 0 29066 800 29096
rect 3969 29066 4035 29069
rect 0 29064 4035 29066
rect 0 29008 3974 29064
rect 4030 29008 4035 29064
rect 0 29006 4035 29008
rect 0 28976 800 29006
rect 3969 29003 4035 29006
rect 7465 29066 7531 29069
rect 7465 29064 7666 29066
rect 7465 29008 7470 29064
rect 7526 29008 7666 29064
rect 7465 29006 7666 29008
rect 7465 29003 7531 29006
rect 7606 28797 7666 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 7557 28792 7666 28797
rect 7557 28736 7562 28792
rect 7618 28736 7666 28792
rect 7557 28734 7666 28736
rect 7557 28731 7623 28734
rect 0 28522 800 28552
rect 4061 28522 4127 28525
rect 0 28520 4127 28522
rect 0 28464 4066 28520
rect 4122 28464 4127 28520
rect 0 28462 4127 28464
rect 0 28432 800 28462
rect 4061 28459 4127 28462
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 86217 28182 86283 28185
rect 86217 28180 86388 28182
rect 86217 28124 86222 28180
rect 86278 28124 86388 28180
rect 86217 28122 86388 28124
rect 86217 28119 86283 28122
rect 28993 28114 29059 28117
rect 28993 28112 32108 28114
rect 28993 28056 28998 28112
rect 29054 28056 32108 28112
rect 28993 28054 32108 28056
rect 28993 28051 29059 28054
rect 58433 28046 58499 28049
rect 58022 28044 58604 28046
rect 0 27978 800 28008
rect 58022 27988 58438 28044
rect 58494 27988 58604 28044
rect 58022 27986 58604 27988
rect 3509 27978 3575 27981
rect 58022 27978 58082 27986
rect 58433 27983 58499 27986
rect 0 27976 3575 27978
rect 0 27920 3514 27976
rect 3570 27920 3575 27976
rect 0 27918 3575 27920
rect 0 27888 800 27918
rect 3509 27915 3575 27918
rect 55446 27918 58082 27978
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 9121 27570 9187 27573
rect 9254 27570 9260 27572
rect 9121 27568 9260 27570
rect 9121 27512 9126 27568
rect 9182 27512 9260 27568
rect 9121 27510 9260 27512
rect 9121 27507 9187 27510
rect 9254 27508 9260 27510
rect 9324 27508 9330 27572
rect 0 27298 800 27328
rect 4061 27298 4127 27301
rect 55446 27300 55506 27918
rect 0 27296 4127 27298
rect 0 27240 4066 27296
rect 4122 27240 4127 27296
rect 0 27238 4127 27240
rect 0 27208 800 27238
rect 4061 27235 4127 27238
rect 55438 27236 55444 27300
rect 55508 27236 55514 27300
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 55254 27100 55260 27164
rect 55324 27162 55330 27164
rect 56409 27162 56475 27165
rect 57421 27162 57487 27165
rect 55324 27160 57487 27162
rect 55324 27104 56414 27160
rect 56470 27104 57426 27160
rect 57482 27104 57487 27160
rect 55324 27102 57487 27104
rect 55324 27100 55330 27102
rect 56409 27099 56475 27102
rect 57421 27099 57487 27102
rect 58433 26822 58499 26825
rect 58433 26820 58604 26822
rect 0 26754 800 26784
rect 58433 26764 58438 26820
rect 58494 26764 58604 26820
rect 58433 26762 58604 26764
rect 58433 26759 58499 26762
rect 3509 26754 3575 26757
rect 0 26752 3575 26754
rect 0 26696 3514 26752
rect 3570 26696 3575 26752
rect 0 26694 3575 26696
rect 0 26664 800 26694
rect 3509 26691 3575 26694
rect 28901 26754 28967 26757
rect 28901 26752 32108 26754
rect 28901 26696 28906 26752
rect 28962 26696 32108 26752
rect 28901 26694 32108 26696
rect 28901 26691 28967 26694
rect 83406 26692 83412 26756
rect 83476 26754 83482 26756
rect 86217 26754 86283 26757
rect 83476 26752 86388 26754
rect 83476 26696 86222 26752
rect 86278 26696 86388 26752
rect 83476 26694 86388 26696
rect 83476 26692 83482 26694
rect 86217 26691 86283 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 4208 26144 4528 26145
rect 0 26074 800 26104
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 3509 26074 3575 26077
rect 0 26072 3575 26074
rect 0 26016 3514 26072
rect 3570 26016 3575 26072
rect 0 26014 3575 26016
rect 0 25984 800 26014
rect 3509 26011 3575 26014
rect 19568 25600 19888 25601
rect 0 25530 800 25560
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 58433 25598 58499 25601
rect 86217 25598 86283 25601
rect 58433 25596 58604 25598
rect 58433 25540 58438 25596
rect 58494 25540 58604 25596
rect 58433 25538 58604 25540
rect 86217 25596 86388 25598
rect 86217 25540 86222 25596
rect 86278 25540 86388 25596
rect 86217 25538 86388 25540
rect 58433 25535 58499 25538
rect 86217 25535 86283 25538
rect 3969 25530 4035 25533
rect 0 25528 4035 25530
rect 0 25472 3974 25528
rect 4030 25472 4035 25528
rect 0 25470 4035 25472
rect 0 25440 800 25470
rect 3969 25467 4035 25470
rect 28993 25530 29059 25533
rect 28993 25528 32108 25530
rect 28993 25472 28998 25528
rect 29054 25472 32108 25528
rect 28993 25470 32108 25472
rect 28993 25467 29059 25470
rect 4208 25056 4528 25057
rect 0 24986 800 25016
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 3969 24986 4035 24989
rect 0 24984 4035 24986
rect 0 24928 3974 24984
rect 4030 24928 4035 24984
rect 0 24926 4035 24928
rect 0 24896 800 24926
rect 3969 24923 4035 24926
rect 13353 24850 13419 24853
rect 14273 24850 14339 24853
rect 13353 24848 14339 24850
rect 13353 24792 13358 24848
rect 13414 24792 14278 24848
rect 14334 24792 14339 24848
rect 13353 24790 14339 24792
rect 13353 24787 13419 24790
rect 14273 24787 14339 24790
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 0 24306 800 24336
rect 3969 24306 4035 24309
rect 0 24304 4035 24306
rect 0 24248 3974 24304
rect 4030 24248 4035 24304
rect 0 24246 4035 24248
rect 0 24216 800 24246
rect 3969 24243 4035 24246
rect 86217 24238 86283 24241
rect 85806 24236 86388 24238
rect 85806 24180 86222 24236
rect 86278 24180 86388 24236
rect 85806 24178 86388 24180
rect 28993 24170 29059 24173
rect 28993 24168 32108 24170
rect 28993 24112 28998 24168
rect 29054 24112 32108 24168
rect 28993 24110 32108 24112
rect 28993 24107 29059 24110
rect 52678 24108 52684 24172
rect 52748 24170 52754 24172
rect 55254 24170 55260 24172
rect 52748 24110 55260 24170
rect 52748 24108 52754 24110
rect 55254 24108 55260 24110
rect 55324 24108 55330 24172
rect 58065 24170 58131 24173
rect 58433 24170 58499 24173
rect 58065 24168 58604 24170
rect 58065 24112 58070 24168
rect 58126 24112 58438 24168
rect 58494 24112 58604 24168
rect 58065 24110 58604 24112
rect 58065 24107 58131 24110
rect 58433 24107 58499 24110
rect 83038 24108 83044 24172
rect 83108 24170 83114 24172
rect 85806 24170 85866 24178
rect 86217 24175 86283 24178
rect 83108 24110 85866 24170
rect 83108 24108 83114 24110
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 53046 23836 53052 23900
rect 53116 23898 53122 23900
rect 55438 23898 55444 23900
rect 53116 23838 55444 23898
rect 53116 23836 53122 23838
rect 55438 23836 55444 23838
rect 55508 23836 55514 23900
rect 0 23762 800 23792
rect 4061 23762 4127 23765
rect 0 23760 4127 23762
rect 0 23704 4066 23760
rect 4122 23704 4127 23760
rect 0 23702 4127 23704
rect 0 23672 800 23702
rect 4061 23699 4127 23702
rect 15837 23492 15903 23493
rect 15837 23490 15884 23492
rect 15792 23488 15884 23490
rect 15792 23432 15842 23488
rect 15792 23430 15884 23432
rect 15837 23428 15884 23430
rect 15948 23428 15954 23492
rect 22553 23490 22619 23493
rect 31886 23490 31892 23492
rect 22553 23488 31892 23490
rect 22553 23432 22558 23488
rect 22614 23432 31892 23488
rect 22553 23430 31892 23432
rect 15837 23427 15903 23428
rect 22553 23427 22619 23430
rect 31886 23428 31892 23430
rect 31956 23428 31962 23492
rect 52310 23428 52316 23492
rect 52380 23490 52386 23492
rect 58341 23490 58407 23493
rect 52380 23488 58407 23490
rect 52380 23432 58346 23488
rect 58402 23432 58407 23488
rect 52380 23430 58407 23432
rect 52380 23428 52386 23430
rect 58341 23427 58407 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 55254 23292 55260 23356
rect 55324 23354 55330 23356
rect 58065 23354 58131 23357
rect 55324 23352 58131 23354
rect 55324 23296 58070 23352
rect 58126 23296 58131 23352
rect 55324 23294 58131 23296
rect 55324 23292 55330 23294
rect 58065 23291 58131 23294
rect 108297 23218 108363 23221
rect 111440 23218 112240 23248
rect 108297 23216 112240 23218
rect 108297 23160 108302 23216
rect 108358 23160 112240 23216
rect 108297 23158 112240 23160
rect 108297 23155 108363 23158
rect 111440 23128 112240 23158
rect 0 23082 800 23112
rect 4061 23082 4127 23085
rect 0 23080 4127 23082
rect 0 23024 4066 23080
rect 4122 23024 4127 23080
rect 0 23022 4127 23024
rect 0 22992 800 23022
rect 4061 23019 4127 23022
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 86033 22878 86099 22881
rect 4208 22815 4528 22816
rect 85806 22876 86388 22878
rect 85806 22820 86038 22876
rect 86094 22820 86388 22876
rect 85806 22818 86388 22820
rect 9949 22812 10015 22813
rect 9949 22810 9996 22812
rect 9904 22808 9996 22810
rect 9904 22752 9954 22808
rect 9904 22750 9996 22752
rect 9949 22748 9996 22750
rect 10060 22748 10066 22812
rect 29085 22810 29151 22813
rect 29085 22808 32108 22810
rect 29085 22752 29090 22808
rect 29146 22752 32108 22808
rect 29085 22750 32108 22752
rect 9949 22747 10015 22748
rect 29085 22747 29151 22750
rect 54518 22748 54524 22812
rect 54588 22810 54594 22812
rect 58433 22810 58499 22813
rect 54588 22808 58604 22810
rect 54588 22752 58438 22808
rect 58494 22752 58604 22808
rect 54588 22750 58604 22752
rect 54588 22748 54594 22750
rect 58433 22747 58499 22750
rect 83958 22748 83964 22812
rect 84028 22810 84034 22812
rect 85806 22810 85866 22818
rect 86033 22815 86099 22818
rect 84028 22750 85866 22810
rect 84028 22748 84034 22750
rect 0 22538 800 22568
rect 3325 22538 3391 22541
rect 0 22536 3391 22538
rect 0 22480 3330 22536
rect 3386 22480 3391 22536
rect 0 22478 3391 22480
rect 0 22448 800 22478
rect 3325 22475 3391 22478
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 18597 22130 18663 22133
rect 19190 22130 19196 22132
rect 18597 22128 19196 22130
rect 18597 22072 18602 22128
rect 18658 22072 19196 22128
rect 18597 22070 19196 22072
rect 18597 22067 18663 22070
rect 19190 22068 19196 22070
rect 19260 22068 19266 22132
rect 52310 22068 52316 22132
rect 52380 22130 52386 22132
rect 55622 22130 55628 22132
rect 52380 22070 55628 22130
rect 52380 22068 52386 22070
rect 55622 22068 55628 22070
rect 55692 22068 55698 22132
rect 19374 21932 19380 21996
rect 19444 21994 19450 21996
rect 31886 21994 31892 21996
rect 19444 21934 31892 21994
rect 19444 21932 19450 21934
rect 31886 21932 31892 21934
rect 31956 21932 31962 21996
rect 0 21858 800 21888
rect 4061 21858 4127 21861
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 800 21798
rect 4061 21795 4127 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 14457 21450 14523 21453
rect 14590 21450 14596 21452
rect 14457 21448 14596 21450
rect 14457 21392 14462 21448
rect 14518 21392 14596 21448
rect 14457 21390 14596 21392
rect 14457 21387 14523 21390
rect 14590 21388 14596 21390
rect 14660 21388 14666 21452
rect 0 21314 800 21344
rect 3969 21314 4035 21317
rect 0 21312 4035 21314
rect 0 21256 3974 21312
rect 4030 21256 4035 21312
rect 0 21254 4035 21256
rect 0 21224 800 21254
rect 3969 21251 4035 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 0 20770 800 20800
rect 4061 20770 4127 20773
rect 0 20768 4127 20770
rect 0 20712 4066 20768
rect 4122 20712 4127 20768
rect 0 20710 4127 20712
rect 0 20680 800 20710
rect 4061 20707 4127 20710
rect 23933 20770 23999 20773
rect 24158 20770 24164 20772
rect 23933 20768 24164 20770
rect 23933 20712 23938 20768
rect 23994 20712 24164 20768
rect 23933 20710 24164 20712
rect 23933 20707 23999 20710
rect 24158 20708 24164 20710
rect 24228 20708 24234 20772
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 19568 20160 19888 20161
rect 0 20090 800 20120
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 85941 20158 86007 20161
rect 19568 20095 19888 20096
rect 85806 20156 86388 20158
rect 85806 20100 85946 20156
rect 86002 20100 86388 20156
rect 85806 20098 86388 20100
rect 2865 20090 2931 20093
rect 0 20088 2931 20090
rect 0 20032 2870 20088
rect 2926 20032 2931 20088
rect 0 20030 2931 20032
rect 0 20000 800 20030
rect 2865 20027 2931 20030
rect 29085 20090 29151 20093
rect 29085 20088 32108 20090
rect 29085 20032 29090 20088
rect 29146 20032 32108 20088
rect 29085 20030 32108 20032
rect 29085 20027 29151 20030
rect 56174 20028 56180 20092
rect 56244 20090 56250 20092
rect 58433 20090 58499 20093
rect 56244 20088 58604 20090
rect 56244 20032 58438 20088
rect 58494 20032 58604 20088
rect 56244 20030 58604 20032
rect 56244 20028 56250 20030
rect 58433 20027 58499 20030
rect 83222 20028 83228 20092
rect 83292 20090 83298 20092
rect 85806 20090 85866 20098
rect 85941 20095 86007 20098
rect 83292 20030 85866 20090
rect 83292 20028 83298 20030
rect 4208 19616 4528 19617
rect 0 19546 800 19576
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 3693 19546 3759 19549
rect 0 19544 3759 19546
rect 0 19488 3698 19544
rect 3754 19488 3759 19544
rect 0 19486 3759 19488
rect 0 19456 800 19486
rect 3693 19483 3759 19486
rect 25037 19274 25103 19277
rect 25405 19274 25471 19277
rect 25037 19272 25471 19274
rect 25037 19216 25042 19272
rect 25098 19216 25410 19272
rect 25466 19216 25471 19272
rect 25037 19214 25471 19216
rect 25037 19211 25103 19214
rect 25405 19211 25471 19214
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 0 18866 800 18896
rect 3969 18866 4035 18869
rect 0 18864 4035 18866
rect 0 18808 3974 18864
rect 4030 18808 4035 18864
rect 0 18806 4035 18808
rect 0 18776 800 18806
rect 3969 18803 4035 18806
rect 27705 18730 27771 18733
rect 27838 18730 27844 18732
rect 27705 18728 27844 18730
rect 27705 18672 27710 18728
rect 27766 18672 27844 18728
rect 27705 18670 27844 18672
rect 27705 18667 27771 18670
rect 27838 18668 27844 18670
rect 27908 18668 27914 18732
rect 14457 18594 14523 18597
rect 17125 18594 17191 18597
rect 14457 18592 17191 18594
rect 14457 18536 14462 18592
rect 14518 18536 17130 18592
rect 17186 18536 17191 18592
rect 14457 18534 17191 18536
rect 14457 18531 14523 18534
rect 17125 18531 17191 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 0 18322 800 18352
rect 3417 18322 3483 18325
rect 0 18320 3483 18322
rect 0 18264 3422 18320
rect 3478 18264 3483 18320
rect 0 18262 3483 18264
rect 0 18232 800 18262
rect 3417 18259 3483 18262
rect 8109 18050 8175 18053
rect 9581 18050 9647 18053
rect 8109 18048 9647 18050
rect 8109 17992 8114 18048
rect 8170 17992 9586 18048
rect 9642 17992 9647 18048
rect 8109 17990 9647 17992
rect 8109 17987 8175 17990
rect 9581 17987 9647 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 0 17778 800 17808
rect 3325 17778 3391 17781
rect 0 17776 3391 17778
rect 0 17720 3330 17776
rect 3386 17720 3391 17776
rect 0 17718 3391 17720
rect 0 17688 800 17718
rect 3325 17715 3391 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 22553 17370 22619 17373
rect 22686 17370 22692 17372
rect 22553 17368 22692 17370
rect 22553 17312 22558 17368
rect 22614 17312 22692 17368
rect 22553 17310 22692 17312
rect 22553 17307 22619 17310
rect 22686 17308 22692 17310
rect 22756 17308 22762 17372
rect 82854 17172 82860 17236
rect 82924 17234 82930 17236
rect 83222 17234 83228 17236
rect 82924 17174 83228 17234
rect 82924 17172 82930 17174
rect 83222 17172 83228 17174
rect 83292 17172 83298 17236
rect 0 17098 800 17128
rect 4061 17098 4127 17101
rect 0 17096 4127 17098
rect 0 17040 4066 17096
rect 4122 17040 4127 17096
rect 0 17038 4127 17040
rect 0 17008 800 17038
rect 4061 17035 4127 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 10501 16692 10567 16693
rect 10501 16690 10548 16692
rect 10456 16688 10548 16690
rect 10456 16632 10506 16688
rect 10456 16630 10548 16632
rect 10501 16628 10548 16630
rect 10612 16628 10618 16692
rect 10501 16627 10567 16628
rect 0 16554 800 16584
rect 4061 16554 4127 16557
rect 0 16552 4127 16554
rect 0 16496 4066 16552
rect 4122 16496 4127 16552
rect 0 16494 4127 16496
rect 0 16464 800 16494
rect 4061 16491 4127 16494
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 21909 16012 21975 16013
rect 21909 16010 21956 16012
rect 21864 16008 21956 16010
rect 21864 15952 21914 16008
rect 21864 15950 21956 15952
rect 21909 15948 21956 15950
rect 22020 15948 22026 16012
rect 21909 15947 21975 15948
rect 0 15874 800 15904
rect 3877 15874 3943 15877
rect 0 15872 3943 15874
rect 0 15816 3882 15872
rect 3938 15816 3943 15872
rect 0 15814 3943 15816
rect 0 15784 800 15814
rect 3877 15811 3943 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 0 15330 800 15360
rect 3969 15330 4035 15333
rect 24853 15332 24919 15333
rect 24853 15330 24900 15332
rect 0 15328 4035 15330
rect 0 15272 3974 15328
rect 4030 15272 4035 15328
rect 0 15270 4035 15272
rect 24808 15328 24900 15330
rect 24808 15272 24858 15328
rect 24808 15270 24900 15272
rect 0 15240 800 15270
rect 3969 15267 4035 15270
rect 24853 15268 24900 15270
rect 24964 15268 24970 15332
rect 24853 15267 24919 15268
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 58433 14854 58499 14857
rect 86217 14854 86283 14857
rect 58433 14852 58604 14854
rect 58433 14796 58438 14852
rect 58494 14796 58604 14852
rect 58433 14794 58604 14796
rect 85806 14852 86388 14854
rect 85806 14796 86222 14852
rect 86278 14796 86388 14852
rect 85806 14794 86388 14796
rect 58433 14791 58499 14794
rect 28993 14786 29059 14789
rect 28993 14784 32108 14786
rect 28993 14728 28998 14784
rect 29054 14728 32108 14784
rect 28993 14726 32108 14728
rect 28993 14723 29059 14726
rect 82854 14724 82860 14788
rect 82924 14786 82930 14788
rect 85806 14786 85866 14794
rect 86217 14791 86283 14794
rect 82924 14726 85866 14786
rect 82924 14724 82930 14726
rect 19568 14720 19888 14721
rect 0 14650 800 14680
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 4889 14650 4955 14653
rect 0 14648 4955 14650
rect 0 14592 4894 14648
rect 4950 14592 4955 14648
rect 0 14590 4955 14592
rect 0 14560 800 14590
rect 4889 14587 4955 14590
rect 4208 14176 4528 14177
rect 0 14106 800 14136
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 3969 14106 4035 14109
rect 0 14104 4035 14106
rect 0 14048 3974 14104
rect 4030 14048 4035 14104
rect 0 14046 4035 14048
rect 0 14016 800 14046
rect 3969 14043 4035 14046
rect 24025 13970 24091 13973
rect 24158 13970 24164 13972
rect 24025 13968 24164 13970
rect 24025 13912 24030 13968
rect 24086 13912 24164 13968
rect 24025 13910 24164 13912
rect 24025 13907 24091 13910
rect 24158 13908 24164 13910
rect 24228 13908 24234 13972
rect 19568 13632 19888 13633
rect 0 13562 800 13592
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 4061 13562 4127 13565
rect 0 13560 4127 13562
rect 0 13504 4066 13560
rect 4122 13504 4127 13560
rect 0 13502 4127 13504
rect 0 13472 800 13502
rect 4061 13499 4127 13502
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 0 12882 800 12912
rect 3969 12882 4035 12885
rect 0 12880 4035 12882
rect 0 12824 3974 12880
rect 4030 12824 4035 12880
rect 0 12822 4035 12824
rect 0 12792 800 12822
rect 3969 12819 4035 12822
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 0 12338 800 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 0 11658 800 11688
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11568 800 11598
rect 4061 11595 4127 11598
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 0 11114 800 11144
rect 3969 11114 4035 11117
rect 0 11112 4035 11114
rect 0 11056 3974 11112
rect 4030 11056 4035 11112
rect 0 11054 4035 11056
rect 0 11024 800 11054
rect 3969 11051 4035 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 0 10570 800 10600
rect 4061 10570 4127 10573
rect 0 10568 4127 10570
rect 0 10512 4066 10568
rect 4122 10512 4127 10568
rect 0 10510 4127 10512
rect 0 10480 800 10510
rect 4061 10507 4127 10510
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 0 9890 800 9920
rect 3969 9890 4035 9893
rect 0 9888 4035 9890
rect 0 9832 3974 9888
rect 4030 9832 4035 9888
rect 0 9830 4035 9832
rect 0 9800 800 9830
rect 3969 9827 4035 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 0 9346 800 9376
rect 4061 9346 4127 9349
rect 0 9344 4127 9346
rect 0 9288 4066 9344
rect 4122 9288 4127 9344
rect 0 9286 4127 9288
rect 0 9256 800 9286
rect 4061 9283 4127 9286
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 4208 8736 4528 8737
rect 0 8666 800 8696
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 4061 8666 4127 8669
rect 0 8664 4127 8666
rect 0 8608 4066 8664
rect 4122 8608 4127 8664
rect 0 8606 4127 8608
rect 0 8576 800 8606
rect 4061 8603 4127 8606
rect 19568 8192 19888 8193
rect 0 8122 800 8152
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 3969 8122 4035 8125
rect 0 8120 4035 8122
rect 0 8064 3974 8120
rect 4030 8064 4035 8120
rect 0 8062 4035 8064
rect 0 8032 800 8062
rect 3969 8059 4035 8062
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 0 7442 800 7472
rect 4061 7442 4127 7445
rect 0 7440 4127 7442
rect 0 7384 4066 7440
rect 4122 7384 4127 7440
rect 0 7382 4127 7384
rect 0 7352 800 7382
rect 4061 7379 4127 7382
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 0 6898 800 6928
rect 3325 6898 3391 6901
rect 0 6896 3391 6898
rect 0 6840 3330 6896
rect 3386 6840 3391 6896
rect 0 6838 3391 6840
rect 0 6808 800 6838
rect 3325 6835 3391 6838
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 0 6354 800 6384
rect 3693 6354 3759 6357
rect 0 6352 3759 6354
rect 0 6296 3698 6352
rect 3754 6296 3759 6352
rect 0 6294 3759 6296
rect 0 6264 800 6294
rect 3693 6291 3759 6294
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 0 5674 800 5704
rect 3969 5674 4035 5677
rect 0 5672 4035 5674
rect 0 5616 3974 5672
rect 4030 5616 4035 5672
rect 0 5614 4035 5616
rect 0 5584 800 5614
rect 3969 5611 4035 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 0 5130 800 5160
rect 4061 5130 4127 5133
rect 0 5128 4127 5130
rect 0 5072 4066 5128
rect 4122 5072 4127 5128
rect 0 5070 4127 5072
rect 0 5040 800 5070
rect 4061 5067 4127 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 29913 4858 29979 4861
rect 56409 4858 56475 4861
rect 84009 4858 84075 4861
rect 29913 4856 32108 4858
rect 29913 4800 29918 4856
rect 29974 4800 32108 4856
rect 29913 4798 32108 4800
rect 56409 4856 58604 4858
rect 56409 4800 56414 4856
rect 56470 4800 58604 4856
rect 56409 4798 58604 4800
rect 84009 4856 86388 4858
rect 84009 4800 84014 4856
rect 84070 4800 86388 4856
rect 84009 4798 86388 4800
rect 29913 4795 29979 4798
rect 56409 4795 56475 4798
rect 84009 4795 84075 4798
rect 0 4450 800 4480
rect 3969 4450 4035 4453
rect 0 4448 4035 4450
rect 0 4392 3974 4448
rect 4030 4392 4035 4448
rect 0 4390 4035 4392
rect 0 4360 800 4390
rect 3969 4387 4035 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 0 3906 800 3936
rect 4061 3906 4127 3909
rect 0 3904 4127 3906
rect 0 3848 4066 3904
rect 4122 3848 4127 3904
rect 0 3846 4127 3848
rect 0 3816 800 3846
rect 4061 3843 4127 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 0 3362 800 3392
rect 3969 3362 4035 3365
rect 0 3360 4035 3362
rect 0 3304 3974 3360
rect 4030 3304 4035 3360
rect 0 3302 4035 3304
rect 0 3272 800 3302
rect 3969 3299 4035 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 19568 2752 19888 2753
rect 0 2682 800 2712
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 2681 2682 2747 2685
rect 0 2680 2747 2682
rect 0 2624 2686 2680
rect 2742 2624 2747 2680
rect 0 2622 2747 2624
rect 0 2592 800 2622
rect 2681 2619 2747 2622
rect 4208 2208 4528 2209
rect 0 2138 800 2168
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 4061 2138 4127 2141
rect 0 2136 4127 2138
rect 0 2080 4066 2136
rect 4122 2080 4127 2136
rect 0 2078 4127 2080
rect 0 2048 800 2078
rect 4061 2075 4127 2078
rect 0 1458 800 1488
rect 3785 1458 3851 1461
rect 0 1456 3851 1458
rect 0 1400 3790 1456
rect 3846 1400 3851 1456
rect 0 1398 3851 1400
rect 0 1368 800 1398
rect 3785 1395 3851 1398
rect 0 914 800 944
rect 2773 914 2839 917
rect 0 912 2839 914
rect 0 856 2778 912
rect 2834 856 2839 912
rect 0 854 2839 856
rect 0 824 800 854
rect 2773 851 2839 854
rect 0 370 800 400
rect 3049 370 3115 373
rect 0 368 3115 370
rect 0 312 3054 368
rect 3110 312 3115 368
rect 0 310 3115 312
rect 0 280 800 310
rect 3049 307 3115 310
<< via3 >>
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 50296 44092 50360 44096
rect 50296 44036 50300 44092
rect 50300 44036 50356 44092
rect 50356 44036 50360 44092
rect 50296 44032 50360 44036
rect 50376 44092 50440 44096
rect 50376 44036 50380 44092
rect 50380 44036 50436 44092
rect 50436 44036 50440 44092
rect 50376 44032 50440 44036
rect 50456 44092 50520 44096
rect 50456 44036 50460 44092
rect 50460 44036 50516 44092
rect 50516 44036 50520 44092
rect 50456 44032 50520 44036
rect 50536 44092 50600 44096
rect 50536 44036 50540 44092
rect 50540 44036 50596 44092
rect 50596 44036 50600 44092
rect 50536 44032 50600 44036
rect 81016 44092 81080 44096
rect 81016 44036 81020 44092
rect 81020 44036 81076 44092
rect 81076 44036 81080 44092
rect 81016 44032 81080 44036
rect 81096 44092 81160 44096
rect 81096 44036 81100 44092
rect 81100 44036 81156 44092
rect 81156 44036 81160 44092
rect 81096 44032 81160 44036
rect 81176 44092 81240 44096
rect 81176 44036 81180 44092
rect 81180 44036 81236 44092
rect 81236 44036 81240 44092
rect 81176 44032 81240 44036
rect 81256 44092 81320 44096
rect 81256 44036 81260 44092
rect 81260 44036 81316 44092
rect 81316 44036 81320 44092
rect 81256 44032 81320 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 65656 43548 65720 43552
rect 65656 43492 65660 43548
rect 65660 43492 65716 43548
rect 65716 43492 65720 43548
rect 65656 43488 65720 43492
rect 65736 43548 65800 43552
rect 65736 43492 65740 43548
rect 65740 43492 65796 43548
rect 65796 43492 65800 43548
rect 65736 43488 65800 43492
rect 65816 43548 65880 43552
rect 65816 43492 65820 43548
rect 65820 43492 65876 43548
rect 65876 43492 65880 43548
rect 65816 43488 65880 43492
rect 65896 43548 65960 43552
rect 65896 43492 65900 43548
rect 65900 43492 65956 43548
rect 65956 43492 65960 43548
rect 65896 43488 65960 43492
rect 96376 43548 96440 43552
rect 96376 43492 96380 43548
rect 96380 43492 96436 43548
rect 96436 43492 96440 43548
rect 96376 43488 96440 43492
rect 96456 43548 96520 43552
rect 96456 43492 96460 43548
rect 96460 43492 96516 43548
rect 96516 43492 96520 43548
rect 96456 43488 96520 43492
rect 96536 43548 96600 43552
rect 96536 43492 96540 43548
rect 96540 43492 96596 43548
rect 96596 43492 96600 43548
rect 96536 43488 96600 43492
rect 96616 43548 96680 43552
rect 96616 43492 96620 43548
rect 96620 43492 96676 43548
rect 96676 43492 96680 43548
rect 96616 43488 96680 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 50296 43004 50360 43008
rect 50296 42948 50300 43004
rect 50300 42948 50356 43004
rect 50356 42948 50360 43004
rect 50296 42944 50360 42948
rect 50376 43004 50440 43008
rect 50376 42948 50380 43004
rect 50380 42948 50436 43004
rect 50436 42948 50440 43004
rect 50376 42944 50440 42948
rect 50456 43004 50520 43008
rect 50456 42948 50460 43004
rect 50460 42948 50516 43004
rect 50516 42948 50520 43004
rect 50456 42944 50520 42948
rect 50536 43004 50600 43008
rect 50536 42948 50540 43004
rect 50540 42948 50596 43004
rect 50596 42948 50600 43004
rect 50536 42944 50600 42948
rect 81016 43004 81080 43008
rect 81016 42948 81020 43004
rect 81020 42948 81076 43004
rect 81076 42948 81080 43004
rect 81016 42944 81080 42948
rect 81096 43004 81160 43008
rect 81096 42948 81100 43004
rect 81100 42948 81156 43004
rect 81156 42948 81160 43004
rect 81096 42944 81160 42948
rect 81176 43004 81240 43008
rect 81176 42948 81180 43004
rect 81180 42948 81236 43004
rect 81236 42948 81240 43004
rect 81176 42944 81240 42948
rect 81256 43004 81320 43008
rect 81256 42948 81260 43004
rect 81260 42948 81316 43004
rect 81316 42948 81320 43004
rect 81256 42944 81320 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 65656 42460 65720 42464
rect 65656 42404 65660 42460
rect 65660 42404 65716 42460
rect 65716 42404 65720 42460
rect 65656 42400 65720 42404
rect 65736 42460 65800 42464
rect 65736 42404 65740 42460
rect 65740 42404 65796 42460
rect 65796 42404 65800 42460
rect 65736 42400 65800 42404
rect 65816 42460 65880 42464
rect 65816 42404 65820 42460
rect 65820 42404 65876 42460
rect 65876 42404 65880 42460
rect 65816 42400 65880 42404
rect 65896 42460 65960 42464
rect 65896 42404 65900 42460
rect 65900 42404 65956 42460
rect 65956 42404 65960 42460
rect 65896 42400 65960 42404
rect 96376 42460 96440 42464
rect 96376 42404 96380 42460
rect 96380 42404 96436 42460
rect 96436 42404 96440 42460
rect 96376 42400 96440 42404
rect 96456 42460 96520 42464
rect 96456 42404 96460 42460
rect 96460 42404 96516 42460
rect 96516 42404 96520 42460
rect 96456 42400 96520 42404
rect 96536 42460 96600 42464
rect 96536 42404 96540 42460
rect 96540 42404 96596 42460
rect 96596 42404 96600 42460
rect 96536 42400 96600 42404
rect 96616 42460 96680 42464
rect 96616 42404 96620 42460
rect 96620 42404 96676 42460
rect 96676 42404 96680 42460
rect 96616 42400 96680 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 50296 41916 50360 41920
rect 50296 41860 50300 41916
rect 50300 41860 50356 41916
rect 50356 41860 50360 41916
rect 50296 41856 50360 41860
rect 50376 41916 50440 41920
rect 50376 41860 50380 41916
rect 50380 41860 50436 41916
rect 50436 41860 50440 41916
rect 50376 41856 50440 41860
rect 50456 41916 50520 41920
rect 50456 41860 50460 41916
rect 50460 41860 50516 41916
rect 50516 41860 50520 41916
rect 50456 41856 50520 41860
rect 50536 41916 50600 41920
rect 50536 41860 50540 41916
rect 50540 41860 50596 41916
rect 50596 41860 50600 41916
rect 50536 41856 50600 41860
rect 81016 41916 81080 41920
rect 81016 41860 81020 41916
rect 81020 41860 81076 41916
rect 81076 41860 81080 41916
rect 81016 41856 81080 41860
rect 81096 41916 81160 41920
rect 81096 41860 81100 41916
rect 81100 41860 81156 41916
rect 81156 41860 81160 41916
rect 81096 41856 81160 41860
rect 81176 41916 81240 41920
rect 81176 41860 81180 41916
rect 81180 41860 81236 41916
rect 81236 41860 81240 41916
rect 81176 41856 81240 41860
rect 81256 41916 81320 41920
rect 81256 41860 81260 41916
rect 81260 41860 81316 41916
rect 81316 41860 81320 41916
rect 81256 41856 81320 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 65656 41372 65720 41376
rect 65656 41316 65660 41372
rect 65660 41316 65716 41372
rect 65716 41316 65720 41372
rect 65656 41312 65720 41316
rect 65736 41372 65800 41376
rect 65736 41316 65740 41372
rect 65740 41316 65796 41372
rect 65796 41316 65800 41372
rect 65736 41312 65800 41316
rect 65816 41372 65880 41376
rect 65816 41316 65820 41372
rect 65820 41316 65876 41372
rect 65876 41316 65880 41372
rect 65816 41312 65880 41316
rect 65896 41372 65960 41376
rect 65896 41316 65900 41372
rect 65900 41316 65956 41372
rect 65956 41316 65960 41372
rect 65896 41312 65960 41316
rect 96376 41372 96440 41376
rect 96376 41316 96380 41372
rect 96380 41316 96436 41372
rect 96436 41316 96440 41372
rect 96376 41312 96440 41316
rect 96456 41372 96520 41376
rect 96456 41316 96460 41372
rect 96460 41316 96516 41372
rect 96516 41316 96520 41372
rect 96456 41312 96520 41316
rect 96536 41372 96600 41376
rect 96536 41316 96540 41372
rect 96540 41316 96596 41372
rect 96596 41316 96600 41372
rect 96536 41312 96600 41316
rect 96616 41372 96680 41376
rect 96616 41316 96620 41372
rect 96620 41316 96676 41372
rect 96676 41316 96680 41372
rect 96616 41312 96680 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 50296 40828 50360 40832
rect 50296 40772 50300 40828
rect 50300 40772 50356 40828
rect 50356 40772 50360 40828
rect 50296 40768 50360 40772
rect 50376 40828 50440 40832
rect 50376 40772 50380 40828
rect 50380 40772 50436 40828
rect 50436 40772 50440 40828
rect 50376 40768 50440 40772
rect 50456 40828 50520 40832
rect 50456 40772 50460 40828
rect 50460 40772 50516 40828
rect 50516 40772 50520 40828
rect 50456 40768 50520 40772
rect 50536 40828 50600 40832
rect 50536 40772 50540 40828
rect 50540 40772 50596 40828
rect 50596 40772 50600 40828
rect 50536 40768 50600 40772
rect 81016 40828 81080 40832
rect 81016 40772 81020 40828
rect 81020 40772 81076 40828
rect 81076 40772 81080 40828
rect 81016 40768 81080 40772
rect 81096 40828 81160 40832
rect 81096 40772 81100 40828
rect 81100 40772 81156 40828
rect 81156 40772 81160 40828
rect 81096 40768 81160 40772
rect 81176 40828 81240 40832
rect 81176 40772 81180 40828
rect 81180 40772 81236 40828
rect 81236 40772 81240 40828
rect 81176 40768 81240 40772
rect 81256 40828 81320 40832
rect 81256 40772 81260 40828
rect 81260 40772 81316 40828
rect 81316 40772 81320 40828
rect 81256 40768 81320 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 65656 40284 65720 40288
rect 65656 40228 65660 40284
rect 65660 40228 65716 40284
rect 65716 40228 65720 40284
rect 65656 40224 65720 40228
rect 65736 40284 65800 40288
rect 65736 40228 65740 40284
rect 65740 40228 65796 40284
rect 65796 40228 65800 40284
rect 65736 40224 65800 40228
rect 65816 40284 65880 40288
rect 65816 40228 65820 40284
rect 65820 40228 65876 40284
rect 65876 40228 65880 40284
rect 65816 40224 65880 40228
rect 65896 40284 65960 40288
rect 65896 40228 65900 40284
rect 65900 40228 65956 40284
rect 65956 40228 65960 40284
rect 65896 40224 65960 40228
rect 96376 40284 96440 40288
rect 96376 40228 96380 40284
rect 96380 40228 96436 40284
rect 96436 40228 96440 40284
rect 96376 40224 96440 40228
rect 96456 40284 96520 40288
rect 96456 40228 96460 40284
rect 96460 40228 96516 40284
rect 96516 40228 96520 40284
rect 96456 40224 96520 40228
rect 96536 40284 96600 40288
rect 96536 40228 96540 40284
rect 96540 40228 96596 40284
rect 96596 40228 96600 40284
rect 96536 40224 96600 40228
rect 96616 40284 96680 40288
rect 96616 40228 96620 40284
rect 96620 40228 96676 40284
rect 96676 40228 96680 40284
rect 96616 40224 96680 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 50296 39740 50360 39744
rect 50296 39684 50300 39740
rect 50300 39684 50356 39740
rect 50356 39684 50360 39740
rect 50296 39680 50360 39684
rect 50376 39740 50440 39744
rect 50376 39684 50380 39740
rect 50380 39684 50436 39740
rect 50436 39684 50440 39740
rect 50376 39680 50440 39684
rect 50456 39740 50520 39744
rect 50456 39684 50460 39740
rect 50460 39684 50516 39740
rect 50516 39684 50520 39740
rect 50456 39680 50520 39684
rect 50536 39740 50600 39744
rect 50536 39684 50540 39740
rect 50540 39684 50596 39740
rect 50596 39684 50600 39740
rect 50536 39680 50600 39684
rect 81016 39740 81080 39744
rect 81016 39684 81020 39740
rect 81020 39684 81076 39740
rect 81076 39684 81080 39740
rect 81016 39680 81080 39684
rect 81096 39740 81160 39744
rect 81096 39684 81100 39740
rect 81100 39684 81156 39740
rect 81156 39684 81160 39740
rect 81096 39680 81160 39684
rect 81176 39740 81240 39744
rect 81176 39684 81180 39740
rect 81180 39684 81236 39740
rect 81236 39684 81240 39740
rect 81176 39680 81240 39684
rect 81256 39740 81320 39744
rect 81256 39684 81260 39740
rect 81260 39684 81316 39740
rect 81316 39684 81320 39740
rect 81256 39680 81320 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 65656 39196 65720 39200
rect 65656 39140 65660 39196
rect 65660 39140 65716 39196
rect 65716 39140 65720 39196
rect 65656 39136 65720 39140
rect 65736 39196 65800 39200
rect 65736 39140 65740 39196
rect 65740 39140 65796 39196
rect 65796 39140 65800 39196
rect 65736 39136 65800 39140
rect 65816 39196 65880 39200
rect 65816 39140 65820 39196
rect 65820 39140 65876 39196
rect 65876 39140 65880 39196
rect 65816 39136 65880 39140
rect 65896 39196 65960 39200
rect 65896 39140 65900 39196
rect 65900 39140 65956 39196
rect 65956 39140 65960 39196
rect 65896 39136 65960 39140
rect 96376 39196 96440 39200
rect 96376 39140 96380 39196
rect 96380 39140 96436 39196
rect 96436 39140 96440 39196
rect 96376 39136 96440 39140
rect 96456 39196 96520 39200
rect 96456 39140 96460 39196
rect 96460 39140 96516 39196
rect 96516 39140 96520 39196
rect 96456 39136 96520 39140
rect 96536 39196 96600 39200
rect 96536 39140 96540 39196
rect 96540 39140 96596 39196
rect 96596 39140 96600 39196
rect 96536 39136 96600 39140
rect 96616 39196 96680 39200
rect 96616 39140 96620 39196
rect 96620 39140 96676 39196
rect 96676 39140 96680 39196
rect 96616 39136 96680 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 50296 38652 50360 38656
rect 50296 38596 50300 38652
rect 50300 38596 50356 38652
rect 50356 38596 50360 38652
rect 50296 38592 50360 38596
rect 50376 38652 50440 38656
rect 50376 38596 50380 38652
rect 50380 38596 50436 38652
rect 50436 38596 50440 38652
rect 50376 38592 50440 38596
rect 50456 38652 50520 38656
rect 50456 38596 50460 38652
rect 50460 38596 50516 38652
rect 50516 38596 50520 38652
rect 50456 38592 50520 38596
rect 50536 38652 50600 38656
rect 50536 38596 50540 38652
rect 50540 38596 50596 38652
rect 50596 38596 50600 38652
rect 50536 38592 50600 38596
rect 81016 38652 81080 38656
rect 81016 38596 81020 38652
rect 81020 38596 81076 38652
rect 81076 38596 81080 38652
rect 81016 38592 81080 38596
rect 81096 38652 81160 38656
rect 81096 38596 81100 38652
rect 81100 38596 81156 38652
rect 81156 38596 81160 38652
rect 81096 38592 81160 38596
rect 81176 38652 81240 38656
rect 81176 38596 81180 38652
rect 81180 38596 81236 38652
rect 81236 38596 81240 38652
rect 81176 38592 81240 38596
rect 81256 38652 81320 38656
rect 81256 38596 81260 38652
rect 81260 38596 81316 38652
rect 81316 38596 81320 38652
rect 81256 38592 81320 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 65656 38108 65720 38112
rect 65656 38052 65660 38108
rect 65660 38052 65716 38108
rect 65716 38052 65720 38108
rect 65656 38048 65720 38052
rect 65736 38108 65800 38112
rect 65736 38052 65740 38108
rect 65740 38052 65796 38108
rect 65796 38052 65800 38108
rect 65736 38048 65800 38052
rect 65816 38108 65880 38112
rect 65816 38052 65820 38108
rect 65820 38052 65876 38108
rect 65876 38052 65880 38108
rect 65816 38048 65880 38052
rect 65896 38108 65960 38112
rect 65896 38052 65900 38108
rect 65900 38052 65956 38108
rect 65956 38052 65960 38108
rect 65896 38048 65960 38052
rect 96376 38108 96440 38112
rect 96376 38052 96380 38108
rect 96380 38052 96436 38108
rect 96436 38052 96440 38108
rect 96376 38048 96440 38052
rect 96456 38108 96520 38112
rect 96456 38052 96460 38108
rect 96460 38052 96516 38108
rect 96516 38052 96520 38108
rect 96456 38048 96520 38052
rect 96536 38108 96600 38112
rect 96536 38052 96540 38108
rect 96540 38052 96596 38108
rect 96596 38052 96600 38108
rect 96536 38048 96600 38052
rect 96616 38108 96680 38112
rect 96616 38052 96620 38108
rect 96620 38052 96676 38108
rect 96676 38052 96680 38108
rect 96616 38048 96680 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 81016 37564 81080 37568
rect 81016 37508 81020 37564
rect 81020 37508 81076 37564
rect 81076 37508 81080 37564
rect 81016 37504 81080 37508
rect 81096 37564 81160 37568
rect 81096 37508 81100 37564
rect 81100 37508 81156 37564
rect 81156 37508 81160 37564
rect 81096 37504 81160 37508
rect 81176 37564 81240 37568
rect 81176 37508 81180 37564
rect 81180 37508 81236 37564
rect 81236 37508 81240 37564
rect 81176 37504 81240 37508
rect 81256 37564 81320 37568
rect 81256 37508 81260 37564
rect 81260 37508 81316 37564
rect 81316 37508 81320 37564
rect 81256 37504 81320 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 65656 37020 65720 37024
rect 65656 36964 65660 37020
rect 65660 36964 65716 37020
rect 65716 36964 65720 37020
rect 65656 36960 65720 36964
rect 65736 37020 65800 37024
rect 65736 36964 65740 37020
rect 65740 36964 65796 37020
rect 65796 36964 65800 37020
rect 65736 36960 65800 36964
rect 65816 37020 65880 37024
rect 65816 36964 65820 37020
rect 65820 36964 65876 37020
rect 65876 36964 65880 37020
rect 65816 36960 65880 36964
rect 65896 37020 65960 37024
rect 65896 36964 65900 37020
rect 65900 36964 65956 37020
rect 65956 36964 65960 37020
rect 65896 36960 65960 36964
rect 96376 37020 96440 37024
rect 96376 36964 96380 37020
rect 96380 36964 96436 37020
rect 96436 36964 96440 37020
rect 96376 36960 96440 36964
rect 96456 37020 96520 37024
rect 96456 36964 96460 37020
rect 96460 36964 96516 37020
rect 96516 36964 96520 37020
rect 96456 36960 96520 36964
rect 96536 37020 96600 37024
rect 96536 36964 96540 37020
rect 96540 36964 96596 37020
rect 96596 36964 96600 37020
rect 96536 36960 96600 36964
rect 96616 37020 96680 37024
rect 96616 36964 96620 37020
rect 96620 36964 96676 37020
rect 96676 36964 96680 37020
rect 96616 36960 96680 36964
rect 17908 36620 17972 36684
rect 26188 36484 26252 36548
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 81016 36476 81080 36480
rect 81016 36420 81020 36476
rect 81020 36420 81076 36476
rect 81076 36420 81080 36476
rect 81016 36416 81080 36420
rect 81096 36476 81160 36480
rect 81096 36420 81100 36476
rect 81100 36420 81156 36476
rect 81156 36420 81160 36476
rect 81096 36416 81160 36420
rect 81176 36476 81240 36480
rect 81176 36420 81180 36476
rect 81180 36420 81236 36476
rect 81236 36420 81240 36476
rect 81176 36416 81240 36420
rect 81256 36476 81320 36480
rect 81256 36420 81260 36476
rect 81260 36420 81316 36476
rect 81316 36420 81320 36476
rect 81256 36416 81320 36420
rect 17908 36212 17972 36276
rect 26188 36212 26252 36276
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 65656 35932 65720 35936
rect 65656 35876 65660 35932
rect 65660 35876 65716 35932
rect 65716 35876 65720 35932
rect 65656 35872 65720 35876
rect 65736 35932 65800 35936
rect 65736 35876 65740 35932
rect 65740 35876 65796 35932
rect 65796 35876 65800 35932
rect 65736 35872 65800 35876
rect 65816 35932 65880 35936
rect 65816 35876 65820 35932
rect 65820 35876 65876 35932
rect 65876 35876 65880 35932
rect 65816 35872 65880 35876
rect 65896 35932 65960 35936
rect 65896 35876 65900 35932
rect 65900 35876 65956 35932
rect 65956 35876 65960 35932
rect 65896 35872 65960 35876
rect 96376 35932 96440 35936
rect 96376 35876 96380 35932
rect 96380 35876 96436 35932
rect 96436 35876 96440 35932
rect 96376 35872 96440 35876
rect 96456 35932 96520 35936
rect 96456 35876 96460 35932
rect 96460 35876 96516 35932
rect 96516 35876 96520 35932
rect 96456 35872 96520 35876
rect 96536 35932 96600 35936
rect 96536 35876 96540 35932
rect 96540 35876 96596 35932
rect 96596 35876 96600 35932
rect 96536 35872 96600 35876
rect 96616 35932 96680 35936
rect 96616 35876 96620 35932
rect 96620 35876 96676 35932
rect 96676 35876 96680 35932
rect 96616 35872 96680 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 81016 35388 81080 35392
rect 81016 35332 81020 35388
rect 81020 35332 81076 35388
rect 81076 35332 81080 35388
rect 81016 35328 81080 35332
rect 81096 35388 81160 35392
rect 81096 35332 81100 35388
rect 81100 35332 81156 35388
rect 81156 35332 81160 35388
rect 81096 35328 81160 35332
rect 81176 35388 81240 35392
rect 81176 35332 81180 35388
rect 81180 35332 81236 35388
rect 81236 35332 81240 35388
rect 81176 35328 81240 35332
rect 81256 35388 81320 35392
rect 81256 35332 81260 35388
rect 81260 35332 81316 35388
rect 81316 35332 81320 35388
rect 81256 35328 81320 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 65656 34844 65720 34848
rect 65656 34788 65660 34844
rect 65660 34788 65716 34844
rect 65716 34788 65720 34844
rect 65656 34784 65720 34788
rect 65736 34844 65800 34848
rect 65736 34788 65740 34844
rect 65740 34788 65796 34844
rect 65796 34788 65800 34844
rect 65736 34784 65800 34788
rect 65816 34844 65880 34848
rect 65816 34788 65820 34844
rect 65820 34788 65876 34844
rect 65876 34788 65880 34844
rect 65816 34784 65880 34788
rect 65896 34844 65960 34848
rect 65896 34788 65900 34844
rect 65900 34788 65956 34844
rect 65956 34788 65960 34844
rect 65896 34784 65960 34788
rect 96376 34844 96440 34848
rect 96376 34788 96380 34844
rect 96380 34788 96436 34844
rect 96436 34788 96440 34844
rect 96376 34784 96440 34788
rect 96456 34844 96520 34848
rect 96456 34788 96460 34844
rect 96460 34788 96516 34844
rect 96516 34788 96520 34844
rect 96456 34784 96520 34788
rect 96536 34844 96600 34848
rect 96536 34788 96540 34844
rect 96540 34788 96596 34844
rect 96596 34788 96600 34844
rect 96536 34784 96600 34788
rect 96616 34844 96680 34848
rect 96616 34788 96620 34844
rect 96620 34788 96676 34844
rect 96676 34788 96680 34844
rect 96616 34784 96680 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 81016 34300 81080 34304
rect 81016 34244 81020 34300
rect 81020 34244 81076 34300
rect 81076 34244 81080 34300
rect 81016 34240 81080 34244
rect 81096 34300 81160 34304
rect 81096 34244 81100 34300
rect 81100 34244 81156 34300
rect 81156 34244 81160 34300
rect 81096 34240 81160 34244
rect 81176 34300 81240 34304
rect 81176 34244 81180 34300
rect 81180 34244 81236 34300
rect 81236 34244 81240 34300
rect 81176 34240 81240 34244
rect 81256 34300 81320 34304
rect 81256 34244 81260 34300
rect 81260 34244 81316 34300
rect 81316 34244 81320 34300
rect 81256 34240 81320 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 55628 30092 55692 30156
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 55812 29412 55876 29476
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 9260 27508 9324 27572
rect 55444 27236 55508 27300
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 55260 27100 55324 27164
rect 83412 26692 83476 26756
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 52684 24108 52748 24172
rect 55260 24108 55324 24172
rect 83044 24108 83108 24172
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 53052 23836 53116 23900
rect 55444 23836 55508 23900
rect 15884 23488 15948 23492
rect 15884 23432 15898 23488
rect 15898 23432 15948 23488
rect 15884 23428 15948 23432
rect 31892 23428 31956 23492
rect 52316 23428 52380 23492
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 55260 23292 55324 23356
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 9996 22808 10060 22812
rect 9996 22752 10010 22808
rect 10010 22752 10060 22808
rect 9996 22748 10060 22752
rect 54524 22748 54588 22812
rect 83964 22748 84028 22812
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 19196 22068 19260 22132
rect 52316 22068 52380 22132
rect 55628 22068 55692 22132
rect 19380 21932 19444 21996
rect 31892 21932 31956 21996
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 14596 21388 14660 21452
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 24164 20708 24228 20772
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 56180 20028 56244 20092
rect 83228 20028 83292 20092
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 27844 18668 27908 18732
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 22692 17308 22756 17372
rect 82860 17172 82924 17236
rect 83228 17172 83292 17236
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 10548 16688 10612 16692
rect 10548 16632 10562 16688
rect 10562 16632 10612 16688
rect 10548 16628 10612 16632
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 21956 16008 22020 16012
rect 21956 15952 21970 16008
rect 21970 15952 22020 16008
rect 21956 15948 22020 15952
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 24900 15328 24964 15332
rect 24900 15272 24914 15328
rect 24914 15272 24964 15328
rect 24900 15268 24964 15272
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 82860 14724 82924 14788
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 24164 13908 24228 13972
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
<< metal4 >>
rect 4208 43552 4528 44112
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43014 4528 43488
rect 4208 42778 4250 43014
rect 4486 42778 4528 43014
rect 4208 42694 4528 42778
rect 4208 42464 4250 42694
rect 4486 42464 4528 42694
rect 4208 42400 4216 42464
rect 4280 42400 4296 42458
rect 4360 42400 4376 42458
rect 4440 42400 4456 42458
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 19568 44096 19888 44112
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 17907 36684 17973 36685
rect 17907 36620 17908 36684
rect 17972 36620 17973 36684
rect 17907 36619 17973 36620
rect 17910 36277 17970 36619
rect 19568 36480 19888 37504
rect 34928 43552 35248 44112
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43014 35248 43488
rect 34928 42778 34970 43014
rect 35206 42778 35248 43014
rect 34928 42694 35248 42778
rect 34928 42464 34970 42694
rect 35206 42464 35248 42694
rect 34928 42400 34936 42464
rect 35000 42400 35016 42458
rect 35080 42400 35096 42458
rect 35160 42400 35176 42458
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 26187 36548 26253 36549
rect 26187 36484 26188 36548
rect 26252 36484 26253 36548
rect 26187 36483 26253 36484
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 17907 36276 17973 36277
rect 17907 36212 17908 36276
rect 17972 36212 17973 36276
rect 17907 36211 17973 36212
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 19568 35392 19888 36416
rect 26190 36277 26250 36483
rect 26187 36276 26253 36277
rect 26187 36212 26188 36276
rect 26252 36212 26253 36276
rect 26187 36211 26253 36212
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33880 35248 34784
rect 50288 44096 50608 44112
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 43008 50608 44032
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 41920 50608 42944
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 40832 50608 41856
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 39744 50608 40768
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 38656 50608 39680
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 37568 50608 38592
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33880 50608 34240
rect 65648 43552 65968 44112
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43014 65968 43488
rect 65648 42778 65690 43014
rect 65926 42778 65968 43014
rect 65648 42694 65968 42778
rect 65648 42464 65690 42694
rect 65926 42464 65968 42694
rect 65648 42400 65656 42464
rect 65720 42400 65736 42458
rect 65800 42400 65816 42458
rect 65880 42400 65896 42458
rect 65960 42400 65968 42464
rect 65648 41376 65968 42400
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 40288 65968 41312
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 39200 65968 40224
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 38112 65968 39136
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 37024 65968 38048
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 35936 65968 36960
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 34848 65968 35872
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 33880 65968 34784
rect 81008 44096 81328 44112
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 43008 81328 44032
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 41920 81328 42944
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 40832 81328 41856
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 39744 81328 40768
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 38656 81328 39680
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 37568 81328 38592
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 36480 81328 37504
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 35392 81328 36416
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 34304 81328 35328
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 33880 81328 34240
rect 96368 43552 96688 44112
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43014 96688 43488
rect 96368 42778 96410 43014
rect 96646 42778 96688 43014
rect 96368 42694 96688 42778
rect 96368 42464 96410 42694
rect 96646 42464 96688 42694
rect 96368 42400 96376 42464
rect 96440 42400 96456 42458
rect 96520 42400 96536 42458
rect 96600 42400 96616 42458
rect 96680 42400 96688 42464
rect 96368 41376 96688 42400
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 40288 96688 41312
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 39200 96688 40224
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 38112 96688 39136
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 37024 96688 38048
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 35936 96688 36960
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 34848 96688 35872
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 33880 96688 34784
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 55627 30156 55693 30157
rect 55627 30092 55628 30156
rect 55692 30092 55693 30156
rect 55627 30091 55693 30092
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 19568 26688 19888 27712
rect 55262 27165 55322 27422
rect 55443 27300 55509 27301
rect 55443 27236 55444 27300
rect 55508 27236 55509 27300
rect 55443 27235 55509 27236
rect 55259 27164 55325 27165
rect 55259 27100 55260 27164
rect 55324 27100 55325 27164
rect 55259 27099 55325 27100
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25014 19888 25536
rect 19568 24778 19610 25014
rect 19846 24778 19888 25014
rect 19568 24694 19888 24778
rect 19568 24512 19610 24694
rect 19846 24512 19888 24694
rect 19568 24448 19576 24512
rect 19640 24448 19656 24458
rect 19720 24448 19736 24458
rect 19800 24448 19816 24458
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 52683 24172 52749 24173
rect 52683 24108 52684 24172
rect 52748 24108 52749 24172
rect 52683 24107 52749 24108
rect 55259 24172 55325 24173
rect 55259 24108 55260 24172
rect 55324 24108 55325 24172
rect 55259 24107 55325 24108
rect 31891 23492 31957 23493
rect 31891 23428 31892 23492
rect 31956 23428 31957 23492
rect 31891 23427 31957 23428
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 19568 22336 19888 23360
rect 31894 22898 31954 23427
rect 52686 22898 52746 24107
rect 53051 23900 53117 23901
rect 53051 23836 53052 23900
rect 53116 23836 53117 23900
rect 53051 23835 53117 23836
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19195 22132 19261 22133
rect 19195 22068 19196 22132
rect 19260 22130 19261 22132
rect 19260 22070 19442 22130
rect 19260 22068 19261 22070
rect 19195 22067 19261 22068
rect 19382 21997 19442 22070
rect 19379 21996 19445 21997
rect 19379 21932 19380 21996
rect 19444 21932 19445 21996
rect 19379 21931 19445 21932
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 30974 19498 31034 22662
rect 31891 21996 31957 21997
rect 31891 21932 31892 21996
rect 31956 21932 31957 21996
rect 31891 21931 31957 21932
rect 31894 20090 31954 21931
rect 34470 20090 34530 21982
rect 31894 20030 34530 20090
rect 53054 19498 53114 23835
rect 55262 23357 55322 24107
rect 55446 23901 55506 27235
rect 55443 23900 55509 23901
rect 55443 23836 55444 23900
rect 55508 23836 55509 23900
rect 55443 23835 55509 23836
rect 55259 23356 55325 23357
rect 55259 23292 55260 23356
rect 55324 23292 55325 23356
rect 55259 23291 55325 23292
rect 54523 22812 54589 22813
rect 54523 22748 54524 22812
rect 54588 22748 54589 22812
rect 54523 22747 54589 22748
rect 54526 20178 54586 22747
rect 55630 22133 55690 30091
rect 55811 29476 55877 29477
rect 55811 29412 55812 29476
rect 55876 29412 55877 29476
rect 55811 29411 55877 29412
rect 55627 22132 55693 22133
rect 55627 22068 55628 22132
rect 55692 22068 55693 22132
rect 55627 22067 55693 22068
rect 55814 21538 55874 29411
rect 83411 26756 83477 26757
rect 83411 26692 83412 26756
rect 83476 26692 83477 26756
rect 83411 26691 83477 26692
rect 83043 24172 83109 24173
rect 83043 24108 83044 24172
rect 83108 24108 83109 24172
rect 83043 24107 83109 24108
rect 56179 20092 56245 20093
rect 56179 20028 56180 20092
rect 56244 20028 56245 20092
rect 56179 20027 56245 20028
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 56182 18818 56242 20027
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 83046 17370 83106 24107
rect 83227 20092 83293 20093
rect 83227 20028 83228 20092
rect 83292 20028 83293 20092
rect 83227 20027 83293 20028
rect 82642 17310 83106 17370
rect 83230 17237 83290 20027
rect 82859 17236 82925 17237
rect 82859 17172 82860 17236
rect 82924 17172 82925 17236
rect 82859 17171 82925 17172
rect 83227 17236 83293 17237
rect 83227 17172 83228 17236
rect 83292 17172 83293 17236
rect 83227 17171 83293 17172
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7014 4528 7584
rect 4208 6778 4250 7014
rect 4486 6778 4528 7014
rect 4208 6694 4528 6778
rect 4208 6560 4250 6694
rect 4486 6560 4528 6694
rect 4208 6496 4216 6560
rect 4520 6496 4528 6560
rect 4208 6458 4250 6496
rect 4486 6458 4528 6496
rect 4208 5472 4528 6458
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 82862 15418 82922 17171
rect 83414 16778 83474 26691
rect 83963 22812 84029 22813
rect 83963 22748 83964 22812
rect 84028 22748 84029 22812
rect 83963 22747 84029 22748
rect 83966 16098 84026 22747
rect 82859 14788 82925 14789
rect 82859 14724 82860 14788
rect 82924 14724 82925 14788
rect 82859 14723 82925 14724
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 82862 14058 82922 14723
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
<< via4 >>
rect 4250 42778 4486 43014
rect 4250 42464 4486 42694
rect 4250 42458 4280 42464
rect 4280 42458 4296 42464
rect 4296 42458 4360 42464
rect 4360 42458 4376 42464
rect 4376 42458 4440 42464
rect 4440 42458 4456 42464
rect 4456 42458 4486 42464
rect 34970 42778 35206 43014
rect 34970 42464 35206 42694
rect 34970 42458 35000 42464
rect 35000 42458 35016 42464
rect 35016 42458 35080 42464
rect 35080 42458 35096 42464
rect 35096 42458 35160 42464
rect 35160 42458 35176 42464
rect 35176 42458 35206 42464
rect 65690 42778 65926 43014
rect 65690 42464 65926 42694
rect 65690 42458 65720 42464
rect 65720 42458 65736 42464
rect 65736 42458 65800 42464
rect 65800 42458 65816 42464
rect 65816 42458 65880 42464
rect 65880 42458 65896 42464
rect 65896 42458 65926 42464
rect 96410 42778 96646 43014
rect 96410 42464 96646 42694
rect 96410 42458 96440 42464
rect 96440 42458 96456 42464
rect 96456 42458 96520 42464
rect 96520 42458 96536 42464
rect 96536 42458 96600 42464
rect 96600 42458 96616 42464
rect 96616 42458 96646 42464
rect 9174 27572 9410 27658
rect 9174 27508 9260 27572
rect 9260 27508 9324 27572
rect 9324 27508 9410 27572
rect 9174 27422 9410 27508
rect 55174 27422 55410 27658
rect 19610 24778 19846 25014
rect 19610 24512 19846 24694
rect 19610 24458 19640 24512
rect 19640 24458 19656 24512
rect 19656 24458 19720 24512
rect 19720 24458 19736 24512
rect 19736 24458 19800 24512
rect 19800 24458 19816 24512
rect 19816 24458 19846 24512
rect 15798 23492 16034 23578
rect 15798 23428 15884 23492
rect 15884 23428 15948 23492
rect 15948 23428 16034 23492
rect 15798 23342 16034 23428
rect 52230 23492 52466 23578
rect 52230 23428 52316 23492
rect 52316 23428 52380 23492
rect 52380 23428 52466 23492
rect 9910 22812 10146 22898
rect 9910 22748 9996 22812
rect 9996 22748 10060 22812
rect 10060 22748 10146 22812
rect 9910 22662 10146 22748
rect 52230 23342 52466 23428
rect 30886 22662 31122 22898
rect 31806 22662 32042 22898
rect 52598 22662 52834 22898
rect 14510 21452 14746 21538
rect 14510 21388 14596 21452
rect 14596 21388 14660 21452
rect 14660 21388 14746 21452
rect 14510 21302 14746 21388
rect 24078 20772 24314 20858
rect 24078 20708 24164 20772
rect 24164 20708 24228 20772
rect 24228 20708 24314 20772
rect 24078 20622 24314 20708
rect 34382 21982 34618 22218
rect 52230 22132 52466 22218
rect 52230 22068 52316 22132
rect 52316 22068 52380 22132
rect 52380 22068 52466 22132
rect 52230 21982 52466 22068
rect 55726 21302 55962 21538
rect 54438 19942 54674 20178
rect 30886 19262 31122 19498
rect 52966 19262 53202 19498
rect 27758 18732 27994 18818
rect 27758 18668 27844 18732
rect 27844 18668 27908 18732
rect 27908 18668 27994 18732
rect 27758 18582 27994 18668
rect 56094 18582 56330 18818
rect 22606 17372 22842 17458
rect 22606 17308 22692 17372
rect 22692 17308 22756 17372
rect 22756 17308 22842 17372
rect 22606 17222 22842 17308
rect 82406 17222 82642 17458
rect 10462 16692 10698 16778
rect 10462 16628 10548 16692
rect 10548 16628 10612 16692
rect 10612 16628 10698 16692
rect 10462 16542 10698 16628
rect 4250 6778 4486 7014
rect 4250 6560 4486 6694
rect 4250 6496 4280 6560
rect 4280 6496 4296 6560
rect 4296 6496 4360 6560
rect 4360 6496 4376 6560
rect 4376 6496 4440 6560
rect 4440 6496 4456 6560
rect 4456 6496 4486 6560
rect 4250 6458 4486 6496
rect 21870 16012 22106 16098
rect 21870 15948 21956 16012
rect 21956 15948 22020 16012
rect 22020 15948 22106 16012
rect 21870 15862 22106 15948
rect 83326 16542 83562 16778
rect 83878 15862 84114 16098
rect 24814 15332 25050 15418
rect 24814 15268 24900 15332
rect 24900 15268 24964 15332
rect 24964 15268 25050 15332
rect 24814 15182 25050 15268
rect 82774 15182 83010 15418
rect 24078 13972 24314 14058
rect 24078 13908 24164 13972
rect 24164 13908 24228 13972
rect 24228 13908 24314 13972
rect 24078 13822 24314 13908
rect 82774 13822 83010 14058
<< metal5 >>
rect 4208 43036 4528 43038
rect 34928 43036 35248 43038
rect 65648 43036 65968 43038
rect 96368 43036 96688 43038
rect 1104 43014 111136 43036
rect 1104 42778 4250 43014
rect 4486 42778 34970 43014
rect 35206 42778 65690 43014
rect 65926 42778 96410 43014
rect 96646 42778 111136 43014
rect 1104 42694 111136 42778
rect 1104 42458 4250 42694
rect 4486 42458 34970 42694
rect 35206 42458 65690 42694
rect 65926 42458 96410 42694
rect 96646 42458 111136 42694
rect 1104 42436 111136 42458
rect 4208 42434 4528 42436
rect 34928 42434 35248 42436
rect 65648 42434 65968 42436
rect 96368 42434 96688 42436
rect 9132 27658 55452 27700
rect 9132 27422 9174 27658
rect 9410 27422 55174 27658
rect 55410 27422 55452 27658
rect 9132 27380 55452 27422
rect 19568 25036 19888 25038
rect 1104 25014 111136 25036
rect 1104 24778 19610 25014
rect 19846 24778 111136 25014
rect 1104 24694 111136 24778
rect 1104 24458 19610 24694
rect 19846 24458 111136 24694
rect 1104 24436 111136 24458
rect 19568 24434 19888 24436
rect 34340 23708 38892 24028
rect 34340 23620 34660 23708
rect 15756 23578 34660 23620
rect 15756 23342 15798 23578
rect 16034 23342 34660 23578
rect 15756 23300 34660 23342
rect 38572 23620 38892 23708
rect 38572 23578 52508 23620
rect 38572 23342 52230 23578
rect 52466 23342 52508 23578
rect 38572 23300 52508 23342
rect 9868 22898 31164 22940
rect 9868 22662 9910 22898
rect 10146 22662 30886 22898
rect 31122 22662 31164 22898
rect 9868 22620 31164 22662
rect 31764 22898 52876 22940
rect 31764 22662 31806 22898
rect 32042 22662 52598 22898
rect 52834 22662 52876 22898
rect 31764 22620 52876 22662
rect 34340 22218 52508 22260
rect 34340 21982 34382 22218
rect 34618 21982 52230 22218
rect 52466 21982 52508 22218
rect 34340 21940 52508 21982
rect 14468 21538 56004 21580
rect 14468 21302 14510 21538
rect 14746 21302 55726 21538
rect 55962 21302 56004 21538
rect 14468 21260 56004 21302
rect 24036 20858 43308 20900
rect 24036 20622 24078 20858
rect 24314 20622 43308 20858
rect 24036 20580 43308 20622
rect 42988 20220 43308 20580
rect 42988 20178 54716 20220
rect 42988 19942 54438 20178
rect 54674 19942 54716 20178
rect 42988 19900 54716 19942
rect 30844 19498 53244 19540
rect 30844 19262 30886 19498
rect 31122 19262 52966 19498
rect 53202 19262 53244 19498
rect 30844 19220 53244 19262
rect 27716 18818 56372 18860
rect 27716 18582 27758 18818
rect 27994 18582 56094 18818
rect 56330 18582 56372 18818
rect 27716 18540 56372 18582
rect 22564 17458 82684 17500
rect 22564 17222 22606 17458
rect 22842 17222 82406 17458
rect 82642 17222 82684 17458
rect 22564 17180 82684 17222
rect 10420 16778 83604 16820
rect 10420 16542 10462 16778
rect 10698 16542 83326 16778
rect 83562 16542 83604 16778
rect 10420 16500 83604 16542
rect 21828 16098 84156 16140
rect 21828 15862 21870 16098
rect 22106 15862 83878 16098
rect 84114 15862 84156 16098
rect 21828 15820 84156 15862
rect 24772 15418 83052 15460
rect 24772 15182 24814 15418
rect 25050 15182 82774 15418
rect 83010 15182 83052 15418
rect 24772 15140 83052 15182
rect 24036 14058 83052 14100
rect 24036 13822 24078 14058
rect 24314 13822 82774 14058
rect 83010 13822 83052 14058
rect 24036 13780 83052 13822
rect 4208 7036 4528 7038
rect 1104 7014 111136 7036
rect 1104 6778 4250 7014
rect 4486 6778 111136 7014
rect 1104 6694 111136 6778
rect 1104 6458 4250 6694
rect 4486 6458 111136 6694
rect 1104 6436 111136 6458
rect 4208 6434 4528 6436
use sky130_fd_sc_hd__decap_8  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2484 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607194113
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607194113
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1607194113
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607194113
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1483_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3312 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_47
timestamp 1607194113
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607194113
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__D
timestamp 1607194113
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1607194113
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607194113
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1607194113
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1607194113
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1607194113
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607194113
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1607194113
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1607194113
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607194113
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1607194113
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607194113
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1607194113
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1607194113
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607194113
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1607194113
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1607194113
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1607194113
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1607194113
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1607194113
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607194113
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1607194113
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1607194113
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1607194113
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607194113
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1607194113
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1607194113
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1607194113
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1607194113
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1607194113
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1607194113
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1607194113
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1607194113
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607194113
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1607194113
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1607194113
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1607194113
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1607194113
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607194113
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1607194113
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1607194113
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1607194113
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1607194113
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1607194113
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607194113
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607194113
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607194113
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607194113
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607194113
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1607194113
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607194113
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607194113
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607194113
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607194113
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1607194113
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1607194113
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1607194113
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1607194113
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1607194113
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1607194113
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1607194113
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1607194113
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1607194113
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1607194113
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1607194113
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1607194113
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1607194113
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1607194113
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1607194113
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1607194113
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1607194113
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607194113
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607194113
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1484_
timestamp 1607194113
transform 1 0 2852 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__D
timestamp 1607194113
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_54
timestamp 1607194113
transform 1 0 6072 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_42
timestamp 1607194113
transform 1 0 4968 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__CLK
timestamp 1607194113
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1607194113
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1607194113
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1607194113
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1607194113
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1607194113
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1607194113
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1607194113
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1607194113
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1607194113
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1607194113
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1607194113
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1607194113
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1607194113
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1607194113
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1607194113
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1607194113
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1607194113
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1607194113
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1607194113
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1607194113
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607194113
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607194113
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607194113
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607194113
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607194113
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1607194113
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_44
timestamp 1607194113
transform 1 0 5152 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1485_
timestamp 1607194113
transform 1 0 5888 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_73
timestamp 1607194113
transform 1 0 7820 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__CLK
timestamp 1607194113
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1607194113
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1607194113
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1607194113
transform 1 0 8924 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1607194113
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1607194113
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1607194113
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1607194113
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1607194113
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1607194113
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1607194113
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1607194113
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1607194113
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1607194113
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1607194113
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1607194113
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1607194113
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1607194113
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1607194113
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1607194113
transform 1 0 2484 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607194113
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607194113
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1486_
timestamp 1607194113
transform 1 0 2576 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_5_37
timestamp 1607194113
transform 1 0 4508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__CLK
timestamp 1607194113
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_49
timestamp 1607194113
transform 1 0 5612 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1607194113
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1607194113
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607194113
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1607194113
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1607194113
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1607194113
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1607194113
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1607194113
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607194113
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1607194113
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1607194113
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1607194113
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1607194113
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1607194113
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607194113
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1607194113
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1607194113
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1607194113
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607194113
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1607194113
transform 1 0 2484 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607194113
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1607194113
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607194113
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607194113
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607194113
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1487_
timestamp 1607194113
transform 1 0 2576 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_7_37
timestamp 1607194113
transform 1 0 4508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1607194113
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1607194113
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__CLK
timestamp 1607194113
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607194113
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_49
timestamp 1607194113
transform 1 0 5612 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1607194113
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1607194113
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1607194113
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607194113
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1342_
timestamp 1607194113
transform 1 0 6808 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_7_83
timestamp 1607194113
transform 1 0 8740 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1607194113
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1607194113
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__CLK
timestamp 1607194113
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607194113
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1341_
timestamp 1607194113
transform 1 0 9844 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_7_116
timestamp 1607194113
transform 1 0 11776 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1607194113
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1607194113
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__CLK
timestamp 1607194113
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1607194113
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1607194113
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1607194113
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607194113
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:4.inst.g_clkdly15_2.dly $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13708 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_158
timestamp 1607194113
transform 1 0 15640 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_146
timestamp 1607194113
transform 1 0 14536 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1607194113
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1607194113
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607194113
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_170
timestamp 1607194113
transform 1 0 16744 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1607194113
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1607194113
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1607194113
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1607194113
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1607194113
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1607194113
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607194113
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1607194113
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1607194113
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1607194113
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607194113
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1607194113
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1607194113
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1607194113
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1607194113
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607194113
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1607194113
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607194113
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607194113
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1607194113
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607194113
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:6.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_59
timestamp 1607194113
transform 1 0 6532 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1607194113
transform 1 0 5980 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1607194113
transform 1 0 4876 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_69
timestamp 1607194113
transform 1 0 7452 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:5.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 6624 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1607194113
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1607194113
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_81
timestamp 1607194113
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607194113
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_105
timestamp 1607194113
transform 1 0 10764 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1333_
timestamp 1607194113
transform 1 0 11316 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_8_132
timestamp 1607194113
transform 1 0 13248 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__CLK
timestamp 1607194113
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1607194113
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1607194113
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_144
timestamp 1607194113
transform 1 0 14352 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607194113
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_166
timestamp 1607194113
transform 1 0 16376 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1332_
timestamp 1607194113
transform 1 0 16652 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1607194113
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__CLK
timestamp 1607194113
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1607194113
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1607194113
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607194113
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1607194113
transform 1 0 21988 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__CLK
timestamp 1607194113
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1339_
timestamp 1607194113
transform 1 0 22540 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_9_15
timestamp 1607194113
transform 1 0 2484 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607194113
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607194113
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1343_
timestamp 1607194113
transform 1 0 3036 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_9_54
timestamp 1607194113
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1607194113
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__CLK
timestamp 1607194113
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp 1607194113
transform 1 0 7544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1607194113
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1607194113
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607194113
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1334_
timestamp 1607194113
transform 1 0 7636 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_92
timestamp 1607194113
transform 1 0 9568 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__CLK
timestamp 1607194113
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1607194113
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_104
timestamp 1607194113
transform 1 0 10672 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1607194113
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1607194113
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607194113
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_153
timestamp 1607194113
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_147
timestamp 1607194113
transform 1 0 14628 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1607194113
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1340_
timestamp 1607194113
transform 1 0 15456 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1607194113
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1607194113
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1607194113
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607194113
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1607194113
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_233
timestamp 1607194113
transform 1 0 22540 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1607194113
transform 1 0 21344 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:3.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 21712 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_241
timestamp 1607194113
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607194113
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1607194113
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607194113
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607194113
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1607194113
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1607194113
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607194113
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1335_
timestamp 1607194113
transform 1 0 4140 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1607194113
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__CLK
timestamp 1607194113
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_78
timestamp 1607194113
transform 1 0 8280 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1607194113
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1607194113
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1607194113
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607194113
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_105
timestamp 1607194113
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1446_
timestamp 1607194113
transform 1 0 10856 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_127
timestamp 1607194113
transform 1 0 12788 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__CLK
timestamp 1607194113
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_154
timestamp 1607194113
transform 1 0 15272 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1607194113
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_139
timestamp 1607194113
transform 1 0 13892 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607194113
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_162
timestamp 1607194113
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1445_
timestamp 1607194113
transform 1 0 16100 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_196
timestamp 1607194113
transform 1 0 19136 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1607194113
transform 1 0 18032 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__CLK
timestamp 1607194113
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1607194113
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1607194113
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607194113
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_237
timestamp 1607194113
transform 1 0 22908 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_227
timestamp 1607194113
transform 1 0 21988 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:2.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 22080 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__CLK
timestamp 1607194113
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1607194113
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607194113
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607194113
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1488_
timestamp 1607194113
transform 1 0 2576 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1607194113
transform 1 0 4508 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__CLK
timestamp 1607194113
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_49
timestamp 1607194113
transform 1 0 5612 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1607194113
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607194113
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1447_
timestamp 1607194113
transform 1 0 7544 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_11_91
timestamp 1607194113
transform 1 0 9476 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__CLK
timestamp 1607194113
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 10028 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1607194113
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_111
timestamp 1607194113
transform 1 0 11316 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_130
timestamp 1607194113
transform 1 0 13064 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607194113
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 12420 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_11_154
timestamp 1607194113
transform 1 0 15272 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_142
timestamp 1607194113
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1607194113
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 1607194113
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1166_
timestamp 1607194113
transform 1 0 15916 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_11_198
timestamp 1607194113
transform 1 0 19320 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607194113
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1167_
timestamp 1607194113
transform 1 0 18032 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_11_216
timestamp 1607194113
transform 1 0 20976 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_210
timestamp 1607194113
transform 1 0 20424 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1338_
timestamp 1607194113
transform 1 0 21068 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_11_238
timestamp 1607194113
transform 1 0 23000 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__CLK
timestamp 1607194113
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607194113
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1607194113
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607194113
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607194113
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1607194113
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1607194113
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607194113
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1607194113
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1607194113
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1607194113
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1607194113
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1607194113
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607194113
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_111
timestamp 1607194113
transform 1 0 11316 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_105
timestamp 1607194113
transform 1 0 10764 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _1165_
timestamp 1607194113
transform 1 0 11408 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_12_126
timestamp 1607194113
transform 1 0 12696 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0983_
timestamp 1607194113
transform 1 0 13432 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1607194113
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1607194113
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A
timestamp 1607194113
transform 1 0 15640 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607194113
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_160
timestamp 1607194113
transform 1 0 15824 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1444_
timestamp 1607194113
transform 1 0 16560 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_12_189
timestamp 1607194113
transform 1 0 18492 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__CLK
timestamp 1607194113
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1607194113
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1607194113
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1607194113
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607194113
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_231
timestamp 1607194113
transform 1 0 22356 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_227
timestamp 1607194113
transform 1 0 21988 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__CLK
timestamp 1607194113
transform 1 0 22632 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 22080 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1330_
timestamp 1607194113
transform 1 0 22816 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607194113
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607194113
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_15
timestamp 1607194113
transform 1 0 2484 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607194113
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607194113
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607194113
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1489_
timestamp 1607194113
transform 1 0 2576 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1607194113
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607194113
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_37
timestamp 1607194113
transform 1 0 4508 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__CLK
timestamp 1607194113
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607194113
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_44
timestamp 1607194113
transform 1 0 5152 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_49
timestamp 1607194113
transform 1 0 5612 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1448_
timestamp 1607194113
transform 1 0 5704 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_14_71
timestamp 1607194113
transform 1 0 7636 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_78
timestamp 1607194113
transform 1 0 8280 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__CLK
timestamp 1607194113
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A2
timestamp 1607194113
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607194113
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1162_
timestamp 1607194113
transform 1 0 6808 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _0960_
timestamp 1607194113
transform 1 0 8188 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1607194113
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1607194113
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_91
timestamp 1607194113
transform 1 0 9476 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607194113
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 10212 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0969_
timestamp 1607194113
transform 1 0 8832 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_14_105
timestamp 1607194113
transform 1 0 10764 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_117
timestamp 1607194113
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_105
timestamp 1607194113
transform 1 0 10764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A
timestamp 1607194113
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1607194113
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 11500 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_136
timestamp 1607194113
transform 1 0 13616 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_124
timestamp 1607194113
transform 1 0 12512 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_132
timestamp 1607194113
transform 1 0 13248 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1607194113
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A
timestamp 1607194113
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607194113
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0990_
timestamp 1607194113
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_148
timestamp 1607194113
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1607194113
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_144
timestamp 1607194113
transform 1 0 14352 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__CLK
timestamp 1607194113
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607194113
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1443_
timestamp 1607194113
transform 1 0 15272 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _1168_
timestamp 1607194113
transform 1 0 15640 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_14_173
timestamp 1607194113
transform 1 0 17020 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_172
timestamp 1607194113
transform 1 0 16928 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1607194113
transform 1 0 19228 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_185
timestamp 1607194113
transform 1 0 18124 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1607194113
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1607194113
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1607194113
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607194113
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1607194113
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1607194113
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1607194113
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607194113
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_238
timestamp 1607194113
transform 1 0 23000 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_226
timestamp 1607194113
transform 1 0 21896 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1607194113
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1607194113
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly_A
timestamp 1607194113
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:1.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 21620 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607194113
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1607194113
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607194113
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607194113
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1490_
timestamp 1607194113
transform 1 0 2576 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1607194113
transform 1 0 4508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__CLK
timestamp 1607194113
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_49
timestamp 1607194113
transform 1 0 5612 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_79
timestamp 1607194113
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1607194113
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__C
timestamp 1607194113
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607194113
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0968_
timestamp 1607194113
transform 1 0 7360 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_91
timestamp 1607194113
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1607194113
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_103
timestamp 1607194113
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_135
timestamp 1607194113
transform 1 0 13524 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1607194113
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1607194113
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607194113
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1169_
timestamp 1607194113
transform 1 0 13800 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_15_154
timestamp 1607194113
transform 1 0 15272 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B1
timestamp 1607194113
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_176
timestamp 1607194113
transform 1 0 17296 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_164
timestamp 1607194113
transform 1 0 16192 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1161_
timestamp 1607194113
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1607194113
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1607194113
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1607194113
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607194113
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_216
timestamp 1607194113
transform 1 0 20976 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_208
timestamp 1607194113
transform 1 0 20240 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1337_
timestamp 1607194113
transform 1 0 21068 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_15_238
timestamp 1607194113
transform 1 0 23000 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__CLK
timestamp 1607194113
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607194113
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1607194113
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607194113
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607194113
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1607194113
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1607194113
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607194113
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_50
timestamp 1607194113
transform 1 0 5704 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1607194113
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6440 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1607194113
transform 1 0 5336 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1607194113
transform 1 0 7084 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0975_
timestamp 1607194113
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1607194113
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_84
timestamp 1607194113
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__C
timestamp 1607194113
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607194113
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_117
timestamp 1607194113
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1607194113
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_123
timestamp 1607194113
transform 1 0 12420 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1442_
timestamp 1607194113
transform 1 0 12696 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1607194113
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607194113
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1170_
timestamp 1607194113
transform 1 0 15272 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_16_170
timestamp 1607194113
transform 1 0 16744 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__B1
timestamp 1607194113
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 1607194113
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_182
timestamp 1607194113
transform 1 0 17848 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1328_
timestamp 1607194113
transform 1 0 18308 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1607194113
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_208
timestamp 1607194113
transform 1 0 20240 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__CLK
timestamp 1607194113
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607194113
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1329_
timestamp 1607194113
transform 1 0 21988 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_17_15
timestamp 1607194113
transform 1 0 2484 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607194113
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607194113
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1491_
timestamp 1607194113
transform 1 0 2576 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1607194113
transform 1 0 4508 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__CLK
timestamp 1607194113
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_49
timestamp 1607194113
transform 1 0 5612 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_71
timestamp 1607194113
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__B
timestamp 1607194113
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607194113
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1002_
timestamp 1607194113
transform 1 0 8188 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0956_
timestamp 1607194113
transform 1 0 6808 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_96
timestamp 1607194113
transform 1 0 9936 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_84
timestamp 1607194113
transform 1 0 8832 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_108
timestamp 1607194113
transform 1 0 11040 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1607194113
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1607194113
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__CLK
timestamp 1607194113
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607194113
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1441_
timestamp 1607194113
transform 1 0 12880 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1607194113
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1607194113
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1607194113
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1607194113
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607194113
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1336_
timestamp 1607194113
transform 1 0 18584 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_213
timestamp 1607194113
transform 1 0 20700 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__CLK
timestamp 1607194113
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__D
timestamp 1607194113
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1607194113
transform 1 0 22908 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1607194113
transform 1 0 21804 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1607194113
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607194113
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607194113
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607194113
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607194113
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1607194113
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607194113
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607194113
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_56
timestamp 1607194113
transform 1 0 6256 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1607194113
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1360_
timestamp 1607194113
transform 1 0 6348 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_78
timestamp 1607194113
transform 1 0 8280 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__CLK
timestamp 1607194113
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1607194113
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1607194113
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607194113
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1607194113
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 1607194113
transform 1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_138
timestamp 1607194113
transform 1 0 13800 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1607194113
transform 1 0 13156 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_122
timestamp 1607194113
transform 1 0 12328 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1607194113
transform 1 0 12144 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk_i
timestamp 1607194113
transform 1 0 12880 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1607194113
transform 1 0 13524 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_154
timestamp 1607194113
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1607194113
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607194113
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_162
timestamp 1607194113
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__B1
timestamp 1607194113
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 16284 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_193
timestamp 1607194113
transform 1 0 18860 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_181
timestamp 1607194113
transform 1 0 17756 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1607194113
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1607194113
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_205
timestamp 1607194113
transform 1 0 19964 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607194113
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_235
timestamp 1607194113
transform 1 0 22724 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_227
timestamp 1607194113
transform 1 0 21988 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1607194113
transform 1 0 22816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_241
timestamp 1607194113
transform 1 0 23276 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A
timestamp 1607194113
transform 1 0 23092 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607194113
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607194113
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_15
timestamp 1607194113
transform 1 0 2484 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607194113
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607194113
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607194113
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1492_
timestamp 1607194113
transform 1 0 2576 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1607194113
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607194113
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1607194113
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__CLK
timestamp 1607194113
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__D
timestamp 1607194113
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607194113
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_54
timestamp 1607194113
transform 1 0 6072 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_44
timestamp 1607194113
transform 1 0 5152 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1607194113
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__B1
timestamp 1607194113
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1296_
timestamp 1607194113
transform 1 0 5704 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_78
timestamp 1607194113
transform 1 0 8280 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_78
timestamp 1607194113
transform 1 0 8280 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B1
timestamp 1607194113
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607194113
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1301_
timestamp 1607194113
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1299_
timestamp 1607194113
transform 1 0 6808 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1607194113
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1607194113
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_95
timestamp 1607194113
transform 1 0 9844 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_89
timestamp 1607194113
transform 1 0 9292 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1607194113
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__B1
timestamp 1607194113
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607194113
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1303_
timestamp 1607194113
transform 1 0 10120 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1607194113
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1607194113
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1607194113
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1359_
timestamp 1607194113
transform 1 0 10948 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_134
timestamp 1607194113
transform 1 0 13432 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_128
timestamp 1607194113
transform 1 0 12880 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1607194113
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1607194113
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_i_A
timestamp 1607194113
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk_i
timestamp 1607194113
transform 1 0 13524 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607194113
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1284_
timestamp 1607194113
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1607194113
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1607194113
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_140
timestamp 1607194113
transform 1 0 13984 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1607194113
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1607194113
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607194113
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_166
timestamp 1607194113
transform 1 0 16376 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1607194113
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_163
timestamp 1607194113
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__CLK
timestamp 1607194113
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1365_
timestamp 1607194113
transform 1 0 16836 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1607194113
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_189
timestamp 1607194113
transform 1 0 18492 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A
timestamp 1607194113
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607194113
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1607194113
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1607194113
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1607194113
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_217
timestamp 1607194113
transform 1 0 21068 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_213
timestamp 1607194113
transform 1 0 20700 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_201
timestamp 1607194113
transform 1 0 19596 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B1
timestamp 1607194113
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607194113
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1607194113
transform 1 0 21988 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_236
timestamp 1607194113
transform 1 0 22816 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1367_
timestamp 1607194113
transform 1 0 22356 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1287_
timestamp 1607194113
transform 1 0 21344 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607194113
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1607194113
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607194113
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607194113
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1493_
timestamp 1607194113
transform 1 0 2576 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1607194113
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__CLK
timestamp 1607194113
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__D
timestamp 1607194113
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1607194113
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1607194113
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_70
timestamp 1607194113
transform 1 0 7544 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1607194113
transform 1 0 6808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607194113
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1362_
timestamp 1607194113
transform 1 0 7820 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1607194113
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__CLK
timestamp 1607194113
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1607194113
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_106
timestamp 1607194113
transform 1 0 10856 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1607194113
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1607194113
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607194113
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1607194113
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__CLK
timestamp 1607194113
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1363_
timestamp 1607194113
transform 1 0 14720 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_21_167
timestamp 1607194113
transform 1 0 16468 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1607194113
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1607194113
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__B1
timestamp 1607194113
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607194113
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1292_
timestamp 1607194113
transform 1 0 18124 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_217
timestamp 1607194113
transform 1 0 21068 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_213
timestamp 1607194113
transform 1 0 20700 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1607194113
transform 1 0 19596 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__B1
timestamp 1607194113
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_236
timestamp 1607194113
transform 1 0 22816 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1285_
timestamp 1607194113
transform 1 0 21344 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607194113
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607194113
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607194113
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607194113
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607194113
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607194113
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607194113
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1607194113
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1607194113
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B1
timestamp 1607194113
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1297_
timestamp 1607194113
transform 1 0 6992 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_98
timestamp 1607194113
transform 1 0 10120 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1607194113
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1607194113
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607194113
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1295_
timestamp 1607194113
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_117
timestamp 1607194113
transform 1 0 11868 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_110
timestamp 1607194113
transform 1 0 11224 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1283_
timestamp 1607194113
transform 1 0 11500 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1607194113
transform 1 0 13064 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1607194113
transform 1 0 12604 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1289_
timestamp 1607194113
transform 1 0 12696 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1005_
timestamp 1607194113
transform 1 0 13800 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1607194113
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1607194113
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607194113
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1607194113
transform 1 0 15548 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_174
timestamp 1607194113
transform 1 0 17112 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_162
timestamp 1607194113
transform 1 0 16008 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A
timestamp 1607194113
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_198
timestamp 1607194113
transform 1 0 19320 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_186
timestamp 1607194113
transform 1 0 18216 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1607194113
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1607194113
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_202
timestamp 1607194113
transform 1 0 19688 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A
timestamp 1607194113
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A2
timestamp 1607194113
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607194113
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1607194113
transform 1 0 19780 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_235
timestamp 1607194113
transform 1 0 22724 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1607194113
transform 1 0 22540 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 21252 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_23_15
timestamp 1607194113
transform 1 0 2484 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607194113
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607194113
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1494_
timestamp 1607194113
transform 1 0 2576 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1607194113
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__CLK
timestamp 1607194113
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__D
timestamp 1607194113
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1607194113
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1607194113
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1607194113
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607194113
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1361_
timestamp 1607194113
transform 1 0 7544 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_91
timestamp 1607194113
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__CLK
timestamp 1607194113
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_115
timestamp 1607194113
transform 1 0 11684 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_103
timestamp 1607194113
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk_i
timestamp 1607194113
transform 1 0 11960 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_134
timestamp 1607194113
transform 1 0 13432 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1607194113
transform 1 0 12972 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_123
timestamp 1607194113
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1607194113
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607194113
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0958_
timestamp 1607194113
transform 1 0 13064 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_158
timestamp 1607194113
transform 1 0 15640 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__B1
timestamp 1607194113
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1294_
timestamp 1607194113
transform 1 0 14168 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_170
timestamp 1607194113
transform 1 0 16744 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_196
timestamp 1607194113
transform 1 0 19136 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1607194113
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1607194113
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__CLK
timestamp 1607194113
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607194113
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_218
timestamp 1607194113
transform 1 0 21160 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1364_
timestamp 1607194113
transform 1 0 19412 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_230
timestamp 1607194113
transform 1 0 22264 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_242
timestamp 1607194113
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607194113
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607194113
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607194113
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607194113
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607194113
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607194113
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1496_
timestamp 1607194113
transform 1 0 4048 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1607194113
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__CLK
timestamp 1607194113
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1607194113
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__D
timestamp 1607194113
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1011_
timestamp 1607194113
transform 1 0 6532 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_76
timestamp 1607194113
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_68
timestamp 1607194113
transform 1 0 7360 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 1607194113
transform 1 0 8372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1607194113
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_84
timestamp 1607194113
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A
timestamp 1607194113
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1607194113
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607194113
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1607194113
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1607194113
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_128
timestamp 1607194113
transform 1 0 12880 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1607194113
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1607194113
transform 1 0 12604 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1607194113
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A2
timestamp 1607194113
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607194113
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15456 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_24_175
timestamp 1607194113
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1607194113
transform 1 0 17020 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_187
timestamp 1607194113
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_218
timestamp 1607194113
transform 1 0 21160 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_215
timestamp 1607194113
transform 1 0 20884 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1607194113
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_199
timestamp 1607194113
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A2
timestamp 1607194113
transform 1 0 20976 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607194113
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A2
timestamp 1607194113
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _0967_
timestamp 1607194113
transform 1 0 21620 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_24_242
timestamp 1607194113
transform 1 0 23368 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1607194113
transform 1 0 23184 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1607194113
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607194113
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607194113
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1495_
timestamp 1607194113
transform 1 0 2576 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_25_37
timestamp 1607194113
transform 1 0 4508 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__CLK
timestamp 1607194113
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1607194113
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_47
timestamp 1607194113
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1607194113
transform 1 0 5060 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1607194113
transform 1 0 7452 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607194113
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1004_
timestamp 1607194113
transform 1 0 6808 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_25_85
timestamp 1607194113
transform 1 0 8924 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1607194113
transform 1 0 8556 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A1
timestamp 1607194113
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _1001_
timestamp 1607194113
transform 1 0 9200 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1607194113
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_107
timestamp 1607194113
transform 1 0 10948 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A2
timestamp 1607194113
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1607194113
transform 1 0 12972 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_123
timestamp 1607194113
transform 1 0 12420 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607194113
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1020_
timestamp 1607194113
transform 1 0 13064 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_25_144
timestamp 1607194113
transform 1 0 14352 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0957_
timestamp 1607194113
transform 1 0 15088 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1607194113
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1607194113
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1607194113
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1607194113
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607194113
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1607194113
transform 1 0 21068 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_208
timestamp 1607194113
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_i_A
timestamp 1607194113
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1
timestamp 1607194113
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk_i
timestamp 1607194113
transform 1 0 20792 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_4  _0974_
timestamp 1607194113
transform 1 0 21160 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_25_235
timestamp 1607194113
transform 1 0 22724 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1607194113
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607194113
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1607194113
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607194113
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1607194113
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607194113
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1607194113
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1607194113
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607194113
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607194113
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0680_
timestamp 1607194113
transform 1 0 2852 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_25
timestamp 1607194113
transform 1 0 3404 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_38
timestamp 1607194113
transform 1 0 4600 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1607194113
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1607194113
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607194113
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1003_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 4140 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0679_
timestamp 1607194113
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0667_
timestamp 1607194113
transform 1 0 3036 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_53
timestamp 1607194113
transform 1 0 5980 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_42
timestamp 1607194113
transform 1 0 4968 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_48
timestamp 1607194113
transform 1 0 5520 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1607194113
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0905_
timestamp 1607194113
transform 1 0 5152 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1607194113
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_74
timestamp 1607194113
transform 1 0 7912 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1607194113
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_72
timestamp 1607194113
transform 1 0 7728 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_60
timestamp 1607194113
transform 1 0 6624 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607194113
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_98
timestamp 1607194113
transform 1 0 10120 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1607194113
transform 1 0 8464 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_84
timestamp 1607194113
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1607194113
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607194113
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0995_
timestamp 1607194113
transform 1 0 9660 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__a32o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8556 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1607194113
transform 1 0 11500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_112
timestamp 1607194113
transform 1 0 11408 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A2
timestamp 1607194113
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0941_
timestamp 1607194113
transform 1 0 10856 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1607194113
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1607194113
transform 1 0 12512 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1607194113
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607194113
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1607194113
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_136
timestamp 1607194113
transform 1 0 13616 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_128
timestamp 1607194113
transform 1 0 12880 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1607194113
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B
timestamp 1607194113
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1007_
timestamp 1607194113
transform 1 0 13248 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1607194113
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_148
timestamp 1607194113
transform 1 0 14720 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_154
timestamp 1607194113
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1607194113
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_139
timestamp 1607194113
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1607194113
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607194113
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1017_
timestamp 1607194113
transform 1 0 14076 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1607194113
transform 1 0 15456 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_177
timestamp 1607194113
transform 1 0 17388 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1607194113
transform 1 0 16468 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1607194113
transform 1 0 15732 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1607194113
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B1
timestamp 1607194113
transform 1 0 17388 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1000_
timestamp 1607194113
transform 1 0 15824 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_4  _0984_
timestamp 1607194113
transform 1 0 16560 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1607194113
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1607194113
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_191
timestamp 1607194113
transform 1 0 18676 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_179
timestamp 1607194113
transform 1 0 17572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607194113
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_216
timestamp 1607194113
transform 1 0 20976 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_204
timestamp 1607194113
transform 1 0 19872 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_206
timestamp 1607194113
transform 1 0 20056 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1607194113
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A2
timestamp 1607194113
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607194113
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0981_
timestamp 1607194113
transform 1 0 20884 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_4  _0977_
timestamp 1607194113
transform 1 0 20148 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1607194113
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1607194113
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_234
timestamp 1607194113
transform 1 0 22632 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A1
timestamp 1607194113
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1607194113
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0962_
timestamp 1607194113
transform 1 0 21528 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_27_241
timestamp 1607194113
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_243
timestamp 1607194113
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607194113
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1607194113
transform 1 0 23184 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_15
timestamp 1607194113
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607194113
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1607194113
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607194113
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_23
timestamp 1607194113
transform 1 0 3220 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B
timestamp 1607194113
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607194113
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0669_
timestamp 1607194113
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1607194113
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1607194113
transform 1 0 4876 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _0907_
timestamp 1607194113
transform 1 0 5980 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_78
timestamp 1607194113
transform 1 0 8280 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1607194113
transform 1 0 7912 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1607194113
transform 1 0 6808 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1607194113
transform 1 0 8372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_93
timestamp 1607194113
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1607194113
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_83
timestamp 1607194113
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607194113
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_110
timestamp 1607194113
transform 1 0 11224 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1607194113
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1282_
timestamp 1607194113
transform 1 0 11776 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_137
timestamp 1607194113
transform 1 0 13708 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_125
timestamp 1607194113
transform 1 0 12604 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_154
timestamp 1607194113
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1607194113
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607194113
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0994_
timestamp 1607194113
transform 1 0 16008 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_28_191
timestamp 1607194113
transform 1 0 18676 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_179
timestamp 1607194113
transform 1 0 17572 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1607194113
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607194113
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1607194113
transform 1 0 19780 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0946_
timestamp 1607194113
transform 1 0 20884 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_28_224
timestamp 1607194113
transform 1 0 21712 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1607194113
transform 1 0 21528 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1607194113
transform 1 0 22908 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0970_
timestamp 1607194113
transform 1 0 22264 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_28_239
timestamp 1607194113
transform 1 0 23092 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1607194113
transform 1 0 2852 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_11
timestamp 1607194113
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1607194113
transform 1 0 1380 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1607194113
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607194113
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1607194113
transform 1 0 2576 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_36
timestamp 1607194113
transform 1 0 4416 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__C
timestamp 1607194113
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1607194113
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0866_
timestamp 1607194113
transform 1 0 3588 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1607194113
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0948_
timestamp 1607194113
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_78
timestamp 1607194113
transform 1 0 8280 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_66
timestamp 1607194113
transform 1 0 7176 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607194113
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0908_
timestamp 1607194113
transform 1 0 7912 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1607194113
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_90
timestamp 1607194113
transform 1 0 9384 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0993_
timestamp 1607194113
transform 1 0 9476 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_112
timestamp 1607194113
transform 1 0 11408 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_100
timestamp 1607194113
transform 1 0 10304 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp 1607194113
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1607194113
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1607194113
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607194113
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 12880 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1607194113
transform 1 0 15640 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_141
timestamp 1607194113
transform 1 0 14076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1021_
timestamp 1607194113
transform 1 0 14812 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_170
timestamp 1607194113
transform 1 0 16744 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0961_
timestamp 1607194113
transform 1 0 16376 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1607194113
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1607194113
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1607194113
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607194113
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_200
timestamp 1607194113
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__CLK
timestamp 1607194113
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1375_
timestamp 1607194113
transform 1 0 19780 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_234
timestamp 1607194113
transform 1 0 22632 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_222
timestamp 1607194113
transform 1 0 21528 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_242
timestamp 1607194113
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607194113
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1607194113
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607194113
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607194113
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_32
timestamp 1607194113
transform 1 0 4048 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1607194113
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1607194113
transform 1 0 4140 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607194113
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1022_
timestamp 1607194113
transform 1 0 4324 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1607194113
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1607194113
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1607194113
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1607194113
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607194113
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0999_
timestamp 1607194113
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_119
timestamp 1607194113
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_104
timestamp 1607194113
transform 1 0 10672 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__D
timestamp 1607194113
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1158_
timestamp 1607194113
transform 1 0 11224 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_131
timestamp 1607194113
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1607194113
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1607194113
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_143
timestamp 1607194113
transform 1 0 14260 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607194113
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1013_
timestamp 1607194113
transform 1 0 15456 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_30_175
timestamp 1607194113
transform 1 0 17204 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_165
timestamp 1607194113
transform 1 0 16284 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1607194113
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1607194113
transform 1 0 16836 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1607194113
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A2
timestamp 1607194113
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A3
timestamp 1607194113
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1272_
timestamp 1607194113
transform 1 0 18492 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1607194113
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1607194113
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__B1
timestamp 1607194113
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607194113
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1607194113
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_239
timestamp 1607194113
transform 1 0 23092 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 1607194113
transform 1 0 2484 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607194113
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607194113
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1498_
timestamp 1607194113
transform 1 0 2576 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_31_37
timestamp 1607194113
transform 1 0 4508 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__CLK
timestamp 1607194113
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_52
timestamp 1607194113
transform 1 0 5888 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1607194113
transform 1 0 5704 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1012_
timestamp 1607194113
transform 1 0 5060 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_31_75
timestamp 1607194113
transform 1 0 8004 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1607194113
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1607194113
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__D
timestamp 1607194113
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607194113
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0682_
timestamp 1607194113
transform 1 0 7176 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_83
timestamp 1607194113
transform 1 0 8740 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A2
timestamp 1607194113
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B1
timestamp 1607194113
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0992_
timestamp 1607194113
transform 1 0 9016 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1607194113
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_111
timestamp 1607194113
transform 1 0 11316 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_101
timestamp 1607194113
transform 1 0 10396 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1025_
timestamp 1607194113
transform 1 0 10948 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1607194113
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1607194113
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607194113
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1607194113
transform 1 0 14628 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__CLK
timestamp 1607194113
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1372_
timestamp 1607194113
transform 1 0 15180 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1607194113
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1607194113
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1607194113
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__CLK
timestamp 1607194113
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607194113
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1376_
timestamp 1607194113
transform 1 0 19320 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_31_217
timestamp 1607194113
transform 1 0 21068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1607194113
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1607194113
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607194113
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_15
timestamp 1607194113
transform 1 0 2484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1607194113
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1607194113
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607194113
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0939_
timestamp 1607194113
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp 1607194113
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1607194113
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607194113
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0670_
timestamp 1607194113
transform 1 0 4600 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_55
timestamp 1607194113
transform 1 0 6164 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_50
timestamp 1607194113
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_42
timestamp 1607194113
transform 1 0 4968 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0949_
timestamp 1607194113
transform 1 0 5796 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_79
timestamp 1607194113
transform 1 0 8372 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_67
timestamp 1607194113
transform 1 0 7268 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_87
timestamp 1607194113
transform 1 0 9108 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B1
timestamp 1607194113
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607194113
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0998_
timestamp 1607194113
transform 1 0 9660 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_32_118
timestamp 1607194113
transform 1 0 11960 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_108
timestamp 1607194113
transform 1 0 11040 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A2
timestamp 1607194113
transform 1 0 10856 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1607194113
transform 1 0 11408 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0950_
timestamp 1607194113
transform 1 0 11592 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_130
timestamp 1607194113
transform 1 0 13064 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1224_
timestamp 1607194113
transform 1 0 12696 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1607194113
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_150
timestamp 1607194113
transform 1 0 14904 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_142
timestamp 1607194113
transform 1 0 14168 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A2
timestamp 1607194113
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A3
timestamp 1607194113
transform 1 0 15364 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607194113
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1275_
timestamp 1607194113
transform 1 0 15548 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_32_176
timestamp 1607194113
transform 1 0 17296 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B1
timestamp 1607194113
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_188
timestamp 1607194113
transform 1 0 18400 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1607194113
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1607194113
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_200
timestamp 1607194113
transform 1 0 19504 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607194113
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1607194113
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_239
timestamp 1607194113
transform 1 0 23092 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607194113
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607194113
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_15
timestamp 1607194113
transform 1 0 2484 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607194113
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607194113
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607194113
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1497_
timestamp 1607194113
transform 1 0 2576 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1607194113
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1607194113
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_37
timestamp 1607194113
transform 1 0 4508 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__CLK
timestamp 1607194113
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607194113
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1607194113
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1607194113
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_49
timestamp 1607194113
transform 1 0 5612 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1607194113
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1607194113
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1607194113
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607194113
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_98
timestamp 1607194113
transform 1 0 10120 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1607194113
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_98
timestamp 1607194113
transform 1 0 10120 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1607194113
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1607194113
transform 1 0 9936 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607194113
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1607194113
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_107
timestamp 1607194113
transform 1 0 10948 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1607194113
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_111
timestamp 1607194113
transform 1 0 11316 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__B1
timestamp 1607194113
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1233_
timestamp 1607194113
transform 1 0 10672 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1231_
timestamp 1607194113
transform 1 0 11684 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1607194113
transform 1 0 10672 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1607194113
transform 1 0 13156 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1607194113
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607194113
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1220_
timestamp 1607194113
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_148
timestamp 1607194113
transform 1 0 14720 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1607194113
transform 1 0 14352 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_147
timestamp 1607194113
transform 1 0 14628 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_139
timestamp 1607194113
transform 1 0 13892 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1607194113
transform 1 0 14168 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1607194113
transform 1 0 14720 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1607194113
transform 1 0 13892 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A2
timestamp 1607194113
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B2
timestamp 1607194113
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607194113
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1607194113
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1015_
timestamp 1607194113
transform 1 0 15272 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1607194113
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_175
timestamp 1607194113
transform 1 0 17204 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_163
timestamp 1607194113
transform 1 0 16100 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_184
timestamp 1607194113
transform 1 0 18032 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607194113
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_196
timestamp 1607194113
transform 1 0 19136 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1607194113
transform 1 0 18768 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_192
timestamp 1607194113
transform 1 0 18768 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A2
timestamp 1607194113
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A3
timestamp 1607194113
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1221_
timestamp 1607194113
transform 1 0 19228 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1607194113
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _1271_
timestamp 1607194113
transform 1 0 19228 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1607194113
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1607194113
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1607194113
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_216
timestamp 1607194113
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__B1
timestamp 1607194113
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A2
timestamp 1607194113
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607194113
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_227
timestamp 1607194113
transform 1 0 21988 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1607194113
transform 1 0 23000 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B2
timestamp 1607194113
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1607194113
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1406_
timestamp 1607194113
transform 1 0 22356 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _0972_
timestamp 1607194113
transform 1 0 21528 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607194113
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_15
timestamp 1607194113
transform 1 0 2484 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1607194113
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607194113
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1482_
timestamp 1607194113
transform 1 0 2576 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1607194113
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__CLK
timestamp 1607194113
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__D
timestamp 1607194113
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1607194113
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1607194113
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_70
timestamp 1607194113
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_62
timestamp 1607194113
transform 1 0 6808 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__B1
timestamp 1607194113
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607194113
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1229_
timestamp 1607194113
transform 1 0 7912 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_35_90
timestamp 1607194113
transform 1 0 9384 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0867_
timestamp 1607194113
transform 1 0 10120 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_114
timestamp 1607194113
transform 1 0 11592 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1607194113
transform 1 0 10488 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1228_
timestamp 1607194113
transform 1 0 11224 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1607194113
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__CLK
timestamp 1607194113
transform 1 0 12604 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607194113
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1401_
timestamp 1607194113
transform 1 0 12788 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_35_154
timestamp 1607194113
transform 1 0 15272 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_146
timestamp 1607194113
transform 1 0 14536 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B1
timestamp 1607194113
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_175
timestamp 1607194113
transform 1 0 17204 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1232_
timestamp 1607194113
transform 1 0 15732 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_196
timestamp 1607194113
transform 1 0 19136 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1607194113
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607194113
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1234_
timestamp 1607194113
transform 1 0 19228 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_216
timestamp 1607194113
transform 1 0 20976 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_212
timestamp 1607194113
transform 1 0 20608 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_200
timestamp 1607194113
transform 1 0 19504 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B1
timestamp 1607194113
transform 1 0 21068 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_235
timestamp 1607194113
transform 1 0 22724 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1225_
timestamp 1607194113
transform 1 0 21252 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_243
timestamp 1607194113
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607194113
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1607194113
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1607194113
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607194113
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1607194113
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1607194113
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607194113
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_56
timestamp 1607194113
transform 1 0 6256 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1607194113
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_64
timestamp 1607194113
transform 1 0 6992 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B1
timestamp 1607194113
transform 1 0 7176 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1230_
timestamp 1607194113
transform 1 0 7360 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_36_98
timestamp 1607194113
transform 1 0 10120 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_84
timestamp 1607194113
transform 1 0 8832 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1607194113
transform 1 0 9936 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607194113
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1607194113
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_110
timestamp 1607194113
transform 1 0 11224 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1607194113
transform 1 0 11960 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_136
timestamp 1607194113
transform 1 0 13616 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_124
timestamp 1607194113
transform 1 0 12512 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1607194113
transform 1 0 12144 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1607194113
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1607194113
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_148
timestamp 1607194113
transform 1 0 14720 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607194113
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_166
timestamp 1607194113
transform 1 0 16376 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__CLK
timestamp 1607194113
transform 1 0 16744 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1400_
timestamp 1607194113
transform 1 0 16928 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_36_191
timestamp 1607194113
transform 1 0 18676 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_209
timestamp 1607194113
transform 1 0 20332 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_203
timestamp 1607194113
transform 1 0 19780 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A2
timestamp 1607194113
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B2
timestamp 1607194113
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607194113
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0979_
timestamp 1607194113
transform 1 0 20884 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_36_231
timestamp 1607194113
transform 1 0 22356 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A1
timestamp 1607194113
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_243
timestamp 1607194113
transform 1 0 23460 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_15
timestamp 1607194113
transform 1 0 2484 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1607194113
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607194113
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1499_
timestamp 1607194113
transform 1 0 2576 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1607194113
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__CLK
timestamp 1607194113
transform 1 0 4508 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__D
timestamp 1607194113
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1607194113
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1607194113
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_74
timestamp 1607194113
transform 1 0 7912 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1607194113
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607194113
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1402_
timestamp 1607194113
transform 1 0 8280 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_37_99
timestamp 1607194113
transform 1 0 10212 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__CLK
timestamp 1607194113
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_119
timestamp 1607194113
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_111
timestamp 1607194113
transform 1 0 11316 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1607194113
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B1
timestamp 1607194113
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607194113
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1227_
timestamp 1607194113
transform 1 0 13708 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_37_153
timestamp 1607194113
transform 1 0 15180 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_177
timestamp 1607194113
transform 1 0 17388 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_165
timestamp 1607194113
transform 1 0 16284 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_189
timestamp 1607194113
transform 1 0 18492 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1607194113
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607194113
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1607194113
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_201
timestamp 1607194113
transform 1 0 19596 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B1
timestamp 1607194113
transform 1 0 19872 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1226_
timestamp 1607194113
transform 1 0 20056 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_37_234
timestamp 1607194113
transform 1 0 22632 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_222
timestamp 1607194113
transform 1 0 21528 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_242
timestamp 1607194113
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607194113
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1607194113
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1607194113
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607194113
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1607194113
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1607194113
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607194113
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1607194113
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1607194113
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1607194113
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1607194113
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1607194113
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607194113
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_109
timestamp 1607194113
transform 1 0 11132 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_105
timestamp 1607194113
transform 1 0 10764 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1607194113
transform 1 0 12052 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 11224 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1607194113
transform 1 0 13340 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1607194113
transform 1 0 12236 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_145
timestamp 1607194113
transform 1 0 14444 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1607194113
transform 1 0 13892 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B2
timestamp 1607194113
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1607194113
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A2
timestamp 1607194113
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607194113
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0987_
timestamp 1607194113
transform 1 0 15272 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1607194113
transform 1 0 14168 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1607194113
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_192
timestamp 1607194113
transform 1 0 18768 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1607194113
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_204
timestamp 1607194113
transform 1 0 19872 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607194113
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1405_
timestamp 1607194113
transform 1 0 20884 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_38_234
timestamp 1607194113
transform 1 0 22632 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1607194113
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1607194113
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_15
timestamp 1607194113
transform 1 0 2484 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1607194113
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607194113
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607194113
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1500_
timestamp 1607194113
transform 1 0 2576 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1607194113
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1607194113
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_37
timestamp 1607194113
transform 1 0 4508 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__CLK
timestamp 1607194113
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607194113
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_44
timestamp 1607194113
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_53
timestamp 1607194113
transform 1 0 5980 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_49
timestamp 1607194113
transform 1 0 5612 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1517_
timestamp 1607194113
transform 1 0 5336 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1607194113
transform 1 0 5704 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_79
timestamp 1607194113
transform 1 0 8372 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_67
timestamp 1607194113
transform 1 0 7268 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_73
timestamp 1607194113
transform 1 0 7820 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__CLK
timestamp 1607194113
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1607194113
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607194113
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0683_
timestamp 1607194113
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_87
timestamp 1607194113
transform 1 0 9108 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__CLK
timestamp 1607194113
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607194113
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1412_
timestamp 1607194113
transform 1 0 9660 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1403_
timestamp 1607194113
transform 1 0 8556 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_40_112
timestamp 1607194113
transform 1 0 11408 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_112
timestamp 1607194113
transform 1 0 11408 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_102
timestamp 1607194113
transform 1 0 10488 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__CLK
timestamp 1607194113
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1607194113
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1607194113
transform 1 0 11040 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_136
timestamp 1607194113
transform 1 0 13616 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_124
timestamp 1607194113
transform 1 0 12512 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1607194113
transform 1 0 13524 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1607194113
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_120
timestamp 1607194113
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607194113
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1607194113
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1607194113
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_148
timestamp 1607194113
transform 1 0 14720 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_139
timestamp 1607194113
transform 1 0 13892 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__CLK
timestamp 1607194113
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607194113
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1404_
timestamp 1607194113
transform 1 0 14168 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1607194113
transform 1 0 15456 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_167
timestamp 1607194113
transform 1 0 16468 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_161
timestamp 1607194113
transform 1 0 15916 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_173
timestamp 1607194113
transform 1 0 17020 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_161
timestamp 1607194113
transform 1 0 15916 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1607194113
transform 1 0 15732 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1371_
timestamp 1607194113
transform 1 0 16560 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1607194113
transform 1 0 19228 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_189
timestamp 1607194113
transform 1 0 18492 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_189
timestamp 1607194113
transform 1 0 18492 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_181
timestamp 1607194113
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__CLK
timestamp 1607194113
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1607194113
transform 1 0 18308 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607194113
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1607194113
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1607194113
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1607194113
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_205
timestamp 1607194113
transform 1 0 19964 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_213
timestamp 1607194113
transform 1 0 20700 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_201
timestamp 1607194113
transform 1 0 19596 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_i_A
timestamp 1607194113
transform 1 0 19780 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk_i
timestamp 1607194113
transform 1 0 19504 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607194113
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_233
timestamp 1607194113
transform 1 0 22540 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_230
timestamp 1607194113
transform 1 0 22264 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1607194113
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1607194113
transform 1 0 21988 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1315_
timestamp 1607194113
transform 1 0 22172 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1607194113
transform 1 0 21804 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_242
timestamp 1607194113
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__B1
timestamp 1607194113
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607194113
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1316_
timestamp 1607194113
transform 1 0 23276 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_41_15
timestamp 1607194113
transform 1 0 2484 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1607194113
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607194113
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1501_
timestamp 1607194113
transform 1 0 2576 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_41_37
timestamp 1607194113
transform 1 0 4508 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__CLK
timestamp 1607194113
transform 1 0 4324 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_49
timestamp 1607194113
transform 1 0 5612 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A1
timestamp 1607194113
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B1
timestamp 1607194113
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607194113
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0684_
timestamp 1607194113
transform 1 0 6808 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_41_91
timestamp 1607194113
transform 1 0 9476 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_80
timestamp 1607194113
transform 1 0 8464 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B1
timestamp 1607194113
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk_i
timestamp 1607194113
transform 1 0 9200 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1215_
timestamp 1607194113
transform 1 0 10028 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_41_115
timestamp 1607194113
transform 1 0 11684 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1_N
timestamp 1607194113
transform 1 0 11500 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_130
timestamp 1607194113
transform 1 0 13064 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1607194113
transform 1 0 12696 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1607194113
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A1_N
timestamp 1607194113
transform 1 0 13156 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A2_N
timestamp 1607194113
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607194113
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1006_
timestamp 1607194113
transform 1 0 13524 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1607194113
transform 1 0 12420 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_151
timestamp 1607194113
transform 1 0 14996 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__B1
timestamp 1607194113
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1607194113
transform 1 0 17388 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A1_N
timestamp 1607194113
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1277_
timestamp 1607194113
transform 1 0 15732 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__CLK
timestamp 1607194113
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607194113
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1413_
timestamp 1607194113
transform 1 0 18032 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_41_215
timestamp 1607194113
transform 1 0 20884 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_203
timestamp 1607194113
transform 1 0 19780 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_227
timestamp 1607194113
transform 1 0 21988 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1607194113
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1607194113
transform 1 0 23092 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607194113
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1607194113
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1607194113
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607194113
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1607194113
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1607194113
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607194113
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_44
timestamp 1607194113
transform 1 0 5152 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1518_
timestamp 1607194113
transform 1 0 5244 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1607194113
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_66
timestamp 1607194113
transform 1 0 7176 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__CLK
timestamp 1607194113
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1607194113
transform 1 0 7728 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1607194113
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1607194113
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_87
timestamp 1607194113
transform 1 0 9108 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607194113
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_113
timestamp 1607194113
transform 1 0 11500 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_105
timestamp 1607194113
transform 1 0 10764 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1213_
timestamp 1607194113
transform 1 0 11776 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_132
timestamp 1607194113
transform 1 0 13248 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_120
timestamp 1607194113
transform 1 0 12144 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_154
timestamp 1607194113
transform 1 0 15272 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_152
timestamp 1607194113
transform 1 0 15088 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_144
timestamp 1607194113
transform 1 0 14352 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607194113
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B1
timestamp 1607194113
transform 1 0 16376 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1214_
timestamp 1607194113
transform 1 0 16560 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_196
timestamp 1607194113
transform 1 0 19136 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_184
timestamp 1607194113
transform 1 0 18032 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1607194113
transform 1 0 20884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_208
timestamp 1607194113
transform 1 0 20240 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607194113
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1607194113
transform 1 0 21988 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_239
timestamp 1607194113
transform 1 0 23092 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1607194113
transform 1 0 2484 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1607194113
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607194113
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1502_
timestamp 1607194113
transform 1 0 2576 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_43_37
timestamp 1607194113
transform 1 0 4508 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__CLK
timestamp 1607194113
transform 1 0 4324 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_49
timestamp 1607194113
transform 1 0 5612 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_71
timestamp 1607194113
transform 1 0 7636 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_62
timestamp 1607194113
transform 1 0 6808 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607194113
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0674_
timestamp 1607194113
transform 1 0 8372 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1607194113
transform 1 0 7360 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_92
timestamp 1607194113
transform 1 0 9568 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B
timestamp 1607194113
transform 1 0 9384 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1607194113
transform 1 0 9200 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_110
timestamp 1607194113
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_104
timestamp 1607194113
transform 1 0 10672 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_i_A
timestamp 1607194113
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk_i
timestamp 1607194113
transform 1 0 10764 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_135
timestamp 1607194113
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1607194113
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607194113
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_147
timestamp 1607194113
transform 1 0 14628 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B1
timestamp 1607194113
transform 1 0 15364 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1216_
timestamp 1607194113
transform 1 0 15548 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_43_175
timestamp 1607194113
transform 1 0 17204 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1_N
timestamp 1607194113
transform 1 0 17020 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_187
timestamp 1607194113
transform 1 0 18308 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607194113
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1607194113
transform 1 0 18032 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_211
timestamp 1607194113
transform 1 0 20516 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_199
timestamp 1607194113
transform 1 0 19412 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_235
timestamp 1607194113
transform 1 0 22724 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_223
timestamp 1607194113
transform 1 0 21620 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_243
timestamp 1607194113
transform 1 0 23460 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607194113
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1607194113
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1607194113
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1607194113
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1607194113
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607194113
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1504_
timestamp 1607194113
transform 1 0 4048 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_44_53
timestamp 1607194113
transform 1 0 5980 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1519_
timestamp 1607194113
transform 1 0 6532 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__CLK
timestamp 1607194113
transform 1 0 8280 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1607194113
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_80
timestamp 1607194113
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607194113
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1607194113
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1607194113
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1607194113
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_154
timestamp 1607194113
transform 1 0 15272 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1607194113
transform 1 0 14076 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607194113
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_162
timestamp 1607194113
transform 1 0 16008 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1411_
timestamp 1607194113
transform 1 0 16192 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1607194113
transform 1 0 19228 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_185
timestamp 1607194113
transform 1 0 18124 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__CLK
timestamp 1607194113
transform 1 0 17940 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_215
timestamp 1607194113
transform 1 0 20884 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1607194113
transform 1 0 20700 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1607194113
transform 1 0 20332 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__CLK
timestamp 1607194113
transform 1 0 21068 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607194113
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_238
timestamp 1607194113
transform 1 0 23000 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1414_
timestamp 1607194113
transform 1 0 21252 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp 1607194113
transform 1 0 2484 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1607194113
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1607194113
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1503_
timestamp 1607194113
transform 1 0 2576 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_45_37
timestamp 1607194113
transform 1 0 4508 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__CLK
timestamp 1607194113
transform 1 0 4324 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_49
timestamp 1607194113
transform 1 0 5612 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_74
timestamp 1607194113
transform 1 0 7912 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_68
timestamp 1607194113
transform 1 0 7360 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_62
timestamp 1607194113
transform 1 0 6808 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1607194113
transform 1 0 7452 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607194113
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1607194113
transform 1 0 7636 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_96
timestamp 1607194113
transform 1 0 9936 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B1
timestamp 1607194113
transform 1 0 8464 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A2
timestamp 1607194113
transform 1 0 9752 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_119
timestamp 1607194113
transform 1 0 12052 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_111
timestamp 1607194113
transform 1 0 11316 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1607194113
transform 1 0 11132 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1023_
timestamp 1607194113
transform 1 0 10488 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_45_133
timestamp 1607194113
transform 1 0 13340 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_129
timestamp 1607194113
transform 1 0 12972 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_123
timestamp 1607194113
transform 1 0 12420 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607194113
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1607194113
transform 1 0 13064 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__CLK
timestamp 1607194113
transform 1 0 14076 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1369_
timestamp 1607194113
transform 1 0 14260 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_45_173
timestamp 1607194113
transform 1 0 17020 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_162
timestamp 1607194113
transform 1 0 16008 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1607194113
transform 1 0 16744 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1607194113
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1607194113
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1607194113
transform 1 0 17756 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607194113
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_208
timestamp 1607194113
transform 1 0 20240 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B1
timestamp 1607194113
transform 1 0 20516 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1212_
timestamp 1607194113
transform 1 0 20700 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_231
timestamp 1607194113
transform 1 0 22356 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A1_N
timestamp 1607194113
transform 1 0 22172 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1607194113
transform 1 0 23460 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607194113
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_15
timestamp 1607194113
transform 1 0 2484 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1607194113
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1607194113
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1607194113
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1607194113
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1607194113
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1505_
timestamp 1607194113
transform 1 0 2576 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_47_37
timestamp 1607194113
transform 1 0 4508 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1607194113
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__CLK
timestamp 1607194113
transform 1 0 4324 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607194113
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0901_
timestamp 1607194113
transform 1 0 4048 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_47_52
timestamp 1607194113
transform 1 0 5888 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_55
timestamp 1607194113
transform 1 0 6164 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_43
timestamp 1607194113
transform 1 0 5060 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1607194113
transform 1 0 4876 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0912_
timestamp 1607194113
transform 1 0 5060 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_47_73
timestamp 1607194113
transform 1 0 7820 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_62
timestamp 1607194113
transform 1 0 6808 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_60
timestamp 1607194113
transform 1 0 6624 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_67
timestamp 1607194113
transform 1 0 7268 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607194113
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1607194113
transform 1 0 7544 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1326_
timestamp 1607194113
transform 1 0 8004 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_47_97
timestamp 1607194113
transform 1 0 10028 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_81
timestamp 1607194113
transform 1 0 8556 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_93
timestamp 1607194113
transform 1 0 9660 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1607194113
transform 1 0 9200 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__B
timestamp 1607194113
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A2
timestamp 1607194113
transform 1 0 9844 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A
timestamp 1607194113
transform 1 0 8832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607194113
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1325_
timestamp 1607194113
transform 1 0 8740 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_105
timestamp 1607194113
transform 1 0 10764 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_104
timestamp 1607194113
transform 1 0 10672 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk_i
timestamp 1607194113
transform 1 0 10396 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0665_
timestamp 1607194113
transform 1 0 10948 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_119
timestamp 1607194113
transform 1 0 12052 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1607194113
transform 1 0 11500 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_110
timestamp 1607194113
transform 1 0 11224 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__CLK
timestamp 1607194113
transform 1 0 11316 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A
timestamp 1607194113
transform 1 0 11316 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1410_
timestamp 1607194113
transform 1 0 11500 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_46_132
timestamp 1607194113
transform 1 0 13248 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B1
timestamp 1607194113
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607194113
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1218_
timestamp 1607194113
transform 1 0 12420 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_151
timestamp 1607194113
transform 1 0 14996 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_139
timestamp 1607194113
transform 1 0 13892 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_154
timestamp 1607194113
transform 1 0 15272 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_152
timestamp 1607194113
transform 1 0 15088 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_144
timestamp 1607194113
transform 1 0 14352 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B1
timestamp 1607194113
transform 1 0 15456 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607194113
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1279_
timestamp 1607194113
transform 1 0 15640 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_47_175
timestamp 1607194113
transform 1 0 17204 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_163
timestamp 1607194113
transform 1 0 16100 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_178
timestamp 1607194113
transform 1 0 17480 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B2
timestamp 1607194113
transform 1 0 17296 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1_N
timestamp 1607194113
transform 1 0 17112 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_196
timestamp 1607194113
transform 1 0 19136 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1607194113
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_190
timestamp 1607194113
transform 1 0 18584 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607194113
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_218
timestamp 1607194113
transform 1 0 21160 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_210
timestamp 1607194113
transform 1 0 20424 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_202
timestamp 1607194113
transform 1 0 19688 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__B1
timestamp 1607194113
transform 1 0 19504 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607194113
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1370_
timestamp 1607194113
transform 1 0 20884 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1278_
timestamp 1607194113
transform 1 0 19688 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_230
timestamp 1607194113
transform 1 0 22264 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_234
timestamp 1607194113
transform 1 0 22632 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_242
timestamp 1607194113
transform 1 0 23368 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_240
timestamp 1607194113
transform 1 0 23184 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1607194113
transform 1 0 23276 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607194113
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1607194113
transform 1 0 23460 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1607194113
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1607194113
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1607194113
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1607194113
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607194113
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0899_
timestamp 1607194113
transform 1 0 4048 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_48_55
timestamp 1607194113
transform 1 0 6164 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_43
timestamp 1607194113
transform 1 0 5060 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1607194113
transform 1 0 4876 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_75
timestamp 1607194113
transform 1 0 8004 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_67
timestamp 1607194113
transform 1 0 7268 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A
timestamp 1607194113
transform 1 0 8188 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1607194113
transform 1 0 8372 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1607194113
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_90
timestamp 1607194113
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_82
timestamp 1607194113
transform 1 0 8648 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607194113
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_105
timestamp 1607194113
transform 1 0 10764 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B1
timestamp 1607194113
transform 1 0 11316 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1217_
timestamp 1607194113
transform 1 0 11500 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_48_131
timestamp 1607194113
transform 1 0 13156 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1_N
timestamp 1607194113
transform 1 0 12972 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1172_
timestamp 1607194113
transform 1 0 13708 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_154
timestamp 1607194113
transform 1 0 15272 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1607194113
transform 1 0 14076 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607194113
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_172
timestamp 1607194113
transform 1 0 16928 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_166
timestamp 1607194113
transform 1 0 16376 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__CLK
timestamp 1607194113
transform 1 0 17020 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1368_
timestamp 1607194113
transform 1 0 17204 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_48_194
timestamp 1607194113
transform 1 0 18952 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1607194113
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_206
timestamp 1607194113
transform 1 0 20056 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A
timestamp 1607194113
transform 1 0 19504 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607194113
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1276_
timestamp 1607194113
transform 1 0 19688 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1607194113
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1607194113
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1607194113
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1607194113
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1607194113
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_38
timestamp 1607194113
transform 1 0 4600 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_27
timestamp 1607194113
transform 1 0 3588 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0914_
timestamp 1607194113
transform 1 0 3772 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_49_58
timestamp 1607194113
transform 1 0 6440 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_50
timestamp 1607194113
transform 1 0 5704 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0895_
timestamp 1607194113
transform 1 0 5336 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_74
timestamp 1607194113
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1607194113
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607194113
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_98
timestamp 1607194113
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_86
timestamp 1607194113
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_110
timestamp 1607194113
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607194113
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1409_
timestamp 1607194113
transform 1 0 12420 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_49_153
timestamp 1607194113
transform 1 0 15180 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_144
timestamp 1607194113
transform 1 0 14352 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__CLK
timestamp 1607194113
transform 1 0 14168 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1607194113
transform 1 0 14904 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_172
timestamp 1607194113
transform 1 0 16928 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_165
timestamp 1607194113
transform 1 0 16284 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk_i
timestamp 1607194113
transform 1 0 16652 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_197
timestamp 1607194113
transform 1 0 19228 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_189
timestamp 1607194113
transform 1 0 18492 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_180
timestamp 1607194113
transform 1 0 17664 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A
timestamp 1607194113
transform 1 0 18308 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607194113
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1607194113
transform 1 0 18032 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_215
timestamp 1607194113
transform 1 0 20884 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_203
timestamp 1607194113
transform 1 0 19780 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1240_
timestamp 1607194113
transform 1 0 19412 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_227
timestamp 1607194113
transform 1 0 21988 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_243
timestamp 1607194113
transform 1 0 23460 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_239
timestamp 1607194113
transform 1 0 23092 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607194113
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_11
timestamp 1607194113
transform 1 0 2116 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1607194113
transform 1 0 1380 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1607194113
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0932_
timestamp 1607194113
transform 1 0 2392 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_50_25
timestamp 1607194113
transform 1 0 3404 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__B
timestamp 1607194113
transform 1 0 3220 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607194113
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0921_
timestamp 1607194113
transform 1 0 4048 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_50_43
timestamp 1607194113
transform 1 0 5060 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1607194113
transform 1 0 4876 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1506_
timestamp 1607194113
transform 1 0 5796 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_72
timestamp 1607194113
transform 1 0 7728 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__CLK
timestamp 1607194113
transform 1 0 7544 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_99
timestamp 1607194113
transform 1 0 10212 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_93
timestamp 1607194113
transform 1 0 9660 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_84
timestamp 1607194113
transform 1 0 8832 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607194113
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__CLK
timestamp 1607194113
transform 1 0 10304 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1426_
timestamp 1607194113
transform 1 0 10488 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1607194113
transform 1 0 13340 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1607194113
transform 1 0 12236 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_154
timestamp 1607194113
transform 1 0 15272 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_151
timestamp 1607194113
transform 1 0 14996 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_143
timestamp 1607194113
transform 1 0 14260 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607194113
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1173_
timestamp 1607194113
transform 1 0 13892 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B1
timestamp 1607194113
transform 1 0 16376 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1280_
timestamp 1607194113
transform 1 0 16560 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_50_188
timestamp 1607194113
transform 1 0 18400 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1607194113
transform 1 0 18584 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A2_N
timestamp 1607194113
transform 1 0 18216 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B2
timestamp 1607194113
transform 1 0 18032 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0804_
timestamp 1607194113
transform 1 0 18768 0 -1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_50_215
timestamp 1607194113
transform 1 0 20884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1607194113
transform 1 0 20424 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1607194113
transform 1 0 20240 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B2
timestamp 1607194113
transform 1 0 20056 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607194113
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1607194113
transform 1 0 21988 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__CLK
timestamp 1607194113
transform 1 0 23092 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1373_
timestamp 1607194113
transform 1 0 23276 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_51_11
timestamp 1607194113
transform 1 0 2116 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1607194113
transform 1 0 1380 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1607194113
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0934_
timestamp 1607194113
transform 1 0 2392 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_51_25
timestamp 1607194113
transform 1 0 3404 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B
timestamp 1607194113
transform 1 0 3220 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0926_
timestamp 1607194113
transform 1 0 3956 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_51_52
timestamp 1607194113
transform 1 0 5888 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_42
timestamp 1607194113
transform 1 0 4968 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B
timestamp 1607194113
transform 1 0 4784 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0922_
timestamp 1607194113
transform 1 0 5520 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_74
timestamp 1607194113
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_62
timestamp 1607194113
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_60
timestamp 1607194113
transform 1 0 6624 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607194113
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_92
timestamp 1607194113
transform 1 0 9568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_86
timestamp 1607194113
transform 1 0 9016 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B1
timestamp 1607194113
transform 1 0 9660 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1258_
timestamp 1607194113
transform 1 0 9844 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1607194113
transform 1 0 11500 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A1_N
timestamp 1607194113
transform 1 0 11316 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1607194113
transform 1 0 13708 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_126
timestamp 1607194113
transform 1 0 12696 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_121
timestamp 1607194113
transform 1 0 12236 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607194113
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1607194113
transform 1 0 13432 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1607194113
transform 1 0 12420 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_156
timestamp 1607194113
transform 1 0 15456 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_149
timestamp 1607194113
transform 1 0 14812 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_i_A
timestamp 1607194113
transform 1 0 15272 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk_i
timestamp 1607194113
transform 1 0 14996 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_160
timestamp 1607194113
transform 1 0 15824 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp 1607194113
transform 1 0 17388 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B2
timestamp 1607194113
transform 1 0 17204 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0706_
timestamp 1607194113
transform 1 0 15916 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_51_193
timestamp 1607194113
transform 1 0 18860 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_179
timestamp 1607194113
transform 1 0 17572 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B
timestamp 1607194113
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607194113
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0805_
timestamp 1607194113
transform 1 0 18032 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_51_217
timestamp 1607194113
transform 1 0 21068 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1607194113
transform 1 0 19964 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B1
timestamp 1607194113
transform 1 0 21160 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1235_
timestamp 1607194113
transform 1 0 19596 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_238
timestamp 1607194113
transform 1 0 23000 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A1_N
timestamp 1607194113
transform 1 0 22816 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1211_
timestamp 1607194113
transform 1 0 21344 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607194113
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_15
timestamp 1607194113
transform 1 0 2484 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1607194113
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_15
timestamp 1607194113
transform 1 0 2484 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1607194113
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1607194113
transform 1 0 2760 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1607194113
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1607194113
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1507_
timestamp 1607194113
transform 1 0 2576 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_53_37
timestamp 1607194113
transform 1 0 4508 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_23
timestamp 1607194113
transform 1 0 3220 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__CLK
timestamp 1607194113
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607194113
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0928_
timestamp 1607194113
transform 1 0 4048 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1607194113
transform 1 0 2944 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_49
timestamp 1607194113
transform 1 0 5612 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_43
timestamp 1607194113
transform 1 0 5060 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B
timestamp 1607194113
transform 1 0 6440 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B
timestamp 1607194113
transform 1 0 4876 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0936_
timestamp 1607194113
transform 1 0 5612 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_52_72
timestamp 1607194113
transform 1 0 7728 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_60
timestamp 1607194113
transform 1 0 6624 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1_N
timestamp 1607194113
transform 1 0 8280 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607194113
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1257_
timestamp 1607194113
transform 1 0 6808 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_53_92
timestamp 1607194113
transform 1 0 9568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_80
timestamp 1607194113
transform 1 0 8464 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_93
timestamp 1607194113
transform 1 0 9660 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_84
timestamp 1607194113
transform 1 0 8832 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B1
timestamp 1607194113
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607194113
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1195_
timestamp 1607194113
transform 1 0 9844 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1607194113
transform 1 0 11500 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_101
timestamp 1607194113
transform 1 0 10396 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A1_N
timestamp 1607194113
transform 1 0 11316 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1385_
timestamp 1607194113
transform 1 0 10488 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_53_127
timestamp 1607194113
transform 1 0 12788 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_123
timestamp 1607194113
transform 1 0 12420 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_121
timestamp 1607194113
transform 1 0 12236 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_123
timestamp 1607194113
transform 1 0 12420 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__CLK
timestamp 1607194113
transform 1 0 12236 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607194113
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_132
timestamp 1607194113
transform 1 0 13248 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_135
timestamp 1607194113
transform 1 0 13524 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_131
timestamp 1607194113
transform 1 0 13156 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk_i
timestamp 1607194113
transform 1 0 13248 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1176_
timestamp 1607194113
transform 1 0 12880 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1181_
timestamp 1607194113
transform 1 0 13708 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_158
timestamp 1607194113
transform 1 0 15640 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_146
timestamp 1607194113
transform 1 0 14536 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_154
timestamp 1607194113
transform 1 0 15272 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1607194113
transform 1 0 14076 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A
timestamp 1607194113
transform 1 0 14352 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607194113
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1255_
timestamp 1607194113
transform 1 0 13984 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_170
timestamp 1607194113
transform 1 0 16744 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_176
timestamp 1607194113
transform 1 0 17296 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_162
timestamp 1607194113
transform 1 0 16008 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A
timestamp 1607194113
transform 1 0 16100 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B
timestamp 1607194113
transform 1 0 16284 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0707_
timestamp 1607194113
transform 1 0 16468 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_53_191
timestamp 1607194113
transform 1 0 18676 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_184
timestamp 1607194113
transform 1 0 18032 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_182
timestamp 1607194113
transform 1 0 17848 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1607194113
transform 1 0 19320 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607194113
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1210_
timestamp 1607194113
transform 1 0 18308 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _0900_
timestamp 1607194113
transform 1 0 18032 0 -1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_53_199
timestamp 1607194113
transform 1 0 19412 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1607194113
transform 1 0 20884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_202
timestamp 1607194113
transform 1 0 19688 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__CLK
timestamp 1607194113
transform 1 0 19688 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1607194113
transform 1 0 19504 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607194113
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1388_
timestamp 1607194113
transform 1 0 19872 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_53_235
timestamp 1607194113
transform 1 0 22724 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_223
timestamp 1607194113
transform 1 0 21620 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1607194113
transform 1 0 21988 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_243
timestamp 1607194113
transform 1 0 23460 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_239
timestamp 1607194113
transform 1 0 23092 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607194113
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1607194113
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1607194113
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1607194113
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_36
timestamp 1607194113
transform 1 0 4416 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1607194113
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607194113
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0861_
timestamp 1607194113
transform 1 0 4048 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_48
timestamp 1607194113
transform 1 0 5520 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1194_
timestamp 1607194113
transform 1 0 5796 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_54_78
timestamp 1607194113
transform 1 0 8280 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_69
timestamp 1607194113
transform 1 0 7452 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A1_N
timestamp 1607194113
transform 1 0 7268 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1607194113
transform 1 0 8004 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1607194113
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_90
timestamp 1607194113
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607194113
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_117
timestamp 1607194113
transform 1 0 11868 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_105
timestamp 1607194113
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_138
timestamp 1607194113
transform 1 0 13800 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1607194113
transform 1 0 13616 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1607194113
transform 1 0 13432 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0913_
timestamp 1607194113
transform 1 0 12144 0 -1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_54_154
timestamp 1607194113
transform 1 0 15272 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_150
timestamp 1607194113
transform 1 0 14904 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607194113
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_178
timestamp 1607194113
transform 1 0 17480 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_166
timestamp 1607194113
transform 1 0 16376 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1607194113
transform 1 0 18032 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1191_
timestamp 1607194113
transform 1 0 18216 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_54_215
timestamp 1607194113
transform 1 0 20884 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_212
timestamp 1607194113
transform 1 0 20608 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_204
timestamp 1607194113
transform 1 0 19872 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1_N
timestamp 1607194113
transform 1 0 19688 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607194113
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1607194113
transform 1 0 20976 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_230
timestamp 1607194113
transform 1 0 22264 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_219
timestamp 1607194113
transform 1 0 21252 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1607194113
transform 1 0 21988 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_242
timestamp 1607194113
transform 1 0 23368 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_15
timestamp 1607194113
transform 1 0 2484 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1607194113
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1607194113
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1508_
timestamp 1607194113
transform 1 0 2576 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_55_37
timestamp 1607194113
transform 1 0 4508 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__CLK
timestamp 1607194113
transform 1 0 4324 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_49
timestamp 1607194113
transform 1 0 5612 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607194113
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1386_
timestamp 1607194113
transform 1 0 6808 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_55_95
timestamp 1607194113
transform 1 0 9844 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_83
timestamp 1607194113
transform 1 0 8740 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__CLK
timestamp 1607194113
transform 1 0 8556 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_115
timestamp 1607194113
transform 1 0 11684 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_107
timestamp 1607194113
transform 1 0 10948 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1
timestamp 1607194113
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_137
timestamp 1607194113
transform 1 0 13708 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1607194113
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607194113
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0911_
timestamp 1607194113
transform 1 0 12420 0 1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_55_151
timestamp 1607194113
transform 1 0 14996 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_145
timestamp 1607194113
transform 1 0 14444 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1189_
timestamp 1607194113
transform 1 0 14628 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_175
timestamp 1607194113
transform 1 0 17204 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_163
timestamp 1607194113
transform 1 0 16100 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_196
timestamp 1607194113
transform 1 0 19136 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1607194113
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1607194113
transform 1 0 19228 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607194113
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_218
timestamp 1607194113
transform 1 0 21160 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1429_
timestamp 1607194113
transform 1 0 19412 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_55_230
timestamp 1607194113
transform 1 0 22264 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_242
timestamp 1607194113
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607194113
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1607194113
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1607194113
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1607194113
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1607194113
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607194113
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0938_
timestamp 1607194113
transform 1 0 4048 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_56_49
timestamp 1607194113
transform 1 0 5612 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 1607194113
transform 1 0 4876 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1427_
timestamp 1607194113
transform 1 0 5704 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_56_71
timestamp 1607194113
transform 1 0 7636 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__CLK
timestamp 1607194113
transform 1 0 7452 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1607194113
transform 1 0 8188 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1607194113
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_80
timestamp 1607194113
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607194113
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_117
timestamp 1607194113
transform 1 0 11868 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_105
timestamp 1607194113
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_134
timestamp 1607194113
transform 1 0 13432 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_130
timestamp 1607194113
transform 1 0 13064 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_123
timestamp 1607194113
transform 1 0 12420 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1607194113
transform 1 0 12880 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1607194113
transform 1 0 13524 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1192_
timestamp 1607194113
transform 1 0 12512 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0896_
timestamp 1607194113
transform 1 0 13708 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_154
timestamp 1607194113
transform 1 0 15272 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1607194113
transform 1 0 14076 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607194113
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_178
timestamp 1607194113
transform 1 0 17480 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_166
timestamp 1607194113
transform 1 0 16376 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_184
timestamp 1607194113
transform 1 0 18032 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__B1
timestamp 1607194113
transform 1 0 18124 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1254_
timestamp 1607194113
transform 1 0 18308 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_56_213
timestamp 1607194113
transform 1 0 20700 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_205
timestamp 1607194113
transform 1 0 19964 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A1_N
timestamp 1607194113
transform 1 0 19780 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607194113
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0920_
timestamp 1607194113
transform 1 0 20884 0 -1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_56_229
timestamp 1607194113
transform 1 0 22172 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_241
timestamp 1607194113
transform 1 0 23276 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_15
timestamp 1607194113
transform 1 0 2484 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1607194113
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1607194113
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1509_
timestamp 1607194113
transform 1 0 2576 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_57_37
timestamp 1607194113
transform 1 0 4508 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__CLK
timestamp 1607194113
transform 1 0 4324 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1607194113
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_47
timestamp 1607194113
transform 1 0 5428 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0880_
timestamp 1607194113
transform 1 0 5060 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_74
timestamp 1607194113
transform 1 0 7912 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1607194113
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607194113
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8004 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_57_88
timestamp 1607194113
transform 1 0 9200 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_108
timestamp 1607194113
transform 1 0 11040 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_100
timestamp 1607194113
transform 1 0 10304 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0903_
timestamp 1607194113
transform 1 0 10396 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__B1
timestamp 1607194113
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607194113
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1193_
timestamp 1607194113
transform 1 0 12420 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1607194113
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_139
timestamp 1607194113
transform 1 0 13892 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1607194113
transform 1 0 14444 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0897_
timestamp 1607194113
transform 1 0 14628 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_175
timestamp 1607194113
transform 1 0 17204 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_163
timestamp 1607194113
transform 1 0 16100 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_192
timestamp 1607194113
transform 1 0 18768 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_184
timestamp 1607194113
transform 1 0 18032 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1607194113
transform 1 0 19228 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607194113
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1252_
timestamp 1607194113
transform 1 0 18860 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_199
timestamp 1607194113
transform 1 0 19412 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B1
timestamp 1607194113
transform 1 0 19780 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1190_
timestamp 1607194113
transform 1 0 19964 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_57_235
timestamp 1607194113
transform 1 0 22724 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_223
timestamp 1607194113
transform 1 0 21620 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A1_N
timestamp 1607194113
transform 1 0 21436 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1607194113
transform 1 0 23460 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607194113
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1607194113
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1607194113
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1607194113
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_32
timestamp 1607194113
transform 1 0 4048 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1607194113
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607194113
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_49
timestamp 1607194113
transform 1 0 5612 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _0894_
timestamp 1607194113
transform 1 0 4784 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_73
timestamp 1607194113
transform 1 0 7820 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_61
timestamp 1607194113
transform 1 0 6716 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1607194113
transform 1 0 9292 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1607194113
transform 1 0 8924 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1607194113
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607194113
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _0909_
timestamp 1607194113
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_117
timestamp 1607194113
transform 1 0 11868 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_105
timestamp 1607194113
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_125
timestamp 1607194113
transform 1 0 12604 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B1
timestamp 1607194113
transform 1 0 12788 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1256_
timestamp 1607194113
transform 1 0 12972 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_58_145
timestamp 1607194113
transform 1 0 14444 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1607194113
transform 1 0 15548 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607194113
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1607194113
transform 1 0 15272 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_171
timestamp 1607194113
transform 1 0 16836 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_159
timestamp 1607194113
transform 1 0 15732 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_191
timestamp 1607194113
transform 1 0 18676 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_183
timestamp 1607194113
transform 1 0 17940 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0898_
timestamp 1607194113
transform 1 0 18768 0 -1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_58_210
timestamp 1607194113
transform 1 0 20424 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1
timestamp 1607194113
transform 1 0 20240 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1607194113
transform 1 0 20056 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__B1
timestamp 1607194113
transform 1 0 20608 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607194113
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1253_
timestamp 1607194113
transform 1 0 20884 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1607194113
transform 1 0 22540 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A1_N
timestamp 1607194113
transform 1 0 22356 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1607194113
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1607194113
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_15
timestamp 1607194113
transform 1 0 2484 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1607194113
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1607194113
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1607194113
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1510_
timestamp 1607194113
transform 1 0 2576 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_60_32
timestamp 1607194113
transform 1 0 4048 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1607194113
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_37
timestamp 1607194113
transform 1 0 4508 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__CLK
timestamp 1607194113
transform 1 0 4324 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607194113
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0884_
timestamp 1607194113
transform 1 0 4416 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_60_45
timestamp 1607194113
transform 1 0 5244 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_52
timestamp 1607194113
transform 1 0 5888 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0888_
timestamp 1607194113
transform 1 0 5980 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0886_
timestamp 1607194113
transform 1 0 5060 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_74
timestamp 1607194113
transform 1 0 7912 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_62
timestamp 1607194113
transform 1 0 6808 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_74
timestamp 1607194113
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_62
timestamp 1607194113
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_60
timestamp 1607194113
transform 1 0 6624 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607194113
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_86
timestamp 1607194113
transform 1 0 9016 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_94
timestamp 1607194113
transform 1 0 9752 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_86
timestamp 1607194113
transform 1 0 9016 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1607194113
transform 1 0 9568 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607194113
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0917_
timestamp 1607194113
transform 1 0 9660 0 -1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0868_
timestamp 1607194113
transform 1 0 9200 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_118
timestamp 1607194113
transform 1 0 11960 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_106
timestamp 1607194113
transform 1 0 10856 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_118
timestamp 1607194113
transform 1 0 11960 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1
timestamp 1607194113
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1607194113
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1607194113
transform 1 0 11408 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0937_
timestamp 1607194113
transform 1 0 10304 0 1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1607194113
transform 1 0 11592 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_130
timestamp 1607194113
transform 1 0 13064 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_135
timestamp 1607194113
transform 1 0 13524 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1607194113
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__CLK
timestamp 1607194113
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607194113
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1607194113
transform 1 0 13800 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_151
timestamp 1607194113
transform 1 0 14996 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_143
timestamp 1607194113
transform 1 0 14260 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1607194113
transform 1 0 14076 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1607194113
transform 1 0 15640 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607194113
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1387_
timestamp 1607194113
transform 1 0 13984 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0923_
timestamp 1607194113
transform 1 0 15272 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_172
timestamp 1607194113
transform 1 0 16928 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_160
timestamp 1607194113
transform 1 0 15824 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_171
timestamp 1607194113
transform 1 0 16836 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_159
timestamp 1607194113
transform 1 0 15732 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A
timestamp 1607194113
transform 1 0 16744 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1236_
timestamp 1607194113
transform 1 0 16376 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_196
timestamp 1607194113
transform 1 0 19136 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_184
timestamp 1607194113
transform 1 0 18032 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_196
timestamp 1607194113
transform 1 0 19136 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1607194113
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607194113
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_208
timestamp 1607194113
transform 1 0 20240 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_202
timestamp 1607194113
transform 1 0 19688 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__B1
timestamp 1607194113
transform 1 0 19780 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607194113
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1198_
timestamp 1607194113
transform 1 0 19964 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1196_
timestamp 1607194113
transform 1 0 20884 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_237
timestamp 1607194113
transform 1 0 22908 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_219
timestamp 1607194113
transform 1 0 21252 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_233
timestamp 1607194113
transform 1 0 22540 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_221
timestamp 1607194113
transform 1 0 21436 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1607194113
transform 1 0 22356 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1266_
timestamp 1607194113
transform 1 0 22540 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1203_
timestamp 1607194113
transform 1 0 22172 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_241
timestamp 1607194113
transform 1 0 23276 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607194113
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1607194113
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1607194113
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1607194113
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1511_
timestamp 1607194113
transform 1 0 3588 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_61_48
timestamp 1607194113
transform 1 0 5520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__CLK
timestamp 1607194113
transform 1 0 5336 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_71
timestamp 1607194113
transform 1 0 7636 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_60
timestamp 1607194113
transform 1 0 6624 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607194113
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0892_
timestamp 1607194113
transform 1 0 6808 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_61_95
timestamp 1607194113
transform 1 0 9844 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_83
timestamp 1607194113
transform 1 0 8740 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B1
timestamp 1607194113
transform 1 0 10120 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_114
timestamp 1607194113
transform 1 0 11592 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A1
timestamp 1607194113
transform 1 0 11408 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0916_
timestamp 1607194113
transform 1 0 10304 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_123
timestamp 1607194113
transform 1 0 12420 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1607194113
transform 1 0 13156 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607194113
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1428_
timestamp 1607194113
transform 1 0 13340 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_61_152
timestamp 1607194113
transform 1 0 15088 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1607194113
transform 1 0 15640 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_176
timestamp 1607194113
transform 1 0 17296 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_164
timestamp 1607194113
transform 1 0 16192 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0924_
timestamp 1607194113
transform 1 0 15824 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1607194113
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1607194113
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_182
timestamp 1607194113
transform 1 0 17848 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607194113
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_208
timestamp 1607194113
transform 1 0 20240 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1383_
timestamp 1607194113
transform 1 0 20332 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_61_230
timestamp 1607194113
transform 1 0 22264 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__CLK
timestamp 1607194113
transform 1 0 22080 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_242
timestamp 1607194113
transform 1 0 23368 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607194113
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1607194113
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1607194113
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1607194113
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_32
timestamp 1607194113
transform 1 0 4048 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1607194113
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607194113
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_50
timestamp 1607194113
transform 1 0 5704 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_40
timestamp 1607194113
transform 1 0 4784 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0879_
timestamp 1607194113
transform 1 0 4876 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0862_
timestamp 1607194113
transform 1 0 6440 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_74
timestamp 1607194113
transform 1 0 7912 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_62
timestamp 1607194113
transform 1 0 6808 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_93
timestamp 1607194113
transform 1 0 9660 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_86
timestamp 1607194113
transform 1 0 9016 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607194113
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_112
timestamp 1607194113
transform 1 0 11408 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_101
timestamp 1607194113
transform 1 0 10396 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1607194113
transform 1 0 11224 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0915_
timestamp 1607194113
transform 1 0 10580 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_136
timestamp 1607194113
transform 1 0 13616 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_124
timestamp 1607194113
transform 1 0 12512 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_158
timestamp 1607194113
transform 1 0 15640 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_152
timestamp 1607194113
transform 1 0 15088 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_148
timestamp 1607194113
transform 1 0 14720 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607194113
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1182_
timestamp 1607194113
transform 1 0 15272 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_176
timestamp 1607194113
transform 1 0 17296 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_166
timestamp 1607194113
transform 1 0 16376 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1607194113
transform 1 0 17112 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0703_
timestamp 1607194113
transform 1 0 16468 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_188
timestamp 1607194113
transform 1 0 18400 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_215
timestamp 1607194113
transform 1 0 20884 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_212
timestamp 1607194113
transform 1 0 20608 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_200
timestamp 1607194113
transform 1 0 19504 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607194113
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1424_
timestamp 1607194113
transform 1 0 20976 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1607194113
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__CLK
timestamp 1607194113
transform 1 0 22724 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1607194113
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1607194113
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1607194113
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_39
timestamp 1607194113
transform 1 0 4692 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1607194113
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_52
timestamp 1607194113
transform 1 0 5888 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0877_
timestamp 1607194113
transform 1 0 5060 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1607194113
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1607194113
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_60
timestamp 1607194113
transform 1 0 6624 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607194113
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_98
timestamp 1607194113
transform 1 0 10120 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1607194113
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_109
timestamp 1607194113
transform 1 0 11132 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_104
timestamp 1607194113
transform 1 0 10672 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1607194113
transform 1 0 10764 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_135
timestamp 1607194113
transform 1 0 13524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1607194113
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_121
timestamp 1607194113
transform 1 0 12236 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607194113
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_147
timestamp 1607194113
transform 1 0 14628 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__B1
timestamp 1607194113
transform 1 0 14904 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1183_
timestamp 1607194113
transform 1 0 15088 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_168
timestamp 1607194113
transform 1 0 16560 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_197
timestamp 1607194113
transform 1 0 19228 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_193
timestamp 1607194113
transform 1 0 18860 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_180
timestamp 1607194113
transform 1 0 17664 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B
timestamp 1607194113
transform 1 0 18676 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__B1
timestamp 1607194113
transform 1 0 19320 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607194113
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0802_
timestamp 1607194113
transform 1 0 18032 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_63_216
timestamp 1607194113
transform 1 0 20976 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1261_
timestamp 1607194113
transform 1 0 19504 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_227
timestamp 1607194113
transform 1 0 21988 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1607194113
transform 1 0 21712 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_243
timestamp 1607194113
transform 1 0 23460 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_239
timestamp 1607194113
transform 1 0 23092 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607194113
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1607194113
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1607194113
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1607194113
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_32
timestamp 1607194113
transform 1 0 4048 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1607194113
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1607194113
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_40
timestamp 1607194113
transform 1 0 4784 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1512_
timestamp 1607194113
transform 1 0 4968 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1607194113
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1607194113
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__CLK
timestamp 1607194113
transform 1 0 6716 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_99
timestamp 1607194113
transform 1 0 10212 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1607194113
transform 1 0 9660 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_91
timestamp 1607194113
transform 1 0 9476 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_87
timestamp 1607194113
transform 1 0 9108 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1607194113
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0882_
timestamp 1607194113
transform 1 0 9844 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _0883_
timestamp 1607194113
transform 1 0 10948 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_64_133
timestamp 1607194113
transform 1 0 13340 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1607194113
transform 1 0 12236 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_145
timestamp 1607194113
transform 1 0 14444 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__B1
timestamp 1607194113
transform 1 0 14996 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1607194113
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1184_
timestamp 1607194113
transform 1 0 15272 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1607194113
transform 1 0 16928 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1_N
timestamp 1607194113
transform 1 0 16744 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B1
timestamp 1607194113
transform 1 0 17296 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1246_
timestamp 1607194113
transform 1 0 17480 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_194
timestamp 1607194113
transform 1 0 18952 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_206
timestamp 1607194113
transform 1 0 20056 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_202
timestamp 1607194113
transform 1 0 19688 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1607194113
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1259_
timestamp 1607194113
transform 1 0 20884 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1607194113
transform 1 0 19780 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1607194113
transform 1 0 22540 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1607194113
transform 1 0 21436 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A
timestamp 1607194113
transform 1 0 21252 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_15
timestamp 1607194113
transform 1 0 2484 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1607194113
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1607194113
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1344_
timestamp 1607194113
transform 1 0 2576 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_65_39
timestamp 1607194113
transform 1 0 4692 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__CLK
timestamp 1607194113
transform 1 0 4508 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__D
timestamp 1607194113
transform 1 0 4324 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_55
timestamp 1607194113
transform 1 0 6164 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_43
timestamp 1607194113
transform 1 0 5060 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B
timestamp 1607194113
transform 1 0 5980 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0873_
timestamp 1607194113
transform 1 0 5152 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_71
timestamp 1607194113
transform 1 0 7636 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1607194113
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0875_
timestamp 1607194113
transform 1 0 6808 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_65_95
timestamp 1607194113
transform 1 0 9844 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_83
timestamp 1607194113
transform 1 0 8740 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0891_
timestamp 1607194113
transform 1 0 10120 0 1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_65_112
timestamp 1607194113
transform 1 0 11408 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_135
timestamp 1607194113
transform 1 0 13524 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_123
timestamp 1607194113
transform 1 0 12420 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_120
timestamp 1607194113
transform 1 0 12144 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1607194113
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_154
timestamp 1607194113
transform 1 0 15272 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_146
timestamp 1607194113
transform 1 0 14536 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_139
timestamp 1607194113
transform 1 0 13892 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1607194113
transform 1 0 14352 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B1
timestamp 1607194113
transform 1 0 15548 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1248_
timestamp 1607194113
transform 1 0 13984 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_177
timestamp 1607194113
transform 1 0 17388 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1_N
timestamp 1607194113
transform 1 0 17204 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1247_
timestamp 1607194113
transform 1 0 15732 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_65_192
timestamp 1607194113
transform 1 0 18768 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_184
timestamp 1607194113
transform 1 0 18032 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1607194113
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1394_
timestamp 1607194113
transform 1 0 18952 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_215
timestamp 1607194113
transform 1 0 20884 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__CLK
timestamp 1607194113
transform 1 0 20700 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_227
timestamp 1607194113
transform 1 0 21988 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_243
timestamp 1607194113
transform 1 0 23460 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_239
timestamp 1607194113
transform 1 0 23092 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1607194113
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_15
timestamp 1607194113
transform 1 0 2484 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1607194113
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1607194113
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1607194113
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1607194113
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1607194113
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1514_
timestamp 1607194113
transform 1 0 2668 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_67_38
timestamp 1607194113
transform 1 0 4600 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_66_32
timestamp 1607194113
transform 1 0 4048 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1607194113
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__CLK
timestamp 1607194113
transform 1 0 4416 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1607194113
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1513_
timestamp 1607194113
transform 1 0 4324 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_67_53
timestamp 1607194113
transform 1 0 5980 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_56
timestamp 1607194113
transform 1 0 6256 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__CLK
timestamp 1607194113
transform 1 0 6072 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0871_
timestamp 1607194113
transform 1 0 5152 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_67_74
timestamp 1607194113
transform 1 0 7912 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1607194113
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_64
timestamp 1607194113
transform 1 0 6992 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B1
timestamp 1607194113
transform 1 0 7176 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A1
timestamp 1607194113
transform 1 0 7360 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1607194113
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0893_
timestamp 1607194113
transform 1 0 7544 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_67_98
timestamp 1607194113
transform 1 0 10120 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_86
timestamp 1607194113
transform 1 0 9016 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_98
timestamp 1607194113
transform 1 0 10120 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_93
timestamp 1607194113
transform 1 0 9660 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_84
timestamp 1607194113
transform 1 0 8832 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1607194113
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0864_
timestamp 1607194113
transform 1 0 9752 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_118
timestamp 1607194113
transform 1 0 11960 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B1
timestamp 1607194113
transform 1 0 11776 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A1
timestamp 1607194113
transform 1 0 11592 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0887_
timestamp 1607194113
transform 1 0 10304 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _0885_
timestamp 1607194113
transform 1 0 10856 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_67_135
timestamp 1607194113
transform 1 0 13524 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_123
timestamp 1607194113
transform 1 0 12420 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_132
timestamp 1607194113
transform 1 0 13248 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_124
timestamp 1607194113
transform 1 0 12512 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B1
timestamp 1607194113
transform 1 0 12328 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A1
timestamp 1607194113
transform 1 0 12144 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1607194113
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0869_
timestamp 1607194113
transform 1 0 12880 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_152
timestamp 1607194113
transform 1 0 15088 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_144
timestamp 1607194113
transform 1 0 14352 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__B2
timestamp 1607194113
transform 1 0 14904 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__B1
timestamp 1607194113
transform 1 0 14076 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__B1
timestamp 1607194113
transform 1 0 14720 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1607194113
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1249_
timestamp 1607194113
transform 1 0 15272 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1186_
timestamp 1607194113
transform 1 0 14260 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_67_174
timestamp 1607194113
transform 1 0 17112 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1607194113
transform 1 0 16468 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1607194113
transform 1 0 15916 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_172
timestamp 1607194113
transform 1 0 16928 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A
timestamp 1607194113
transform 1 0 16928 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A1_N
timestamp 1607194113
transform 1 0 16744 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1_N
timestamp 1607194113
transform 1 0 15732 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1245_
timestamp 1607194113
transform 1 0 16560 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_187
timestamp 1607194113
transform 1 0 18308 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1607194113
transform 1 0 17848 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_196
timestamp 1607194113
transform 1 0 19136 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_184
timestamp 1607194113
transform 1 0 18032 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1607194113
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1607194113
transform 1 0 18032 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_215
timestamp 1607194113
transform 1 0 20884 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_213
timestamp 1607194113
transform 1 0 20700 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_205
timestamp 1607194113
transform 1 0 19964 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__CLK
timestamp 1607194113
transform 1 0 21160 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1607194113
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1435_
timestamp 1607194113
transform 1 0 19412 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1607194113
transform 1 0 19688 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_232
timestamp 1607194113
transform 1 0 22448 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_220
timestamp 1607194113
transform 1 0 21344 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_227
timestamp 1607194113
transform 1 0 21988 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_240
timestamp 1607194113
transform 1 0 23184 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_239
timestamp 1607194113
transform 1 0 23092 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A1_N
timestamp 1607194113
transform 1 0 23460 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A1_N
timestamp 1607194113
transform 1 0 23368 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1607194113
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1607194113
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1607194113
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1607194113
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_32
timestamp 1607194113
transform 1 0 4048 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1607194113
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B1
timestamp 1607194113
transform 1 0 4232 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1607194113
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1188_
timestamp 1607194113
transform 1 0 4416 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_54
timestamp 1607194113
transform 1 0 6072 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1_N
timestamp 1607194113
transform 1 0 5888 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_78
timestamp 1607194113
transform 1 0 8280 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_66
timestamp 1607194113
transform 1 0 7176 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_93
timestamp 1607194113
transform 1 0 9660 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_90
timestamp 1607194113
transform 1 0 9384 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1607194113
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_101
timestamp 1607194113
transform 1 0 10396 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B1
timestamp 1607194113
transform 1 0 10488 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1187_
timestamp 1607194113
transform 1 0 10672 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_131
timestamp 1607194113
transform 1 0 13156 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_120
timestamp 1607194113
transform 1 0 12144 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1607194113
transform 1 0 12696 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1607194113
transform 1 0 12880 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_154
timestamp 1607194113
transform 1 0 15272 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_151
timestamp 1607194113
transform 1 0 14996 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_143
timestamp 1607194113
transform 1 0 14260 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1607194113
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1433_
timestamp 1607194113
transform 1 0 16376 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_196
timestamp 1607194113
transform 1 0 19136 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_187
timestamp 1607194113
transform 1 0 18308 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__CLK
timestamp 1607194113
transform 1 0 18124 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1607194113
transform 1 0 18860 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_215
timestamp 1607194113
transform 1 0 20884 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_208
timestamp 1607194113
transform 1 0 20240 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1607194113
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_235
timestamp 1607194113
transform 1 0 22724 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_227
timestamp 1607194113
transform 1 0 21988 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B1
timestamp 1607194113
transform 1 0 22908 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1_N
timestamp 1607194113
transform 1 0 23092 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0784_
timestamp 1607194113
transform 1 0 23276 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_15
timestamp 1607194113
transform 1 0 2484 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1607194113
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1607194113
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1390_
timestamp 1607194113
transform 1 0 2852 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__CLK
timestamp 1607194113
transform 1 0 4600 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_53
timestamp 1607194113
transform 1 0 5980 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_48
timestamp 1607194113
transform 1 0 5520 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_40
timestamp 1607194113
transform 1 0 4784 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1607194113
transform 1 0 5704 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_68
timestamp 1607194113
transform 1 0 7360 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_62
timestamp 1607194113
transform 1 0 6808 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1607194113
transform 1 0 6900 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1607194113
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1607194113
transform 1 0 7084 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_92
timestamp 1607194113
transform 1 0 9568 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_80
timestamp 1607194113
transform 1 0 8464 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B1
timestamp 1607194113
transform 1 0 9752 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1250_
timestamp 1607194113
transform 1 0 9936 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_69_116
timestamp 1607194113
transform 1 0 11776 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__A2_N
timestamp 1607194113
transform 1 0 11592 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B2
timestamp 1607194113
transform 1 0 11408 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_136
timestamp 1607194113
transform 1 0 13616 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_129
timestamp 1607194113
transform 1 0 12972 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_123
timestamp 1607194113
transform 1 0 12420 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1607194113
transform 1 0 13432 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1607194113
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1185_
timestamp 1607194113
transform 1 0 13064 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_148
timestamp 1607194113
transform 1 0 14720 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_178
timestamp 1607194113
transform 1 0 17480 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_172
timestamp 1607194113
transform 1 0 16928 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_160
timestamp 1607194113
transform 1 0 15824 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B2
timestamp 1607194113
transform 1 0 17572 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A2
timestamp 1607194113
transform 1 0 17756 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1607194113
transform 1 0 19320 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1607194113
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0870_
timestamp 1607194113
transform 1 0 18032 0 1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_69_214
timestamp 1607194113
transform 1 0 20792 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_202
timestamp 1607194113
transform 1 0 19688 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1607194113
transform 1 0 19504 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_238
timestamp 1607194113
transform 1 0 23000 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_226
timestamp 1607194113
transform 1 0 21896 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_243
timestamp 1607194113
transform 1 0 23460 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A1_N
timestamp 1607194113
transform 1 0 23276 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B1
timestamp 1607194113
transform 1 0 23092 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1607194113
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1607194113
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1607194113
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1607194113
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_32
timestamp 1607194113
transform 1 0 4048 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_27
timestamp 1607194113
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1607194113
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__CLK
timestamp 1607194113
transform 1 0 6532 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1431_
timestamp 1607194113
transform 1 0 4784 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_73
timestamp 1607194113
transform 1 0 7820 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_61
timestamp 1607194113
transform 1 0 6716 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_93
timestamp 1607194113
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1607194113
transform 1 0 9476 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_85
timestamp 1607194113
transform 1 0 8924 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1607194113
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_105
timestamp 1607194113
transform 1 0 10764 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1391_
timestamp 1607194113
transform 1 0 10856 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_138
timestamp 1607194113
transform 1 0 13800 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_127
timestamp 1607194113
transform 1 0 12788 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__CLK
timestamp 1607194113
transform 1 0 12604 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1607194113
transform 1 0 13616 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1607194113
transform 1 0 13340 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_154
timestamp 1607194113
transform 1 0 15272 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_150
timestamp 1607194113
transform 1 0 14904 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1607194113
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_166
timestamp 1607194113
transform 1 0 16376 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1392_
timestamp 1607194113
transform 1 0 16652 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_190
timestamp 1607194113
transform 1 0 18584 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__CLK
timestamp 1607194113
transform 1 0 18400 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_215
timestamp 1607194113
transform 1 0 20884 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_202
timestamp 1607194113
transform 1 0 19688 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1607194113
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_227
timestamp 1607194113
transform 1 0 21988 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_239
timestamp 1607194113
transform 1 0 23092 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_71_15
timestamp 1607194113
transform 1 0 2484 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1607194113
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1607194113
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A1_N
timestamp 1607194113
transform 1 0 4692 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B1
timestamp 1607194113
transform 1 0 3036 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1251_
timestamp 1607194113
transform 1 0 3220 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_71_58
timestamp 1607194113
transform 1 0 6440 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_50
timestamp 1607194113
transform 1 0 5704 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_45
timestamp 1607194113
transform 1 0 5244 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A2_N
timestamp 1607194113
transform 1 0 5060 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B2
timestamp 1607194113
transform 1 0 4876 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1607194113
transform 1 0 5428 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_74
timestamp 1607194113
transform 1 0 7912 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_62
timestamp 1607194113
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1607194113
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_82
timestamp 1607194113
transform 1 0 8648 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A1
timestamp 1607194113
transform 1 0 10120 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0876_
timestamp 1607194113
transform 1 0 8832 0 1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_71_118
timestamp 1607194113
transform 1 0 11960 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_106
timestamp 1607194113
transform 1 0 10856 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B2
timestamp 1607194113
transform 1 0 10672 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A2
timestamp 1607194113
transform 1 0 10488 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B1
timestamp 1607194113
transform 1 0 10304 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1607194113
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1432_
timestamp 1607194113
transform 1 0 12420 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_156
timestamp 1607194113
transform 1 0 15456 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_144
timestamp 1607194113
transform 1 0 14352 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1607194113
transform 1 0 14168 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_168
timestamp 1607194113
transform 1 0 16560 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_190
timestamp 1607194113
transform 1 0 18584 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_71_180
timestamp 1607194113
transform 1 0 17664 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A
timestamp 1607194113
transform 1 0 18400 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1607194113
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1241_
timestamp 1607194113
transform 1 0 19136 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1237_
timestamp 1607194113
transform 1 0 18032 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_214
timestamp 1607194113
transform 1 0 20792 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_202
timestamp 1607194113
transform 1 0 19688 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A
timestamp 1607194113
transform 1 0 19504 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_238
timestamp 1607194113
transform 1 0 23000 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_226
timestamp 1607194113
transform 1 0 21896 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1607194113
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_11
timestamp 1607194113
transform 1 0 2116 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_3
timestamp 1607194113
transform 1 0 1380 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1607194113
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1607194113
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__D
timestamp 1607194113
transform 1 0 2392 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1607194113
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1607194113
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1345_
timestamp 1607194113
transform 1 0 2576 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_73_37
timestamp 1607194113
transform 1 0 4508 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1607194113
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__CLK
timestamp 1607194113
transform 1 0 4324 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1607194113
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1180_
timestamp 1607194113
transform 1 0 4048 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_48
timestamp 1607194113
transform 1 0 5520 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_50
timestamp 1607194113
transform 1 0 5704 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A1_N
timestamp 1607194113
transform 1 0 5520 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1607194113
transform 1 0 5244 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_74
timestamp 1607194113
transform 1 0 7912 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_62
timestamp 1607194113
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_60
timestamp 1607194113
transform 1 0 6624 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_62
timestamp 1607194113
transform 1 0 6808 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B1
timestamp 1607194113
transform 1 0 7176 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1607194113
transform 1 0 7360 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1607194113
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0878_
timestamp 1607194113
transform 1 0 7544 0 -1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_73_86
timestamp 1607194113
transform 1 0 9016 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_88
timestamp 1607194113
transform 1 0 9200 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B2
timestamp 1607194113
transform 1 0 9016 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1607194113
transform 1 0 8832 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_90
timestamp 1607194113
transform 1 0 9384 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B1
timestamp 1607194113
transform 1 0 9476 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B1
timestamp 1607194113
transform 1 0 9384 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1607194113
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1243_
timestamp 1607194113
transform 1 0 9660 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1179_
timestamp 1607194113
transform 1 0 9660 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_73_119
timestamp 1607194113
transform 1 0 12052 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_111
timestamp 1607194113
transform 1 0 11316 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_115
timestamp 1607194113
transform 1 0 11684 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A2_N
timestamp 1607194113
transform 1 0 11500 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B2
timestamp 1607194113
transform 1 0 11316 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A1_N
timestamp 1607194113
transform 1 0 11132 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1_N
timestamp 1607194113
transform 1 0 11132 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_138
timestamp 1607194113
transform 1 0 13800 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_126
timestamp 1607194113
transform 1 0 12696 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_135
timestamp 1607194113
transform 1 0 13524 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_127
timestamp 1607194113
transform 1 0 12788 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1607194113
transform 1 0 13800 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1607194113
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1607194113
transform 1 0 12420 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_156
timestamp 1607194113
transform 1 0 15456 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_150
timestamp 1607194113
transform 1 0 14904 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_154
timestamp 1607194113
transform 1 0 15272 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_152
timestamp 1607194113
transform 1 0 15088 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_144
timestamp 1607194113
transform 1 0 14352 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B2
timestamp 1607194113
transform 1 0 15548 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1607194113
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1177_
timestamp 1607194113
transform 1 0 13984 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_166
timestamp 1607194113
transform 1 0 16376 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A2
timestamp 1607194113
transform 1 0 15732 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1607194113
transform 1 0 17388 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1607194113
transform 1 0 17204 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B1
timestamp 1607194113
transform 1 0 16560 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1242_
timestamp 1607194113
transform 1 0 16744 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0874_
timestamp 1607194113
transform 1 0 15916 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_72_190
timestamp 1607194113
transform 1 0 18584 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B2
timestamp 1607194113
transform 1 0 18400 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B2
timestamp 1607194113
transform 1 0 17572 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A2
timestamp 1607194113
transform 1 0 17756 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1_N
timestamp 1607194113
transform 1 0 18216 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A1
timestamp 1607194113
transform 1 0 19320 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1607194113
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0872_
timestamp 1607194113
transform 1 0 18032 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_73_209
timestamp 1607194113
transform 1 0 20332 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_202
timestamp 1607194113
transform 1 0 19688 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_215
timestamp 1607194113
transform 1 0 20884 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_202
timestamp 1607194113
transform 1 0 19688 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B1
timestamp 1607194113
transform 1 0 19504 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1607194113
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1607194113
transform 1 0 20056 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_233
timestamp 1607194113
transform 1 0 22540 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_221
timestamp 1607194113
transform 1 0 21436 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_227
timestamp 1607194113
transform 1 0 21988 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B1
timestamp 1607194113
transform 1 0 22908 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_243
timestamp 1607194113
transform 1 0 23460 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_239
timestamp 1607194113
transform 1 0 23092 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A1_N
timestamp 1607194113
transform 1 0 23460 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A2_N
timestamp 1607194113
transform 1 0 23092 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B2
timestamp 1607194113
transform 1 0 23276 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1607194113
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1607194113
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1607194113
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1607194113
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_32
timestamp 1607194113
transform 1 0 4048 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1607194113
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1607194113
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__CLK
timestamp 1607194113
transform 1 0 6532 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1395_
timestamp 1607194113
transform 1 0 4784 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_73
timestamp 1607194113
transform 1 0 7820 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_61
timestamp 1607194113
transform 1 0 6716 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_93
timestamp 1607194113
transform 1 0 9660 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1607194113
transform 1 0 9476 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1607194113
transform 1 0 8924 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1607194113
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1396_
timestamp 1607194113
transform 1 0 10396 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_131
timestamp 1607194113
transform 1 0 13156 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_122
timestamp 1607194113
transform 1 0 12328 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__CLK
timestamp 1607194113
transform 1 0 12144 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1607194113
transform 1 0 12880 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_143
timestamp 1607194113
transform 1 0 14260 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A2_N
timestamp 1607194113
transform 1 0 15272 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B1
timestamp 1607194113
transform 1 0 14996 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1607194113
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1178_
timestamp 1607194113
transform 1 0 15456 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_74_174
timestamp 1607194113
transform 1 0 17112 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A1_N
timestamp 1607194113
transform 1 0 16928 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1397_
timestamp 1607194113
transform 1 0 17664 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_215
timestamp 1607194113
transform 1 0 20884 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_213
timestamp 1607194113
transform 1 0 20700 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_201
timestamp 1607194113
transform 1 0 19596 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__CLK
timestamp 1607194113
transform 1 0 19412 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1607194113
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_227
timestamp 1607194113
transform 1 0 21988 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_239
timestamp 1607194113
transform 1 0 23092 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A2_N
timestamp 1607194113
transform 1 0 23184 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B2
timestamp 1607194113
transform 1 0 23368 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B1
timestamp 1607194113
transform 1 0 23552 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1607194113
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1607194113
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1607194113
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_27
timestamp 1607194113
transform 1 0 3588 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1436_
timestamp 1607194113
transform 1 0 3680 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_49
timestamp 1607194113
transform 1 0 5612 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__CLK
timestamp 1607194113
transform 1 0 5428 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_77
timestamp 1607194113
transform 1 0 8188 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_65
timestamp 1607194113
transform 1 0 7084 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1607194113
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1607194113
transform 1 0 6808 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_89
timestamp 1607194113
transform 1 0 9292 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1437_
timestamp 1607194113
transform 1 0 9844 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_75_116
timestamp 1607194113
transform 1 0 11776 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__CLK
timestamp 1607194113
transform 1 0 11592 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_135
timestamp 1607194113
transform 1 0 13524 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_123
timestamp 1607194113
transform 1 0 12420 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1607194113
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_147
timestamp 1607194113
transform 1 0 14628 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_171
timestamp 1607194113
transform 1 0 16836 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_159
timestamp 1607194113
transform 1 0 15732 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1607194113
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1438_
timestamp 1607194113
transform 1 0 18032 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_217
timestamp 1607194113
transform 1 0 21068 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1607194113
transform 1 0 19964 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__CLK
timestamp 1607194113
transform 1 0 19780 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_229
timestamp 1607194113
transform 1 0 22172 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_241
timestamp 1607194113
transform 1 0 23276 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B1
timestamp 1607194113
transform 1 0 23368 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1607194113
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1607194113
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1607194113
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1607194113
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_32
timestamp 1607194113
transform 1 0 4048 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1607194113
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1607194113
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1244_
timestamp 1607194113
transform 1 0 4416 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_58
timestamp 1607194113
transform 1 0 6440 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A2_N
timestamp 1607194113
transform 1 0 6256 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B2
timestamp 1607194113
transform 1 0 6072 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A1_N
timestamp 1607194113
transform 1 0 5888 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_75
timestamp 1607194113
transform 1 0 8004 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_63
timestamp 1607194113
transform 1 0 6900 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1607194113
transform 1 0 6808 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_94
timestamp 1607194113
transform 1 0 9752 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_87
timestamp 1607194113
transform 1 0 9108 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1607194113
transform 1 0 9660 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_118
timestamp 1607194113
transform 1 0 11960 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_106
timestamp 1607194113
transform 1 0 10856 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_137
timestamp 1607194113
transform 1 0 13708 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_125
timestamp 1607194113
transform 1 0 12604 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1607194113
transform 1 0 12512 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_156
timestamp 1607194113
transform 1 0 15456 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_149
timestamp 1607194113
transform 1 0 14812 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1607194113
transform 1 0 15364 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_168
timestamp 1607194113
transform 1 0 16560 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_196
timestamp 1607194113
transform 1 0 19136 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_187
timestamp 1607194113
transform 1 0 18308 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_76_180
timestamp 1607194113
transform 1 0 17664 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1607194113
transform 1 0 18216 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1607194113
transform 1 0 18860 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_218
timestamp 1607194113
transform 1 0 21160 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_216
timestamp 1607194113
transform 1 0 20976 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_208
timestamp 1607194113
transform 1 0 20240 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1607194113
transform 1 0 21068 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_230
timestamp 1607194113
transform 1 0 22264 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_242
timestamp 1607194113
transform 1 0 23368 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1607194113
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1607194113
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1607194113
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1607194113
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607194113
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1607194113
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1607194113
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1607194113
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1607194113
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607194113
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_301
timestamp 1607194113
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1607194113
transform 1 0 28060 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_300
timestamp 1607194113
transform 1 0 28704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_292
timestamp 1607194113
transform 1 0 27968 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1607194113
transform -1 0 29256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1607194113
transform -1 0 29256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1607194113
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1607194113
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1607194113
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1607194113
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1607194113
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1607194113
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1607194113
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1607194113
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_301
timestamp 1607194113
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_293
timestamp 1607194113
transform 1 0 28060 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_300
timestamp 1607194113
transform 1 0 28704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1607194113
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607194113
transform -1 0 29256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607194113
transform -1 0 29256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1607194113
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1607194113
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1607194113
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1607194113
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_300
timestamp 1607194113
transform 1 0 28704 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1607194113
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607194113
transform -1 0 29256 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_263
timestamp 1607194113
transform 1 0 25300 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1607194113
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1607194113
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1607194113
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1607194113
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1607194113
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__CLK
timestamp 1607194113
transform 1 0 26036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__D
timestamp 1607194113
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607194113
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1346_
timestamp 1607194113
transform 1 0 26496 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_6_295
timestamp 1607194113
transform 1 0 28244 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_301
timestamp 1607194113
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_293
timestamp 1607194113
transform 1 0 28060 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607194113
transform -1 0 29256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607194113
transform -1 0 29256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1607194113
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1607194113
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1607194113
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1607194113
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_301
timestamp 1607194113
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_293
timestamp 1607194113
transform 1 0 28060 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607194113
transform -1 0 29256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1607194113
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1607194113
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_264
timestamp 1607194113
transform 1 0 25392 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_252
timestamp 1607194113
transform 1 0 24288 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1607194113
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1607194113
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1607194113
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1607194113
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607194113
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_301
timestamp 1607194113
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_293
timestamp 1607194113
transform 1 0 28060 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_300
timestamp 1607194113
transform 1 0 28704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_288
timestamp 1607194113
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607194113
transform -1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607194113
transform -1 0 29256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_264
timestamp 1607194113
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1331_
timestamp 1607194113
transform 1 0 23644 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1607194113
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_272
timestamp 1607194113
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607194113
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_300
timestamp 1607194113
transform 1 0 28704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_288
timestamp 1607194113
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607194113
transform -1 0 29256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_255
timestamp 1607194113
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1607194113
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1607194113
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1607194113
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_267
timestamp 1607194113
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1607194113
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1607194113
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607194113
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_300
timestamp 1607194113
transform 1 0 28704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_288
timestamp 1607194113
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_301
timestamp 1607194113
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1607194113
transform 1 0 28060 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607194113
transform -1 0 29256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607194113
transform -1 0 29256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_256
timestamp 1607194113
transform 1 0 24656 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_245
timestamp 1607194113
transform 1 0 23644 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_i_A
timestamp 1607194113
transform 1 0 24196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk_i
timestamp 1607194113
transform 1 0 24380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_268
timestamp 1607194113
transform 1 0 25760 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__CLK
timestamp 1607194113
transform 1 0 26128 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1347_
timestamp 1607194113
transform 1 0 26312 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_301
timestamp 1607194113
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_293
timestamp 1607194113
transform 1 0 28060 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607194113
transform -1 0 29256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_263
timestamp 1607194113
transform 1 0 25300 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_257
timestamp 1607194113
transform 1 0 24748 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1607194113
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_262
timestamp 1607194113
transform 1 0 25208 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_250
timestamp 1607194113
transform 1 0 24104 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__CLK
timestamp 1607194113
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_270
timestamp 1607194113
transform 1 0 25944 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607194113
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1349_
timestamp 1607194113
transform 1 0 25576 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1348_
timestamp 1607194113
transform 1 0 26496 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_15_297
timestamp 1607194113
transform 1 0 28428 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_285
timestamp 1607194113
transform 1 0 27324 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_295
timestamp 1607194113
transform 1 0 28244 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607194113
transform -1 0 29256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607194113
transform -1 0 29256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_260
timestamp 1607194113
transform 1 0 25024 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_248
timestamp 1607194113
transform 1 0 23920 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__CLK
timestamp 1607194113
transform 1 0 23736 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1607194113
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_272
timestamp 1607194113
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607194113
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_300
timestamp 1607194113
transform 1 0 28704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_288
timestamp 1607194113
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607194113
transform -1 0 29256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1607194113
transform 1 0 24380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_257
timestamp 1607194113
transform 1 0 24748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_251
timestamp 1607194113
transform 1 0 24196 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_245
timestamp 1607194113
transform 1 0 23644 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__CLK
timestamp 1607194113
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk_i
timestamp 1607194113
transform 1 0 24472 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1449_
timestamp 1607194113
transform 1 0 24840 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1607194113
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1607194113
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1607194113
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_277
timestamp 1607194113
transform 1 0 26588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607194113
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_300
timestamp 1607194113
transform 1 0 28704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_288
timestamp 1607194113
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_301
timestamp 1607194113
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_289
timestamp 1607194113
transform 1 0 27692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607194113
transform -1 0 29256 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607194113
transform -1 0 29256 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_264
timestamp 1607194113
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_252
timestamp 1607194113
transform 1 0 24288 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__CLK
timestamp 1607194113
transform 1 0 24104 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__CLK
timestamp 1607194113
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1366_
timestamp 1607194113
transform 1 0 23644 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_272
timestamp 1607194113
transform 1 0 26128 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_266
timestamp 1607194113
transform 1 0 25576 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__CLK
timestamp 1607194113
transform 1 0 26312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__B1
timestamp 1607194113
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607194113
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1358_
timestamp 1607194113
transform 1 0 26496 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1305_
timestamp 1607194113
transform 1 0 26496 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_20_300
timestamp 1607194113
transform 1 0 28704 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_292
timestamp 1607194113
transform 1 0 27968 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_295
timestamp 1607194113
transform 1 0 28244 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607194113
transform -1 0 29256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607194113
transform -1 0 29256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_262
timestamp 1607194113
transform 1 0 25208 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_250
timestamp 1607194113
transform 1 0 24104 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A
timestamp 1607194113
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1281_
timestamp 1607194113
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_274
timestamp 1607194113
transform 1 0 26312 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_291
timestamp 1607194113
transform 1 0 27876 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_286
timestamp 1607194113
transform 1 0 27416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607194113
transform -1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1607194113
transform 1 0 27600 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_257
timestamp 1607194113
transform 1 0 24748 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1607194113
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_259
timestamp 1607194113
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_247
timestamp 1607194113
transform 1 0 23828 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__B1
timestamp 1607194113
transform 1 0 25300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1607194113
transform 1 0 26956 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_271
timestamp 1607194113
transform 1 0 26036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607194113
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1357_
timestamp 1607194113
transform 1 0 26496 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1307_
timestamp 1607194113
transform 1 0 25484 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_300
timestamp 1607194113
transform 1 0 28704 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_292
timestamp 1607194113
transform 1 0 27968 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_295
timestamp 1607194113
transform 1 0 28244 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607194113
transform -1 0 29256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607194113
transform -1 0 29256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1306_
timestamp 1607194113
transform 1 0 27692 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_262
timestamp 1607194113
transform 1 0 25208 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_254
timestamp 1607194113
transform 1 0 24472 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1607194113
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1159_
timestamp 1607194113
transform 1 0 24840 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_270
timestamp 1607194113
transform 1 0 25944 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607194113
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1408_
timestamp 1607194113
transform 1 0 26496 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_24_295
timestamp 1607194113
transform 1 0 28244 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607194113
transform -1 0 29256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_255
timestamp 1607194113
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_260
timestamp 1607194113
transform 1 0 25024 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_248
timestamp 1607194113
transform 1 0 23920 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1607194113
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1607194113
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_267
timestamp 1607194113
transform 1 0 25668 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_280
timestamp 1607194113
transform 1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 1607194113
transform 1 0 26128 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607194113
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1607194113
transform 1 0 27140 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_300
timestamp 1607194113
transform 1 0 28704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_288
timestamp 1607194113
transform 1 0 27600 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_300
timestamp 1607194113
transform 1 0 28704 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_288
timestamp 1607194113
transform 1 0 27600 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1607194113
transform 1 0 27416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607194113
transform -1 0 29256 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607194113
transform -1 0 29256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_261
timestamp 1607194113
transform 1 0 25116 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_257
timestamp 1607194113
transform 1 0 24748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1607194113
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B1
timestamp 1607194113
transform 1 0 25208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1222_
timestamp 1607194113
transform 1 0 25392 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_280
timestamp 1607194113
transform 1 0 26864 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_300
timestamp 1607194113
transform 1 0 28704 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_292
timestamp 1607194113
transform 1 0 27968 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607194113
transform -1 0 29256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_257
timestamp 1607194113
transform 1 0 24748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1607194113
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_247
timestamp 1607194113
transform 1 0 23828 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__B2
timestamp 1607194113
transform 1 0 23920 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A2
timestamp 1607194113
transform 1 0 24104 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B1
timestamp 1607194113
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1223_
timestamp 1607194113
transform 1 0 25116 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0953_
timestamp 1607194113
transform 1 0 24288 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_29_277
timestamp 1607194113
transform 1 0 26588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_272
timestamp 1607194113
transform 1 0 26128 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_266
timestamp 1607194113
transform 1 0 25576 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607194113
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1407_
timestamp 1607194113
transform 1 0 26496 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_29_302
timestamp 1607194113
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_290
timestamp 1607194113
transform 1 0 27784 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_295
timestamp 1607194113
transform 1 0 28244 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1607194113
transform 1 0 27600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607194113
transform -1 0 29256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607194113
transform -1 0 29256 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1607194113
transform 1 0 27324 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A2
timestamp 1607194113
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B2
timestamp 1607194113
transform 1 0 24012 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0965_
timestamp 1607194113
transform 1 0 24196 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1607194113
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_273
timestamp 1607194113
transform 1 0 26220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1607194113
transform 1 0 25484 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607194113
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_300
timestamp 1607194113
transform 1 0 28704 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_288
timestamp 1607194113
transform 1 0 27600 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607194113
transform -1 0 29256 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_247
timestamp 1607194113
transform 1 0 23828 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_257
timestamp 1607194113
transform 1 0 24748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1607194113
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B1
timestamp 1607194113
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B1
timestamp 1607194113
transform 1 0 24012 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1209_
timestamp 1607194113
transform 1 0 24196 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1208_
timestamp 1607194113
transform 1 0 25024 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1607194113
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A2_N
timestamp 1607194113
transform 1 0 25852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B2
timestamp 1607194113
transform 1 0 25668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_282
timestamp 1607194113
transform 1 0 27048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1607194113
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1607194113
transform 1 0 26864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A2_N
timestamp 1607194113
transform 1 0 26680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B2
timestamp 1607194113
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607194113
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1607194113
transform 1 0 26588 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_280
timestamp 1607194113
transform 1 0 26864 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_291
timestamp 1607194113
transform 1 0 27876 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_300
timestamp 1607194113
transform 1 0 28704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_292
timestamp 1607194113
transform 1 0 27968 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1607194113
transform 1 0 27416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607194113
transform -1 0 29256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607194113
transform -1 0 29256 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1607194113
transform 1 0 27600 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_257
timestamp 1607194113
transform 1 0 24748 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1607194113
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_265
timestamp 1607194113
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__CLK
timestamp 1607194113
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1416_
timestamp 1607194113
transform 1 0 25852 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_33_300
timestamp 1607194113
transform 1 0 28704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_288
timestamp 1607194113
transform 1 0 27600 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607194113
transform -1 0 29256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_262
timestamp 1607194113
transform 1 0 25208 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_250
timestamp 1607194113
transform 1 0 24104 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_264
timestamp 1607194113
transform 1 0 25392 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_252
timestamp 1607194113
transform 1 0 24288 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__CLK
timestamp 1607194113
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1607194113
transform 1 0 23920 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1607194113
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_274
timestamp 1607194113
transform 1 0 26312 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_272
timestamp 1607194113
transform 1 0 26128 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607194113
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1417_
timestamp 1607194113
transform 1 0 26496 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_35_302
timestamp 1607194113
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_298
timestamp 1607194113
transform 1 0 28520 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1607194113
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_295
timestamp 1607194113
transform 1 0 28244 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607194113
transform -1 0 29256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607194113
transform -1 0 29256 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1607194113
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1607194113
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_255
timestamp 1607194113
transform 1 0 24564 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_273
timestamp 1607194113
transform 1 0 26220 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_269
timestamp 1607194113
transform 1 0 25852 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1607194113
transform 1 0 26496 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_267
timestamp 1607194113
transform 1 0 25668 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__CLK
timestamp 1607194113
transform 1 0 26312 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607194113
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1356_
timestamp 1607194113
transform 1 0 26496 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_37_295
timestamp 1607194113
transform 1 0 28244 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_291
timestamp 1607194113
transform 1 0 27876 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607194113
transform -1 0 29256 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607194113
transform -1 0 29256 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1607194113
transform 1 0 27600 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_246
timestamp 1607194113
transform 1 0 23736 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__B1
timestamp 1607194113
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1313_
timestamp 1607194113
transform 1 0 24104 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_38_272
timestamp 1607194113
transform 1 0 26128 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_266
timestamp 1607194113
transform 1 0 25576 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__B1
timestamp 1607194113
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607194113
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1311_
timestamp 1607194113
transform 1 0 26496 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_38_300
timestamp 1607194113
transform 1 0 28704 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_292
timestamp 1607194113
transform 1 0 27968 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607194113
transform -1 0 29256 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_252
timestamp 1607194113
transform 1 0 24288 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_245
timestamp 1607194113
transform 1 0 23644 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__CLK
timestamp 1607194113
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1607194113
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1355_
timestamp 1607194113
transform 1 0 24656 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1309_
timestamp 1607194113
transform 1 0 23736 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_275
timestamp 1607194113
transform 1 0 26404 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1607194113
transform 1 0 26956 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 27140 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607194113
transform -1 0 29256 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_257
timestamp 1607194113
transform 1 0 24748 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_284
timestamp 1607194113
transform 1 0 27232 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1607194113
transform 1 0 26864 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_269
timestamp 1607194113
transform 1 0 25852 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607194113
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1312_
timestamp 1607194113
transform 1 0 27324 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1310_
timestamp 1607194113
transform 1 0 26496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_296
timestamp 1607194113
transform 1 0 28336 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_288
timestamp 1607194113
transform 1 0 27600 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_i_A
timestamp 1607194113
transform 1 0 28520 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk_i
timestamp 1607194113
transform 1 0 28704 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607194113
transform -1 0 29256 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_247
timestamp 1607194113
transform 1 0 23828 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1607194113
transform 1 0 23644 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__B1
timestamp 1607194113
transform 1 0 24012 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1354_
timestamp 1607194113
transform 1 0 23828 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1318_
timestamp 1607194113
transform 1 0 24196 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_276
timestamp 1607194113
transform 1 0 26496 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_267
timestamp 1607194113
transform 1 0 25668 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_277
timestamp 1607194113
transform 1 0 26588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_266
timestamp 1607194113
transform 1 0 25576 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607194113
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1607194113
transform 1 0 26312 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_300
timestamp 1607194113
transform 1 0 28704 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_288
timestamp 1607194113
transform 1 0 27600 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_301
timestamp 1607194113
transform 1 0 28796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_289
timestamp 1607194113
transform 1 0 27692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607194113
transform -1 0 29256 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607194113
transform -1 0 29256 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_264
timestamp 1607194113
transform 1 0 25392 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_245
timestamp 1607194113
transform 1 0 23644 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__B1
timestamp 1607194113
transform 1 0 23736 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1320_
timestamp 1607194113
transform 1 0 23920 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_43_270
timestamp 1607194113
transform 1 0 25944 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__CLK
timestamp 1607194113
transform 1 0 26036 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1353_
timestamp 1607194113
transform 1 0 26220 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_43_300
timestamp 1607194113
transform 1 0 28704 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_292
timestamp 1607194113
transform 1 0 27968 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607194113
transform -1 0 29256 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_261
timestamp 1607194113
transform 1 0 25116 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_249
timestamp 1607194113
transform 1 0 24012 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1319_
timestamp 1607194113
transform 1 0 25392 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1607194113
transform 1 0 23736 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_281
timestamp 1607194113
transform 1 0 26956 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_276
timestamp 1607194113
transform 1 0 26496 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_267
timestamp 1607194113
transform 1 0 25668 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607194113
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1317_
timestamp 1607194113
transform 1 0 26680 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_301
timestamp 1607194113
transform 1 0 28796 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_293
timestamp 1607194113
transform 1 0 28060 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1607194113
transform -1 0 29256 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_257
timestamp 1607194113
transform 1 0 24748 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1607194113
transform 1 0 23644 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__CLK
timestamp 1607194113
transform 1 0 24840 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1352_
timestamp 1607194113
transform 1 0 25024 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_45_279
timestamp 1607194113
transform 1 0 26772 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_291
timestamp 1607194113
transform 1 0 27876 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1607194113
transform -1 0 29256 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1607194113
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_246
timestamp 1607194113
transform 1 0 23736 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_270
timestamp 1607194113
transform 1 0 25944 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__B1
timestamp 1607194113
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607194113
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1322_
timestamp 1607194113
transform 1 0 26496 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_46_300
timestamp 1607194113
transform 1 0 28704 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_292
timestamp 1607194113
transform 1 0 27968 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1607194113
transform -1 0 29256 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_263
timestamp 1607194113
transform 1 0 25300 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_251
timestamp 1607194113
transform 1 0 24196 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_249
timestamp 1607194113
transform 1 0 24012 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1607194113
transform 1 0 23644 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__B1
timestamp 1607194113
transform 1 0 24104 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1324_
timestamp 1607194113
transform 1 0 24288 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1323_
timestamp 1607194113
transform 1 0 25392 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_284
timestamp 1607194113
transform 1 0 27232 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_276
timestamp 1607194113
transform 1 0 26496 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_267
timestamp 1607194113
transform 1 0 25668 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_268
timestamp 1607194113
transform 1 0 25760 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607194113
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1351_
timestamp 1607194113
transform 1 0 26496 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1321_
timestamp 1607194113
transform 1 0 27324 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_300
timestamp 1607194113
transform 1 0 28704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_288
timestamp 1607194113
transform 1 0 27600 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_297
timestamp 1607194113
transform 1 0 28428 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__CLK
timestamp 1607194113
transform 1 0 28244 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1607194113
transform -1 0 29256 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1607194113
transform -1 0 29256 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_255
timestamp 1607194113
transform 1 0 24564 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_249
timestamp 1607194113
transform 1 0 24012 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_245
timestamp 1607194113
transform 1 0 23644 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1607194113
transform 1 0 24380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1350_
timestamp 1607194113
transform 1 0 25116 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1607194113
transform 1 0 24104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_282
timestamp 1607194113
transform 1 0 27048 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__CLK
timestamp 1607194113
transform 1 0 26864 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_302
timestamp 1607194113
transform 1 0 28888 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_294
timestamp 1607194113
transform 1 0 28152 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1607194113
transform -1 0 29256 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_260
timestamp 1607194113
transform 1 0 25024 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_276
timestamp 1607194113
transform 1 0 26496 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_272
timestamp 1607194113
transform 1 0 26128 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607194113
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_300
timestamp 1607194113
transform 1 0 28704 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_288
timestamp 1607194113
transform 1 0 27600 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1607194113
transform -1 0 29256 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1607194113
transform 1 0 25484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1_N
timestamp 1607194113
transform 1 0 25300 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B1
timestamp 1607194113
transform 1 0 23644 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1274_
timestamp 1607194113
transform 1 0 23828 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_277
timestamp 1607194113
transform 1 0 26588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_301
timestamp 1607194113
transform 1 0 28796 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_289
timestamp 1607194113
transform 1 0 27692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1607194113
transform -1 0 29256 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_247
timestamp 1607194113
transform 1 0 23828 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1415_
timestamp 1607194113
transform 1 0 23920 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_52_269
timestamp 1607194113
transform 1 0 25852 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__CLK
timestamp 1607194113
transform 1 0 25668 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607194113
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1374_
timestamp 1607194113
transform 1 0 26496 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_52_297
timestamp 1607194113
transform 1 0 28428 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__CLK
timestamp 1607194113
transform 1 0 28244 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1607194113
transform -1 0 29256 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_262
timestamp 1607194113
transform 1 0 25208 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_250
timestamp 1607194113
transform 1 0 24104 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A
timestamp 1607194113
transform 1 0 23644 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1607194113
transform 1 0 23828 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B1
timestamp 1607194113
transform 1 0 25760 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1273_
timestamp 1607194113
transform 1 0 25944 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_53_300
timestamp 1607194113
transform 1 0 28704 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_288
timestamp 1607194113
transform 1 0 27600 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A1_N
timestamp 1607194113
transform 1 0 27416 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1607194113
transform -1 0 29256 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_263
timestamp 1607194113
transform 1 0 25300 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_245
timestamp 1607194113
transform 1 0 23644 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_264
timestamp 1607194113
transform 1 0 25392 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_254
timestamp 1607194113
transform 1 0 24472 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A
timestamp 1607194113
transform 1 0 24840 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A
timestamp 1607194113
transform 1 0 24748 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1607194113
transform 1 0 25024 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1206_
timestamp 1607194113
transform 1 0 24932 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_274
timestamp 1607194113
transform 1 0 26312 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_284
timestamp 1607194113
transform 1 0 27232 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_276
timestamp 1607194113
transform 1 0 26496 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_272
timestamp 1607194113
transform 1 0 26128 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607194113
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1607194113
transform 1 0 26036 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_302
timestamp 1607194113
transform 1 0 28888 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_298
timestamp 1607194113
transform 1 0 28520 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1607194113
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_300
timestamp 1607194113
transform 1 0 28704 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_292
timestamp 1607194113
transform 1 0 27968 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1607194113
transform 1 0 27784 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1607194113
transform -1 0 29256 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1607194113
transform -1 0 29256 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1607194113
transform 1 0 27508 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_249
timestamp 1607194113
transform 1 0 24012 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0854_
timestamp 1607194113
transform 1 0 24196 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_276
timestamp 1607194113
transform 1 0 26496 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_273
timestamp 1607194113
transform 1 0 26220 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2_N
timestamp 1607194113
transform 1 0 26036 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B1
timestamp 1607194113
transform 1 0 25852 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B2
timestamp 1607194113
transform 1 0 25668 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607194113
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_300
timestamp 1607194113
transform 1 0 28704 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_288
timestamp 1607194113
transform 1 0 27600 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1607194113
transform -1 0 29256 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_253
timestamp 1607194113
transform 1 0 24380 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_245
timestamp 1607194113
transform 1 0 23644 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A1_N
timestamp 1607194113
transform 1 0 24472 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0783_
timestamp 1607194113
transform 1 0 24656 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_276
timestamp 1607194113
transform 1 0 26496 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A2_N
timestamp 1607194113
transform 1 0 26312 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B2
timestamp 1607194113
transform 1 0 26128 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_300
timestamp 1607194113
transform 1 0 28704 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_288
timestamp 1607194113
transform 1 0 27600 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1607194113
transform -1 0 29256 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_257
timestamp 1607194113
transform 1 0 24748 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_245
timestamp 1607194113
transform 1 0 23644 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_269
timestamp 1607194113
transform 1 0 25852 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607194113
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1418_
timestamp 1607194113
transform 1 0 26496 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_58_297
timestamp 1607194113
transform 1 0 28428 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__CLK
timestamp 1607194113
transform 1 0 28244 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1607194113
transform -1 0 29256 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_257
timestamp 1607194113
transform 1 0 24748 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_245
timestamp 1607194113
transform 1 0 23644 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B2
timestamp 1607194113
transform 1 0 25024 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A2_N
timestamp 1607194113
transform 1 0 25208 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B1
timestamp 1607194113
transform 1 0 25392 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_284
timestamp 1607194113
transform 1 0 27232 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A1_N
timestamp 1607194113
transform 1 0 27048 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1207_
timestamp 1607194113
transform 1 0 25576 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_59_304
timestamp 1607194113
transform 1 0 29072 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_296
timestamp 1607194113
transform 1 0 28336 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607194113
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1377_
timestamp 1607194113
transform 1 0 29256 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_327
timestamp 1607194113
transform 1 0 31188 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__CLK
timestamp 1607194113
transform 1 0 31004 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_339
timestamp 1607194113
transform 1 0 32292 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1607194113
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_363
timestamp 1607194113
transform 1 0 34500 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_351
timestamp 1607194113
transform 1 0 33396 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607194113
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1607194113
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_391
timestamp 1607194113
transform 1 0 37076 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A1_N
timestamp 1607194113
transform 1 0 37812 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1607194113
transform 1 0 37996 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0740_
timestamp 1607194113
transform 1 0 38180 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_428
timestamp 1607194113
transform 1 0 40480 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_423
timestamp 1607194113
transform 1 0 40020 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B2
timestamp 1607194113
transform 1 0 39836 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A2_N
timestamp 1607194113
transform 1 0 39652 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607194113
transform 1 0 40388 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_444
timestamp 1607194113
transform 1 0 41952 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_440
timestamp 1607194113
transform 1 0 41584 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A1_N
timestamp 1607194113
transform 1 0 42044 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B1
timestamp 1607194113
transform 1 0 42228 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0727_
timestamp 1607194113
transform 1 0 42412 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_469
timestamp 1607194113
transform 1 0 44252 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A2_N
timestamp 1607194113
transform 1 0 44068 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B2
timestamp 1607194113
transform 1 0 43884 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_487
timestamp 1607194113
transform 1 0 45908 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_481
timestamp 1607194113
transform 1 0 45356 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607194113
transform 1 0 46000 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_260
timestamp 1607194113
transform 1 0 25024 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_248
timestamp 1607194113
transform 1 0 23920 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1607194113
transform 1 0 23644 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_274
timestamp 1607194113
transform 1 0 26312 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_268
timestamp 1607194113
transform 1 0 25760 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A2_N
timestamp 1607194113
transform 1 0 26128 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__B1
timestamp 1607194113
transform 1 0 25944 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607194113
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1270_
timestamp 1607194113
transform 1 0 26496 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_304
timestamp 1607194113
transform 1 0 29072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_300
timestamp 1607194113
transform 1 0 28704 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_294
timestamp 1607194113
transform 1 0 28152 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A1_N
timestamp 1607194113
transform 1 0 27968 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1607194113
transform 1 0 28796 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1607194113
transform 1 0 30636 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_316
timestamp 1607194113
transform 1 0 30176 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1607194113
transform 1 0 30360 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_345
timestamp 1607194113
transform 1 0 32844 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_337
timestamp 1607194113
transform 1 0 32108 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_333
timestamp 1607194113
transform 1 0 31740 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__CLK
timestamp 1607194113
transform 1 0 32936 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607194113
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1425_
timestamp 1607194113
transform 1 0 33120 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_60_367
timestamp 1607194113
transform 1 0 34868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_379
timestamp 1607194113
transform 1 0 35972 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_398
timestamp 1607194113
transform 1 0 37720 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_391
timestamp 1607194113
transform 1 0 37076 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1607194113
transform 1 0 38088 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1_N
timestamp 1607194113
transform 1 0 38272 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607194113
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0759_
timestamp 1607194113
transform 1 0 38456 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B2
timestamp 1607194113
transform 1 0 40112 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2_N
timestamp 1607194113
transform 1 0 39928 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B1
timestamp 1607194113
transform 1 0 40296 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A1_N
timestamp 1607194113
transform 1 0 40480 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0732_
timestamp 1607194113
transform 1 0 40664 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_450
timestamp 1607194113
transform 1 0 42504 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B2
timestamp 1607194113
transform 1 0 42320 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A2_N
timestamp 1607194113
transform 1 0 42136 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_471
timestamp 1607194113
transform 1 0 44436 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_459
timestamp 1607194113
transform 1 0 43332 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607194113
transform 1 0 43240 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_483
timestamp 1607194113
transform 1 0 45540 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_257
timestamp 1607194113
transform 1 0 24748 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1607194113
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_263
timestamp 1607194113
transform 1 0 25300 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_257
timestamp 1607194113
transform 1 0 24748 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_245
timestamp 1607194113
transform 1 0 23644 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1607194113
transform 1 0 25024 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__B1
timestamp 1607194113
transform 1 0 25392 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1262_
timestamp 1607194113
transform 1 0 25208 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_270
timestamp 1607194113
transform 1 0 25944 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_266
timestamp 1607194113
transform 1 0 25576 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_284
timestamp 1607194113
transform 1 0 27232 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B2
timestamp 1607194113
transform 1 0 26036 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A2
timestamp 1607194113
transform 1 0 26220 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1_N
timestamp 1607194113
transform 1 0 27048 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607194113
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1197_
timestamp 1607194113
transform 1 0 25576 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0925_
timestamp 1607194113
transform 1 0 26496 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_62_302
timestamp 1607194113
transform 1 0 28888 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_290
timestamp 1607194113
transform 1 0 27784 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_300
timestamp 1607194113
transform 1 0 28704 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_296
timestamp 1607194113
transform 1 0 28336 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A1_N
timestamp 1607194113
transform 1 0 28796 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B1
timestamp 1607194113
transform 1 0 28980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607194113
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0701_
timestamp 1607194113
transform 1 0 29256 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_316
timestamp 1607194113
transform 1 0 30176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_310
timestamp 1607194113
transform 1 0 29624 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A1_N
timestamp 1607194113
transform 1 0 31096 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A2_N
timestamp 1607194113
transform 1 0 30912 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B2
timestamp 1607194113
transform 1 0 30728 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk_i
timestamp 1607194113
transform 1 0 29900 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_328
timestamp 1607194113
transform 1 0 31280 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__CLK
timestamp 1607194113
transform 1 0 31832 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B1
timestamp 1607194113
transform 1 0 31280 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A2_N
timestamp 1607194113
transform 1 0 33120 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B2
timestamp 1607194113
transform 1 0 32936 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607194113
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1384_
timestamp 1607194113
transform 1 0 32108 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _0799_
timestamp 1607194113
transform 1 0 31464 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_62_356
timestamp 1607194113
transform 1 0 33856 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A2_N
timestamp 1607194113
transform 1 0 34040 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B2
timestamp 1607194113
transform 1 0 34224 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B2
timestamp 1607194113
transform 1 0 34408 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A2
timestamp 1607194113
transform 1 0 34592 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B1
timestamp 1607194113
transform 1 0 34408 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607194113
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_350
timestamp 1607194113
transform 1 0 33304 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1205_
timestamp 1607194113
transform 1 0 34592 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0935_
timestamp 1607194113
transform 1 0 34868 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_380
timestamp 1607194113
transform 1 0 36064 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_381
timestamp 1607194113
transform 1 0 36156 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_410
timestamp 1607194113
transform 1 0 38824 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_398
timestamp 1607194113
transform 1 0 37720 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_396
timestamp 1607194113
transform 1 0 37536 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_392
timestamp 1607194113
transform 1 0 37168 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_393
timestamp 1607194113
transform 1 0 37260 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1607194113
transform 1 0 37812 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1_N
timestamp 1607194113
transform 1 0 37996 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607194113
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0760_
timestamp 1607194113
transform 1 0 38180 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_62_416
timestamp 1607194113
transform 1 0 39376 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2_N
timestamp 1607194113
transform 1 0 39836 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B2
timestamp 1607194113
transform 1 0 39744 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1607194113
transform 1 0 39652 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1607194113
transform 1 0 39468 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_422
timestamp 1607194113
transform 1 0 39928 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_426
timestamp 1607194113
transform 1 0 40296 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_423
timestamp 1607194113
transform 1 0 40020 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A1_N
timestamp 1607194113
transform 1 0 40112 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B1
timestamp 1607194113
transform 1 0 40296 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607194113
transform 1 0 40388 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0758_
timestamp 1607194113
transform 1 0 40480 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0736_
timestamp 1607194113
transform 1 0 40480 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_448
timestamp 1607194113
transform 1 0 42320 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_448
timestamp 1607194113
transform 1 0 42320 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B2
timestamp 1607194113
transform 1 0 42136 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A2_N
timestamp 1607194113
transform 1 0 42136 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2_N
timestamp 1607194113
transform 1 0 41952 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B2
timestamp 1607194113
transform 1 0 41952 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0741_
timestamp 1607194113
transform 1 0 42688 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1607194113
transform 1 0 44620 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1607194113
transform 1 0 43516 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B1
timestamp 1607194113
transform 1 0 43056 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607194113
transform 1 0 43240 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0836_
timestamp 1607194113
transform 1 0 43332 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_62_483
timestamp 1607194113
transform 1 0 45540 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_479
timestamp 1607194113
transform 1 0 45172 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_485
timestamp 1607194113
transform 1 0 45724 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B2
timestamp 1607194113
transform 1 0 45632 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A2
timestamp 1607194113
transform 1 0 45816 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A2_N
timestamp 1607194113
transform 1 0 44988 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B2
timestamp 1607194113
transform 1 0 44804 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607194113
transform 1 0 46000 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0931_
timestamp 1607194113
transform 1 0 46000 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_63_257
timestamp 1607194113
transform 1 0 24748 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1607194113
transform 1 0 23644 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B1
timestamp 1607194113
transform 1 0 25116 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1260_
timestamp 1607194113
transform 1 0 25300 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1607194113
transform 1 0 26956 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A1_N
timestamp 1607194113
transform 1 0 26772 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1607194113
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1607194113
transform 1 0 28060 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607194113
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1607194113
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_342
timestamp 1607194113
transform 1 0 32568 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_330
timestamp 1607194113
transform 1 0 31464 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_365
timestamp 1607194113
transform 1 0 34684 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_360
timestamp 1607194113
transform 1 0 34224 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_354
timestamp 1607194113
transform 1 0 33672 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A2_N
timestamp 1607194113
transform 1 0 34316 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B2
timestamp 1607194113
transform 1 0 34500 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607194113
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1268_
timestamp 1607194113
transform 1 0 34868 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_383
timestamp 1607194113
transform 1 0 36340 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_407
timestamp 1607194113
transform 1 0 38548 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_395
timestamp 1607194113
transform 1 0 37444 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_428
timestamp 1607194113
transform 1 0 40480 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_419
timestamp 1607194113
transform 1 0 39652 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607194113
transform 1 0 40388 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_452
timestamp 1607194113
transform 1 0 42688 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_441
timestamp 1607194113
transform 1 0 41676 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1607194113
transform 1 0 42412 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0764_
timestamp 1607194113
transform 1 0 40848 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_63_464
timestamp 1607194113
transform 1 0 43792 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0841_
timestamp 1607194113
transform 1 0 44160 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_487
timestamp 1607194113
transform 1 0 45908 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_477
timestamp 1607194113
transform 1 0 44988 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A2_N
timestamp 1607194113
transform 1 0 45540 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B2
timestamp 1607194113
transform 1 0 45724 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607194113
transform 1 0 46000 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_257
timestamp 1607194113
transform 1 0 24748 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_245
timestamp 1607194113
transform 1 0 23644 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1607194113
transform 1 0 25024 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1199_
timestamp 1607194113
transform 1 0 25208 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_274
timestamp 1607194113
transform 1 0 26312 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_266
timestamp 1607194113
transform 1 0 25576 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B2
timestamp 1607194113
transform 1 0 26128 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B1
timestamp 1607194113
transform 1 0 25944 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1607194113
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1200_
timestamp 1607194113
transform 1 0 26496 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_304
timestamp 1607194113
transform 1 0 29072 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_292
timestamp 1607194113
transform 1 0 27968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_321
timestamp 1607194113
transform 1 0 30636 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__C
timestamp 1607194113
transform 1 0 29624 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0720_
timestamp 1607194113
transform 1 0 29808 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1607194113
transform 1 0 32108 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1607194113
transform 1 0 31924 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_329
timestamp 1607194113
transform 1 0 31372 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_i_A
timestamp 1607194113
transform 1 0 31740 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk_i
timestamp 1607194113
transform 1 0 31464 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1607194113
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_367
timestamp 1607194113
transform 1 0 34868 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_361
timestamp 1607194113
transform 1 0 34316 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1607194113
transform 1 0 33212 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__CLK
timestamp 1607194113
transform 1 0 34960 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B1
timestamp 1607194113
transform 1 0 34684 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_389
timestamp 1607194113
transform 1 0 36892 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1419_
timestamp 1607194113
transform 1 0 35144 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_410
timestamp 1607194113
transform 1 0 38824 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_398
timestamp 1607194113
transform 1 0 37720 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1607194113
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_422
timestamp 1607194113
transform 1 0 39928 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A1_N
timestamp 1607194113
transform 1 0 40020 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B1
timestamp 1607194113
transform 1 0 40204 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0763_
timestamp 1607194113
transform 1 0 40388 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1607194113
transform 1 0 42044 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A2_N
timestamp 1607194113
transform 1 0 41860 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_471
timestamp 1607194113
transform 1 0 44436 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_459
timestamp 1607194113
transform 1 0 43332 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_457
timestamp 1607194113
transform 1 0 43148 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1607194113
transform 1 0 43240 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_483
timestamp 1607194113
transform 1 0 45540 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B1
timestamp 1607194113
transform 1 0 45908 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_263
timestamp 1607194113
transform 1 0 25300 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_257
timestamp 1607194113
transform 1 0 24748 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_245
timestamp 1607194113
transform 1 0 23644 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B2
timestamp 1607194113
transform 1 0 25392 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_284
timestamp 1607194113
transform 1 0 27232 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B1
timestamp 1607194113
transform 1 0 25576 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1263_
timestamp 1607194113
transform 1 0 25760 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_65_304
timestamp 1607194113
transform 1 0 29072 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_296
timestamp 1607194113
transform 1 0 28336 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1607194113
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1382_
timestamp 1607194113
transform 1 0 29256 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_65_327
timestamp 1607194113
transform 1 0 31188 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__CLK
timestamp 1607194113
transform 1 0 31004 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_342
timestamp 1607194113
transform 1 0 32568 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__C
timestamp 1607194113
transform 1 0 31556 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0815_
timestamp 1607194113
transform 1 0 31740 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_65_367
timestamp 1607194113
transform 1 0 34868 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_354
timestamp 1607194113
transform 1 0 33672 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1607194113
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_371
timestamp 1607194113
transform 1 0 35236 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__CLK
timestamp 1607194113
transform 1 0 35328 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1378_
timestamp 1607194113
transform 1 0 35512 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_404
timestamp 1607194113
transform 1 0 38272 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_393
timestamp 1607194113
transform 1 0 37260 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1607194113
transform 1 0 37996 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_428
timestamp 1607194113
transform 1 0 40480 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_424
timestamp 1607194113
transform 1 0 40112 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_416
timestamp 1607194113
transform 1 0 39376 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1607194113
transform 1 0 40388 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_436
timestamp 1607194113
transform 1 0 41216 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1_N
timestamp 1607194113
transform 1 0 41400 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B1
timestamp 1607194113
transform 1 0 41584 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0840_
timestamp 1607194113
transform 1 0 41768 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_472
timestamp 1607194113
transform 1 0 44528 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_460
timestamp 1607194113
transform 1 0 43424 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A2_N
timestamp 1607194113
transform 1 0 43240 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_484
timestamp 1607194113
transform 1 0 45632 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A2_N
timestamp 1607194113
transform 1 0 45816 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1607194113
transform 1 0 46000 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_265
timestamp 1607194113
transform 1 0 25484 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A2_N
timestamp 1607194113
transform 1 0 25300 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B2
timestamp 1607194113
transform 1 0 25116 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0851_
timestamp 1607194113
transform 1 0 23644 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_276
timestamp 1607194113
transform 1 0 26496 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_273
timestamp 1607194113
transform 1 0 26220 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1607194113
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_288
timestamp 1607194113
transform 1 0 27600 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__CLK
timestamp 1607194113
transform 1 0 27876 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1423_
timestamp 1607194113
transform 1 0 28060 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_324
timestamp 1607194113
transform 1 0 30912 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_320
timestamp 1607194113
transform 1 0 30544 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_312
timestamp 1607194113
transform 1 0 29808 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1607194113
transform 1 0 30636 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_345
timestamp 1607194113
transform 1 0 32844 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_337
timestamp 1607194113
transform 1 0 32108 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk_i
timestamp 1607194113
transform 1 0 33028 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1607194113
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_362
timestamp 1607194113
transform 1 0 34408 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_350
timestamp 1607194113
transform 1 0 33304 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_388
timestamp 1607194113
transform 1 0 36800 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_382
timestamp 1607194113
transform 1 0 36248 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_374
timestamp 1607194113
transform 1 0 35512 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1607194113
transform 1 0 36524 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_396
timestamp 1607194113
transform 1 0 37536 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1607194113
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0828_
timestamp 1607194113
transform 1 0 37720 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_418
timestamp 1607194113
transform 1 0 39560 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__D
timestamp 1607194113
transform 1 0 40664 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B2
timestamp 1607194113
transform 1 0 39376 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A2_N
timestamp 1607194113
transform 1 0 39192 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_441
timestamp 1607194113
transform 1 0 41676 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0786_
timestamp 1607194113
transform 1 0 40848 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_471
timestamp 1607194113
transform 1 0 44436 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_459
timestamp 1607194113
transform 1 0 43332 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_457
timestamp 1607194113
transform 1 0 43148 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_453
timestamp 1607194113
transform 1 0 42780 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1607194113
transform 1 0 43240 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_483
timestamp 1607194113
transform 1 0 45540 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_261
timestamp 1607194113
transform 1 0 25116 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_265
timestamp 1607194113
transform 1 0 25484 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A2_N
timestamp 1607194113
transform 1 0 25300 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2_N
timestamp 1607194113
transform 1 0 24932 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B2
timestamp 1607194113
transform 1 0 24748 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B2
timestamp 1607194113
transform 1 0 25116 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0777_
timestamp 1607194113
transform 1 0 23644 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_285
timestamp 1607194113
transform 1 0 27324 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_273
timestamp 1607194113
transform 1 0 26220 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_278
timestamp 1607194113
transform 1 0 26680 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1607194113
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0856_
timestamp 1607194113
transform 1 0 26496 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0785_
timestamp 1607194113
transform 1 0 25852 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_68_297
timestamp 1607194113
transform 1 0 28428 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_306
timestamp 1607194113
transform 1 0 29256 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_302
timestamp 1607194113
transform 1 0 28888 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_290
timestamp 1607194113
transform 1 0 27784 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1607194113
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_309
timestamp 1607194113
transform 1 0 29532 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_325
timestamp 1607194113
transform 1 0 31004 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_313
timestamp 1607194113
transform 1 0 29900 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A2_N
timestamp 1607194113
transform 1 0 31096 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0698_
timestamp 1607194113
transform 1 0 29624 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1607194113
transform 1 0 29624 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1607194113
transform 1 0 32108 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_330
timestamp 1607194113
transform 1 0 31464 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1607194113
transform 1 0 32108 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B2
timestamp 1607194113
transform 1 0 31280 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1607194113
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_365
timestamp 1607194113
transform 1 0 34684 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_361
timestamp 1607194113
transform 1 0 34316 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_365
timestamp 1607194113
transform 1 0 34684 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_361
timestamp 1607194113
transform 1 0 34316 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B1
timestamp 1607194113
transform 1 0 34776 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A1_N
timestamp 1607194113
transform 1 0 34960 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1607194113
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_349
timestamp 1607194113
transform 1 0 33212 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1607194113
transform 1 0 34868 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1607194113
transform 1 0 33212 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_390
timestamp 1607194113
transform 1 0 36984 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_383
timestamp 1607194113
transform 1 0 36340 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_379
timestamp 1607194113
transform 1 0 35972 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A2_N
timestamp 1607194113
transform 1 0 36800 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B2
timestamp 1607194113
transform 1 0 36616 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0845_
timestamp 1607194113
transform 1 0 35144 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0746_
timestamp 1607194113
transform 1 0 36432 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_410
timestamp 1607194113
transform 1 0 38824 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_398
timestamp 1607194113
transform 1 0 37720 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_396
timestamp 1607194113
transform 1 0 37536 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_404
timestamp 1607194113
transform 1 0 38272 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B2
timestamp 1607194113
transform 1 0 38088 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2_N
timestamp 1607194113
transform 1 0 37904 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1607194113
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_430
timestamp 1607194113
transform 1 0 40664 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_422
timestamp 1607194113
transform 1 0 39928 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_428
timestamp 1607194113
transform 1 0 40480 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_67_424
timestamp 1607194113
transform 1 0 40112 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_416
timestamp 1607194113
transform 1 0 39376 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1607194113
transform 1 0 40388 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_434
timestamp 1607194113
transform 1 0 41032 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A2_N
timestamp 1607194113
transform 1 0 42688 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A1_N
timestamp 1607194113
transform 1 0 42504 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B1
timestamp 1607194113
transform 1 0 40848 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A1_N
timestamp 1607194113
transform 1 0 41124 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B1
timestamp 1607194113
transform 1 0 41308 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0834_
timestamp 1607194113
transform 1 0 41032 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0755_
timestamp 1607194113
transform 1 0 41492 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_67_459
timestamp 1607194113
transform 1 0 43332 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B2
timestamp 1607194113
transform 1 0 43148 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B2
timestamp 1607194113
transform 1 0 42872 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A2_N
timestamp 1607194113
transform 1 0 42964 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__D
timestamp 1607194113
transform 1 0 43516 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B1
timestamp 1607194113
transform 1 0 43056 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1607194113
transform 1 0 43240 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0857_
timestamp 1607194113
transform 1 0 43700 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_67_472
timestamp 1607194113
transform 1 0 44528 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _0830_
timestamp 1607194113
transform 1 0 43332 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_479
timestamp 1607194113
transform 1 0 45172 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_484
timestamp 1607194113
transform 1 0 45632 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A2_N
timestamp 1607194113
transform 1 0 44988 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B2
timestamp 1607194113
transform 1 0 44804 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1607194113
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B2
timestamp 1607194113
transform 1 0 25300 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1607194113
transform 1 0 25484 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A2_N
timestamp 1607194113
transform 1 0 25116 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0780_
timestamp 1607194113
transform 1 0 23644 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1_N
timestamp 1607194113
transform 1 0 25668 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B2
timestamp 1607194113
transform 1 0 27324 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0855_
timestamp 1607194113
transform 1 0 25852 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_306
timestamp 1607194113
transform 1 0 29256 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_301
timestamp 1607194113
transform 1 0 28796 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_289
timestamp 1607194113
transform 1 0 27692 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2_N
timestamp 1607194113
transform 1 0 27508 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1607194113
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0797_
timestamp 1607194113
transform 1 0 30360 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_338
timestamp 1607194113
transform 1 0 32200 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B2
timestamp 1607194113
transform 1 0 32016 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A2_N
timestamp 1607194113
transform 1 0 31832 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0814_
timestamp 1607194113
transform 1 0 32568 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_69_367
timestamp 1607194113
transform 1 0 34868 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_365
timestamp 1607194113
transform 1 0 34684 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_353
timestamp 1607194113
transform 1 0 33580 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B
timestamp 1607194113
transform 1 0 33396 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1607194113
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A1_N
timestamp 1607194113
transform 1 0 35604 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B1
timestamp 1607194113
transform 1 0 35788 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0753_
timestamp 1607194113
transform 1 0 35972 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B2
timestamp 1607194113
transform 1 0 37628 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A1_N
timestamp 1607194113
transform 1 0 37812 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B1
timestamp 1607194113
transform 1 0 37996 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2_N
timestamp 1607194113
transform 1 0 37444 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0832_
timestamp 1607194113
transform 1 0 38180 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_69_428
timestamp 1607194113
transform 1 0 40480 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_423
timestamp 1607194113
transform 1 0 40020 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B2
timestamp 1607194113
transform 1 0 39836 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A2_N
timestamp 1607194113
transform 1 0 39652 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1607194113
transform 1 0 40388 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_434
timestamp 1607194113
transform 1 0 41032 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1_N
timestamp 1607194113
transform 1 0 41124 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1607194113
transform 1 0 41308 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0749_
timestamp 1607194113
transform 1 0 41492 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_472
timestamp 1607194113
transform 1 0 44528 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_461
timestamp 1607194113
transform 1 0 43516 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A1_N
timestamp 1607194113
transform 1 0 42964 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2_N
timestamp 1607194113
transform 1 0 43332 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B2
timestamp 1607194113
transform 1 0 43148 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0835_
timestamp 1607194113
transform 1 0 43700 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_69_484
timestamp 1607194113
transform 1 0 45632 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1607194113
transform 1 0 46000 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B2
timestamp 1607194113
transform 1 0 25484 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B1
timestamp 1607194113
transform 1 0 23644 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A2_N
timestamp 1607194113
transform 1 0 25300 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0711_
timestamp 1607194113
transform 1 0 23828 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_70_284
timestamp 1607194113
transform 1 0 27232 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_276
timestamp 1607194113
transform 1 0 26496 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_267
timestamp 1607194113
transform 1 0 25668 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1607194113
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0719_
timestamp 1607194113
transform 1 0 27324 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_70_304
timestamp 1607194113
transform 1 0 29072 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_296
timestamp 1607194113
transform 1 0 28336 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1607194113
transform 1 0 29164 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B
timestamp 1607194113
transform 1 0 28152 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_327
timestamp 1607194113
transform 1 0 31188 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B2
timestamp 1607194113
transform 1 0 31004 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A2_N
timestamp 1607194113
transform 1 0 30820 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0807_
timestamp 1607194113
transform 1 0 29348 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_337
timestamp 1607194113
transform 1 0 32108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_335
timestamp 1607194113
transform 1 0 31924 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1607194113
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_361
timestamp 1607194113
transform 1 0 34316 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_349
timestamp 1607194113
transform 1 0 33212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B1
timestamp 1607194113
transform 1 0 34592 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A1_N
timestamp 1607194113
transform 1 0 34776 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0769_
timestamp 1607194113
transform 1 0 34960 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_70_388
timestamp 1607194113
transform 1 0 36800 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A2_N
timestamp 1607194113
transform 1 0 36616 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B2
timestamp 1607194113
transform 1 0 36432 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_398
timestamp 1607194113
transform 1 0 37720 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_396
timestamp 1607194113
transform 1 0 37536 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1607194113
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0850_
timestamp 1607194113
transform 1 0 38272 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_425
timestamp 1607194113
transform 1 0 40204 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_413
timestamp 1607194113
transform 1 0 39100 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_443
timestamp 1607194113
transform 1 0 41860 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_433
timestamp 1607194113
transform 1 0 40940 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0756_
timestamp 1607194113
transform 1 0 41032 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_70_473
timestamp 1607194113
transform 1 0 44620 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_465
timestamp 1607194113
transform 1 0 43884 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_459
timestamp 1607194113
transform 1 0 43332 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_455
timestamp 1607194113
transform 1 0 42964 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1607194113
transform 1 0 43240 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1607194113
transform 1 0 43608 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_482
timestamp 1607194113
transform 1 0 45448 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1054_
timestamp 1607194113
transform 1 0 44804 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_71_245
timestamp 1607194113
transform 1 0 23644 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1_N
timestamp 1607194113
transform 1 0 23736 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B2
timestamp 1607194113
transform 1 0 25392 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0716_
timestamp 1607194113
transform 1 0 23920 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_71_283
timestamp 1607194113
transform 1 0 27140 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_275
timestamp 1607194113
transform 1 0 26404 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_268
timestamp 1607194113
transform 1 0 25760 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A2_N
timestamp 1607194113
transform 1 0 25576 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk_i
timestamp 1607194113
transform 1 0 26128 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk_i
timestamp 1607194113
transform 1 0 27232 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_71_306
timestamp 1607194113
transform 1 0 29256 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_301
timestamp 1607194113
transform 1 0 28796 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_289
timestamp 1607194113
transform 1 0 27692 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_i_A
timestamp 1607194113
transform 1 0 27508 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1607194113
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1_N
timestamp 1607194113
transform 1 0 29808 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0811_
timestamp 1607194113
transform 1 0 29992 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_346
timestamp 1607194113
transform 1 0 32936 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_334
timestamp 1607194113
transform 1 0 31832 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A2_N
timestamp 1607194113
transform 1 0 31648 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B2
timestamp 1607194113
transform 1 0 31464 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_367
timestamp 1607194113
transform 1 0 34868 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_358
timestamp 1607194113
transform 1 0 34040 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1607194113
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_375
timestamp 1607194113
transform 1 0 35604 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0772_
timestamp 1607194113
transform 1 0 35880 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_71_396
timestamp 1607194113
transform 1 0 37536 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2_N
timestamp 1607194113
transform 1 0 37352 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0775_
timestamp 1607194113
transform 1 0 38088 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_428
timestamp 1607194113
transform 1 0 40480 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_423
timestamp 1607194113
transform 1 0 40020 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_411
timestamp 1607194113
transform 1 0 38916 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1607194113
transform 1 0 40388 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_452
timestamp 1607194113
transform 1 0 42688 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_440
timestamp 1607194113
transform 1 0 41584 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_468
timestamp 1607194113
transform 1 0 44160 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_460
timestamp 1607194113
transform 1 0 43424 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_456
timestamp 1607194113
transform 1 0 43056 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A
timestamp 1607194113
transform 1 0 44436 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1052_
timestamp 1607194113
transform 1 0 44620 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1607194113
transform 1 0 43148 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_480
timestamp 1607194113
transform 1 0 45264 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1607194113
transform 1 0 46000 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B2
timestamp 1607194113
transform 1 0 25484 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B1
timestamp 1607194113
transform 1 0 23644 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A2_N
timestamp 1607194113
transform 1 0 25300 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0852_
timestamp 1607194113
transform 1 0 23828 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_276
timestamp 1607194113
transform 1 0 26496 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_274
timestamp 1607194113
transform 1 0 26312 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_267
timestamp 1607194113
transform 1 0 25668 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk_i
timestamp 1607194113
transform 1 0 26036 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1607194113
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_300
timestamp 1607194113
transform 1 0 28704 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_288
timestamp 1607194113
transform 1 0 27600 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_326
timestamp 1607194113
transform 1 0 31096 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_315
timestamp 1607194113
transform 1 0 30084 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1607194113
transform 1 0 30820 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1607194113
transform 1 0 29808 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_337
timestamp 1607194113
transform 1 0 32108 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_334
timestamp 1607194113
transform 1 0 31832 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1607194113
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_361
timestamp 1607194113
transform 1 0 34316 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_349
timestamp 1607194113
transform 1 0 33212 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2_N
timestamp 1607194113
transform 1 0 36892 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0847_
timestamp 1607194113
transform 1 0 35420 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_72_396
timestamp 1607194113
transform 1 0 37536 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_391
timestamp 1607194113
transform 1 0 37076 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B1
timestamp 1607194113
transform 1 0 37352 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1_N
timestamp 1607194113
transform 1 0 37168 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1607194113
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0849_
timestamp 1607194113
transform 1 0 37720 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_428
timestamp 1607194113
transform 1 0 40480 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_416
timestamp 1607194113
transform 1 0 39376 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B2
timestamp 1607194113
transform 1 0 39192 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_452
timestamp 1607194113
transform 1 0 42688 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_440
timestamp 1607194113
transform 1 0 41584 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_466
timestamp 1607194113
transform 1 0 43976 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__CLK
timestamp 1607194113
transform 1 0 44528 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1607194113
transform 1 0 43240 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1055_
timestamp 1607194113
transform 1 0 43332 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1481_
timestamp 1607194113
transform 1 0 44712 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_73_263
timestamp 1607194113
transform 1 0 25300 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A1_N
timestamp 1607194113
transform 1 0 25116 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1174_
timestamp 1607194113
transform 1 0 23644 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A1_N
timestamp 1607194113
transform 1 0 25576 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B1
timestamp 1607194113
transform 1 0 25760 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0718_
timestamp 1607194113
transform 1 0 25944 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_73_306
timestamp 1607194113
transform 1 0 29256 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_302
timestamp 1607194113
transform 1 0 28888 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_290
timestamp 1607194113
transform 1 0 27784 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A2_N
timestamp 1607194113
transform 1 0 27600 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B2
timestamp 1607194113
transform 1 0 27416 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1607194113
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A1_N
timestamp 1607194113
transform 1 0 29440 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B1
timestamp 1607194113
transform 1 0 29624 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0813_
timestamp 1607194113
transform 1 0 29808 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_344
timestamp 1607194113
transform 1 0 32752 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_332
timestamp 1607194113
transform 1 0 31648 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A2_N
timestamp 1607194113
transform 1 0 31464 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B2
timestamp 1607194113
transform 1 0 31280 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_364
timestamp 1607194113
transform 1 0 34592 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_356
timestamp 1607194113
transform 1 0 33856 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1607194113
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1607194113
transform 1 0 34868 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_378
timestamp 1607194113
transform 1 0 35880 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_370
timestamp 1607194113
transform 1 0 35144 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1
timestamp 1607194113
transform 1 0 36064 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1_N
timestamp 1607194113
transform 1 0 36248 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0774_
timestamp 1607194113
transform 1 0 36432 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_402
timestamp 1607194113
transform 1 0 38088 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B2
timestamp 1607194113
transform 1 0 37904 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_428
timestamp 1607194113
transform 1 0 40480 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_426
timestamp 1607194113
transform 1 0 40296 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_414
timestamp 1607194113
transform 1 0 39192 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1607194113
transform 1 0 40388 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_452
timestamp 1607194113
transform 1 0 42688 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_440
timestamp 1607194113
transform 1 0 41584 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A1
timestamp 1607194113
transform 1 0 43792 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1059_
timestamp 1607194113
transform 1 0 43976 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_73_482
timestamp 1607194113
transform 1 0 45448 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B1
timestamp 1607194113
transform 1 0 45264 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1607194113
transform 1 0 46000 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_263
timestamp 1607194113
transform 1 0 25300 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_264
timestamp 1607194113
transform 1 0 25392 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A1_N
timestamp 1607194113
transform 1 0 25116 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1_N
timestamp 1607194113
transform 1 0 25208 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1238_
timestamp 1607194113
transform 1 0 23644 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1175_
timestamp 1607194113
transform 1 0 23736 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_75_275
timestamp 1607194113
transform 1 0 26404 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_276
timestamp 1607194113
transform 1 0 26496 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_272
timestamp 1607194113
transform 1 0 26128 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__CLK
timestamp 1607194113
transform 1 0 26496 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1607194113
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1439_
timestamp 1607194113
transform 1 0 26680 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_306
timestamp 1607194113
transform 1 0 29256 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_297
timestamp 1607194113
transform 1 0 28428 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_296
timestamp 1607194113
transform 1 0 28336 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_288
timestamp 1607194113
transform 1 0 27600 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__CLK
timestamp 1607194113
transform 1 0 28520 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1607194113
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1398_
timestamp 1607194113
transform 1 0 28704 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_318
timestamp 1607194113
transform 1 0 30360 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_319
timestamp 1607194113
transform 1 0 30452 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_338
timestamp 1607194113
transform 1 0 32200 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_330
timestamp 1607194113
transform 1 0 31464 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_337
timestamp 1607194113
transform 1 0 32108 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_335
timestamp 1607194113
transform 1 0 31924 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_331
timestamp 1607194113
transform 1 0 31556 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1607194113
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1440_
timestamp 1607194113
transform 1 0 32292 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1399_
timestamp 1607194113
transform 1 0 32660 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1607194113
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_360
timestamp 1607194113
transform 1 0 34224 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_364
timestamp 1607194113
transform 1 0 34592 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__CLK
timestamp 1607194113
transform 1 0 34040 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__CLK
timestamp 1607194113
transform 1 0 34408 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1607194113
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_387
timestamp 1607194113
transform 1 0 36708 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_379
timestamp 1607194113
transform 1 0 35972 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_385
timestamp 1607194113
transform 1 0 36524 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_373
timestamp 1607194113
transform 1 0 35420 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1_N
timestamp 1607194113
transform 1 0 36800 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1607194113
transform 1 0 36984 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1607194113
transform 1 0 35144 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_408
timestamp 1607194113
transform 1 0 38640 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_408
timestamp 1607194113
transform 1 0 38640 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_400
timestamp 1607194113
transform 1 0 37904 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_396
timestamp 1607194113
transform 1 0 37536 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__CLK
timestamp 1607194113
transform 1 0 38824 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_i_A
timestamp 1607194113
transform 1 0 37720 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk_i
timestamp 1607194113
transform 1 0 37260 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1607194113
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0767_
timestamp 1607194113
transform 1 0 37168 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_75_426
timestamp 1607194113
transform 1 0 40296 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_420
timestamp 1607194113
transform 1 0 39744 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_431
timestamp 1607194113
transform 1 0 40756 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1607194113
transform 1 0 40388 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1479_
timestamp 1607194113
transform 1 0 39008 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0766_
timestamp 1607194113
transform 1 0 40480 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_444
timestamp 1607194113
transform 1 0 41952 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_432
timestamp 1607194113
transform 1 0 40848 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_443
timestamp 1607194113
transform 1 0 41860 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__CLK
timestamp 1607194113
transform 1 0 42136 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1480_
timestamp 1607194113
transform 1 0 42320 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_467
timestamp 1607194113
transform 1 0 44068 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_462
timestamp 1607194113
transform 1 0 43608 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_455
timestamp 1607194113
transform 1 0 42964 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1607194113
transform 1 0 43240 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1607194113
transform 1 0 43332 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_487
timestamp 1607194113
transform 1 0 45908 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_479
timestamp 1607194113
transform 1 0 45172 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_474
timestamp 1607194113
transform 1 0 44712 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1607194113
transform 1 0 45908 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1607194113
transform 1 0 46000 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1056_
timestamp 1607194113
transform 1 0 45080 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1_N
timestamp 1607194113
transform 1 0 25484 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B1
timestamp 1607194113
transform 1 0 23736 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1607194113
transform 1 0 23920 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1239_
timestamp 1607194113
transform 1 0 24012 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_280
timestamp 1607194113
transform 1 0 26864 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_267
timestamp 1607194113
transform 1 0 25668 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1607194113
transform 1 0 26772 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_304
timestamp 1607194113
transform 1 0 29072 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_292
timestamp 1607194113
transform 1 0 27968 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_323
timestamp 1607194113
transform 1 0 30820 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_311
timestamp 1607194113
transform 1 0 29716 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1607194113
transform 1 0 29624 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_342
timestamp 1607194113
transform 1 0 32568 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_335
timestamp 1607194113
transform 1 0 31924 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1607194113
transform 1 0 32476 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_366
timestamp 1607194113
transform 1 0 34776 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_354
timestamp 1607194113
transform 1 0 33672 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_385
timestamp 1607194113
transform 1 0 36524 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_373
timestamp 1607194113
transform 1 0 35420 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1607194113
transform 1 0 35328 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_397
timestamp 1607194113
transform 1 0 37628 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A1_N
timestamp 1607194113
transform 1 0 37812 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__B1
timestamp 1607194113
transform 1 0 37996 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1607194113
transform 1 0 38180 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0843_
timestamp 1607194113
transform 1 0 38272 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_420
timestamp 1607194113
transform 1 0 39744 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_447
timestamp 1607194113
transform 1 0 42228 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_435
timestamp 1607194113
transform 1 0 41124 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_432
timestamp 1607194113
transform 1 0 40848 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1607194113
transform 1 0 41032 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_466
timestamp 1607194113
transform 1 0 43976 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_459
timestamp 1607194113
transform 1 0 43332 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1607194113
transform 1 0 43884 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_478
timestamp 1607194113
transform 1 0 45080 0 -1 44064
box -38 -48 1142 592
use delayline_9_hs  inst_tdelay_line
timestamp 1607276359
transform 1 0 31280 0 1 3761
box 800 801 23264 27367
use sky130_fd_sc_hd__decap_12  FILLER_59_500
timestamp 1607194113
transform 1 0 47104 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_489
timestamp 1607194113
transform 1 0 46092 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_i_A
timestamp 1607194113
transform 1 0 46644 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk_i
timestamp 1607194113
transform 1 0 46828 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_512
timestamp 1607194113
transform 1 0 48208 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A1_N
timestamp 1607194113
transform 1 0 48300 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B1
timestamp 1607194113
transform 1 0 48484 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0825_
timestamp 1607194113
transform 1 0 48668 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_537
timestamp 1607194113
transform 1 0 50508 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B2
timestamp 1607194113
transform 1 0 50324 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A2_N
timestamp 1607194113
transform 1 0 50140 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_562
timestamp 1607194113
transform 1 0 52808 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_550
timestamp 1607194113
transform 1 0 51704 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607194113
transform 1 0 51612 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1516_
timestamp 1607194113
transform 1 0 53544 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_59_600
timestamp 1607194113
transform 1 0 56304 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_591
timestamp 1607194113
transform 1 0 55476 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__CLK
timestamp 1607194113
transform 1 0 55292 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A2_N
timestamp 1607194113
transform 1 0 56764 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B2
timestamp 1607194113
transform 1 0 56948 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B1
timestamp 1607194113
transform 1 0 56580 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1607194113
transform 1 0 56028 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_609
timestamp 1607194113
transform 1 0 57132 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_inp_i
timestamp 1607194113
transform 1 0 58788 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607194113
transform 1 0 57224 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1267_
timestamp 1607194113
transform 1 0 57316 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_642
timestamp 1607194113
transform 1 0 60168 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[8]
timestamp 1607194113
transform 1 0 59340 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[7]
timestamp 1607194113
transform 1 0 59156 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[6]
timestamp 1607194113
transform 1 0 58972 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[4]
timestamp 1607194113
transform 1 0 59984 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[2]
timestamp 1607194113
transform 1 0 59800 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk_i
timestamp 1607194113
transform 1 0 59524 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_663
timestamp 1607194113
transform 1 0 62100 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_654
timestamp 1607194113
transform 1 0 61272 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1607194113
transform 1 0 61824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__D
timestamp 1607194113
transform 1 0 62652 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607194113
transform 1 0 62836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1389_
timestamp 1607194113
transform 1 0 62928 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_703
timestamp 1607194113
transform 1 0 65780 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_691
timestamp 1607194113
transform 1 0 64676 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_715
timestamp 1607194113
transform 1 0 66884 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_731
timestamp 1607194113
transform 1 0 68356 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_727
timestamp 1607194113
transform 1 0 67988 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607194113
transform 1 0 68448 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_507
timestamp 1607194113
transform 1 0 47748 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_495
timestamp 1607194113
transform 1 0 46644 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_520
timestamp 1607194113
transform 1 0 48944 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B1
timestamp 1607194113
transform 1 0 49312 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1_N
timestamp 1607194113
transform 1 0 49496 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607194113
transform 1 0 48852 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0821_
timestamp 1607194113
transform 1 0 49680 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B2
timestamp 1607194113
transform 1 0 51336 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A2_N
timestamp 1607194113
transform 1 0 51152 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1_N
timestamp 1607194113
transform 1 0 51520 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B1
timestamp 1607194113
transform 1 0 51704 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0818_
timestamp 1607194113
transform 1 0 51888 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_581
timestamp 1607194113
transform 1 0 54556 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_572
timestamp 1607194113
transform 1 0 53728 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2_N
timestamp 1607194113
transform 1 0 53544 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B2
timestamp 1607194113
transform 1 0 53360 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607194113
transform 1 0 54464 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_595
timestamp 1607194113
transform 1 0 55844 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_589
timestamp 1607194113
transform 1 0 55292 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk_i
timestamp 1607194113
transform 1 0 55568 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1515_
timestamp 1607194113
transform 1 0 56028 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_60_616
timestamp 1607194113
transform 1 0 57776 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_i_A
timestamp 1607194113
transform 1 0 58328 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[5]
timestamp 1607194113
transform 1 0 58788 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk_i
timestamp 1607194113
transform 1 0 58512 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_642
timestamp 1607194113
transform 1 0 60168 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_635
timestamp 1607194113
transform 1 0 59524 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[3]
timestamp 1607194113
transform 1 0 59340 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[1]
timestamp 1607194113
transform 1 0 59156 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[0]
timestamp 1607194113
transform 1 0 58972 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607194113
transform 1 0 60076 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_654
timestamp 1607194113
transform 1 0 61272 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1379_
timestamp 1607194113
transform 1 0 62008 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_60_681
timestamp 1607194113
transform 1 0 63756 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_706
timestamp 1607194113
transform 1 0 66056 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_700
timestamp 1607194113
transform 1 0 65504 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_692
timestamp 1607194113
transform 1 0 64768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607194113
transform 1 0 65688 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1607194113
transform 1 0 65780 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1607194113
transform 1 0 64492 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_718
timestamp 1607194113
transform 1 0 67160 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_730
timestamp 1607194113
transform 1 0 68264 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_502
timestamp 1607194113
transform 1 0 47288 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_501
timestamp 1607194113
transform 1 0 47196 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_489
timestamp 1607194113
transform 1 0 46092 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_518
timestamp 1607194113
transform 1 0 48760 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_514
timestamp 1607194113
transform 1 0 48392 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_513
timestamp 1607194113
transform 1 0 48300 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_520
timestamp 1607194113
transform 1 0 48944 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A1_N
timestamp 1607194113
transform 1 0 49036 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B1
timestamp 1607194113
transform 1 0 49496 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B1
timestamp 1607194113
transform 1 0 49220 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A1_N
timestamp 1607194113
transform 1 0 49680 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607194113
transform 1 0 48852 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0823_
timestamp 1607194113
transform 1 0 49404 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_545
timestamp 1607194113
transform 1 0 51244 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B2
timestamp 1607194113
transform 1 0 51060 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A2_N
timestamp 1607194113
transform 1 0 50876 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A2_N
timestamp 1607194113
transform 1 0 51336 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0837_
timestamp 1607194113
transform 1 0 49864 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_563
timestamp 1607194113
transform 1 0 52900 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_550
timestamp 1607194113
transform 1 0 51704 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_559
timestamp 1607194113
transform 1 0 52532 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B2
timestamp 1607194113
transform 1 0 51520 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B
timestamp 1607194113
transform 1 0 51888 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607194113
transform 1 0 51612 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0826_
timestamp 1607194113
transform 1 0 51704 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1607194113
transform 1 0 53268 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0787_
timestamp 1607194113
transform 1 0 52072 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_581
timestamp 1607194113
transform 1 0 54556 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_579
timestamp 1607194113
transform 1 0 54372 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_575
timestamp 1607194113
transform 1 0 54004 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_582
timestamp 1607194113
transform 1 0 54648 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_570
timestamp 1607194113
transform 1 0 53544 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B2
timestamp 1607194113
transform 1 0 54832 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1607194113
transform 1 0 55016 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607194113
transform 1 0 54464 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_593
timestamp 1607194113
transform 1 0 55660 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_601
timestamp 1607194113
transform 1 0 56396 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_602
timestamp 1607194113
transform 1 0 56488 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A2_N
timestamp 1607194113
transform 1 0 56764 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B2
timestamp 1607194113
transform 1 0 56948 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B2
timestamp 1607194113
transform 1 0 56488 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1607194113
transform 1 0 56672 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B1
timestamp 1607194113
transform 1 0 56580 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0933_
timestamp 1607194113
transform 1 0 55200 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _0927_
timestamp 1607194113
transform 1 0 56856 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_620
timestamp 1607194113
transform 1 0 58144 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_627
timestamp 1607194113
transform 1 0 58788 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_609
timestamp 1607194113
transform 1 0 57132 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607194113
transform 1 0 57224 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1204_
timestamp 1607194113
transform 1 0 57316 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_642
timestamp 1607194113
transform 1 0 60168 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_640
timestamp 1607194113
transform 1 0 59984 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_632
timestamp 1607194113
transform 1 0 59248 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_639
timestamp 1607194113
transform 1 0 59892 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607194113
transform 1 0 60076 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_662
timestamp 1607194113
transform 1 0 62008 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_654
timestamp 1607194113
transform 1 0 61272 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_663
timestamp 1607194113
transform 1 0 62100 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_651
timestamp 1607194113
transform 1 0 60996 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__D
timestamp 1607194113
transform 1 0 62192 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1430_
timestamp 1607194113
transform 1 0 62376 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_685
timestamp 1607194113
transform 1 0 64124 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_680
timestamp 1607194113
transform 1 0 63664 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_672
timestamp 1607194113
transform 1 0 62928 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607194113
transform 1 0 62836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1420_
timestamp 1607194113
transform 1 0 63756 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_62_701
timestamp 1607194113
transform 1 0 65596 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_697
timestamp 1607194113
transform 1 0 65228 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_700
timestamp 1607194113
transform 1 0 65504 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607194113
transform 1 0 65688 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0795_
timestamp 1607194113
transform 1 0 65780 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_724
timestamp 1607194113
transform 1 0 67712 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_712
timestamp 1607194113
transform 1 0 66608 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_723
timestamp 1607194113
transform 1 0 67620 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_711
timestamp 1607194113
transform 1 0 66516 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1607194113
transform 1 0 66240 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_731
timestamp 1607194113
transform 1 0 68356 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607194113
transform 1 0 68448 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1607194113
transform 1 0 47564 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1265_
timestamp 1607194113
transform 1 0 46092 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1607194113
transform 1 0 48300 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1
timestamp 1607194113
transform 1 0 48576 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1_N
timestamp 1607194113
transform 1 0 48760 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0838_
timestamp 1607194113
transform 1 0 48944 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_63_540
timestamp 1607194113
transform 1 0 50784 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A2_N
timestamp 1607194113
transform 1 0 50600 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B2
timestamp 1607194113
transform 1 0 50416 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_561
timestamp 1607194113
transform 1 0 52716 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_553
timestamp 1607194113
transform 1 0 51980 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_548
timestamp 1607194113
transform 1 0 51520 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1607194113
transform 1 0 51612 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0827_
timestamp 1607194113
transform 1 0 52992 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1607194113
transform 1 0 51704 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_578
timestamp 1607194113
transform 1 0 54280 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_602
timestamp 1607194113
transform 1 0 56488 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_590
timestamp 1607194113
transform 1 0 55384 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_623
timestamp 1607194113
transform 1 0 58420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_611
timestamp 1607194113
transform 1 0 57316 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1607194113
transform 1 0 57224 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_647
timestamp 1607194113
transform 1 0 60628 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_635
timestamp 1607194113
transform 1 0 59524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_663
timestamp 1607194113
transform 1 0 62100 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_653
timestamp 1607194113
transform 1 0 61180 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0695_
timestamp 1607194113
transform 1 0 61272 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_672
timestamp 1607194113
transform 1 0 62928 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1607194113
transform 1 0 62836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0688_
timestamp 1607194113
transform 1 0 63020 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_63_689
timestamp 1607194113
transform 1 0 64492 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B1
timestamp 1607194113
transform 1 0 64308 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0694_
timestamp 1607194113
transform 1 0 65044 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_63_725
timestamp 1607194113
transform 1 0 67804 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_713
timestamp 1607194113
transform 1 0 66700 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A2
timestamp 1607194113
transform 1 0 66516 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B2
timestamp 1607194113
transform 1 0 66332 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_731
timestamp 1607194113
transform 1 0 68356 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1607194113
transform 1 0 68448 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_489
timestamp 1607194113
transform 1 0 46092 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1380_
timestamp 1607194113
transform 1 0 46276 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_64_520
timestamp 1607194113
transform 1 0 48944 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_518
timestamp 1607194113
transform 1 0 48760 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_512
timestamp 1607194113
transform 1 0 48208 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__CLK
timestamp 1607194113
transform 1 0 48024 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__D
timestamp 1607194113
transform 1 0 49680 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1607194113
transform 1 0 48852 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1434_
timestamp 1607194113
transform 1 0 49864 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_64_551
timestamp 1607194113
transform 1 0 51796 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__CLK
timestamp 1607194113
transform 1 0 51612 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0742_
timestamp 1607194113
transform 1 0 52348 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_64_577
timestamp 1607194113
transform 1 0 54188 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_571
timestamp 1607194113
transform 1 0 53636 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1607194113
transform 1 0 54280 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1607194113
transform 1 0 54464 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0858_
timestamp 1607194113
transform 1 0 54556 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_64_602
timestamp 1607194113
transform 1 0 56488 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_590
timestamp 1607194113
transform 1 0 55384 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A2_N
timestamp 1607194113
transform 1 0 57224 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B2
timestamp 1607194113
transform 1 0 57408 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B1
timestamp 1607194113
transform 1 0 57592 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1201_
timestamp 1607194113
transform 1 0 57776 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_642
timestamp 1607194113
transform 1 0 60168 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_640
timestamp 1607194113
transform 1 0 59984 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_632
timestamp 1607194113
transform 1 0 59248 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1607194113
transform 1 0 60076 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_662
timestamp 1607194113
transform 1 0 62008 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_658
timestamp 1607194113
transform 1 0 61640 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_654
timestamp 1607194113
transform 1 0 61272 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1607194113
transform 1 0 61732 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_684
timestamp 1607194113
transform 1 0 64032 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1607194113
transform 1 0 62560 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0790_
timestamp 1607194113
transform 1 0 62744 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_64_696
timestamp 1607194113
transform 1 0 65136 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1607194113
transform 1 0 65688 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0794_
timestamp 1607194113
transform 1 0 65780 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_64_721
timestamp 1607194113
transform 1 0 67436 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A2
timestamp 1607194113
transform 1 0 67252 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B2
timestamp 1607194113
transform 1 0 67068 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1607194113
transform 1 0 47840 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_491
timestamp 1607194113
transform 1 0 46276 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B2
timestamp 1607194113
transform 1 0 46092 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1202_
timestamp 1607194113
transform 1 0 46368 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_519
timestamp 1607194113
transform 1 0 48852 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1607194113
transform 1 0 48576 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_543
timestamp 1607194113
transform 1 0 51060 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_531
timestamp 1607194113
transform 1 0 49956 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_550
timestamp 1607194113
transform 1 0 51704 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__D
timestamp 1607194113
transform 1 0 52072 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1607194113
transform 1 0 51612 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1393_
timestamp 1607194113
transform 1 0 52256 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_586
timestamp 1607194113
transform 1 0 55016 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_577
timestamp 1607194113
transform 1 0 54188 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__CLK
timestamp 1607194113
transform 1 0 54004 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1607194113
transform 1 0 54740 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_606
timestamp 1607194113
transform 1 0 56856 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_598
timestamp 1607194113
transform 1 0 56120 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A2_N
timestamp 1607194113
transform 1 0 57500 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B2
timestamp 1607194113
transform 1 0 57316 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B1
timestamp 1607194113
transform 1 0 57040 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1607194113
transform 1 0 57224 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1264_
timestamp 1607194113
transform 1 0 57684 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_631
timestamp 1607194113
transform 1 0 59156 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1381_
timestamp 1607194113
transform 1 0 60260 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_662
timestamp 1607194113
transform 1 0 62008 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_678
timestamp 1607194113
transform 1 0 63480 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_672
timestamp 1607194113
transform 1 0 62928 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_670
timestamp 1607194113
transform 1 0 62744 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1607194113
transform 1 0 62836 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0691_
timestamp 1607194113
transform 1 0 63572 0 1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_65_704
timestamp 1607194113
transform 1 0 65872 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_697
timestamp 1607194113
transform 1 0 65228 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A2
timestamp 1607194113
transform 1 0 65044 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B2
timestamp 1607194113
transform 1 0 64860 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1607194113
transform 1 0 65596 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_716
timestamp 1607194113
transform 1 0 66976 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_728
timestamp 1607194113
transform 1 0 68080 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1607194113
transform 1 0 68448 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_508
timestamp 1607194113
transform 1 0 47840 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_504
timestamp 1607194113
transform 1 0 47472 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_492
timestamp 1607194113
transform 1 0 46368 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_489
timestamp 1607194113
transform 1 0 46092 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B1
timestamp 1607194113
transform 1 0 46184 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1607194113
transform 1 0 47564 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_520
timestamp 1607194113
transform 1 0 48944 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_516
timestamp 1607194113
transform 1 0 48576 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1607194113
transform 1 0 48852 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_544
timestamp 1607194113
transform 1 0 51152 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_532
timestamp 1607194113
transform 1 0 50048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A2_N
timestamp 1607194113
transform 1 0 53176 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0724_
timestamp 1607194113
transform 1 0 51704 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_581
timestamp 1607194113
transform 1 0 54556 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_578
timestamp 1607194113
transform 1 0 54280 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_570
timestamp 1607194113
transform 1 0 53544 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B1
timestamp 1607194113
transform 1 0 53360 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1607194113
transform 1 0 54464 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_605
timestamp 1607194113
transform 1 0 56764 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_593
timestamp 1607194113
transform 1 0 55660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_617
timestamp 1607194113
transform 1 0 57868 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_646
timestamp 1607194113
transform 1 0 60536 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_642
timestamp 1607194113
transform 1 0 60168 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_629
timestamp 1607194113
transform 1 0 58972 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1607194113
transform 1 0 60076 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1422_
timestamp 1607194113
transform 1 0 60628 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_666
timestamp 1607194113
transform 1 0 62376 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0792_
timestamp 1607194113
transform 1 0 63480 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_66_703
timestamp 1607194113
transform 1 0 65780 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_696
timestamp 1607194113
transform 1 0 65136 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A2
timestamp 1607194113
transform 1 0 64952 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B2
timestamp 1607194113
transform 1 0 64768 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1607194113
transform 1 0 65688 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_715
timestamp 1607194113
transform 1 0 66884 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_727
timestamp 1607194113
transform 1 0 67988 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_503
timestamp 1607194113
transform 1 0 47380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_491
timestamp 1607194113
transform 1 0 46276 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_497
timestamp 1607194113
transform 1 0 46828 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_489
timestamp 1607194113
transform 1 0 46092 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1_N
timestamp 1607194113
transform 1 0 47104 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0809_
timestamp 1607194113
transform 1 0 47288 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_515
timestamp 1607194113
transform 1 0 48484 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_522
timestamp 1607194113
transform 1 0 49128 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2_N
timestamp 1607194113
transform 1 0 48944 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B2
timestamp 1607194113
transform 1 0 48760 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1607194113
transform 1 0 48852 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1421_
timestamp 1607194113
transform 1 0 48944 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_541
timestamp 1607194113
transform 1 0 50876 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_546
timestamp 1607194113
transform 1 0 51336 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_534
timestamp 1607194113
transform 1 0 50232 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__CLK
timestamp 1607194113
transform 1 0 50692 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_557
timestamp 1607194113
transform 1 0 52348 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_553
timestamp 1607194113
transform 1 0 51980 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_558
timestamp 1607194113
transform 1 0 52440 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_550
timestamp 1607194113
transform 1 0 51704 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1607194113
transform 1 0 51612 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1069_
timestamp 1607194113
transform 1 0 53084 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _0817_
timestamp 1607194113
transform 1 0 52624 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1607194113
transform 1 0 52072 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_572
timestamp 1607194113
transform 1 0 53728 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_580
timestamp 1607194113
transform 1 0 54464 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1607194113
transform 1 0 54280 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A2_N
timestamp 1607194113
transform 1 0 54096 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1607194113
transform 1 0 54464 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1078_
timestamp 1607194113
transform 1 0 54556 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_68_592
timestamp 1607194113
transform 1 0 55568 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_598
timestamp 1607194113
transform 1 0 56120 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_592
timestamp 1607194113
transform 1 0 55568 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__CLK
timestamp 1607194113
transform 1 0 55936 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1607194113
transform 1 0 55936 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1607194113
transform 1 0 55384 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1476_
timestamp 1607194113
transform 1 0 56120 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1607194113
transform 1 0 55660 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_617
timestamp 1607194113
transform 1 0 57868 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_623
timestamp 1607194113
transform 1 0 58420 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_611
timestamp 1607194113
transform 1 0 57316 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1607194113
transform 1 0 57224 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_642
timestamp 1607194113
transform 1 0 60168 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_629
timestamp 1607194113
transform 1 0 58972 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_647
timestamp 1607194113
transform 1 0 60628 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_635
timestamp 1607194113
transform 1 0 59524 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1607194113
transform 1 0 60076 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_665
timestamp 1607194113
transform 1 0 62284 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_654
timestamp 1607194113
transform 1 0 61272 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_659
timestamp 1607194113
transform 1 0 61732 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1082_
timestamp 1607194113
transform 1 0 61640 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_68_682
timestamp 1607194113
transform 1 0 63848 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_682
timestamp 1607194113
transform 1 0 63848 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_672
timestamp 1607194113
transform 1 0 62928 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1607194113
transform 1 0 63664 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1607194113
transform 1 0 62836 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1091_
timestamp 1607194113
transform 1 0 63204 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1081_
timestamp 1607194113
transform 1 0 63020 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_68_703
timestamp 1607194113
transform 1 0 65780 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_699
timestamp 1607194113
transform 1 0 65412 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_691
timestamp 1607194113
transform 1 0 64676 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_705
timestamp 1607194113
transform 1 0 65964 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_693
timestamp 1607194113
transform 1 0 64860 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1607194113
transform 1 0 65688 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1607194113
transform 1 0 64400 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1607194113
transform 1 0 64584 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_722
timestamp 1607194113
transform 1 0 67528 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_714
timestamp 1607194113
transform 1 0 66792 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_717
timestamp 1607194113
transform 1 0 67068 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1607194113
transform 1 0 67896 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk_i
timestamp 1607194113
transform 1 0 66516 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1607194113
transform 1 0 67620 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_728
timestamp 1607194113
transform 1 0 68080 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_729
timestamp 1607194113
transform 1 0 68172 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__CLK
timestamp 1607194113
transform 1 0 68448 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1607194113
transform 1 0 68448 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_489
timestamp 1607194113
transform 1 0 46092 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A1_N
timestamp 1607194113
transform 1 0 47196 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0714_
timestamp 1607194113
transform 1 0 47380 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_523
timestamp 1607194113
transform 1 0 49220 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A2_N
timestamp 1607194113
transform 1 0 49036 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B2
timestamp 1607194113
transform 1 0 48852 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_547
timestamp 1607194113
transform 1 0 51428 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_535
timestamp 1607194113
transform 1 0 50324 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_564
timestamp 1607194113
transform 1 0 52992 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_556
timestamp 1607194113
transform 1 0 52256 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_550
timestamp 1607194113
transform 1 0 51704 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1607194113
transform 1 0 51612 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1077_
timestamp 1607194113
transform 1 0 52348 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1475_
timestamp 1607194113
transform 1 0 53728 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_69_605
timestamp 1607194113
transform 1 0 56764 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_593
timestamp 1607194113
transform 1 0 55660 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__CLK
timestamp 1607194113
transform 1 0 55476 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_623
timestamp 1607194113
transform 1 0 58420 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_611
timestamp 1607194113
transform 1 0 57316 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_609
timestamp 1607194113
transform 1 0 57132 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1607194113
transform 1 0 57224 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_641
timestamp 1607194113
transform 1 0 60076 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_635
timestamp 1607194113
transform 1 0 59524 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1470_
timestamp 1607194113
transform 1 0 60168 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_69_663
timestamp 1607194113
transform 1 0 62100 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__CLK
timestamp 1607194113
transform 1 0 61916 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_672
timestamp 1607194113
transform 1 0 62928 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1607194113
transform 1 0 62836 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1471_
timestamp 1607194113
transform 1 0 63664 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_701
timestamp 1607194113
transform 1 0 65596 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__CLK
timestamp 1607194113
transform 1 0 65412 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_724
timestamp 1607194113
transform 1 0 67712 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_713
timestamp 1607194113
transform 1 0 66700 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1607194113
transform 1 0 67252 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1607194113
transform 1 0 67436 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1607194113
transform 1 0 68448 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_506
timestamp 1607194113
transform 1 0 47656 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_494
timestamp 1607194113
transform 1 0 46552 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_520
timestamp 1607194113
transform 1 0 48944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_518
timestamp 1607194113
transform 1 0 48760 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1607194113
transform 1 0 48852 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_544
timestamp 1607194113
transform 1 0 51152 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_532
timestamp 1607194113
transform 1 0 50048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_558
timestamp 1607194113
transform 1 0 52440 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_552
timestamp 1607194113
transform 1 0 51888 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1607194113
transform 1 0 52256 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1068_
timestamp 1607194113
transform 1 0 52992 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1607194113
transform 1 0 51980 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_581
timestamp 1607194113
transform 1 0 54556 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_579
timestamp 1607194113
transform 1 0 54372 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_571
timestamp 1607194113
transform 1 0 53636 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1607194113
transform 1 0 54464 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_600
timestamp 1607194113
transform 1 0 56304 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1607194113
transform 1 0 56120 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1075_
timestamp 1607194113
transform 1 0 56856 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 55292 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_617
timestamp 1607194113
transform 1 0 57868 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1607194113
transform 1 0 57684 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_646
timestamp 1607194113
transform 1 0 60536 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_642
timestamp 1607194113
transform 1 0 60168 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_629
timestamp 1607194113
transform 1 0 58972 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1607194113
transform 1 0 60076 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1607194113
transform 1 0 60628 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_650
timestamp 1607194113
transform 1 0 60904 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1093_
timestamp 1607194113
transform 1 0 61640 0 -1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_70_674
timestamp 1607194113
transform 1 0 63112 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B1
timestamp 1607194113
transform 1 0 62928 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1092_
timestamp 1607194113
transform 1 0 63664 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_703
timestamp 1607194113
transform 1 0 65780 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_699
timestamp 1607194113
transform 1 0 65412 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_691
timestamp 1607194113
transform 1 0 64676 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1607194113
transform 1 0 64492 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1607194113
transform 1 0 65688 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_726
timestamp 1607194113
transform 1 0 67896 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_714
timestamp 1607194113
transform 1 0 66792 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk_i
timestamp 1607194113
transform 1 0 66516 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1607194113
transform 1 0 68448 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_501
timestamp 1607194113
transform 1 0 47196 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_489
timestamp 1607194113
transform 1 0 46092 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_525
timestamp 1607194113
transform 1 0 49404 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_513
timestamp 1607194113
transform 1 0 48300 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_537
timestamp 1607194113
transform 1 0 50508 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_550
timestamp 1607194113
transform 1 0 51704 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B1
timestamp 1607194113
transform 1 0 53176 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1607194113
transform 1 0 51612 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1079_
timestamp 1607194113
transform 1 0 51888 0 1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_71_581
timestamp 1607194113
transform 1 0 54556 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_568
timestamp 1607194113
transform 1 0 53360 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _1032_
timestamp 1607194113
transform 1 0 53912 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_71_598
timestamp 1607194113
transform 1 0 56120 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1607194113
transform 1 0 55936 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1070_
timestamp 1607194113
transform 1 0 55292 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_71_623
timestamp 1607194113
transform 1 0 58420 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_611
timestamp 1607194113
transform 1 0 57316 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1607194113
transform 1 0 57224 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_647
timestamp 1607194113
transform 1 0 60628 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_635
timestamp 1607194113
transform 1 0 59524 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_662
timestamp 1607194113
transform 1 0 62008 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_653
timestamp 1607194113
transform 1 0 61180 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1607194113
transform 1 0 60996 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1607194113
transform 1 0 61548 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1607194113
transform 1 0 60720 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1607194113
transform 1 0 61732 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_683
timestamp 1607194113
transform 1 0 63940 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_670
timestamp 1607194113
transform 1 0 62744 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__C
timestamp 1607194113
transform 1 0 63756 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1607194113
transform 1 0 62836 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1049_
timestamp 1607194113
transform 1 0 62928 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_704
timestamp 1607194113
transform 1 0 65872 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_692
timestamp 1607194113
transform 1 0 64768 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_i_A
timestamp 1607194113
transform 1 0 64308 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk_i
timestamp 1607194113
transform 1 0 64492 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_716
timestamp 1607194113
transform 1 0 66976 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__D
timestamp 1607194113
transform 1 0 68080 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1607194113
transform 1 0 68264 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1607194113
transform 1 0 68448 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_505
timestamp 1607194113
transform 1 0 47564 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_493
timestamp 1607194113
transform 1 0 46460 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_525
timestamp 1607194113
transform 1 0 49404 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_517
timestamp 1607194113
transform 1 0 48668 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1607194113
transform 1 0 49220 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1607194113
transform 1 0 48852 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1607194113
transform 1 0 48944 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_537
timestamp 1607194113
transform 1 0 50508 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_564
timestamp 1607194113
transform 1 0 52992 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_552
timestamp 1607194113
transform 1 0 51888 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1607194113
transform 1 0 51612 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1607194113
transform 1 0 53084 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_574
timestamp 1607194113
transform 1 0 53912 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_568
timestamp 1607194113
transform 1 0 53360 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_i_A
timestamp 1607194113
transform 1 0 54004 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk_i
timestamp 1607194113
transform 1 0 54188 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1607194113
transform 1 0 54464 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1050_
timestamp 1607194113
transform 1 0 54556 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_604
timestamp 1607194113
transform 1 0 56672 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_592
timestamp 1607194113
transform 1 0 55568 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1607194113
transform 1 0 55384 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_616
timestamp 1607194113
transform 1 0 57776 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_635
timestamp 1607194113
transform 1 0 59524 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_628
timestamp 1607194113
transform 1 0 58880 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1607194113
transform 1 0 59892 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1607194113
transform 1 0 59340 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1607194113
transform 1 0 60076 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1086_
timestamp 1607194113
transform 1 0 60168 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0751_
timestamp 1607194113
transform 1 0 58972 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_654
timestamp 1607194113
transform 1 0 61272 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__D
timestamp 1607194113
transform 1 0 61824 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1038_
timestamp 1607194113
transform 1 0 62008 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_686
timestamp 1607194113
transform 1 0 64216 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_671
timestamp 1607194113
transform 1 0 62836 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1083_
timestamp 1607194113
transform 1 0 63572 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_72_698
timestamp 1607194113
transform 1 0 65320 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1607194113
transform 1 0 65688 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0779_
timestamp 1607194113
transform 1 0 65780 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_719
timestamp 1607194113
transform 1 0 67252 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_715
timestamp 1607194113
transform 1 0 66884 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_709
timestamp 1607194113
transform 1 0 66332 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1607194113
transform 1 0 66148 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1607194113
transform 1 0 66976 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_731
timestamp 1607194113
transform 1 0 68356 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1097_
timestamp 1607194113
transform 1 0 68448 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_73_504
timestamp 1607194113
transform 1 0 47472 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_492
timestamp 1607194113
transform 1 0 46368 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1607194113
transform 1 0 46092 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_526
timestamp 1607194113
transform 1 0 49496 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1607194113
transform 1 0 49312 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1066_
timestamp 1607194113
transform 1 0 48024 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_73_546
timestamp 1607194113
transform 1 0 51336 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_538
timestamp 1607194113
transform 1 0 50600 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1607194113
transform 1 0 51612 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1474_
timestamp 1607194113
transform 1 0 51704 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_73_583
timestamp 1607194113
transform 1 0 54740 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_571
timestamp 1607194113
transform 1 0 53636 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__CLK
timestamp 1607194113
transform 1 0 53452 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1607194113
transform 1 0 54924 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_601
timestamp 1607194113
transform 1 0 56396 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_588
timestamp 1607194113
transform 1 0 55200 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1607194113
transform 1 0 56212 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1607194113
transform 1 0 55936 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_623
timestamp 1607194113
transform 1 0 58420 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_611
timestamp 1607194113
transform 1 0 57316 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_609
timestamp 1607194113
transform 1 0 57132 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1607194113
transform 1 0 57224 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_631
timestamp 1607194113
transform 1 0 59156 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A1
timestamp 1607194113
transform 1 0 59340 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1085_
timestamp 1607194113
transform 1 0 59524 0 1 41888
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_73_663
timestamp 1607194113
transform 1 0 62100 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_650
timestamp 1607194113
transform 1 0 60904 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__B1
timestamp 1607194113
transform 1 0 60720 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1084_
timestamp 1607194113
transform 1 0 61456 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_73_681
timestamp 1607194113
transform 1 0 63756 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1607194113
transform 1 0 62836 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1088_
timestamp 1607194113
transform 1 0 62928 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_73_701
timestamp 1607194113
transform 1 0 65596 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_693
timestamp 1607194113
transform 1 0 64860 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1099_
timestamp 1607194113
transform 1 0 65780 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_717
timestamp 1607194113
transform 1 0 67068 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1607194113
transform 1 0 66884 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_729
timestamp 1607194113
transform 1 0 68172 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1607194113
transform 1 0 68448 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_489
timestamp 1607194113
transform 1 0 46092 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_501
timestamp 1607194113
transform 1 0 47196 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_489
timestamp 1607194113
transform 1 0 46092 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1478_
timestamp 1607194113
transform 1 0 46460 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1063_
timestamp 1607194113
transform 1 0 47472 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_75_514
timestamp 1607194113
transform 1 0 48392 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_511
timestamp 1607194113
transform 1 0 48116 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__CLK
timestamp 1607194113
transform 1 0 48208 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1607194113
transform 1 0 48852 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1065_
timestamp 1607194113
transform 1 0 48944 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1051_
timestamp 1607194113
transform 1 0 48944 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_75_540
timestamp 1607194113
transform 1 0 50784 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_75_531
timestamp 1607194113
transform 1 0 49956 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_544
timestamp 1607194113
transform 1 0 51152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_529
timestamp 1607194113
transform 1 0 49772 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1607194113
transform 1 0 49772 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1607194113
transform 1 0 50508 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1061_
timestamp 1607194113
transform 1 0 50508 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_75_562
timestamp 1607194113
transform 1 0 52808 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_550
timestamp 1607194113
transform 1 0 51704 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_548
timestamp 1607194113
transform 1 0 51520 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_556
timestamp 1607194113
transform 1 0 52256 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1607194113
transform 1 0 51612 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_586
timestamp 1607194113
transform 1 0 55016 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_574
timestamp 1607194113
transform 1 0 53912 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_581
timestamp 1607194113
transform 1 0 54556 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_568
timestamp 1607194113
transform 1 0 53360 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1607194113
transform 1 0 54464 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1477_
timestamp 1607194113
transform 1 0 54740 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_75_600
timestamp 1607194113
transform 1 0 56304 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_604
timestamp 1607194113
transform 1 0 56672 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__CLK
timestamp 1607194113
transform 1 0 56488 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1073_
timestamp 1607194113
transform 1 0 55200 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_623
timestamp 1607194113
transform 1 0 58420 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_611
timestamp 1607194113
transform 1 0 57316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_608
timestamp 1607194113
transform 1 0 57040 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_625
timestamp 1607194113
transform 1 0 58604 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B1
timestamp 1607194113
transform 1 0 58420 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1607194113
transform 1 0 57224 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1072_
timestamp 1607194113
transform 1 0 57224 0 -1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_75_631
timestamp 1607194113
transform 1 0 59156 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_646
timestamp 1607194113
transform 1 0 60536 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_642
timestamp 1607194113
transform 1 0 60168 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_637
timestamp 1607194113
transform 1 0 59708 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1607194113
transform 1 0 60076 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1473_
timestamp 1607194113
transform 1 0 59248 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1607194113
transform 1 0 60260 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1607194113
transform 1 0 62284 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_653
timestamp 1607194113
transform 1 0 61180 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__CLK
timestamp 1607194113
transform 1 0 60996 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1472_
timestamp 1607194113
transform 1 0 61272 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_684
timestamp 1607194113
transform 1 0 64032 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_672
timestamp 1607194113
transform 1 0 62928 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_675
timestamp 1607194113
transform 1 0 63204 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__CLK
timestamp 1607194113
transform 1 0 63020 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1607194113
transform 1 0 62836 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_704
timestamp 1607194113
transform 1 0 65872 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_696
timestamp 1607194113
transform 1 0 65136 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_699
timestamp 1607194113
transform 1 0 65412 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_687
timestamp 1607194113
transform 1 0 64308 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1607194113
transform 1 0 65688 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1469_
timestamp 1607194113
transform 1 0 65780 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1098_
timestamp 1607194113
transform 1 0 65964 0 1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_75_722
timestamp 1607194113
transform 1 0 67528 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_724
timestamp 1607194113
transform 1 0 67712 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__CLK
timestamp 1607194113
transform 1 0 67528 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1607194113
transform 1 0 67344 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A1
timestamp 1607194113
transform 1 0 67160 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_730
timestamp 1607194113
transform 1 0 68264 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1607194113
transform 1 0 68448 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_505
timestamp 1607194113
transform 1 0 47564 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_501
timestamp 1607194113
transform 1 0 47196 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_497
timestamp 1607194113
transform 1 0 46828 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_490
timestamp 1607194113
transform 1 0 46184 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1607194113
transform 1 0 46736 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1607194113
transform 1 0 47288 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_526
timestamp 1607194113
transform 1 0 49496 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_518
timestamp 1607194113
transform 1 0 48760 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_513
timestamp 1607194113
transform 1 0 48300 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1607194113
transform 1 0 49588 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1064_
timestamp 1607194113
transform 1 0 49680 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1607194113
transform 1 0 48484 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_547
timestamp 1607194113
transform 1 0 51428 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_535
timestamp 1607194113
transform 1 0 50324 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_559
timestamp 1607194113
transform 1 0 52532 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_555
timestamp 1607194113
transform 1 0 52164 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1607194113
transform 1 0 52440 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_583
timestamp 1607194113
transform 1 0 54740 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_571
timestamp 1607194113
transform 1 0 53636 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_602
timestamp 1607194113
transform 1 0 56488 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_590
timestamp 1607194113
transform 1 0 55384 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1607194113
transform 1 0 55292 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_621
timestamp 1607194113
transform 1 0 58236 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_614
timestamp 1607194113
transform 1 0 57592 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1607194113
transform 1 0 58144 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_645
timestamp 1607194113
transform 1 0 60444 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_633
timestamp 1607194113
transform 1 0 59340 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_658
timestamp 1607194113
transform 1 0 61640 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_652
timestamp 1607194113
transform 1 0 61088 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1607194113
transform 1 0 60996 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1089_
timestamp 1607194113
transform 1 0 61732 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_76_683
timestamp 1607194113
transform 1 0 63940 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_670
timestamp 1607194113
transform 1 0 62744 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A
timestamp 1607194113
transform 1 0 62560 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1607194113
transform 1 0 63848 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_695
timestamp 1607194113
transform 1 0 65044 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_726
timestamp 1607194113
transform 1 0 67896 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_714
timestamp 1607194113
transform 1 0 66792 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_707
timestamp 1607194113
transform 1 0 66148 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1607194113
transform 1 0 66700 0 -1 44064
box -38 -48 130 592
use delayline_9_hs  inst_idelay_line
timestamp 1607276359
transform 1 0 57776 0 1 3761
box 800 801 23264 27367
use sky130_fd_sc_hd__fill_2  FILLER_59_745
timestamp 1607194113
transform 1 0 69644 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_733
timestamp 1607194113
transform 1 0 68540 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__CLK
timestamp 1607194113
transform 1 0 69828 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1450_
timestamp 1607194113
transform 1 0 70012 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_59_768
timestamp 1607194113
transform 1 0 71760 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_791
timestamp 1607194113
transform 1 0 73876 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_779
timestamp 1607194113
transform 1 0 72772 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1607194113
transform 1 0 72312 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1607194113
transform 1 0 72496 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_806
timestamp 1607194113
transform 1 0 75256 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_794
timestamp 1607194113
transform 1 0 74152 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607194113
transform 1 0 74060 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_814
timestamp 1607194113
transform 1 0 75992 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__CLK
timestamp 1607194113
transform 1 0 76176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1456_
timestamp 1607194113
transform 1 0 76360 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_59_849
timestamp 1607194113
transform 1 0 79212 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_837
timestamp 1607194113
transform 1 0 78108 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_864
timestamp 1607194113
transform 1 0 80592 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_853
timestamp 1607194113
transform 1 0 79580 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1607194113
transform 1 0 80408 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607194113
transform 1 0 79672 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1607194113
transform 1 0 81144 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1043_
timestamp 1607194113
transform 1 0 79764 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_59_884
timestamp 1607194113
transform 1 0 82432 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_873
timestamp 1607194113
transform 1 0 81420 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1607194113
transform 1 0 82156 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_911
timestamp 1607194113
transform 1 0 84916 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_899
timestamp 1607194113
transform 1 0 83812 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1141_
timestamp 1607194113
transform 1 0 83168 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_59_916
timestamp 1607194113
transform 1 0 85376 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__CLK
timestamp 1607194113
transform 1 0 85560 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607194113
transform 1 0 85284 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1607194113
transform 1 0 85744 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_950
timestamp 1607194113
transform 1 0 88504 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[5]
timestamp 1607194113
transform 1 0 88044 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[4]
timestamp 1607194113
transform 1 0 87860 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[2]
timestamp 1607194113
transform 1 0 87676 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[0]
timestamp 1607194113
transform 1 0 87492 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1607194113
transform 1 0 88228 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_962
timestamp 1607194113
transform 1 0 89608 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_974
timestamp 1607194113
transform 1 0 90712 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607194113
transform 1 0 90896 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_742
timestamp 1607194113
transform 1 0 69368 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_736
timestamp 1607194113
transform 1 0 68816 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1607194113
transform 1 0 69184 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1155_
timestamp 1607194113
transform 1 0 69920 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1607194113
transform 1 0 68908 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_764
timestamp 1607194113
transform 1 0 71392 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_759
timestamp 1607194113
transform 1 0 70932 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1607194113
transform 1 0 70748 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__B
timestamp 1607194113
transform 1 0 70564 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607194113
transform 1 0 71300 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1156_
timestamp 1607194113
transform 1 0 71668 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_788
timestamp 1607194113
transform 1 0 73600 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_776
timestamp 1607194113
transform 1 0 72496 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_800
timestamp 1607194113
transform 1 0 74704 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_831
timestamp 1607194113
transform 1 0 77556 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_818
timestamp 1607194113
transform 1 0 76360 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_812
timestamp 1607194113
transform 1 0 75808 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1607194113
transform 1 0 76176 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1607194113
transform 1 0 77372 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607194113
transform 1 0 76912 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1607194113
transform 1 0 75900 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0734_
timestamp 1607194113
transform 1 0 77004 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_850
timestamp 1607194113
transform 1 0 79304 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A
timestamp 1607194113
transform 1 0 78292 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1142_
timestamp 1607194113
transform 1 0 78476 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_867
timestamp 1607194113
transform 1 0 80868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _1143_
timestamp 1607194113
transform 1 0 80040 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_886
timestamp 1607194113
transform 1 0 82616 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_879
timestamp 1607194113
transform 1 0 81972 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B
timestamp 1607194113
transform 1 0 82984 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607194113
transform 1 0 82524 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_901
timestamp 1607194113
transform 1 0 83996 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1607194113
transform 1 0 83168 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1146_
timestamp 1607194113
transform 1 0 84732 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1137_
timestamp 1607194113
transform 1 0 83352 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_60_918
timestamp 1607194113
transform 1 0 85560 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[7]
timestamp 1607194113
transform 1 0 85928 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[6]
timestamp 1607194113
transform 1 0 86112 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_inp_i
timestamp 1607194113
transform 1 0 86664 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1607194113
transform 1 0 86296 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_950
timestamp 1607194113
transform 1 0 88504 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_938
timestamp 1607194113
transform 1 0 87400 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[8]
timestamp 1607194113
transform 1 0 86848 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[3]
timestamp 1607194113
transform 1 0 87216 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[1]
timestamp 1607194113
transform 1 0 87032 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607194113
transform 1 0 88136 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1607194113
transform 1 0 88228 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_962
timestamp 1607194113
transform 1 0 89608 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_974
timestamp 1607194113
transform 1 0 90712 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_736
timestamp 1607194113
transform 1 0 68816 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_748
timestamp 1607194113
transform 1 0 69920 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_733
timestamp 1607194113
transform 1 0 68540 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__CLK
timestamp 1607194113
transform 1 0 70104 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A
timestamp 1607194113
transform 1 0 69736 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B
timestamp 1607194113
transform 1 0 69552 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1607194113
transform 1 0 70288 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1157_
timestamp 1607194113
transform 1 0 68908 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1149_
timestamp 1607194113
transform 1 0 69920 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_62_770
timestamp 1607194113
transform 1 0 71944 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_764
timestamp 1607194113
transform 1 0 71392 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_757
timestamp 1607194113
transform 1 0 70748 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_771
timestamp 1607194113
transform 1 0 72036 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__CLK
timestamp 1607194113
transform 1 0 72036 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A
timestamp 1607194113
transform 1 0 70564 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607194113
transform 1 0 71300 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_792
timestamp 1607194113
transform 1 0 73968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_791
timestamp 1607194113
transform 1 0 73876 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_783
timestamp 1607194113
transform 1 0 73140 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1451_
timestamp 1607194113
transform 1 0 72220 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0700_
timestamp 1607194113
transform 1 0 72772 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_804
timestamp 1607194113
transform 1 0 75072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_806
timestamp 1607194113
transform 1 0 75256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_794
timestamp 1607194113
transform 1 0 74152 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607194113
transform 1 0 74060 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_825
timestamp 1607194113
transform 1 0 77004 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_816
timestamp 1607194113
transform 1 0 76176 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_818
timestamp 1607194113
transform 1 0 76360 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__CLK
timestamp 1607194113
transform 1 0 77096 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1607194113
transform 1 0 77096 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607194113
transform 1 0 76912 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1457_
timestamp 1607194113
transform 1 0 77280 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1140_
timestamp 1607194113
transform 1 0 77280 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_847
timestamp 1607194113
transform 1 0 79028 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_848
timestamp 1607194113
transform 1 0 79120 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_840
timestamp 1607194113
transform 1 0 78384 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__D
timestamp 1607194113
transform 1 0 79396 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B
timestamp 1607194113
transform 1 0 79212 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_862
timestamp 1607194113
transform 1 0 80408 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_866
timestamp 1607194113
transform 1 0 80776 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_853
timestamp 1607194113
transform 1 0 79580 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1607194113
transform 1 0 80592 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607194113
transform 1 0 79672 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1138_
timestamp 1607194113
transform 1 0 79764 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1047_
timestamp 1607194113
transform 1 0 79764 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_62_874
timestamp 1607194113
transform 1 0 81512 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_878
timestamp 1607194113
transform 1 0 81880 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_886
timestamp 1607194113
transform 1 0 82616 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_882
timestamp 1607194113
transform 1 0 82248 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B1
timestamp 1607194113
transform 1 0 82708 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A2
timestamp 1607194113
transform 1 0 82892 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1607194113
transform 1 0 82524 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607194113
transform 1 0 82524 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0738_
timestamp 1607194113
transform 1 0 82156 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0726_
timestamp 1607194113
transform 1 0 82800 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A1
timestamp 1607194113
transform 1 0 83076 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_907
timestamp 1607194113
transform 1 0 84548 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_894
timestamp 1607194113
transform 1 0 83352 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_907
timestamp 1607194113
transform 1 0 84548 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1607194113
transform 1 0 83720 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1607194113
transform 1 0 83168 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1147_
timestamp 1607194113
transform 1 0 83260 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _1130_
timestamp 1607194113
transform 1 0 83904 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_62_923
timestamp 1607194113
transform 1 0 86020 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_915
timestamp 1607194113
transform 1 0 85284 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_925
timestamp 1607194113
transform 1 0 86204 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1607194113
transform 1 0 86020 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607194113
transform 1 0 85284 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1145_
timestamp 1607194113
transform 1 0 85376 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1133_
timestamp 1607194113
transform 1 0 85376 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_947
timestamp 1607194113
transform 1 0 88228 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_943
timestamp 1607194113
transform 1 0 87860 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_935
timestamp 1607194113
transform 1 0 87124 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__CLK
timestamp 1607194113
transform 1 0 86940 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607194113
transform 1 0 88136 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1607194113
transform 1 0 87124 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0729_
timestamp 1607194113
transform 1 0 86756 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_959
timestamp 1607194113
transform 1 0 89332 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_966
timestamp 1607194113
transform 1 0 89976 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_954
timestamp 1607194113
transform 1 0 88872 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_971
timestamp 1607194113
transform 1 0 90436 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_974
timestamp 1607194113
transform 1 0 90712 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607194113
transform 1 0 90896 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_739
timestamp 1607194113
transform 1 0 69092 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_733
timestamp 1607194113
transform 1 0 68540 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1607194113
transform 1 0 68908 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1154_
timestamp 1607194113
transform 1 0 69644 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1607194113
transform 1 0 68632 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_754
timestamp 1607194113
transform 1 0 70472 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 1607194113
transform 1 0 71024 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1607194113
transform 1 0 72036 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1046_
timestamp 1607194113
transform 1 0 71208 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_63_790
timestamp 1607194113
transform 1 0 73784 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_782
timestamp 1607194113
transform 1 0 73048 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_773
timestamp 1607194113
transform 1 0 72220 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1607194113
transform 1 0 72772 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_806
timestamp 1607194113
transform 1 0 75256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_794
timestamp 1607194113
transform 1 0 74152 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1607194113
transform 1 0 74060 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_818
timestamp 1607194113
transform 1 0 76360 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B1
timestamp 1607194113
transform 1 0 76912 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1607194113
transform 1 0 77096 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1139_
timestamp 1607194113
transform 1 0 77280 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_63_841
timestamp 1607194113
transform 1 0 78476 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_867
timestamp 1607194113
transform 1 0 80868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_855
timestamp 1607194113
transform 1 0 79764 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_853
timestamp 1607194113
transform 1 0 79580 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1607194113
transform 1 0 79672 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_884
timestamp 1607194113
transform 1 0 82432 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_879
timestamp 1607194113
transform 1 0 81972 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B1
timestamp 1607194113
transform 1 0 82800 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A1
timestamp 1607194113
transform 1 0 82984 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1607194113
transform 1 0 82156 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_906
timestamp 1607194113
transform 1 0 84456 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1135_
timestamp 1607194113
transform 1 0 83168 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_63_925
timestamp 1607194113
transform 1 0 86204 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_914
timestamp 1607194113
transform 1 0 85192 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1607194113
transform 1 0 86020 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1607194113
transform 1 0 85284 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1132_
timestamp 1607194113
transform 1 0 85376 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__CLK
timestamp 1607194113
transform 1 0 86940 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1459_
timestamp 1607194113
transform 1 0 87124 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_63_966
timestamp 1607194113
transform 1 0 89976 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_954
timestamp 1607194113
transform 1 0 88872 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_974
timestamp 1607194113
transform 1 0 90712 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1607194113
transform 1 0 90896 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_741
timestamp 1607194113
transform 1 0 69276 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_733
timestamp 1607194113
transform 1 0 68540 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1152_
timestamp 1607194113
transform 1 0 69460 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_755
timestamp 1607194113
transform 1 0 70564 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1607194113
transform 1 0 71116 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1607194113
transform 1 0 71300 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1153_
timestamp 1607194113
transform 1 0 71392 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_785
timestamp 1607194113
transform 1 0 73324 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_773
timestamp 1607194113
transform 1 0 72220 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_810
timestamp 1607194113
transform 1 0 75624 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_805
timestamp 1607194113
transform 1 0 75164 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_797
timestamp 1607194113
transform 1 0 74428 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1117_
timestamp 1607194113
transform 1 0 75256 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_822
timestamp 1607194113
transform 1 0 76728 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1607194113
transform 1 0 76912 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1120_
timestamp 1607194113
transform 1 0 77004 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_845
timestamp 1607194113
transform 1 0 78844 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_834
timestamp 1607194113
transform 1 0 77832 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1607194113
transform 1 0 78568 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_869
timestamp 1607194113
transform 1 0 81052 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_857
timestamp 1607194113
transform 1 0 79948 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_886
timestamp 1607194113
transform 1 0 82616 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_877
timestamp 1607194113
transform 1 0 81788 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_873
timestamp 1607194113
transform 1 0 81420 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__CLK
timestamp 1607194113
transform 1 0 82892 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1607194113
transform 1 0 82524 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1458_
timestamp 1607194113
transform 1 0 83076 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1607194113
transform 1 0 81512 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_910
timestamp 1607194113
transform 1 0 84824 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _1134_
timestamp 1607194113
transform 1 0 85928 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_947
timestamp 1607194113
transform 1 0 88228 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_943
timestamp 1607194113
transform 1 0 87860 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_931
timestamp 1607194113
transform 1 0 86756 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1607194113
transform 1 0 88136 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_959
timestamp 1607194113
transform 1 0 89332 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_971
timestamp 1607194113
transform 1 0 90436 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_733
timestamp 1607194113
transform 1 0 68540 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__CLK
timestamp 1607194113
transform 1 0 69092 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1607194113
transform 1 0 69276 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_65_760
timestamp 1607194113
transform 1 0 71024 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1607194113
transform 1 0 71576 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1150_
timestamp 1607194113
transform 1 0 71760 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_65_787
timestamp 1607194113
transform 1 0 73508 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_775
timestamp 1607194113
transform 1 0 72404 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_806
timestamp 1607194113
transform 1 0 75256 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_794
timestamp 1607194113
transform 1 0 74152 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1607194113
transform 1 0 74060 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1607194113
transform 1 0 75624 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_815
timestamp 1607194113
transform 1 0 76084 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__CLK
timestamp 1607194113
transform 1 0 76452 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1607194113
transform 1 0 75900 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1463_
timestamp 1607194113
transform 1 0 76636 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_840
timestamp 1607194113
transform 1 0 78384 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_867
timestamp 1607194113
transform 1 0 80868 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_855
timestamp 1607194113
transform 1 0 79764 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_852
timestamp 1607194113
transform 1 0 79488 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1607194113
transform 1 0 79672 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_890
timestamp 1607194113
transform 1 0 82984 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_879
timestamp 1607194113
transform 1 0 81972 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1607194113
transform 1 0 82708 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_903
timestamp 1607194113
transform 1 0 84180 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1607194113
transform 1 0 83996 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1607194113
transform 1 0 83720 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_925
timestamp 1607194113
transform 1 0 86204 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1607194113
transform 1 0 86020 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1607194113
transform 1 0 85284 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1125_
timestamp 1607194113
transform 1 0 85376 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_65_946
timestamp 1607194113
transform 1 0 88136 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_934
timestamp 1607194113
transform 1 0 87032 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1607194113
transform 1 0 86756 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_970
timestamp 1607194113
transform 1 0 90344 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_958
timestamp 1607194113
transform 1 0 89240 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1607194113
transform 1 0 90896 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_739
timestamp 1607194113
transform 1 0 69092 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B1
timestamp 1607194113
transform 1 0 69184 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1151_
timestamp 1607194113
transform 1 0 69368 0 -1 38624
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_66_768
timestamp 1607194113
transform 1 0 71760 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_755
timestamp 1607194113
transform 1 0 70564 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1607194113
transform 1 0 71300 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1607194113
transform 1 0 71392 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_792
timestamp 1607194113
transform 1 0 73968 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_780
timestamp 1607194113
transform 1 0 72864 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_801
timestamp 1607194113
transform 1 0 74796 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1607194113
transform 1 0 74520 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1114_
timestamp 1607194113
transform 1 0 75532 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1607194113
transform 1 0 76360 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__C
timestamp 1607194113
transform 1 0 76544 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1607194113
transform 1 0 76728 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1607194113
transform 1 0 76176 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1607194113
transform 1 0 76912 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1110_
timestamp 1607194113
transform 1 0 77004 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_849
timestamp 1607194113
transform 1 0 79212 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_834
timestamp 1607194113
transform 1 0 77832 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1607194113
transform 1 0 78384 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1119_
timestamp 1607194113
transform 1 0 78568 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_66_861
timestamp 1607194113
transform 1 0 80316 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_886
timestamp 1607194113
transform 1 0 82616 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_873
timestamp 1607194113
transform 1 0 81420 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1607194113
transform 1 0 82524 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_905
timestamp 1607194113
transform 1 0 84364 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1607194113
transform 1 0 83352 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1108_
timestamp 1607194113
transform 1 0 83536 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_928
timestamp 1607194113
transform 1 0 86480 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_917
timestamp 1607194113
transform 1 0 85468 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1127_
timestamp 1607194113
transform 1 0 85652 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_947
timestamp 1607194113
transform 1 0 88228 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_940
timestamp 1607194113
transform 1 0 87584 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1607194113
transform 1 0 88136 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_959
timestamp 1607194113
transform 1 0 89332 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_971
timestamp 1607194113
transform 1 0 90436 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_749
timestamp 1607194113
transform 1 0 70012 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_739
timestamp 1607194113
transform 1 0 69092 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1607194113
transform 1 0 68908 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1607194113
transform 1 0 69460 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1466_
timestamp 1607194113
transform 1 0 68632 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1607194113
transform 1 0 69644 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0722_
timestamp 1607194113
transform 1 0 68540 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_767
timestamp 1607194113
transform 1 0 71668 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_761
timestamp 1607194113
transform 1 0 71116 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_753
timestamp 1607194113
transform 1 0 70380 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_761
timestamp 1607194113
transform 1 0 71116 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1607194113
transform 1 0 71300 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1607194113
transform 1 0 71392 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1607194113
transform 1 0 70748 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_791
timestamp 1607194113
transform 1 0 73876 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_779
timestamp 1607194113
transform 1 0 72772 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_790
timestamp 1607194113
transform 1 0 73784 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_778
timestamp 1607194113
transform 1 0 72680 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1607194113
transform 1 0 72496 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1607194113
transform 1 0 72220 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_811
timestamp 1607194113
transform 1 0 75716 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_803
timestamp 1607194113
transform 1 0 74980 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_794
timestamp 1607194113
transform 1 0 74152 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1607194113
transform 1 0 74888 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1607194113
transform 1 0 74060 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1115_
timestamp 1607194113
transform 1 0 75072 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_68_816
timestamp 1607194113
transform 1 0 76176 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_821
timestamp 1607194113
transform 1 0 76636 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_813
timestamp 1607194113
transform 1 0 75900 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0744_
timestamp 1607194113
transform 1 0 75808 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B1
timestamp 1607194113
transform 1 0 76728 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B
timestamp 1607194113
transform 1 0 76728 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A1
timestamp 1607194113
transform 1 0 76912 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1607194113
transform 1 0 77004 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1607194113
transform 1 0 76912 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1041_
timestamp 1607194113
transform 1 0 77188 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1121_
timestamp 1607194113
transform 1 0 77096 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_68_846
timestamp 1607194113
transform 1 0 78936 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_838
timestamp 1607194113
transform 1 0 78200 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_840
timestamp 1607194113
transform 1 0 78384 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__D
timestamp 1607194113
transform 1 0 78016 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1048_
timestamp 1607194113
transform 1 0 79120 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_68_857
timestamp 1607194113
transform 1 0 79948 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_852
timestamp 1607194113
transform 1 0 79488 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1607194113
transform 1 0 79672 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1040_
timestamp 1607194113
transform 1 0 79764 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1607194113
transform 1 0 80960 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__C
timestamp 1607194113
transform 1 0 80776 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__D
timestamp 1607194113
transform 1 0 80592 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1607194113
transform 1 0 80684 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_868
timestamp 1607194113
transform 1 0 80960 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_870
timestamp 1607194113
transform 1 0 81144 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_886
timestamp 1607194113
transform 1 0 82616 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_884
timestamp 1607194113
transform 1 0 82432 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_880
timestamp 1607194113
transform 1 0 82064 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_882
timestamp 1607194113
transform 1 0 82248 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1607194113
transform 1 0 82524 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_908
timestamp 1607194113
transform 1 0 84640 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_894
timestamp 1607194113
transform 1 0 83352 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B1
timestamp 1607194113
transform 1 0 83352 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1607194113
transform 1 0 83444 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A1
timestamp 1607194113
transform 1 0 83536 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B
timestamp 1607194113
transform 1 0 84456 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1128_
timestamp 1607194113
transform 1 0 83720 0 -1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_4  _1109_
timestamp 1607194113
transform 1 0 83628 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_68_912
timestamp 1607194113
transform 1 0 85008 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_919
timestamp 1607194113
transform 1 0 85652 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_914
timestamp 1607194113
transform 1 0 85192 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1607194113
transform 1 0 85560 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1607194113
transform 1 0 85284 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1607194113
transform 1 0 85376 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1123_
timestamp 1607194113
transform 1 0 85744 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_67_925
timestamp 1607194113
transform 1 0 86204 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__CLK
timestamp 1607194113
transform 1 0 86296 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_927
timestamp 1607194113
transform 1 0 86388 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1461_
timestamp 1607194113
transform 1 0 86480 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_947
timestamp 1607194113
transform 1 0 88228 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_945
timestamp 1607194113
transform 1 0 88044 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_939
timestamp 1607194113
transform 1 0 87492 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_947
timestamp 1607194113
transform 1 0 88228 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1607194113
transform 1 0 88136 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_959
timestamp 1607194113
transform 1 0 89332 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_959
timestamp 1607194113
transform 1 0 89332 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_971
timestamp 1607194113
transform 1 0 90436 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_975
timestamp 1607194113
transform 1 0 90804 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_971
timestamp 1607194113
transform 1 0 90436 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1607194113
transform 1 0 90896 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_739
timestamp 1607194113
transform 1 0 69092 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_733
timestamp 1607194113
transform 1 0 68540 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A1
timestamp 1607194113
transform 1 0 69184 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1106_
timestamp 1607194113
transform 1 0 69368 0 1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_69_768
timestamp 1607194113
transform 1 0 71760 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_760
timestamp 1607194113
transform 1 0 71024 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B1
timestamp 1607194113
transform 1 0 70840 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A2
timestamp 1607194113
transform 1 0 70656 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1607194113
transform 1 0 71392 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_790
timestamp 1607194113
transform 1 0 73784 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_784
timestamp 1607194113
transform 1 0 73232 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A
timestamp 1607194113
transform 1 0 73876 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1087_
timestamp 1607194113
transform 1 0 72864 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_811
timestamp 1607194113
transform 1 0 75716 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_803
timestamp 1607194113
transform 1 0 74980 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1607194113
transform 1 0 74060 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1116_
timestamp 1607194113
transform 1 0 74152 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_69_830
timestamp 1607194113
transform 1 0 77464 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_817
timestamp 1607194113
transform 1 0 76268 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1607194113
transform 1 0 76084 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1607194113
transform 1 0 76636 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1113_
timestamp 1607194113
transform 1 0 76820 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1607194113
transform 1 0 75808 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_844
timestamp 1607194113
transform 1 0 78752 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1607194113
transform 1 0 78568 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0709_
timestamp 1607194113
transform 1 0 78200 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_860
timestamp 1607194113
transform 1 0 80224 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_855
timestamp 1607194113
transform 1 0 79764 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_852
timestamp 1607194113
transform 1 0 79488 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1607194113
transform 1 0 79672 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1607194113
transform 1 0 79948 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_884
timestamp 1607194113
transform 1 0 82432 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_872
timestamp 1607194113
transform 1 0 81328 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_902
timestamp 1607194113
transform 1 0 84088 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_896
timestamp 1607194113
transform 1 0 83536 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1607194113
transform 1 0 83812 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_925
timestamp 1607194113
transform 1 0 86204 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_914
timestamp 1607194113
transform 1 0 85192 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1607194113
transform 1 0 86020 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1607194113
transform 1 0 85284 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1126_
timestamp 1607194113
transform 1 0 85376 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_69_949
timestamp 1607194113
transform 1 0 88412 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_937
timestamp 1607194113
transform 1 0 87308 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_961
timestamp 1607194113
transform 1 0 89516 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_973
timestamp 1607194113
transform 1 0 90620 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1607194113
transform 1 0 90896 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_736
timestamp 1607194113
transform 1 0 68816 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B
timestamp 1607194113
transform 1 0 70196 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1607194113
transform 1 0 69368 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1095_
timestamp 1607194113
transform 1 0 69552 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_70_767
timestamp 1607194113
transform 1 0 71668 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_761
timestamp 1607194113
transform 1 0 71116 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_753
timestamp 1607194113
transform 1 0 70380 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1607194113
transform 1 0 71300 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1607194113
transform 1 0 71392 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__CLK
timestamp 1607194113
transform 1 0 72404 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1464_
timestamp 1607194113
transform 1 0 72588 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_808
timestamp 1607194113
transform 1 0 75440 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_796
timestamp 1607194113
transform 1 0 74336 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_820
timestamp 1607194113
transform 1 0 76544 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1607194113
transform 1 0 76912 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1112_
timestamp 1607194113
transform 1 0 77004 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_839
timestamp 1607194113
transform 1 0 78292 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__CLK
timestamp 1607194113
transform 1 0 78660 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1607194113
transform 1 0 78108 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1462_
timestamp 1607194113
transform 1 0 78844 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_864
timestamp 1607194113
transform 1 0 80592 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_886
timestamp 1607194113
transform 1 0 82616 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_884
timestamp 1607194113
transform 1 0 82432 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_876
timestamp 1607194113
transform 1 0 81696 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1607194113
transform 1 0 82524 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__CLK
timestamp 1607194113
transform 1 0 83168 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1460_
timestamp 1607194113
transform 1 0 83352 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_925
timestamp 1607194113
transform 1 0 86204 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_913
timestamp 1607194113
transform 1 0 85100 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_947
timestamp 1607194113
transform 1 0 88228 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_945
timestamp 1607194113
transform 1 0 88044 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_937
timestamp 1607194113
transform 1 0 87308 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1607194113
transform 1 0 88136 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_959
timestamp 1607194113
transform 1 0 89332 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_971
timestamp 1607194113
transform 1 0 90436 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_750
timestamp 1607194113
transform 1 0 70104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_742
timestamp 1607194113
transform 1 0 69368 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1035_
timestamp 1607194113
transform 1 0 68540 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_71_764
timestamp 1607194113
transform 1 0 71392 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1607194113
transform 1 0 71208 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1607194113
transform 1 0 71760 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1104_
timestamp 1607194113
transform 1 0 70380 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1103_
timestamp 1607194113
transform 1 0 71944 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_71_789
timestamp 1607194113
transform 1 0 73692 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_777
timestamp 1607194113
transform 1 0 72588 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_806
timestamp 1607194113
transform 1 0 75256 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_794
timestamp 1607194113
transform 1 0 74152 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1607194113
transform 1 0 74060 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_818
timestamp 1607194113
transform 1 0 76360 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1607194113
transform 1 0 76912 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1111_
timestamp 1607194113
transform 1 0 77096 0 1 40800
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_71_841
timestamp 1607194113
transform 1 0 78476 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A1
timestamp 1607194113
transform 1 0 78292 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_870
timestamp 1607194113
transform 1 0 81144 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_858
timestamp 1607194113
transform 1 0 80040 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_853
timestamp 1607194113
transform 1 0 79580 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1607194113
transform 1 0 79672 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1607194113
transform 1 0 79764 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_882
timestamp 1607194113
transform 1 0 82248 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_906
timestamp 1607194113
transform 1 0 84456 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_894
timestamp 1607194113
transform 1 0 83352 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_928
timestamp 1607194113
transform 1 0 86480 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_916
timestamp 1607194113
transform 1 0 85376 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_914
timestamp 1607194113
transform 1 0 85192 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1607194113
transform 1 0 85284 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_940
timestamp 1607194113
transform 1 0 87584 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_964
timestamp 1607194113
transform 1 0 89792 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_952
timestamp 1607194113
transform 1 0 88688 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1607194113
transform 1 0 90896 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_739
timestamp 1607194113
transform 1 0 69092 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1096_
timestamp 1607194113
transform 1 0 69828 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_72_768
timestamp 1607194113
transform 1 0 71760 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_762
timestamp 1607194113
transform 1 0 71208 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_754
timestamp 1607194113
transform 1 0 70472 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1607194113
transform 1 0 71300 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0748_
timestamp 1607194113
transform 1 0 71392 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_792
timestamp 1607194113
transform 1 0 73968 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_780
timestamp 1607194113
transform 1 0 72864 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_804
timestamp 1607194113
transform 1 0 75072 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_825
timestamp 1607194113
transform 1 0 77004 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_816
timestamp 1607194113
transform 1 0 76176 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1607194113
transform 1 0 76912 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__CLK
timestamp 1607194113
transform 1 0 77740 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1465_
timestamp 1607194113
transform 1 0 77924 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_72_866
timestamp 1607194113
transform 1 0 80776 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_854
timestamp 1607194113
transform 1 0 79672 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_886
timestamp 1607194113
transform 1 0 82616 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_884
timestamp 1607194113
transform 1 0 82432 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_878
timestamp 1607194113
transform 1 0 81880 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1607194113
transform 1 0 82524 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_910
timestamp 1607194113
transform 1 0 84824 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_898
timestamp 1607194113
transform 1 0 83720 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_922
timestamp 1607194113
transform 1 0 85928 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_947
timestamp 1607194113
transform 1 0 88228 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_934
timestamp 1607194113
transform 1 0 87032 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1607194113
transform 1 0 88136 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_959
timestamp 1607194113
transform 1 0 89332 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_971
timestamp 1607194113
transform 1 0 90436 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_749
timestamp 1607194113
transform 1 0 70012 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_739
timestamp 1607194113
transform 1 0 69092 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_733
timestamp 1607194113
transform 1 0 68540 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1100_
timestamp 1607194113
transform 1 0 69184 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_73_755
timestamp 1607194113
transform 1 0 70564 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__CLK
timestamp 1607194113
transform 1 0 70656 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1467_
timestamp 1607194113
transform 1 0 70840 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_73_789
timestamp 1607194113
transform 1 0 73692 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_777
timestamp 1607194113
transform 1 0 72588 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_806
timestamp 1607194113
transform 1 0 75256 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_794
timestamp 1607194113
transform 1 0 74152 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1607194113
transform 1 0 74060 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_830
timestamp 1607194113
transform 1 0 77464 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_818
timestamp 1607194113
transform 1 0 76360 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_842
timestamp 1607194113
transform 1 0 78568 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_867
timestamp 1607194113
transform 1 0 80868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_855
timestamp 1607194113
transform 1 0 79764 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1607194113
transform 1 0 79672 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_891
timestamp 1607194113
transform 1 0 83076 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_879
timestamp 1607194113
transform 1 0 81972 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_903
timestamp 1607194113
transform 1 0 84180 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_928
timestamp 1607194113
transform 1 0 86480 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_916
timestamp 1607194113
transform 1 0 85376 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1607194113
transform 1 0 85284 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_940
timestamp 1607194113
transform 1 0 87584 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_964
timestamp 1607194113
transform 1 0 89792 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_952
timestamp 1607194113
transform 1 0 88688 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1607194113
transform 1 0 90896 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_733
timestamp 1607194113
transform 1 0 68540 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_749
timestamp 1607194113
transform 1 0 70012 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_736
timestamp 1607194113
transform 1 0 68816 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__CLK
timestamp 1607194113
transform 1 0 68908 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A
timestamp 1607194113
transform 1 0 69828 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1468_
timestamp 1607194113
transform 1 0 69092 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1101_
timestamp 1607194113
transform 1 0 69000 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_770
timestamp 1607194113
transform 1 0 71944 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_758
timestamp 1607194113
transform 1 0 70840 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_767
timestamp 1607194113
transform 1 0 71668 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_761
timestamp 1607194113
transform 1 0 71116 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1607194113
transform 1 0 71300 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1607194113
transform 1 0 71392 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_790
timestamp 1607194113
transform 1 0 73784 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_782
timestamp 1607194113
transform 1 0 73048 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_791
timestamp 1607194113
transform 1 0 73876 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_779
timestamp 1607194113
transform 1 0 72772 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_806
timestamp 1607194113
transform 1 0 75256 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_794
timestamp 1607194113
transform 1 0 74152 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_803
timestamp 1607194113
transform 1 0 74980 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1607194113
transform 1 0 74060 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_830
timestamp 1607194113
transform 1 0 77464 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_818
timestamp 1607194113
transform 1 0 76360 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_825
timestamp 1607194113
transform 1 0 77004 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_823
timestamp 1607194113
transform 1 0 76820 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_815
timestamp 1607194113
transform 1 0 76084 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1607194113
transform 1 0 76912 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_842
timestamp 1607194113
transform 1 0 78568 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_849
timestamp 1607194113
transform 1 0 79212 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_837
timestamp 1607194113
transform 1 0 78108 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_867
timestamp 1607194113
transform 1 0 80868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_855
timestamp 1607194113
transform 1 0 79764 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_861
timestamp 1607194113
transform 1 0 80316 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1607194113
transform 1 0 79672 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_891
timestamp 1607194113
transform 1 0 83076 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_879
timestamp 1607194113
transform 1 0 81972 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_886
timestamp 1607194113
transform 1 0 82616 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_873
timestamp 1607194113
transform 1 0 81420 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1607194113
transform 1 0 82524 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_903
timestamp 1607194113
transform 1 0 84180 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_910
timestamp 1607194113
transform 1 0 84824 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_898
timestamp 1607194113
transform 1 0 83720 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_928
timestamp 1607194113
transform 1 0 86480 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_916
timestamp 1607194113
transform 1 0 85376 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_922
timestamp 1607194113
transform 1 0 85928 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1607194113
transform 1 0 85284 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_940
timestamp 1607194113
transform 1 0 87584 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_947
timestamp 1607194113
transform 1 0 88228 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_934
timestamp 1607194113
transform 1 0 87032 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1607194113
transform 1 0 88136 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_964
timestamp 1607194113
transform 1 0 89792 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_952
timestamp 1607194113
transform 1 0 88688 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_959
timestamp 1607194113
transform 1 0 89332 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_971
timestamp 1607194113
transform 1 0 90436 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1607194113
transform 1 0 90896 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_750
timestamp 1607194113
transform 1 0 70104 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_738
timestamp 1607194113
transform 1 0 69000 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1607194113
transform 1 0 69920 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1607194113
transform 1 0 69552 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1607194113
transform 1 0 69644 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_762
timestamp 1607194113
transform 1 0 71208 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_788
timestamp 1607194113
transform 1 0 73600 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_776
timestamp 1607194113
transform 1 0 72496 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_774
timestamp 1607194113
transform 1 0 72312 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1607194113
transform 1 0 72404 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_807
timestamp 1607194113
transform 1 0 75348 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_800
timestamp 1607194113
transform 1 0 74704 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1607194113
transform 1 0 75256 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_831
timestamp 1607194113
transform 1 0 77556 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_819
timestamp 1607194113
transform 1 0 76452 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_850
timestamp 1607194113
transform 1 0 79304 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_838
timestamp 1607194113
transform 1 0 78200 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1607194113
transform 1 0 78108 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_869
timestamp 1607194113
transform 1 0 81052 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_862
timestamp 1607194113
transform 1 0 80408 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1607194113
transform 1 0 80960 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_881
timestamp 1607194113
transform 1 0 82156 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_900
timestamp 1607194113
transform 1 0 83904 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_893
timestamp 1607194113
transform 1 0 83260 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1607194113
transform 1 0 83812 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_924
timestamp 1607194113
transform 1 0 86112 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_912
timestamp 1607194113
transform 1 0 85008 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1607194113
transform 1 0 86664 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_943
timestamp 1607194113
transform 1 0 87860 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_931
timestamp 1607194113
transform 1 0 86756 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_962
timestamp 1607194113
transform 1 0 89608 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_955
timestamp 1607194113
transform 1 0 88964 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1607194113
transform 1 0 89516 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_974
timestamp 1607194113
transform 1 0 90712 0 -1 44064
box -38 -48 1142 592
use delayline_9_hs  inst_rdelay_line
timestamp 1607276359
transform 1 0 85560 0 1 3761
box 800 801 23264 27367
use sky130_fd_sc_hd__decap_12  FILLER_60_986
timestamp 1607194113
transform 1 0 91816 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_989
timestamp 1607194113
transform 1 0 92092 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_977
timestamp 1607194113
transform 1 0 90988 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1008
timestamp 1607194113
transform 1 0 93840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1006
timestamp 1607194113
transform 1 0 93656 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_998
timestamp 1607194113
transform 1 0 92920 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1001
timestamp 1607194113
transform 1 0 93196 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607194113
transform 1 0 93748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1020
timestamp 1607194113
transform 1 0 94944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1025
timestamp 1607194113
transform 1 0 95404 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1013
timestamp 1607194113
transform 1 0 94300 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1032
timestamp 1607194113
transform 1 0 96048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1038
timestamp 1607194113
transform 1 0 96600 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607194113
transform 1 0 96508 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1056
timestamp 1607194113
transform 1 0 98256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1044
timestamp 1607194113
transform 1 0 97152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1050
timestamp 1607194113
transform 1 0 97704 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1069
timestamp 1607194113
transform 1 0 99452 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1074
timestamp 1607194113
transform 1 0 99912 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1062
timestamp 1607194113
transform 1 0 98808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607194113
transform 1 0 99360 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1081
timestamp 1607194113
transform 1 0 100556 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1086
timestamp 1607194113
transform 1 0 101016 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1105
timestamp 1607194113
transform 1 0 102764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1093
timestamp 1607194113
transform 1 0 101660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1099
timestamp 1607194113
transform 1 0 102212 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607194113
transform 1 0 102120 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1117
timestamp 1607194113
transform 1 0 103868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1123
timestamp 1607194113
transform 1 0 104420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1111
timestamp 1607194113
transform 1 0 103316 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1130
timestamp 1607194113
transform 1 0 105064 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1135
timestamp 1607194113
transform 1 0 105524 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607194113
transform 1 0 104972 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1154
timestamp 1607194113
transform 1 0 107272 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1142
timestamp 1607194113
transform 1 0 106168 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1147
timestamp 1607194113
transform 1 0 106628 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1166
timestamp 1607194113
transform 1 0 108376 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1160
timestamp 1607194113
transform 1 0 107824 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607194113
transform 1 0 107732 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1178
timestamp 1607194113
transform 1 0 109480 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1184
timestamp 1607194113
transform 1 0 110032 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1172
timestamp 1607194113
transform 1 0 108928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_1191
timestamp 1607194113
transform 1 0 110676 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1192
timestamp 1607194113
transform 1 0 110768 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607194113
transform 1 0 110584 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1607194113
transform -1 0 111136 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1607194113
transform -1 0 111136 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_989
timestamp 1607194113
transform 1 0 92092 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_977
timestamp 1607194113
transform 1 0 90988 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_983
timestamp 1607194113
transform 1 0 91540 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_989
timestamp 1607194113
transform 1 0 92092 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_977
timestamp 1607194113
transform 1 0 90988 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1001
timestamp 1607194113
transform 1 0 93196 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1008
timestamp 1607194113
transform 1 0 93840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_995
timestamp 1607194113
transform 1 0 92644 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1001
timestamp 1607194113
transform 1 0 93196 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607194113
transform 1 0 93748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1025
timestamp 1607194113
transform 1 0 95404 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1013
timestamp 1607194113
transform 1 0 94300 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1020
timestamp 1607194113
transform 1 0 94944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1025
timestamp 1607194113
transform 1 0 95404 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1013
timestamp 1607194113
transform 1 0 94300 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1038
timestamp 1607194113
transform 1 0 96600 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1032
timestamp 1607194113
transform 1 0 96048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1038
timestamp 1607194113
transform 1 0 96600 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1607194113
transform 1 0 96508 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607194113
transform 1 0 96508 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1050
timestamp 1607194113
transform 1 0 97704 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1056
timestamp 1607194113
transform 1 0 98256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1044
timestamp 1607194113
transform 1 0 97152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1050
timestamp 1607194113
transform 1 0 97704 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1074
timestamp 1607194113
transform 1 0 99912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1062
timestamp 1607194113
transform 1 0 98808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1069
timestamp 1607194113
transform 1 0 99452 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1074
timestamp 1607194113
transform 1 0 99912 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1062
timestamp 1607194113
transform 1 0 98808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607194113
transform 1 0 99360 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1086
timestamp 1607194113
transform 1 0 101016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1081
timestamp 1607194113
transform 1 0 100556 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1086
timestamp 1607194113
transform 1 0 101016 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1099
timestamp 1607194113
transform 1 0 102212 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1105
timestamp 1607194113
transform 1 0 102764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1093
timestamp 1607194113
transform 1 0 101660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1099
timestamp 1607194113
transform 1 0 102212 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1607194113
transform 1 0 102120 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607194113
transform 1 0 102120 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1123
timestamp 1607194113
transform 1 0 104420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1111
timestamp 1607194113
transform 1 0 103316 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1117
timestamp 1607194113
transform 1 0 103868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1123
timestamp 1607194113
transform 1 0 104420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1111
timestamp 1607194113
transform 1 0 103316 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1135
timestamp 1607194113
transform 1 0 105524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1130
timestamp 1607194113
transform 1 0 105064 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1135
timestamp 1607194113
transform 1 0 105524 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607194113
transform 1 0 104972 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1147
timestamp 1607194113
transform 1 0 106628 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1154
timestamp 1607194113
transform 1 0 107272 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1142
timestamp 1607194113
transform 1 0 106168 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1147
timestamp 1607194113
transform 1 0 106628 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1160
timestamp 1607194113
transform 1 0 107824 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1166
timestamp 1607194113
transform 1 0 108376 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1160
timestamp 1607194113
transform 1 0 107824 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1607194113
transform 1 0 107732 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607194113
transform 1 0 107732 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1184
timestamp 1607194113
transform 1 0 110032 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1172
timestamp 1607194113
transform 1 0 108928 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1178
timestamp 1607194113
transform 1 0 109480 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1184
timestamp 1607194113
transform 1 0 110032 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1172
timestamp 1607194113
transform 1 0 108928 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1192
timestamp 1607194113
transform 1 0 110768 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_1191
timestamp 1607194113
transform 1 0 110676 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1192
timestamp 1607194113
transform 1 0 110768 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607194113
transform 1 0 110584 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1607194113
transform -1 0 111136 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1607194113
transform -1 0 111136 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1607194113
transform -1 0 111136 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_989
timestamp 1607194113
transform 1 0 92092 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_977
timestamp 1607194113
transform 1 0 90988 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_983
timestamp 1607194113
transform 1 0 91540 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1001
timestamp 1607194113
transform 1 0 93196 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1008
timestamp 1607194113
transform 1 0 93840 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_995
timestamp 1607194113
transform 1 0 92644 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1607194113
transform 1 0 93748 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1025
timestamp 1607194113
transform 1 0 95404 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1013
timestamp 1607194113
transform 1 0 94300 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1020
timestamp 1607194113
transform 1 0 94944 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1038
timestamp 1607194113
transform 1 0 96600 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1032
timestamp 1607194113
transform 1 0 96048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1607194113
transform 1 0 96508 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1050
timestamp 1607194113
transform 1 0 97704 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1056
timestamp 1607194113
transform 1 0 98256 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1044
timestamp 1607194113
transform 1 0 97152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1074
timestamp 1607194113
transform 1 0 99912 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1062
timestamp 1607194113
transform 1 0 98808 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1069
timestamp 1607194113
transform 1 0 99452 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1607194113
transform 1 0 99360 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1086
timestamp 1607194113
transform 1 0 101016 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1081
timestamp 1607194113
transform 1 0 100556 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1099
timestamp 1607194113
transform 1 0 102212 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1105
timestamp 1607194113
transform 1 0 102764 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1093
timestamp 1607194113
transform 1 0 101660 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1607194113
transform 1 0 102120 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1123
timestamp 1607194113
transform 1 0 104420 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1111
timestamp 1607194113
transform 1 0 103316 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1117
timestamp 1607194113
transform 1 0 103868 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1135
timestamp 1607194113
transform 1 0 105524 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1130
timestamp 1607194113
transform 1 0 105064 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1607194113
transform 1 0 104972 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1147
timestamp 1607194113
transform 1 0 106628 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1154
timestamp 1607194113
transform 1 0 107272 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1142
timestamp 1607194113
transform 1 0 106168 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1160
timestamp 1607194113
transform 1 0 107824 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1166
timestamp 1607194113
transform 1 0 108376 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1607194113
transform 1 0 107732 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1184
timestamp 1607194113
transform 1 0 110032 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1172
timestamp 1607194113
transform 1 0 108928 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1178
timestamp 1607194113
transform 1 0 109480 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1192
timestamp 1607194113
transform 1 0 110768 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1191
timestamp 1607194113
transform 1 0 110676 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1607194113
transform 1 0 110584 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1607194113
transform -1 0 111136 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1607194113
transform -1 0 111136 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_983
timestamp 1607194113
transform 1 0 91540 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_989
timestamp 1607194113
transform 1 0 92092 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_977
timestamp 1607194113
transform 1 0 90988 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_983
timestamp 1607194113
transform 1 0 91540 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1008
timestamp 1607194113
transform 1 0 93840 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_995
timestamp 1607194113
transform 1 0 92644 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1001
timestamp 1607194113
transform 1 0 93196 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1008
timestamp 1607194113
transform 1 0 93840 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_995
timestamp 1607194113
transform 1 0 92644 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1607194113
transform 1 0 93748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1607194113
transform 1 0 93748 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1020
timestamp 1607194113
transform 1 0 94944 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1025
timestamp 1607194113
transform 1 0 95404 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1013
timestamp 1607194113
transform 1 0 94300 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1020
timestamp 1607194113
transform 1 0 94944 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1032
timestamp 1607194113
transform 1 0 96048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1038
timestamp 1607194113
transform 1 0 96600 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1032
timestamp 1607194113
transform 1 0 96048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1607194113
transform 1 0 96508 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1056
timestamp 1607194113
transform 1 0 98256 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1044
timestamp 1607194113
transform 1 0 97152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1050
timestamp 1607194113
transform 1 0 97704 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1056
timestamp 1607194113
transform 1 0 98256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1044
timestamp 1607194113
transform 1 0 97152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1069
timestamp 1607194113
transform 1 0 99452 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1074
timestamp 1607194113
transform 1 0 99912 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1062
timestamp 1607194113
transform 1 0 98808 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1069
timestamp 1607194113
transform 1 0 99452 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1607194113
transform 1 0 99360 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1607194113
transform 1 0 99360 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1081
timestamp 1607194113
transform 1 0 100556 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1086
timestamp 1607194113
transform 1 0 101016 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1081
timestamp 1607194113
transform 1 0 100556 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1105
timestamp 1607194113
transform 1 0 102764 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1093
timestamp 1607194113
transform 1 0 101660 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1099
timestamp 1607194113
transform 1 0 102212 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1105
timestamp 1607194113
transform 1 0 102764 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1093
timestamp 1607194113
transform 1 0 101660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1607194113
transform 1 0 102120 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1117
timestamp 1607194113
transform 1 0 103868 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1123
timestamp 1607194113
transform 1 0 104420 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1111
timestamp 1607194113
transform 1 0 103316 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1117
timestamp 1607194113
transform 1 0 103868 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1130
timestamp 1607194113
transform 1 0 105064 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1135
timestamp 1607194113
transform 1 0 105524 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1130
timestamp 1607194113
transform 1 0 105064 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1607194113
transform 1 0 104972 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1607194113
transform 1 0 104972 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1154
timestamp 1607194113
transform 1 0 107272 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1142
timestamp 1607194113
transform 1 0 106168 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1147
timestamp 1607194113
transform 1 0 106628 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1154
timestamp 1607194113
transform 1 0 107272 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1142
timestamp 1607194113
transform 1 0 106168 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1166
timestamp 1607194113
transform 1 0 108376 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1160
timestamp 1607194113
transform 1 0 107824 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1166
timestamp 1607194113
transform 1 0 108376 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1607194113
transform 1 0 107732 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1178
timestamp 1607194113
transform 1 0 109480 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1184
timestamp 1607194113
transform 1 0 110032 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1172
timestamp 1607194113
transform 1 0 108928 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1178
timestamp 1607194113
transform 1 0 109480 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_1191
timestamp 1607194113
transform 1 0 110676 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1192
timestamp 1607194113
transform 1 0 110768 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_1191
timestamp 1607194113
transform 1 0 110676 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1607194113
transform 1 0 110584 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1607194113
transform 1 0 110584 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1607194113
transform -1 0 111136 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1607194113
transform -1 0 111136 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1607194113
transform -1 0 111136 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_989
timestamp 1607194113
transform 1 0 92092 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_977
timestamp 1607194113
transform 1 0 90988 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_983
timestamp 1607194113
transform 1 0 91540 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_989
timestamp 1607194113
transform 1 0 92092 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_977
timestamp 1607194113
transform 1 0 90988 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1001
timestamp 1607194113
transform 1 0 93196 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1008
timestamp 1607194113
transform 1 0 93840 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_995
timestamp 1607194113
transform 1 0 92644 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1001
timestamp 1607194113
transform 1 0 93196 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1607194113
transform 1 0 93748 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1025
timestamp 1607194113
transform 1 0 95404 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1013
timestamp 1607194113
transform 1 0 94300 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1020
timestamp 1607194113
transform 1 0 94944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1025
timestamp 1607194113
transform 1 0 95404 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1013
timestamp 1607194113
transform 1 0 94300 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1038
timestamp 1607194113
transform 1 0 96600 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1032
timestamp 1607194113
transform 1 0 96048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1038
timestamp 1607194113
transform 1 0 96600 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1607194113
transform 1 0 96508 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1607194113
transform 1 0 96508 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1050
timestamp 1607194113
transform 1 0 97704 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1056
timestamp 1607194113
transform 1 0 98256 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1044
timestamp 1607194113
transform 1 0 97152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1050
timestamp 1607194113
transform 1 0 97704 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1074
timestamp 1607194113
transform 1 0 99912 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1062
timestamp 1607194113
transform 1 0 98808 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1069
timestamp 1607194113
transform 1 0 99452 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1074
timestamp 1607194113
transform 1 0 99912 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1062
timestamp 1607194113
transform 1 0 98808 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1607194113
transform 1 0 99360 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1086
timestamp 1607194113
transform 1 0 101016 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1081
timestamp 1607194113
transform 1 0 100556 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1086
timestamp 1607194113
transform 1 0 101016 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1099
timestamp 1607194113
transform 1 0 102212 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1105
timestamp 1607194113
transform 1 0 102764 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1093
timestamp 1607194113
transform 1 0 101660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1099
timestamp 1607194113
transform 1 0 102212 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1607194113
transform 1 0 102120 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1607194113
transform 1 0 102120 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1123
timestamp 1607194113
transform 1 0 104420 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1111
timestamp 1607194113
transform 1 0 103316 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1117
timestamp 1607194113
transform 1 0 103868 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1123
timestamp 1607194113
transform 1 0 104420 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1111
timestamp 1607194113
transform 1 0 103316 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1135
timestamp 1607194113
transform 1 0 105524 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1130
timestamp 1607194113
transform 1 0 105064 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1135
timestamp 1607194113
transform 1 0 105524 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1607194113
transform 1 0 104972 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1147
timestamp 1607194113
transform 1 0 106628 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1154
timestamp 1607194113
transform 1 0 107272 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1142
timestamp 1607194113
transform 1 0 106168 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1147
timestamp 1607194113
transform 1 0 106628 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1160
timestamp 1607194113
transform 1 0 107824 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1166
timestamp 1607194113
transform 1 0 108376 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1160
timestamp 1607194113
transform 1 0 107824 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1607194113
transform 1 0 107732 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1607194113
transform 1 0 107732 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_1184
timestamp 1607194113
transform 1 0 110032 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1172
timestamp 1607194113
transform 1 0 108928 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1178
timestamp 1607194113
transform 1 0 109480 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_1184
timestamp 1607194113
transform 1 0 110032 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1172
timestamp 1607194113
transform 1 0 108928 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_1192
timestamp 1607194113
transform 1 0 110768 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_1191
timestamp 1607194113
transform 1 0 110676 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_1192
timestamp 1607194113
transform 1 0 110768 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1607194113
transform 1 0 110584 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1607194113
transform -1 0 111136 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1607194113
transform -1 0 111136 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1607194113
transform -1 0 111136 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_983
timestamp 1607194113
transform 1 0 91540 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_989
timestamp 1607194113
transform 1 0 92092 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_977
timestamp 1607194113
transform 1 0 90988 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_983
timestamp 1607194113
transform 1 0 91540 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1008
timestamp 1607194113
transform 1 0 93840 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_995
timestamp 1607194113
transform 1 0 92644 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1001
timestamp 1607194113
transform 1 0 93196 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1008
timestamp 1607194113
transform 1 0 93840 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_995
timestamp 1607194113
transform 1 0 92644 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1607194113
transform 1 0 93748 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1607194113
transform 1 0 93748 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1020
timestamp 1607194113
transform 1 0 94944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1025
timestamp 1607194113
transform 1 0 95404 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1013
timestamp 1607194113
transform 1 0 94300 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1020
timestamp 1607194113
transform 1 0 94944 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1032
timestamp 1607194113
transform 1 0 96048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1038
timestamp 1607194113
transform 1 0 96600 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1032
timestamp 1607194113
transform 1 0 96048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1607194113
transform 1 0 96508 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1056
timestamp 1607194113
transform 1 0 98256 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1044
timestamp 1607194113
transform 1 0 97152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1050
timestamp 1607194113
transform 1 0 97704 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1056
timestamp 1607194113
transform 1 0 98256 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1044
timestamp 1607194113
transform 1 0 97152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1069
timestamp 1607194113
transform 1 0 99452 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1074
timestamp 1607194113
transform 1 0 99912 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1062
timestamp 1607194113
transform 1 0 98808 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1069
timestamp 1607194113
transform 1 0 99452 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1607194113
transform 1 0 99360 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1607194113
transform 1 0 99360 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1081
timestamp 1607194113
transform 1 0 100556 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1086
timestamp 1607194113
transform 1 0 101016 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1081
timestamp 1607194113
transform 1 0 100556 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1105
timestamp 1607194113
transform 1 0 102764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1093
timestamp 1607194113
transform 1 0 101660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1099
timestamp 1607194113
transform 1 0 102212 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1105
timestamp 1607194113
transform 1 0 102764 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1093
timestamp 1607194113
transform 1 0 101660 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1607194113
transform 1 0 102120 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1117
timestamp 1607194113
transform 1 0 103868 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1123
timestamp 1607194113
transform 1 0 104420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1111
timestamp 1607194113
transform 1 0 103316 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1117
timestamp 1607194113
transform 1 0 103868 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1130
timestamp 1607194113
transform 1 0 105064 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1135
timestamp 1607194113
transform 1 0 105524 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1130
timestamp 1607194113
transform 1 0 105064 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1607194113
transform 1 0 104972 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1607194113
transform 1 0 104972 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1154
timestamp 1607194113
transform 1 0 107272 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1142
timestamp 1607194113
transform 1 0 106168 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1147
timestamp 1607194113
transform 1 0 106628 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1154
timestamp 1607194113
transform 1 0 107272 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1142
timestamp 1607194113
transform 1 0 106168 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1166
timestamp 1607194113
transform 1 0 108376 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1160
timestamp 1607194113
transform 1 0 107824 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1166
timestamp 1607194113
transform 1 0 108376 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1607194113
transform 1 0 107732 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1178
timestamp 1607194113
transform 1 0 109480 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_1184
timestamp 1607194113
transform 1 0 110032 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1172
timestamp 1607194113
transform 1 0 108928 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1178
timestamp 1607194113
transform 1 0 109480 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_1191
timestamp 1607194113
transform 1 0 110676 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_1192
timestamp 1607194113
transform 1 0 110768 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_1191
timestamp 1607194113
transform 1 0 110676 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1607194113
transform 1 0 110584 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1607194113
transform 1 0 110584 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1607194113
transform -1 0 111136 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1607194113
transform -1 0 111136 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1607194113
transform -1 0 111136 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_986
timestamp 1607194113
transform 1 0 91816 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_989
timestamp 1607194113
transform 1 0 92092 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_977
timestamp 1607194113
transform 1 0 90988 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1607194113
transform 1 0 92368 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1005
timestamp 1607194113
transform 1 0 93564 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_993
timestamp 1607194113
transform 1 0 92460 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1001
timestamp 1607194113
transform 1 0 93196 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1024
timestamp 1607194113
transform 1 0 95312 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1017
timestamp 1607194113
transform 1 0 94668 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1025
timestamp 1607194113
transform 1 0 95404 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1013
timestamp 1607194113
transform 1 0 94300 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1607194113
transform 1 0 95220 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1036
timestamp 1607194113
transform 1 0 96416 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1038
timestamp 1607194113
transform 1 0 96600 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1607194113
transform 1 0 96508 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1055
timestamp 1607194113
transform 1 0 98164 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1048
timestamp 1607194113
transform 1 0 97520 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1050
timestamp 1607194113
transform 1 0 97704 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1607194113
transform 1 0 98072 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1067
timestamp 1607194113
transform 1 0 99268 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1074
timestamp 1607194113
transform 1 0 99912 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1062
timestamp 1607194113
transform 1 0 98808 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1086
timestamp 1607194113
transform 1 0 101016 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1079
timestamp 1607194113
transform 1 0 100372 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1086
timestamp 1607194113
transform 1 0 101016 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1607194113
transform 1 0 100924 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1098
timestamp 1607194113
transform 1 0 102120 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1099
timestamp 1607194113
transform 1 0 102212 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1607194113
transform 1 0 102120 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1117
timestamp 1607194113
transform 1 0 103868 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1110
timestamp 1607194113
transform 1 0 103224 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1123
timestamp 1607194113
transform 1 0 104420 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1111
timestamp 1607194113
transform 1 0 103316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1607194113
transform 1 0 103776 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1129
timestamp 1607194113
transform 1 0 104972 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1135
timestamp 1607194113
transform 1 0 105524 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1148
timestamp 1607194113
transform 1 0 106720 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1141
timestamp 1607194113
transform 1 0 106076 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1147
timestamp 1607194113
transform 1 0 106628 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1607194113
transform 1 0 106628 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1160
timestamp 1607194113
transform 1 0 107824 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1160
timestamp 1607194113
transform 1 0 107824 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1607194113
transform 1 0 107732 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1179
timestamp 1607194113
transform 1 0 109572 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1172
timestamp 1607194113
transform 1 0 108928 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1184
timestamp 1607194113
transform 1 0 110032 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1172
timestamp 1607194113
transform 1 0 108928 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1607194113
transform 1 0 109480 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_1191
timestamp 1607194113
transform 1 0 110676 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_1192
timestamp 1607194113
transform 1 0 110768 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1607194113
transform -1 0 111136 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1607194113
transform -1 0 111136 0 1 42976
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 280 800 400 6 bus_in[0]
port 0 nsew default input
rlabel metal3 s 0 12248 800 12368 6 bus_in[10]
port 1 nsew default input
rlabel metal3 s 0 13472 800 13592 6 bus_in[11]
port 2 nsew default input
rlabel metal3 s 0 14560 800 14680 6 bus_in[12]
port 3 nsew default input
rlabel metal3 s 0 15784 800 15904 6 bus_in[13]
port 4 nsew default input
rlabel metal3 s 0 17008 800 17128 6 bus_in[14]
port 5 nsew default input
rlabel metal3 s 0 18232 800 18352 6 bus_in[15]
port 6 nsew default input
rlabel metal3 s 0 19456 800 19576 6 bus_in[16]
port 7 nsew default input
rlabel metal3 s 0 20680 800 20800 6 bus_in[17]
port 8 nsew default input
rlabel metal3 s 0 21768 800 21888 6 bus_in[18]
port 9 nsew default input
rlabel metal3 s 0 22992 800 23112 6 bus_in[19]
port 10 nsew default input
rlabel metal3 s 0 1368 800 1488 6 bus_in[1]
port 11 nsew default input
rlabel metal3 s 0 24216 800 24336 6 bus_in[20]
port 12 nsew default input
rlabel metal3 s 0 25440 800 25560 6 bus_in[21]
port 13 nsew default input
rlabel metal3 s 0 26664 800 26784 6 bus_in[22]
port 14 nsew default input
rlabel metal3 s 0 27888 800 28008 6 bus_in[23]
port 15 nsew default input
rlabel metal3 s 0 28976 800 29096 6 bus_in[24]
port 16 nsew default input
rlabel metal3 s 0 30200 800 30320 6 bus_in[25]
port 17 nsew default input
rlabel metal3 s 0 31424 800 31544 6 bus_in[26]
port 18 nsew default input
rlabel metal3 s 0 32648 800 32768 6 bus_in[27]
port 19 nsew default input
rlabel metal3 s 0 33872 800 33992 6 bus_in[28]
port 20 nsew default input
rlabel metal3 s 0 35096 800 35216 6 bus_in[29]
port 21 nsew default input
rlabel metal3 s 0 2592 800 2712 6 bus_in[2]
port 22 nsew default input
rlabel metal3 s 0 36184 800 36304 6 bus_in[30]
port 23 nsew default input
rlabel metal3 s 0 37408 800 37528 6 bus_in[31]
port 24 nsew default input
rlabel metal3 s 0 38632 800 38752 6 bus_in[32]
port 25 nsew default input
rlabel metal3 s 0 39856 800 39976 6 bus_in[33]
port 26 nsew default input
rlabel metal3 s 0 41080 800 41200 6 bus_in[34]
port 27 nsew default input
rlabel metal3 s 0 42304 800 42424 6 bus_in[35]
port 28 nsew default input
rlabel metal3 s 0 42848 800 42968 6 bus_in[36]
port 29 nsew default input
rlabel metal3 s 0 43392 800 43512 6 bus_in[37]
port 30 nsew default input
rlabel metal3 s 0 44072 800 44192 6 bus_in[38]
port 31 nsew default input
rlabel metal3 s 0 44616 800 44736 6 bus_in[39]
port 32 nsew default input
rlabel metal3 s 0 3816 800 3936 6 bus_in[3]
port 33 nsew default input
rlabel metal3 s 0 45296 800 45416 6 bus_in[40]
port 34 nsew default input
rlabel metal3 s 0 45840 800 45960 6 bus_in[41]
port 35 nsew default input
rlabel metal3 s 0 5040 800 5160 6 bus_in[4]
port 36 nsew default input
rlabel metal3 s 0 6264 800 6384 6 bus_in[5]
port 37 nsew default input
rlabel metal3 s 0 7352 800 7472 6 bus_in[6]
port 38 nsew default input
rlabel metal3 s 0 8576 800 8696 6 bus_in[7]
port 39 nsew default input
rlabel metal3 s 0 9800 800 9920 6 bus_in[8]
port 40 nsew default input
rlabel metal3 s 0 11024 800 11144 6 bus_in[9]
port 41 nsew default input
rlabel metal3 s 0 824 800 944 6 bus_out[0]
port 42 nsew default tristate
rlabel metal3 s 0 12792 800 12912 6 bus_out[10]
port 43 nsew default tristate
rlabel metal3 s 0 14016 800 14136 6 bus_out[11]
port 44 nsew default tristate
rlabel metal3 s 0 15240 800 15360 6 bus_out[12]
port 45 nsew default tristate
rlabel metal3 s 0 16464 800 16584 6 bus_out[13]
port 46 nsew default tristate
rlabel metal3 s 0 17688 800 17808 6 bus_out[14]
port 47 nsew default tristate
rlabel metal3 s 0 18776 800 18896 6 bus_out[15]
port 48 nsew default tristate
rlabel metal3 s 0 20000 800 20120 6 bus_out[16]
port 49 nsew default tristate
rlabel metal3 s 0 21224 800 21344 6 bus_out[17]
port 50 nsew default tristate
rlabel metal3 s 0 22448 800 22568 6 bus_out[18]
port 51 nsew default tristate
rlabel metal3 s 0 23672 800 23792 6 bus_out[19]
port 52 nsew default tristate
rlabel metal3 s 0 2048 800 2168 6 bus_out[1]
port 53 nsew default tristate
rlabel metal3 s 0 24896 800 25016 6 bus_out[20]
port 54 nsew default tristate
rlabel metal3 s 0 25984 800 26104 6 bus_out[21]
port 55 nsew default tristate
rlabel metal3 s 0 27208 800 27328 6 bus_out[22]
port 56 nsew default tristate
rlabel metal3 s 0 28432 800 28552 6 bus_out[23]
port 57 nsew default tristate
rlabel metal3 s 0 29656 800 29776 6 bus_out[24]
port 58 nsew default tristate
rlabel metal3 s 0 30880 800 31000 6 bus_out[25]
port 59 nsew default tristate
rlabel metal3 s 0 32104 800 32224 6 bus_out[26]
port 60 nsew default tristate
rlabel metal3 s 0 33192 800 33312 6 bus_out[27]
port 61 nsew default tristate
rlabel metal3 s 0 34416 800 34536 6 bus_out[28]
port 62 nsew default tristate
rlabel metal3 s 0 35640 800 35760 6 bus_out[29]
port 63 nsew default tristate
rlabel metal3 s 0 3272 800 3392 6 bus_out[2]
port 64 nsew default tristate
rlabel metal3 s 0 36864 800 36984 6 bus_out[30]
port 65 nsew default tristate
rlabel metal3 s 0 38088 800 38208 6 bus_out[31]
port 66 nsew default tristate
rlabel metal3 s 0 39312 800 39432 6 bus_out[32]
port 67 nsew default tristate
rlabel metal3 s 0 40400 800 40520 6 bus_out[33]
port 68 nsew default tristate
rlabel metal3 s 0 41624 800 41744 6 bus_out[34]
port 69 nsew default tristate
rlabel metal3 s 0 4360 800 4480 6 bus_out[3]
port 70 nsew default tristate
rlabel metal3 s 0 5584 800 5704 6 bus_out[4]
port 71 nsew default tristate
rlabel metal3 s 0 6808 800 6928 6 bus_out[5]
port 72 nsew default tristate
rlabel metal3 s 0 8032 800 8152 6 bus_out[6]
port 73 nsew default tristate
rlabel metal3 s 0 9256 800 9376 6 bus_out[7]
port 74 nsew default tristate
rlabel metal3 s 0 10480 800 10600 6 bus_out[8]
port 75 nsew default tristate
rlabel metal3 s 0 11568 800 11688 6 bus_out[9]
port 76 nsew default tristate
rlabel metal2 s 28078 0 28134 800 6 clk_i
port 77 nsew default input
rlabel metal2 s 84198 0 84254 800 6 out1_o
port 78 nsew default tristate
rlabel metal3 s 111440 23128 112240 23248 6 out2_o
port 79 nsew default tristate
rlabel metal2 s 56138 45440 56194 46240 6 rst_n_i
port 80 nsew default input
rlabel metal5 s 1104 6436 111136 7036 6 VPWR
port 81 nsew default input
rlabel metal5 s 1104 24436 111136 25036 6 VGND
port 82 nsew default input
<< properties >>
string FIXED_BBOX 0 0 112240 46240
<< end >>
