magic
tech sky130A
magscale 1 2
timestamp 1607276668
<< locali >>
rect 78951 39879 78985 40049
rect 45371 37703 45405 37805
rect 31939 37227 31973 37465
rect 39207 37227 39241 37329
rect 62391 36615 62425 36921
rect 76007 36751 76041 36921
rect 62391 35187 62425 35289
rect 26051 34575 26085 34745
rect 36999 33895 37033 34133
rect 57515 33555 57549 33657
rect 57055 32807 57089 32909
rect 77019 32807 77053 32909
rect 82631 32875 82665 33113
rect 86035 32263 86069 32501
rect 15287 31379 15321 31481
rect 52271 30631 52305 30801
rect 62207 30087 62241 30393
rect 23107 29203 23141 29305
rect 61195 28455 61229 28693
rect 56135 28047 56169 28149
rect 32951 26823 32985 27061
rect 9031 24647 9065 24885
rect 21543 24647 21577 24681
rect 21485 24613 21577 24647
rect 33963 23355 33997 23729
rect 33963 21723 33997 22573
rect 40403 20431 40437 20601
<< viali >>
rect 66071 41613 66105 41647
rect 66255 41613 66289 41647
rect 66531 41613 66565 41647
rect 88887 41613 88921 41647
rect 89071 41613 89105 41647
rect 89347 41613 89381 41647
rect 67635 41477 67669 41511
rect 90451 41477 90485 41511
rect 3051 41273 3085 41307
rect 3511 41273 3545 41307
rect 18875 41273 18909 41307
rect 24487 41273 24521 41307
rect 27155 41273 27189 41307
rect 30283 41273 30317 41307
rect 48683 41273 48717 41307
rect 52731 41273 52765 41307
rect 74995 41273 75029 41307
rect 82631 41273 82665 41307
rect 1947 41137 1981 41171
rect 5259 41137 5293 41171
rect 6547 41137 6581 41171
rect 12067 41137 12101 41171
rect 23383 41137 23417 41171
rect 24947 41137 24981 41171
rect 43071 41137 43105 41171
rect 54479 41137 54513 41171
rect 55767 41137 55801 41171
rect 57055 41137 57089 41171
rect 60091 41137 60125 41171
rect 61379 41137 61413 41171
rect 62667 41137 62701 41171
rect 80975 41137 81009 41171
rect 86771 41137 86805 41171
rect 1671 41069 1705 41103
rect 3603 41069 3637 41103
rect 4615 41069 4649 41103
rect 6271 41069 6305 41103
rect 12343 41069 12377 41103
rect 17495 41069 17529 41103
rect 17771 41069 17805 41103
rect 23107 41069 23141 41103
rect 25591 41069 25625 41103
rect 25867 41069 25901 41103
rect 28719 41069 28753 41103
rect 28995 41069 29029 41103
rect 32031 41069 32065 41103
rect 33135 41069 33169 41103
rect 33227 41069 33261 41103
rect 36355 41069 36389 41103
rect 37367 41069 37401 41103
rect 37735 41069 37769 41103
rect 38011 41069 38045 41103
rect 43255 41069 43289 41103
rect 43807 41069 43841 41103
rect 47119 41069 47153 41103
rect 47395 41069 47429 41103
rect 51167 41069 51201 41103
rect 51443 41069 51477 41103
rect 54663 41069 54697 41103
rect 55215 41069 55249 41103
rect 55399 41069 55433 41103
rect 56779 41069 56813 41103
rect 60275 41069 60309 41103
rect 60827 41069 60861 41103
rect 61011 41069 61045 41103
rect 62207 41069 62241 41103
rect 62391 41069 62425 41103
rect 73615 41069 73649 41103
rect 73891 41069 73925 41103
rect 80791 41069 80825 41103
rect 81067 41069 81101 41103
rect 81343 41069 81377 41103
rect 85391 41069 85425 41103
rect 85667 41069 85701 41103
rect 43991 41001 44025 41035
rect 7835 40933 7869 40967
rect 8019 40933 8053 40967
rect 13447 40933 13481 40967
rect 13907 40933 13941 40967
rect 17311 40933 17345 40967
rect 22923 40933 22957 40967
rect 27339 40933 27373 40967
rect 30467 40933 30501 40967
rect 32215 40933 32249 40967
rect 32951 40933 32985 40967
rect 36539 40933 36573 40967
rect 37551 40933 37585 40967
rect 48867 40933 48901 40967
rect 52915 40933 52949 40967
rect 56043 40933 56077 40967
rect 58159 40933 58193 40967
rect 58619 40933 58653 40967
rect 61655 40933 61689 40967
rect 63771 40933 63805 40967
rect 75455 40933 75489 40967
rect 85299 40933 85333 40967
rect 5443 40729 5477 40763
rect 28351 40729 28385 40763
rect 47211 40729 47245 40763
rect 81067 40729 81101 40763
rect 82355 40729 82389 40763
rect 88151 40729 88185 40763
rect 16759 40661 16793 40695
rect 28535 40661 28569 40695
rect 51351 40661 51385 40695
rect 57423 40661 57457 40695
rect 2407 40593 2441 40627
rect 3511 40593 3545 40627
rect 6731 40593 6765 40627
rect 8203 40593 8237 40627
rect 26787 40593 26821 40627
rect 31847 40593 31881 40627
rect 33503 40593 33537 40627
rect 35987 40593 36021 40627
rect 37459 40593 37493 40627
rect 38839 40593 38873 40627
rect 41323 40593 41357 40627
rect 43071 40593 43105 40627
rect 45463 40593 45497 40627
rect 49511 40593 49545 40627
rect 51167 40593 51201 40627
rect 55583 40593 55617 40627
rect 58067 40593 58101 40627
rect 61011 40593 61045 40627
rect 61103 40593 61137 40627
rect 63587 40593 63621 40627
rect 66531 40593 66565 40627
rect 68279 40593 68313 40627
rect 71131 40593 71165 40627
rect 78491 40593 78525 40627
rect 79871 40593 79905 40627
rect 80883 40593 80917 40627
rect 82079 40593 82113 40627
rect 82539 40593 82573 40627
rect 83827 40593 83861 40627
rect 83919 40593 83953 40627
rect 3787 40525 3821 40559
rect 4983 40525 5017 40559
rect 6455 40525 6489 40559
rect 11055 40525 11089 40559
rect 11331 40525 11365 40559
rect 14919 40525 14953 40559
rect 15195 40525 15229 40559
rect 17311 40525 17345 40559
rect 17403 40525 17437 40559
rect 17679 40525 17713 40559
rect 18783 40525 18817 40559
rect 20991 40525 21025 40559
rect 21267 40525 21301 40559
rect 22371 40525 22405 40559
rect 27063 40525 27097 40559
rect 32123 40525 32157 40559
rect 33595 40525 33629 40559
rect 34239 40525 34273 40559
rect 34331 40525 34365 40559
rect 34607 40525 34641 40559
rect 37183 40525 37217 40559
rect 39483 40525 39517 40559
rect 39667 40525 39701 40559
rect 39943 40525 39977 40559
rect 42611 40525 42645 40559
rect 42795 40525 42829 40559
rect 44175 40525 44209 40559
rect 45739 40525 45773 40559
rect 46843 40525 46877 40559
rect 49787 40525 49821 40559
rect 55859 40525 55893 40559
rect 58159 40525 58193 40559
rect 61379 40525 61413 40559
rect 63679 40525 63713 40559
rect 66807 40525 66841 40559
rect 70855 40525 70889 40559
rect 73339 40525 73373 40559
rect 73615 40525 73649 40559
rect 77939 40525 77973 40559
rect 78215 40525 78249 40559
rect 84195 40525 84229 40559
rect 88243 40525 88277 40559
rect 88519 40525 88553 40559
rect 90727 40525 90761 40559
rect 91003 40525 91037 40559
rect 92107 40525 92141 40559
rect 2499 40389 2533 40423
rect 5351 40389 5385 40423
rect 8019 40389 8053 40423
rect 12435 40389 12469 40423
rect 12895 40389 12929 40423
rect 16299 40389 16333 40423
rect 20899 40389 20933 40423
rect 36907 40389 36941 40423
rect 56963 40389 56997 40423
rect 62667 40389 62701 40423
rect 67911 40389 67945 40423
rect 72235 40389 72269 40423
rect 72695 40389 72729 40423
rect 74719 40389 74753 40423
rect 75179 40389 75213 40423
rect 78123 40389 78157 40423
rect 80699 40389 80733 40423
rect 85299 40389 85333 40423
rect 89623 40389 89657 40423
rect 90359 40389 90393 40423
rect 90543 40389 90577 40423
rect 12803 40185 12837 40219
rect 14183 40185 14217 40219
rect 20163 40185 20197 40219
rect 41599 40185 41633 40219
rect 46567 40185 46601 40219
rect 49327 40185 49361 40219
rect 55675 40185 55709 40219
rect 61103 40185 61137 40219
rect 82539 40185 82573 40219
rect 8111 40117 8145 40151
rect 21543 40117 21577 40151
rect 6363 40049 6397 40083
rect 6639 40049 6673 40083
rect 9123 40049 9157 40083
rect 12527 40049 12561 40083
rect 18691 40049 18725 40083
rect 18783 40049 18817 40083
rect 26143 40049 26177 40083
rect 27707 40049 27741 40083
rect 32399 40049 32433 40083
rect 41691 40049 41725 40083
rect 47211 40049 47245 40083
rect 50247 40049 50281 40083
rect 68555 40049 68589 40083
rect 75731 40049 75765 40083
rect 78031 40049 78065 40083
rect 78951 40049 78985 40083
rect 81435 40049 81469 40083
rect 89347 40049 89381 40083
rect 8847 39981 8881 40015
rect 10595 39981 10629 40015
rect 12619 39981 12653 40015
rect 13907 39981 13941 40015
rect 13999 39981 14033 40015
rect 19059 39981 19093 40015
rect 21635 39981 21669 40015
rect 25591 39981 25625 40015
rect 25959 39981 25993 40015
rect 27247 39981 27281 40015
rect 27431 39981 27465 40015
rect 28995 39981 29029 40015
rect 29271 39981 29305 40015
rect 31663 39981 31697 40015
rect 32123 39981 32157 40015
rect 37275 39981 37309 40015
rect 37551 39981 37585 40015
rect 41967 39981 42001 40015
rect 46751 39981 46785 40015
rect 47119 39981 47153 40015
rect 49511 39981 49545 40015
rect 50063 39981 50097 40015
rect 54663 39981 54697 40015
rect 54755 39981 54789 40015
rect 55215 39981 55249 40015
rect 55399 39981 55433 40015
rect 57147 39981 57181 40015
rect 59907 39981 59941 40015
rect 60091 39981 60125 40015
rect 60643 39981 60677 40015
rect 60827 39981 60861 40015
rect 62483 39981 62517 40015
rect 68279 39981 68313 40015
rect 68463 39981 68497 40015
rect 71315 39981 71349 40015
rect 71591 39981 71625 40015
rect 73615 39981 73649 40015
rect 74075 39981 74109 40015
rect 75915 39981 75949 40015
rect 76467 39981 76501 40015
rect 76651 39981 76685 40015
rect 77939 39981 77973 40015
rect 8019 39913 8053 39947
rect 10503 39913 10537 39947
rect 62575 39913 62609 39947
rect 77019 39913 77053 39947
rect 81067 39981 81101 40015
rect 81159 39981 81193 40015
rect 85391 39981 85425 40015
rect 85851 39981 85885 40015
rect 88611 39981 88645 40015
rect 89071 39981 89105 40015
rect 21819 39845 21853 39879
rect 28811 39845 28845 39879
rect 37091 39845 37125 39879
rect 37919 39845 37953 39879
rect 43071 39845 43105 39879
rect 57239 39845 57273 39879
rect 71131 39845 71165 39879
rect 73707 39845 73741 39879
rect 75179 39845 75213 39879
rect 75363 39845 75397 39879
rect 75547 39845 75581 39879
rect 78951 39845 78985 39879
rect 85667 39845 85701 39879
rect 4155 39641 4189 39675
rect 37367 39641 37401 39675
rect 41691 39641 41725 39675
rect 49511 39641 49545 39675
rect 49787 39641 49821 39675
rect 54479 39641 54513 39675
rect 55951 39641 55985 39675
rect 84195 39641 84229 39675
rect 88795 39641 88829 39675
rect 21635 39573 21669 39607
rect 32307 39573 32341 39607
rect 73339 39573 73373 39607
rect 77295 39573 77329 39607
rect 12159 39505 12193 39539
rect 12527 39505 12561 39539
rect 17311 39505 17345 39539
rect 17495 39505 17529 39539
rect 17587 39505 17621 39539
rect 21175 39505 21209 39539
rect 27339 39505 27373 39539
rect 27891 39505 27925 39539
rect 28075 39505 28109 39539
rect 31571 39505 31605 39539
rect 32031 39505 32065 39539
rect 33503 39505 33537 39539
rect 34055 39505 34089 39539
rect 34239 39505 34273 39539
rect 37183 39505 37217 39539
rect 40679 39505 40713 39539
rect 41231 39505 41265 39539
rect 41415 39505 41449 39539
rect 42795 39505 42829 39539
rect 49695 39505 49729 39539
rect 50247 39505 50281 39539
rect 54111 39505 54145 39539
rect 55031 39505 55065 39539
rect 55399 39505 55433 39539
rect 57055 39505 57089 39539
rect 68003 39505 68037 39539
rect 68279 39505 68313 39539
rect 70855 39505 70889 39539
rect 72879 39505 72913 39539
rect 73155 39505 73189 39539
rect 77387 39505 77421 39539
rect 77663 39505 77697 39539
rect 83919 39505 83953 39539
rect 84471 39505 84505 39539
rect 88703 39505 88737 39539
rect 89163 39505 89197 39539
rect 3511 39437 3545 39471
rect 11975 39437 12009 39471
rect 12435 39437 12469 39471
rect 21083 39437 21117 39471
rect 27247 39437 27281 39471
rect 33319 39437 33353 39471
rect 40587 39437 40621 39471
rect 42887 39437 42921 39471
rect 55123 39437 55157 39471
rect 55307 39437 55341 39471
rect 55767 39437 55801 39471
rect 65059 39437 65093 39471
rect 65243 39437 65277 39471
rect 65519 39437 65553 39471
rect 68187 39437 68221 39471
rect 21819 39369 21853 39403
rect 27063 39369 27097 39403
rect 28259 39369 28293 39403
rect 43163 39369 43197 39403
rect 56871 39369 56905 39403
rect 71039 39369 71073 39403
rect 11791 39301 11825 39335
rect 17771 39301 17805 39335
rect 18231 39301 18265 39335
rect 34515 39301 34549 39335
rect 34883 39301 34917 39335
rect 54203 39301 54237 39335
rect 66807 39301 66841 39335
rect 71315 39301 71349 39335
rect 78951 39301 78985 39335
rect 19151 39097 19185 39131
rect 20439 39097 20473 39131
rect 26879 39097 26913 39131
rect 32123 39097 32157 39131
rect 34699 39097 34733 39131
rect 42151 39097 42185 39131
rect 50891 39097 50925 39131
rect 54111 39097 54145 39131
rect 65335 39097 65369 39131
rect 68279 39097 68313 39131
rect 74075 39097 74109 39131
rect 76007 39097 76041 39131
rect 90175 39097 90209 39131
rect 33227 39029 33261 39063
rect 47211 39029 47245 39063
rect 2499 38961 2533 38995
rect 8571 38961 8605 38995
rect 9031 38961 9065 38995
rect 12251 38961 12285 38995
rect 16575 38961 16609 38995
rect 32583 38961 32617 38995
rect 35159 38961 35193 38995
rect 40863 38961 40897 38995
rect 41323 38961 41357 38995
rect 43071 38961 43105 38995
rect 45647 38961 45681 38995
rect 48131 38961 48165 38995
rect 51167 38961 51201 38995
rect 53927 38961 53961 38995
rect 55031 38961 55065 38995
rect 74535 38961 74569 38995
rect 76191 38961 76225 38995
rect 77479 38961 77513 38995
rect 79503 38961 79537 38995
rect 90451 38961 90485 38995
rect 2223 38893 2257 38927
rect 8755 38893 8789 38927
rect 9123 38893 9157 38927
rect 11975 38893 12009 38927
rect 13631 38893 13665 38927
rect 16207 38893 16241 38927
rect 18783 38893 18817 38927
rect 18967 38893 19001 38927
rect 19519 38893 19553 38927
rect 20255 38893 20289 38927
rect 27063 38893 27097 38927
rect 27247 38893 27281 38927
rect 27615 38893 27649 38927
rect 27799 38893 27833 38927
rect 32491 38893 32525 38927
rect 32859 38893 32893 38927
rect 33043 38893 33077 38927
rect 34883 38893 34917 38927
rect 41415 38893 41449 38927
rect 41783 38893 41817 38927
rect 41967 38893 42001 38927
rect 43163 38893 43197 38927
rect 43715 38893 43749 38927
rect 43899 38893 43933 38927
rect 45555 38893 45589 38927
rect 45923 38893 45957 38927
rect 47303 38893 47337 38927
rect 48039 38893 48073 38927
rect 51627 38893 51661 38927
rect 51811 38893 51845 38927
rect 52179 38893 52213 38927
rect 52271 38893 52305 38927
rect 54939 38893 54973 38927
rect 55307 38893 55341 38927
rect 55491 38893 55525 38927
rect 60275 38893 60309 38927
rect 60367 38893 60401 38927
rect 64139 38893 64173 38927
rect 64323 38893 64357 38927
rect 64783 38893 64817 38927
rect 64875 38893 64909 38927
rect 66807 38893 66841 38927
rect 68463 38893 68497 38927
rect 68647 38893 68681 38927
rect 69015 38893 69049 38927
rect 69107 38893 69141 38927
rect 74443 38893 74477 38927
rect 74811 38893 74845 38927
rect 74995 38893 75029 38927
rect 76375 38893 76409 38927
rect 76927 38893 76961 38927
rect 77111 38893 77145 38927
rect 79227 38893 79261 38927
rect 90727 38893 90761 38927
rect 3879 38825 3913 38859
rect 8111 38825 8145 38859
rect 16023 38825 16057 38859
rect 18875 38825 18909 38859
rect 36539 38825 36573 38859
rect 44267 38825 44301 38859
rect 54295 38825 54329 38859
rect 63863 38825 63897 38859
rect 64047 38825 64081 38859
rect 4063 38757 4097 38791
rect 8019 38757 8053 38791
rect 13815 38757 13849 38791
rect 33411 38757 33445 38791
rect 42335 38757 42369 38791
rect 47395 38757 47429 38791
rect 50707 38757 50741 38791
rect 60551 38757 60585 38791
rect 66899 38757 66933 38791
rect 69291 38757 69325 38791
rect 78951 38757 78985 38791
rect 80607 38757 80641 38791
rect 91831 38757 91865 38791
rect 2499 38553 2533 38587
rect 11883 38553 11917 38587
rect 29363 38553 29397 38587
rect 32859 38553 32893 38587
rect 33227 38553 33261 38587
rect 41415 38553 41449 38587
rect 48683 38553 48717 38587
rect 51259 38553 51293 38587
rect 54295 38553 54329 38587
rect 60275 38553 60309 38587
rect 63679 38553 63713 38587
rect 72511 38553 72545 38587
rect 80055 38553 80089 38587
rect 88795 38553 88829 38587
rect 90175 38553 90209 38587
rect 16759 38485 16793 38519
rect 23475 38485 23509 38519
rect 54479 38485 54513 38519
rect 54663 38485 54697 38519
rect 73431 38485 73465 38519
rect 91555 38485 91589 38519
rect 4339 38417 4373 38451
rect 10043 38417 10077 38451
rect 16207 38417 16241 38451
rect 16391 38417 16425 38451
rect 17771 38417 17805 38451
rect 17863 38417 17897 38451
rect 23751 38417 23785 38451
rect 23843 38417 23877 38451
rect 24303 38417 24337 38451
rect 24487 38417 24521 38451
rect 27523 38417 27557 38451
rect 27799 38417 27833 38451
rect 33043 38417 33077 38451
rect 33319 38417 33353 38451
rect 39207 38417 39241 38451
rect 39483 38417 39517 38451
rect 40035 38417 40069 38451
rect 41231 38417 41265 38451
rect 44727 38417 44761 38451
rect 48407 38417 48441 38451
rect 48591 38417 48625 38451
rect 51351 38417 51385 38451
rect 51535 38417 51569 38451
rect 51995 38417 52029 38451
rect 52087 38417 52121 38451
rect 55307 38417 55341 38451
rect 55675 38417 55709 38451
rect 55859 38417 55893 38451
rect 55951 38417 55985 38451
rect 60367 38417 60401 38451
rect 63495 38417 63529 38451
rect 66899 38417 66933 38451
rect 67083 38417 67117 38451
rect 67635 38417 67669 38451
rect 67819 38417 67853 38451
rect 68371 38417 68405 38451
rect 69107 38417 69141 38451
rect 72327 38417 72361 38451
rect 74075 38417 74109 38451
rect 74443 38417 74477 38451
rect 74627 38417 74661 38451
rect 77755 38417 77789 38451
rect 79963 38417 79997 38451
rect 83091 38417 83125 38451
rect 83275 38417 83309 38451
rect 83827 38417 83861 38451
rect 84011 38417 84045 38451
rect 85299 38417 85333 38451
rect 88979 38417 89013 38451
rect 89163 38417 89197 38451
rect 89715 38417 89749 38451
rect 89899 38417 89933 38451
rect 91463 38417 91497 38451
rect 1855 38349 1889 38383
rect 4063 38349 4097 38383
rect 5719 38349 5753 38383
rect 10319 38349 10353 38383
rect 29179 38349 29213 38383
rect 33595 38349 33629 38383
rect 40311 38349 40345 38383
rect 44451 38349 44485 38383
rect 55399 38349 55433 38383
rect 60643 38349 60677 38383
rect 69199 38349 69233 38383
rect 74167 38349 74201 38383
rect 77479 38349 77513 38383
rect 84379 38349 84413 38383
rect 24671 38281 24705 38315
rect 39575 38281 39609 38315
rect 52455 38281 52489 38315
rect 5903 38213 5937 38247
rect 11423 38213 11457 38247
rect 17587 38213 17621 38247
rect 18047 38213 18081 38247
rect 18507 38213 18541 38247
rect 25131 38213 25165 38247
rect 25315 38213 25349 38247
rect 34883 38213 34917 38247
rect 41047 38213 41081 38247
rect 46015 38213 46049 38247
rect 46199 38213 46233 38247
rect 48131 38213 48165 38247
rect 49143 38213 49177 38247
rect 56227 38213 56261 38247
rect 61747 38213 61781 38247
rect 63311 38213 63345 38247
rect 68095 38213 68129 38247
rect 72235 38213 72269 38247
rect 77387 38213 77421 38247
rect 79043 38213 79077 38247
rect 84563 38213 84597 38247
rect 85391 38213 85425 38247
rect 9307 38009 9341 38043
rect 17495 38009 17529 38043
rect 20163 38009 20197 38043
rect 27615 38009 27649 38043
rect 33227 38009 33261 38043
rect 40863 38009 40897 38043
rect 42151 38009 42185 38043
rect 69383 38009 69417 38043
rect 86403 38009 86437 38043
rect 90175 38009 90209 38043
rect 8847 37941 8881 37975
rect 47211 37941 47245 37975
rect 72603 37941 72637 37975
rect 7743 37873 7777 37907
rect 16575 37873 16609 37907
rect 18231 37873 18265 37907
rect 20899 37873 20933 37907
rect 22923 37873 22957 37907
rect 23107 37873 23141 37907
rect 23383 37873 23417 37907
rect 25683 37873 25717 37907
rect 29915 37873 29949 37907
rect 32031 37873 32065 37907
rect 36631 37873 36665 37907
rect 47303 37873 47337 37907
rect 47487 37873 47521 37907
rect 50983 37873 51017 37907
rect 51259 37873 51293 37907
rect 58251 37873 58285 37907
rect 59539 37873 59573 37907
rect 68003 37873 68037 37907
rect 68279 37873 68313 37907
rect 69843 37873 69877 37907
rect 74075 37873 74109 37907
rect 79319 37873 79353 37907
rect 82631 37873 82665 37907
rect 85115 37873 85149 37907
rect 88611 37873 88645 37907
rect 89071 37873 89105 37907
rect 90451 37873 90485 37907
rect 2131 37805 2165 37839
rect 2407 37805 2441 37839
rect 7467 37805 7501 37839
rect 12527 37805 12561 37839
rect 12803 37805 12837 37839
rect 16207 37805 16241 37839
rect 17771 37805 17805 37839
rect 20439 37805 20473 37839
rect 24763 37805 24797 37839
rect 25499 37805 25533 37839
rect 25591 37805 25625 37839
rect 27431 37805 27465 37839
rect 28719 37805 28753 37839
rect 29823 37805 29857 37839
rect 31755 37805 31789 37839
rect 31847 37805 31881 37839
rect 32215 37805 32249 37839
rect 32767 37805 32801 37839
rect 32951 37805 32985 37839
rect 34699 37805 34733 37839
rect 34791 37805 34825 37839
rect 36447 37805 36481 37839
rect 36723 37805 36757 37839
rect 37183 37805 37217 37839
rect 37275 37805 37309 37839
rect 40771 37805 40805 37839
rect 41967 37805 42001 37839
rect 45371 37805 45405 37839
rect 45555 37805 45589 37839
rect 48039 37805 48073 37839
rect 48315 37805 48349 37839
rect 48499 37805 48533 37839
rect 51351 37805 51385 37839
rect 51903 37805 51937 37839
rect 52087 37805 52121 37839
rect 54939 37805 54973 37839
rect 55031 37805 55065 37839
rect 56319 37805 56353 37839
rect 57883 37805 57917 37839
rect 58389 37805 58423 37839
rect 58987 37805 59021 37839
rect 59171 37805 59205 37839
rect 61287 37805 61321 37839
rect 62391 37805 62425 37839
rect 62667 37805 62701 37839
rect 72419 37805 72453 37839
rect 73983 37805 74017 37839
rect 74259 37805 74293 37839
rect 74719 37805 74753 37839
rect 74811 37805 74845 37839
rect 76467 37805 76501 37839
rect 79227 37805 79261 37839
rect 82723 37805 82757 37839
rect 83275 37805 83309 37839
rect 83459 37805 83493 37839
rect 84655 37805 84689 37839
rect 84839 37805 84873 37839
rect 88979 37805 89013 37839
rect 89347 37805 89381 37839
rect 89439 37805 89473 37839
rect 90727 37805 90761 37839
rect 3787 37737 3821 37771
rect 14183 37737 14217 37771
rect 16023 37737 16057 37771
rect 17679 37737 17713 37771
rect 18323 37737 18357 37771
rect 20347 37737 20381 37771
rect 29087 37737 29121 37771
rect 37827 37737 37861 37771
rect 40587 37737 40621 37771
rect 75363 37737 75397 37771
rect 83827 37737 83861 37771
rect 3971 37669 4005 37703
rect 14275 37669 14309 37703
rect 27339 37669 27373 37703
rect 28903 37669 28937 37703
rect 29731 37669 29765 37703
rect 33595 37669 33629 37703
rect 34975 37669 35009 37703
rect 38103 37669 38137 37703
rect 40403 37669 40437 37703
rect 41231 37669 41265 37703
rect 41783 37669 41817 37703
rect 45371 37669 45405 37703
rect 45647 37669 45681 37703
rect 52363 37669 52397 37703
rect 55215 37669 55249 37703
rect 56135 37669 56169 37703
rect 57699 37669 57733 37703
rect 58067 37669 58101 37703
rect 59723 37669 59757 37703
rect 61379 37669 61413 37703
rect 62115 37669 62149 37703
rect 63771 37669 63805 37703
rect 72327 37669 72361 37703
rect 76283 37669 76317 37703
rect 84011 37669 84045 37703
rect 91831 37669 91865 37703
rect 5995 37465 6029 37499
rect 10411 37465 10445 37499
rect 12435 37465 12469 37499
rect 27247 37465 27281 37499
rect 31939 37465 31973 37499
rect 32123 37465 32157 37499
rect 33595 37465 33629 37499
rect 75271 37465 75305 37499
rect 82263 37465 82297 37499
rect 88703 37465 88737 37499
rect 90083 37465 90117 37499
rect 15655 37397 15689 37431
rect 16207 37397 16241 37431
rect 4155 37329 4189 37363
rect 4431 37329 4465 37363
rect 10779 37329 10813 37363
rect 11147 37329 11181 37363
rect 11239 37329 11273 37363
rect 12619 37329 12653 37363
rect 12803 37329 12837 37363
rect 13171 37329 13205 37363
rect 15839 37329 15873 37363
rect 17219 37329 17253 37363
rect 17311 37329 17345 37363
rect 20163 37329 20197 37363
rect 20347 37329 20381 37363
rect 27615 37329 27649 37363
rect 27983 37329 28017 37363
rect 28167 37329 28201 37363
rect 29455 37329 29489 37363
rect 10871 37261 10905 37295
rect 13079 37261 13113 37295
rect 20623 37261 20657 37295
rect 27707 37261 27741 37295
rect 29363 37261 29397 37295
rect 40587 37397 40621 37431
rect 58343 37397 58377 37431
rect 60919 37397 60953 37431
rect 72051 37397 72085 37431
rect 32675 37329 32709 37363
rect 33043 37329 33077 37363
rect 33227 37329 33261 37363
rect 37367 37329 37401 37363
rect 37459 37329 37493 37363
rect 37919 37329 37953 37363
rect 38103 37329 38137 37363
rect 39207 37329 39241 37363
rect 39483 37329 39517 37363
rect 40219 37329 40253 37363
rect 41139 37329 41173 37363
rect 41415 37329 41449 37363
rect 42979 37329 43013 37363
rect 43531 37329 43565 37363
rect 43715 37329 43749 37363
rect 44359 37329 44393 37363
rect 45371 37329 45405 37363
rect 46383 37329 46417 37363
rect 46751 37329 46785 37363
rect 50891 37329 50925 37363
rect 55031 37329 55065 37363
rect 55491 37329 55525 37363
rect 55583 37329 55617 37363
rect 57239 37329 57273 37363
rect 57791 37329 57825 37363
rect 57975 37329 58009 37363
rect 58619 37329 58653 37363
rect 59815 37329 59849 37363
rect 60367 37329 60401 37363
rect 60551 37329 60585 37363
rect 62759 37329 62793 37363
rect 67083 37329 67117 37363
rect 67451 37329 67485 37363
rect 67635 37329 67669 37363
rect 68647 37329 68681 37363
rect 69199 37329 69233 37363
rect 69383 37329 69417 37363
rect 72695 37329 72729 37363
rect 73063 37329 73097 37363
rect 73247 37329 73281 37363
rect 74075 37329 74109 37363
rect 74259 37329 74293 37363
rect 74811 37329 74845 37363
rect 74995 37329 75029 37363
rect 77939 37329 77973 37363
rect 80515 37329 80549 37363
rect 82079 37329 82113 37363
rect 82447 37329 82481 37363
rect 84287 37329 84321 37363
rect 85667 37329 85701 37363
rect 86495 37329 86529 37363
rect 88887 37329 88921 37363
rect 89071 37329 89105 37363
rect 89531 37329 89565 37363
rect 89623 37329 89657 37363
rect 91279 37329 91313 37363
rect 32767 37261 32801 37295
rect 40495 37261 40529 37295
rect 41599 37261 41633 37295
rect 41691 37261 41725 37295
rect 42887 37261 42921 37295
rect 46199 37261 46233 37295
rect 46659 37261 46693 37295
rect 50615 37261 50649 37295
rect 54939 37261 54973 37295
rect 56135 37261 56169 37295
rect 57147 37261 57181 37295
rect 59631 37261 59665 37295
rect 62483 37261 62517 37295
rect 67175 37261 67209 37295
rect 68555 37261 68589 37295
rect 72787 37261 72821 37295
rect 77663 37261 77697 37295
rect 84011 37261 84045 37295
rect 5719 37193 5753 37227
rect 17035 37193 17069 37227
rect 31939 37193 31973 37227
rect 33411 37193 33445 37227
rect 38287 37193 38321 37227
rect 38747 37193 38781 37227
rect 39207 37193 39241 37227
rect 66715 37193 66749 37227
rect 69567 37193 69601 37227
rect 91371 37193 91405 37227
rect 17495 37125 17529 37159
rect 21727 37125 21761 37159
rect 29639 37125 29673 37159
rect 39299 37125 39333 37159
rect 39667 37125 39701 37159
rect 43991 37125 44025 37159
rect 45555 37125 45589 37159
rect 46015 37125 46049 37159
rect 52179 37125 52213 37159
rect 52363 37125 52397 37159
rect 61195 37125 61229 37159
rect 62299 37125 62333 37159
rect 64047 37125 64081 37159
rect 77479 37125 77513 37159
rect 79227 37125 79261 37159
rect 80331 37125 80365 37159
rect 80699 37125 80733 37159
rect 83919 37125 83953 37159
rect 86587 37125 86621 37159
rect 2223 36921 2257 36955
rect 16299 36921 16333 36955
rect 17771 36921 17805 36955
rect 21359 36921 21393 36955
rect 57239 36921 57273 36955
rect 62391 36921 62425 36955
rect 64139 36921 64173 36955
rect 73799 36921 73833 36955
rect 76007 36921 76041 36955
rect 88611 36921 88645 36955
rect 40495 36853 40529 36887
rect 43991 36853 44025 36887
rect 45555 36853 45589 36887
rect 50155 36853 50189 36887
rect 58251 36853 58285 36887
rect 3143 36785 3177 36819
rect 18139 36785 18173 36819
rect 19703 36785 19737 36819
rect 20347 36785 20381 36819
rect 31387 36785 31421 36819
rect 32123 36785 32157 36819
rect 51995 36785 52029 36819
rect 53559 36785 53593 36819
rect 1579 36717 1613 36751
rect 3419 36717 3453 36751
rect 9675 36717 9709 36751
rect 16207 36717 16241 36751
rect 17495 36717 17529 36751
rect 17679 36717 17713 36751
rect 19887 36717 19921 36751
rect 20071 36717 20105 36751
rect 21267 36717 21301 36751
rect 28719 36717 28753 36751
rect 31985 36717 32019 36751
rect 32399 36717 32433 36751
rect 32583 36717 32617 36751
rect 32767 36717 32801 36751
rect 37643 36717 37677 36751
rect 40127 36717 40161 36751
rect 40311 36717 40345 36751
rect 42703 36717 42737 36751
rect 42795 36717 42829 36751
rect 43163 36717 43197 36751
rect 43255 36717 43289 36751
rect 46199 36717 46233 36751
rect 46383 36717 46417 36751
rect 46751 36717 46785 36751
rect 46843 36717 46877 36751
rect 50063 36717 50097 36751
rect 51719 36717 51753 36751
rect 56871 36717 56905 36751
rect 57055 36717 57089 36751
rect 58067 36717 58101 36751
rect 58159 36717 58193 36751
rect 4799 36649 4833 36683
rect 20623 36649 20657 36683
rect 43807 36649 43841 36683
rect 62575 36853 62609 36887
rect 68003 36785 68037 36819
rect 69199 36785 69233 36819
rect 80883 36853 80917 36887
rect 79319 36785 79353 36819
rect 84839 36785 84873 36819
rect 85299 36785 85333 36819
rect 86311 36785 86345 36819
rect 62483 36717 62517 36751
rect 64047 36717 64081 36751
rect 68172 36717 68206 36751
rect 68647 36717 68681 36751
rect 68739 36717 68773 36751
rect 73431 36717 73465 36751
rect 73615 36717 73649 36751
rect 74075 36717 74109 36751
rect 76007 36717 76041 36751
rect 76283 36717 76317 36751
rect 79227 36717 79261 36751
rect 80975 36717 81009 36751
rect 85483 36717 85517 36751
rect 85851 36717 85885 36751
rect 85943 36717 85977 36751
rect 88795 36717 88829 36751
rect 88979 36717 89013 36751
rect 89301 36717 89335 36751
rect 89531 36717 89565 36751
rect 73063 36649 73097 36683
rect 4983 36581 5017 36615
rect 9491 36581 9525 36615
rect 9859 36581 9893 36615
rect 16115 36581 16149 36615
rect 28811 36581 28845 36615
rect 32859 36581 32893 36615
rect 37551 36581 37585 36615
rect 37827 36581 37861 36615
rect 46015 36581 46049 36615
rect 53283 36581 53317 36615
rect 62391 36581 62425 36615
rect 73247 36581 73281 36615
rect 76099 36581 76133 36615
rect 81159 36581 81193 36615
rect 86127 36581 86161 36615
rect 2499 36377 2533 36411
rect 7375 36377 7409 36411
rect 9767 36377 9801 36411
rect 15471 36377 15505 36411
rect 17863 36377 17897 36411
rect 29271 36377 29305 36411
rect 65703 36377 65737 36411
rect 66071 36377 66105 36411
rect 80699 36377 80733 36411
rect 82355 36377 82389 36411
rect 88427 36377 88461 36411
rect 7191 36309 7225 36343
rect 37459 36309 37493 36343
rect 39207 36309 39241 36343
rect 40495 36309 40529 36343
rect 5535 36241 5569 36275
rect 5811 36241 5845 36275
rect 9583 36241 9617 36275
rect 11607 36241 11641 36275
rect 11791 36241 11825 36275
rect 12159 36241 12193 36275
rect 15655 36241 15689 36275
rect 18967 36241 19001 36275
rect 21359 36241 21393 36275
rect 21635 36241 21669 36275
rect 23475 36241 23509 36275
rect 24027 36241 24061 36275
rect 24211 36241 24245 36275
rect 27431 36241 27465 36275
rect 32583 36241 32617 36275
rect 32951 36241 32985 36275
rect 33503 36241 33537 36275
rect 33687 36241 33721 36275
rect 34331 36241 34365 36275
rect 37643 36241 37677 36275
rect 39115 36241 39149 36275
rect 39851 36241 39885 36275
rect 40219 36241 40253 36275
rect 45371 36241 45405 36275
rect 45555 36241 45589 36275
rect 45647 36241 45681 36275
rect 51627 36241 51661 36275
rect 51995 36241 52029 36275
rect 54019 36241 54053 36275
rect 56779 36241 56813 36275
rect 61839 36241 61873 36275
rect 62299 36241 62333 36275
rect 62391 36241 62425 36275
rect 65887 36241 65921 36275
rect 67727 36241 67761 36275
rect 73339 36241 73373 36275
rect 73523 36241 73557 36275
rect 73983 36241 74017 36275
rect 74075 36241 74109 36275
rect 80515 36241 80549 36275
rect 82723 36241 82757 36275
rect 83091 36241 83125 36275
rect 88611 36241 88645 36275
rect 88795 36241 88829 36275
rect 89347 36241 89381 36275
rect 89531 36241 89565 36275
rect 91371 36241 91405 36275
rect 1855 36173 1889 36207
rect 12067 36173 12101 36207
rect 16483 36173 16517 36207
rect 16759 36173 16793 36207
rect 23383 36173 23417 36207
rect 27707 36173 27741 36207
rect 32215 36173 32249 36207
rect 32859 36173 32893 36207
rect 34055 36173 34089 36207
rect 38931 36173 38965 36207
rect 39667 36173 39701 36207
rect 40127 36173 40161 36207
rect 50983 36173 51017 36207
rect 51443 36173 51477 36207
rect 51903 36173 51937 36207
rect 54111 36173 54145 36207
rect 56411 36173 56445 36207
rect 56503 36173 56537 36207
rect 61563 36173 61597 36207
rect 61655 36173 61689 36207
rect 67451 36173 67485 36207
rect 82539 36173 82573 36207
rect 82999 36173 83033 36207
rect 23199 36105 23233 36139
rect 37827 36105 37861 36139
rect 58067 36105 58101 36139
rect 69199 36105 69233 36139
rect 80331 36105 80365 36139
rect 91463 36105 91497 36139
rect 11423 36037 11457 36071
rect 16299 36037 16333 36071
rect 19059 36037 19093 36071
rect 21451 36037 21485 36071
rect 24487 36037 24521 36071
rect 28995 36037 29029 36071
rect 32399 36037 32433 36071
rect 40679 36037 40713 36071
rect 52363 36037 52397 36071
rect 52547 36037 52581 36071
rect 62851 36037 62885 36071
rect 63219 36037 63253 36071
rect 69015 36037 69049 36071
rect 74535 36037 74569 36071
rect 88243 36037 88277 36071
rect 89807 36037 89841 36071
rect 16483 35833 16517 35867
rect 21267 35833 21301 35867
rect 28995 35833 29029 35867
rect 48407 35833 48441 35867
rect 54387 35833 54421 35867
rect 85575 35833 85609 35867
rect 91831 35833 91865 35867
rect 17679 35765 17713 35799
rect 34515 35765 34549 35799
rect 34791 35765 34825 35799
rect 40035 35765 40069 35799
rect 56963 35765 56997 35799
rect 68095 35765 68129 35799
rect 76007 35765 76041 35799
rect 2683 35697 2717 35731
rect 10411 35697 10445 35731
rect 12159 35697 12193 35731
rect 18047 35697 18081 35731
rect 23383 35697 23417 35731
rect 29639 35697 29673 35731
rect 32031 35697 32065 35731
rect 37643 35697 37677 35731
rect 43255 35697 43289 35731
rect 48683 35697 48717 35731
rect 49327 35697 49361 35731
rect 57975 35697 58009 35731
rect 58159 35697 58193 35731
rect 59723 35697 59757 35731
rect 63955 35697 63989 35731
rect 69291 35697 69325 35731
rect 70763 35697 70797 35731
rect 73615 35697 73649 35731
rect 86771 35697 86805 35731
rect 88059 35697 88093 35731
rect 88243 35697 88277 35731
rect 90727 35697 90761 35731
rect 2407 35629 2441 35663
rect 10319 35629 10353 35663
rect 10687 35629 10721 35663
rect 10779 35629 10813 35663
rect 11883 35629 11917 35663
rect 13631 35629 13665 35663
rect 14827 35629 14861 35663
rect 16391 35629 16425 35663
rect 17587 35629 17621 35663
rect 17863 35629 17897 35663
rect 20623 35629 20657 35663
rect 20899 35629 20933 35663
rect 21083 35629 21117 35663
rect 23107 35629 23141 35663
rect 24763 35629 24797 35663
rect 25591 35629 25625 35663
rect 25683 35629 25717 35663
rect 29179 35629 29213 35663
rect 29363 35629 29397 35663
rect 29731 35629 29765 35663
rect 32123 35629 32157 35663
rect 32675 35629 32709 35663
rect 32859 35629 32893 35663
rect 34331 35629 34365 35663
rect 37367 35629 37401 35663
rect 39943 35629 39977 35663
rect 42979 35629 43013 35663
rect 45555 35629 45589 35663
rect 46935 35629 46969 35663
rect 48591 35629 48625 35663
rect 48867 35629 48901 35663
rect 52455 35629 52489 35663
rect 52639 35629 52673 35663
rect 52823 35629 52857 35663
rect 53375 35629 53409 35663
rect 53559 35629 53593 35663
rect 56779 35629 56813 35663
rect 57147 35629 57181 35663
rect 58343 35629 58377 35663
rect 58895 35629 58929 35663
rect 59079 35629 59113 35663
rect 62391 35629 62425 35663
rect 62575 35629 62609 35663
rect 63035 35629 63069 35663
rect 63215 35629 63249 35663
rect 68003 35629 68037 35663
rect 69015 35629 69049 35663
rect 73799 35629 73833 35663
rect 74259 35629 74293 35663
rect 74351 35629 74385 35663
rect 75823 35629 75857 35663
rect 79227 35629 79261 35663
rect 79595 35629 79629 35663
rect 82079 35629 82113 35663
rect 82263 35629 82297 35663
rect 82723 35629 82757 35663
rect 82815 35629 82849 35663
rect 85759 35629 85793 35663
rect 85943 35629 85977 35663
rect 86311 35629 86345 35663
rect 86495 35629 86529 35663
rect 88335 35629 88369 35663
rect 88795 35629 88829 35663
rect 88887 35629 88921 35663
rect 90451 35629 90485 35663
rect 20071 35561 20105 35595
rect 24947 35561 24981 35595
rect 33227 35561 33261 35595
rect 39023 35561 39057 35595
rect 44635 35561 44669 35595
rect 45647 35561 45681 35595
rect 59447 35561 59481 35595
rect 70671 35561 70705 35595
rect 83367 35561 83401 35595
rect 89439 35561 89473 35595
rect 3971 35493 4005 35527
rect 4247 35493 4281 35527
rect 9951 35493 9985 35527
rect 13263 35493 13297 35527
rect 14643 35493 14677 35527
rect 17219 35493 17253 35527
rect 18507 35493 18541 35527
rect 30099 35493 30133 35527
rect 33503 35493 33537 35527
rect 37183 35493 37217 35527
rect 42795 35493 42829 35527
rect 47027 35493 47061 35527
rect 53835 35493 53869 35527
rect 54111 35493 54145 35527
rect 62115 35493 62149 35527
rect 63587 35493 63621 35527
rect 64139 35493 64173 35527
rect 74811 35493 74845 35527
rect 75639 35493 75673 35527
rect 79411 35493 79445 35527
rect 81711 35493 81745 35527
rect 81895 35493 81929 35527
rect 86679 35493 86713 35527
rect 90175 35493 90209 35527
rect 2499 35289 2533 35323
rect 6823 35289 6857 35323
rect 13079 35289 13113 35323
rect 15563 35289 15597 35323
rect 19427 35289 19461 35323
rect 24027 35289 24061 35323
rect 28259 35289 28293 35323
rect 29547 35289 29581 35323
rect 39115 35289 39149 35323
rect 43071 35289 43105 35323
rect 47579 35289 47613 35323
rect 49327 35289 49361 35323
rect 62391 35289 62425 35323
rect 80975 35289 81009 35323
rect 89531 35289 89565 35323
rect 15103 35221 15137 35255
rect 18231 35221 18265 35255
rect 23199 35221 23233 35255
rect 23383 35221 23417 35255
rect 50247 35221 50281 35255
rect 54939 35221 54973 35255
rect 68555 35221 68589 35255
rect 1855 35153 1889 35187
rect 5535 35153 5569 35187
rect 10135 35153 10169 35187
rect 11515 35153 11549 35187
rect 13263 35153 13297 35187
rect 13447 35153 13481 35187
rect 14735 35153 14769 35187
rect 14827 35153 14861 35187
rect 18783 35153 18817 35187
rect 19059 35153 19093 35187
rect 19243 35153 19277 35187
rect 21819 35153 21853 35187
rect 22371 35153 22405 35187
rect 22555 35153 22589 35187
rect 23843 35153 23877 35187
rect 24211 35153 24245 35187
rect 26971 35153 27005 35187
rect 27063 35153 27097 35187
rect 27247 35153 27281 35187
rect 27799 35153 27833 35187
rect 27983 35153 28017 35187
rect 29731 35153 29765 35187
rect 29915 35153 29949 35187
rect 30283 35153 30317 35187
rect 30375 35153 30409 35187
rect 33135 35153 33169 35187
rect 33411 35153 33445 35187
rect 34791 35153 34825 35187
rect 35619 35153 35653 35187
rect 35711 35153 35745 35187
rect 37827 35153 37861 35187
rect 40035 35153 40069 35187
rect 43255 35153 43289 35187
rect 43531 35153 43565 35187
rect 44911 35153 44945 35187
rect 46015 35153 46049 35187
rect 49511 35153 49545 35187
rect 49603 35153 49637 35187
rect 49787 35153 49821 35187
rect 51259 35153 51293 35187
rect 51903 35153 51937 35187
rect 52271 35153 52305 35187
rect 52455 35153 52489 35187
rect 54019 35153 54053 35187
rect 62391 35153 62425 35187
rect 62621 35153 62655 35187
rect 62759 35153 62793 35187
rect 63127 35153 63161 35187
rect 63219 35153 63253 35187
rect 65887 35153 65921 35187
rect 66163 35153 66197 35187
rect 69199 35153 69233 35187
rect 69567 35153 69601 35187
rect 70855 35153 70889 35187
rect 73891 35153 73925 35187
rect 74167 35153 74201 35187
rect 79227 35153 79261 35187
rect 79411 35153 79445 35187
rect 79687 35153 79721 35187
rect 83091 35153 83125 35187
rect 83275 35153 83309 35187
rect 83551 35153 83585 35187
rect 89715 35153 89749 35187
rect 89991 35153 90025 35187
rect 5259 35085 5293 35119
rect 9859 35085 9893 35119
rect 15747 35085 15781 35119
rect 16023 35085 16057 35119
rect 21635 35085 21669 35119
rect 30651 35085 30685 35119
rect 37551 35085 37585 35119
rect 45739 35085 45773 35119
rect 51995 35085 52029 35119
rect 54387 35085 54421 35119
rect 54663 35085 54697 35119
rect 69291 35085 69325 35119
rect 69659 35085 69693 35119
rect 69935 35085 69969 35119
rect 75639 35085 75673 35119
rect 22739 35017 22773 35051
rect 34883 35017 34917 35051
rect 37367 35017 37401 35051
rect 70947 35017 70981 35051
rect 7099 34949 7133 34983
rect 11607 34949 11641 34983
rect 13539 34949 13573 34983
rect 17311 34949 17345 34983
rect 21543 34949 21577 34983
rect 40127 34949 40161 34983
rect 47119 34949 47153 34983
rect 52639 34949 52673 34983
rect 52731 34949 52765 34983
rect 54157 34949 54191 34983
rect 54295 34949 54329 34983
rect 63679 34949 63713 34983
rect 65979 34949 66013 34983
rect 68371 34949 68405 34983
rect 75271 34949 75305 34983
rect 84655 34949 84689 34983
rect 91095 34949 91129 34983
rect 4155 34745 4189 34779
rect 12803 34745 12837 34779
rect 17035 34745 17069 34779
rect 18691 34745 18725 34779
rect 26051 34745 26085 34779
rect 26584 34745 26618 34779
rect 27339 34745 27373 34779
rect 33963 34745 33997 34779
rect 34607 34745 34641 34779
rect 91187 34745 91221 34779
rect 2315 34609 2349 34643
rect 21267 34609 21301 34643
rect 24671 34609 24705 34643
rect 26695 34677 26729 34711
rect 29639 34677 29673 34711
rect 29915 34677 29949 34711
rect 48131 34677 48165 34711
rect 51995 34677 52029 34711
rect 54847 34677 54881 34711
rect 68003 34677 68037 34711
rect 69291 34677 69325 34711
rect 81159 34677 81193 34711
rect 26235 34609 26269 34643
rect 26787 34609 26821 34643
rect 40035 34609 40069 34643
rect 47671 34609 47705 34643
rect 52087 34609 52121 34643
rect 53375 34609 53409 34643
rect 58067 34609 58101 34643
rect 59447 34609 59481 34643
rect 59907 34609 59941 34643
rect 62391 34609 62425 34643
rect 74259 34609 74293 34643
rect 74535 34609 74569 34643
rect 80147 34609 80181 34643
rect 2591 34541 2625 34575
rect 6363 34541 6397 34575
rect 6455 34541 6489 34575
rect 12895 34541 12929 34575
rect 17219 34541 17253 34575
rect 18231 34541 18265 34575
rect 20531 34541 20565 34575
rect 20623 34541 20657 34575
rect 20807 34541 20841 34575
rect 24855 34541 24889 34575
rect 25039 34541 25073 34575
rect 25407 34541 25441 34575
rect 25499 34541 25533 34575
rect 26051 34541 26085 34575
rect 29731 34541 29765 34575
rect 34147 34541 34181 34575
rect 34791 34541 34825 34575
rect 35067 34541 35101 34575
rect 36447 34541 36481 34575
rect 38195 34541 38229 34575
rect 40127 34541 40161 34575
rect 40587 34541 40621 34575
rect 40679 34541 40713 34575
rect 46291 34541 46325 34575
rect 46567 34541 46601 34575
rect 48775 34541 48809 34575
rect 51866 34541 51900 34575
rect 53099 34541 53133 34575
rect 53467 34541 53501 34575
rect 54019 34541 54053 34575
rect 54203 34541 54237 34575
rect 58343 34541 58377 34575
rect 58435 34541 58469 34575
rect 58895 34541 58929 34575
rect 59079 34541 59113 34575
rect 59723 34541 59757 34575
rect 62575 34541 62609 34575
rect 63035 34541 63069 34575
rect 63215 34541 63249 34575
rect 67819 34541 67853 34575
rect 68187 34541 68221 34575
rect 68371 34541 68405 34575
rect 68831 34541 68865 34575
rect 68923 34541 68957 34575
rect 76007 34541 76041 34575
rect 80239 34541 80273 34575
rect 80791 34541 80825 34575
rect 80975 34541 81009 34575
rect 82723 34541 82757 34575
rect 82999 34541 83033 34575
rect 85943 34541 85977 34575
rect 86127 34541 86161 34575
rect 86587 34541 86621 34575
rect 86679 34541 86713 34575
rect 91095 34541 91129 34575
rect 6547 34473 6581 34507
rect 20347 34473 20381 34507
rect 26419 34473 26453 34507
rect 41231 34473 41265 34507
rect 48867 34473 48901 34507
rect 51719 34473 51753 34507
rect 52455 34473 52489 34507
rect 87231 34473 87265 34507
rect 3879 34405 3913 34439
rect 13079 34405 13113 34439
rect 17587 34405 17621 34439
rect 18415 34405 18449 34439
rect 21451 34405 21485 34439
rect 25775 34405 25809 34439
rect 25959 34405 25993 34439
rect 27063 34405 27097 34439
rect 38287 34405 38321 34439
rect 51535 34405 51569 34439
rect 54479 34405 54513 34439
rect 55031 34405 55065 34439
rect 63587 34405 63621 34439
rect 69659 34405 69693 34439
rect 75639 34405 75673 34439
rect 82815 34405 82849 34439
rect 85851 34405 85885 34439
rect 87415 34405 87449 34439
rect 15931 34201 15965 34235
rect 17311 34201 17345 34235
rect 17679 34201 17713 34235
rect 52823 34201 52857 34235
rect 81067 34201 81101 34235
rect 6731 34133 6765 34167
rect 36999 34133 37033 34167
rect 45095 34133 45129 34167
rect 46751 34133 46785 34167
rect 54387 34133 54421 34167
rect 60367 34133 60401 34167
rect 63587 34133 63621 34167
rect 67543 34133 67577 34167
rect 69383 34133 69417 34167
rect 74995 34133 75029 34167
rect 80883 34133 80917 34167
rect 5351 34065 5385 34099
rect 8939 34065 8973 34099
rect 9583 34065 9617 34099
rect 9767 34065 9801 34099
rect 10135 34065 10169 34099
rect 10227 34065 10261 34099
rect 16115 34065 16149 34099
rect 16299 34065 16333 34099
rect 16851 34065 16885 34099
rect 17035 34065 17069 34099
rect 22279 34065 22313 34099
rect 23659 34065 23693 34099
rect 25959 34065 25993 34099
rect 28903 34065 28937 34099
rect 31663 34065 31697 34099
rect 32031 34065 32065 34099
rect 33319 34065 33353 34099
rect 33503 34065 33537 34099
rect 34055 34065 34089 34099
rect 34239 34065 34273 34099
rect 34883 34065 34917 34099
rect 5075 33997 5109 34031
rect 21819 33997 21853 34031
rect 22003 33997 22037 34031
rect 26327 33997 26361 34031
rect 26695 33997 26729 34031
rect 6915 33929 6949 33963
rect 17863 33929 17897 33963
rect 25683 33929 25717 33963
rect 26124 33929 26158 33963
rect 26879 33929 26913 33963
rect 29087 33929 29121 33963
rect 34423 33929 34457 33963
rect 39805 34065 39839 34099
rect 39943 34065 39977 34099
rect 40311 34065 40345 34099
rect 40403 34065 40437 34099
rect 45003 34065 45037 34099
rect 46935 34065 46969 34099
rect 51259 34065 51293 34099
rect 51443 34065 51477 34099
rect 51627 34065 51661 34099
rect 51811 34065 51845 34099
rect 52363 34065 52397 34099
rect 52547 34065 52581 34099
rect 55123 34065 55157 34099
rect 59631 34065 59665 34099
rect 60551 34065 60585 34099
rect 63817 34065 63851 34099
rect 67911 34065 67945 34099
rect 68095 34065 68129 34099
rect 68555 34065 68589 34099
rect 68647 34065 68681 34099
rect 73615 34065 73649 34099
rect 74903 34065 74937 34099
rect 77939 34065 77973 34099
rect 78123 34065 78157 34099
rect 78675 34065 78709 34099
rect 78859 34065 78893 34099
rect 80791 34065 80825 34099
rect 90451 34065 90485 34099
rect 91003 34065 91037 34099
rect 91187 34065 91221 34099
rect 40955 33997 40989 34031
rect 54203 33997 54237 34031
rect 54534 33997 54568 34031
rect 54755 33997 54789 34031
rect 59999 33997 60033 34031
rect 63955 33997 63989 34031
rect 64323 33997 64357 34031
rect 73523 33997 73557 34031
rect 74075 33997 74109 34031
rect 90267 33997 90301 34031
rect 59907 33929 59941 33963
rect 63403 33929 63437 33963
rect 67819 33929 67853 33963
rect 69015 33929 69049 33963
rect 79043 33929 79077 33963
rect 91371 33929 91405 33963
rect 9399 33861 9433 33895
rect 26235 33861 26269 33895
rect 31847 33861 31881 33895
rect 35067 33861 35101 33895
rect 36999 33861 37033 33895
rect 47027 33861 47061 33895
rect 53191 33861 53225 33895
rect 53375 33861 53409 33895
rect 54663 33861 54697 33895
rect 59769 33861 59803 33895
rect 63752 33861 63786 33895
rect 64507 33861 64541 33895
rect 74167 33861 74201 33895
rect 2775 33657 2809 33691
rect 17587 33657 17621 33691
rect 23291 33657 23325 33691
rect 29363 33657 29397 33691
rect 53927 33657 53961 33691
rect 57515 33657 57549 33691
rect 58987 33657 59021 33691
rect 60137 33657 60171 33691
rect 60275 33657 60309 33691
rect 60459 33657 60493 33691
rect 63495 33657 63529 33691
rect 64139 33657 64173 33691
rect 75087 33657 75121 33691
rect 85667 33657 85701 33691
rect 85851 33657 85885 33691
rect 13171 33589 13205 33623
rect 26787 33589 26821 33623
rect 63384 33589 63418 33623
rect 65887 33589 65921 33623
rect 91555 33589 91589 33623
rect 2131 33521 2165 33555
rect 9031 33521 9065 33555
rect 12619 33521 12653 33555
rect 12987 33521 13021 33555
rect 24119 33521 24153 33555
rect 24303 33521 24337 33555
rect 30375 33521 30409 33555
rect 57515 33521 57549 33555
rect 59263 33521 59297 33555
rect 63587 33521 63621 33555
rect 65979 33521 66013 33555
rect 68739 33521 68773 33555
rect 73615 33521 73649 33555
rect 74167 33521 74201 33555
rect 81435 33521 81469 33555
rect 90543 33521 90577 33555
rect 3051 33453 3085 33487
rect 4615 33453 4649 33487
rect 4799 33453 4833 33487
rect 5167 33453 5201 33487
rect 5351 33453 5385 33487
rect 8755 33453 8789 33487
rect 10503 33453 10537 33487
rect 12527 33453 12561 33487
rect 12895 33453 12929 33487
rect 13815 33453 13849 33487
rect 13907 33453 13941 33487
rect 17495 33453 17529 33487
rect 18783 33453 18817 33487
rect 20991 33453 21025 33487
rect 23199 33453 23233 33487
rect 24395 33453 24429 33487
rect 24947 33453 24981 33487
rect 25131 33453 25165 33487
rect 26603 33453 26637 33487
rect 29179 33453 29213 33487
rect 30283 33453 30317 33487
rect 31479 33453 31513 33487
rect 31571 33453 31605 33487
rect 32031 33453 32065 33487
rect 32215 33453 32249 33487
rect 35435 33453 35469 33487
rect 35527 33453 35561 33487
rect 40127 33453 40161 33487
rect 40587 33453 40621 33487
rect 44083 33453 44117 33487
rect 47119 33453 47153 33487
rect 51167 33453 51201 33487
rect 52731 33453 52765 33487
rect 52915 33453 52949 33487
rect 53375 33453 53409 33487
rect 53467 33453 53501 33487
rect 54295 33453 54329 33487
rect 54479 33453 54513 33487
rect 57975 33453 58009 33487
rect 58067 33453 58101 33487
rect 58435 33453 58469 33487
rect 58527 33453 58561 33487
rect 60338 33453 60372 33487
rect 60919 33453 60953 33487
rect 63219 33453 63253 33487
rect 63955 33453 63989 33487
rect 65758 33453 65792 33487
rect 68003 33453 68037 33487
rect 68647 33453 68681 33487
rect 69015 33453 69049 33487
rect 69199 33453 69233 33487
rect 73707 33453 73741 33487
rect 74995 33453 75029 33487
rect 79227 33453 79261 33487
rect 79411 33453 79445 33487
rect 79871 33453 79905 33487
rect 79963 33453 79997 33487
rect 81619 33453 81653 33487
rect 82171 33453 82205 33487
rect 82355 33453 82389 33487
rect 86035 33453 86069 33487
rect 86219 33453 86253 33487
rect 86403 33453 86437 33487
rect 86863 33453 86897 33487
rect 86955 33453 86989 33487
rect 90635 33453 90669 33487
rect 91095 33453 91129 33487
rect 91187 33453 91221 33487
rect 3971 33385 4005 33419
rect 10411 33385 10445 33419
rect 11883 33385 11917 33419
rect 13999 33385 14033 33419
rect 18875 33385 18909 33419
rect 39943 33385 39977 33419
rect 46935 33385 46969 33419
rect 47487 33385 47521 33419
rect 51259 33385 51293 33419
rect 59999 33385 60033 33419
rect 63127 33385 63161 33419
rect 65611 33385 65645 33419
rect 66347 33385 66381 33419
rect 80515 33385 80549 33419
rect 82723 33385 82757 33419
rect 87691 33385 87725 33419
rect 4431 33317 4465 33351
rect 20807 33317 20841 33351
rect 21175 33317 21209 33351
rect 25407 33317 25441 33351
rect 32491 33317 32525 33351
rect 32859 33317 32893 33351
rect 40219 33317 40253 33351
rect 43991 33317 44025 33351
rect 44175 33317 44209 33351
rect 52363 33317 52397 33351
rect 52547 33317 52581 33351
rect 57607 33317 57641 33351
rect 59447 33317 59481 33351
rect 65427 33317 65461 33351
rect 67727 33317 67761 33351
rect 69383 33317 69417 33351
rect 74351 33317 74385 33351
rect 87415 33317 87449 33351
rect 6547 33113 6581 33147
rect 13447 33113 13481 33147
rect 18875 33113 18909 33147
rect 22003 33113 22037 33147
rect 28995 33113 29029 33147
rect 33411 33113 33445 33147
rect 33871 33113 33905 33147
rect 35435 33113 35469 33147
rect 39299 33113 39333 33147
rect 43715 33113 43749 33147
rect 58527 33113 58561 33147
rect 60827 33113 60861 33147
rect 61195 33113 61229 33147
rect 65887 33113 65921 33147
rect 66163 33113 66197 33147
rect 82631 33113 82665 33147
rect 82907 33113 82941 33147
rect 18783 33045 18817 33079
rect 25959 33045 25993 33079
rect 46935 33045 46969 33079
rect 4707 32977 4741 33011
rect 4983 32977 5017 33011
rect 10043 32977 10077 33011
rect 11791 32977 11825 33011
rect 12527 32977 12561 33011
rect 13539 32977 13573 33011
rect 17403 32977 17437 33011
rect 17955 32977 17989 33011
rect 18139 32977 18173 33011
rect 20899 32977 20933 33011
rect 22187 32977 22221 33011
rect 25223 32977 25257 33011
rect 26603 32977 26637 33011
rect 26971 32977 27005 33011
rect 28903 32977 28937 33011
rect 31571 32977 31605 33011
rect 31847 32977 31881 33011
rect 34055 32977 34089 33011
rect 34331 32977 34365 33011
rect 37919 32977 37953 33011
rect 41047 32977 41081 33011
rect 41139 32977 41173 33011
rect 41415 32977 41449 33011
rect 43537 32977 43571 33011
rect 44635 32977 44669 33011
rect 44782 32977 44816 33011
rect 47027 32977 47061 33011
rect 48959 32977 48993 33011
rect 49695 32977 49729 33011
rect 54755 32977 54789 33011
rect 57515 32977 57549 33011
rect 58067 32977 58101 33011
rect 58251 32977 58285 33011
rect 59079 32977 59113 33011
rect 59815 32977 59849 33011
rect 60367 32977 60401 33011
rect 60551 32977 60585 33011
rect 62943 32977 62977 33011
rect 63127 32977 63161 33011
rect 63587 32977 63621 33011
rect 63679 32977 63713 33011
rect 65243 32977 65277 33011
rect 66531 32977 66565 33011
rect 67083 32977 67117 33011
rect 67543 32977 67577 33011
rect 67635 32977 67669 33011
rect 69107 32977 69141 33011
rect 74351 32977 74385 33011
rect 74443 32977 74477 33011
rect 74811 32977 74845 33011
rect 74903 32977 74937 33011
rect 77479 32977 77513 33011
rect 77939 32977 77973 33011
rect 78119 32977 78153 33011
rect 10319 32909 10353 32943
rect 12619 32909 12653 32943
rect 17311 32909 17345 32943
rect 20807 32909 20841 32943
rect 26419 32909 26453 32943
rect 26879 32909 26913 32943
rect 38195 32909 38229 32943
rect 41507 32909 41541 32943
rect 45003 32909 45037 32943
rect 49327 32909 49361 32943
rect 57055 32909 57089 32943
rect 57147 32909 57181 32943
rect 57331 32909 57365 32943
rect 59355 32909 59389 32943
rect 59631 32909 59665 32943
rect 64231 32909 64265 32943
rect 65611 32909 65645 32943
rect 66899 32909 66933 32943
rect 75363 32909 75397 32943
rect 77019 32909 77053 32943
rect 77295 32909 77329 32943
rect 22279 32841 22313 32875
rect 25039 32841 25073 32875
rect 37827 32841 37861 32875
rect 41783 32841 41817 32875
rect 41967 32841 42001 32875
rect 44911 32841 44945 32875
rect 45279 32841 45313 32875
rect 54939 32841 54973 32875
rect 64415 32841 64449 32875
rect 64691 32841 64725 32875
rect 65059 32841 65093 32875
rect 65519 32841 65553 32875
rect 68371 32841 68405 32875
rect 68647 32841 68681 32875
rect 74075 32841 74109 32875
rect 82723 32977 82757 33011
rect 83275 32977 83309 33011
rect 83367 32977 83401 33011
rect 83827 32977 83861 33011
rect 84011 32977 84045 33011
rect 86587 32977 86621 33011
rect 87967 32977 88001 33011
rect 87691 32909 87725 32943
rect 82631 32841 82665 32875
rect 6271 32773 6305 32807
rect 11423 32773 11457 32807
rect 13631 32773 13665 32807
rect 18415 32773 18449 32807
rect 21083 32773 21117 32807
rect 25315 32773 25349 32807
rect 27247 32773 27281 32807
rect 27523 32773 27557 32807
rect 33135 32773 33169 32807
rect 40495 32773 40529 32807
rect 44451 32773 44485 32807
rect 46751 32773 46785 32807
rect 47211 32773 47245 32807
rect 47579 32773 47613 32807
rect 57055 32773 57089 32807
rect 58803 32773 58837 32807
rect 61379 32773 61413 32807
rect 64875 32773 64909 32807
rect 65408 32773 65442 32807
rect 66715 32773 66749 32807
rect 68095 32773 68129 32807
rect 69199 32773 69233 32807
rect 75639 32773 75673 32807
rect 77019 32773 77053 32807
rect 77111 32773 77145 32807
rect 78491 32773 78525 32807
rect 84287 32773 84321 32807
rect 86679 32773 86713 32807
rect 87415 32773 87449 32807
rect 89071 32773 89105 32807
rect 4063 32569 4097 32603
rect 16115 32569 16149 32603
rect 16483 32569 16517 32603
rect 18875 32569 18909 32603
rect 21175 32569 21209 32603
rect 26787 32569 26821 32603
rect 33135 32569 33169 32603
rect 34515 32569 34549 32603
rect 35251 32569 35285 32603
rect 40311 32569 40345 32603
rect 43715 32569 43749 32603
rect 64323 32569 64357 32603
rect 65611 32569 65645 32603
rect 65795 32569 65829 32603
rect 77663 32569 77697 32603
rect 83256 32569 83290 32603
rect 4339 32501 4373 32535
rect 5075 32501 5109 32535
rect 7191 32501 7225 32535
rect 17219 32501 17253 32535
rect 20991 32501 21025 32535
rect 35619 32501 35653 32535
rect 41231 32501 41265 32535
rect 43991 32501 44025 32535
rect 44819 32501 44853 32535
rect 48646 32501 48680 32535
rect 49419 32501 49453 32535
rect 52639 32501 52673 32535
rect 58435 32501 58469 32535
rect 59723 32501 59757 32535
rect 65151 32501 65185 32535
rect 65473 32501 65507 32535
rect 71223 32501 71257 32535
rect 77203 32501 77237 32535
rect 83367 32501 83401 32535
rect 83551 32501 83585 32535
rect 86035 32501 86069 32535
rect 2499 32433 2533 32467
rect 14735 32433 14769 32467
rect 16207 32433 16241 32467
rect 21083 32433 21117 32467
rect 25499 32433 25533 32467
rect 41415 32433 41449 32467
rect 47579 32433 47613 32467
rect 48867 32433 48901 32467
rect 51259 32433 51293 32467
rect 58619 32433 58653 32467
rect 60183 32433 60217 32467
rect 64691 32433 64725 32467
rect 65703 32433 65737 32467
rect 70855 32433 70889 32467
rect 75455 32433 75489 32467
rect 75915 32433 75949 32467
rect 76099 32433 76133 32467
rect 80883 32433 80917 32467
rect 82171 32433 82205 32467
rect 83459 32433 83493 32467
rect 2775 32365 2809 32399
rect 5167 32365 5201 32399
rect 5259 32365 5293 32399
rect 7007 32365 7041 32399
rect 12803 32365 12837 32399
rect 12895 32365 12929 32399
rect 13171 32365 13205 32399
rect 13355 32365 13389 32399
rect 14183 32365 14217 32399
rect 14275 32365 14309 32399
rect 15986 32365 16020 32399
rect 17495 32365 17529 32399
rect 17771 32365 17805 32399
rect 20862 32365 20896 32399
rect 25223 32365 25257 32399
rect 33043 32365 33077 32399
rect 34331 32365 34365 32399
rect 34699 32365 34733 32399
rect 35435 32365 35469 32399
rect 38655 32365 38689 32399
rect 39023 32365 39057 32399
rect 40219 32365 40253 32399
rect 40771 32365 40805 32399
rect 41691 32365 41725 32399
rect 43899 32365 43933 32399
rect 44175 32365 44209 32399
rect 44635 32365 44669 32399
rect 47119 32365 47153 32399
rect 47211 32365 47245 32399
rect 47487 32365 47521 32399
rect 48729 32365 48763 32399
rect 49235 32365 49269 32399
rect 51535 32365 51569 32399
rect 53007 32365 53041 32399
rect 58803 32365 58837 32399
rect 59355 32365 59389 32399
rect 59539 32365 59573 32399
rect 60367 32365 60401 32399
rect 63311 32365 63345 32399
rect 63403 32365 63437 32399
rect 63863 32365 63897 32399
rect 64047 32365 64081 32399
rect 69475 32365 69509 32399
rect 69751 32365 69785 32399
rect 73615 32365 73649 32399
rect 73891 32365 73925 32399
rect 76283 32365 76317 32399
rect 76743 32365 76777 32399
rect 76835 32365 76869 32399
rect 81067 32365 81101 32399
rect 81619 32365 81653 32399
rect 81803 32365 81837 32399
rect 83091 32365 83125 32399
rect 12159 32297 12193 32331
rect 15839 32297 15873 32331
rect 20715 32297 20749 32331
rect 38471 32297 38505 32331
rect 40035 32297 40069 32331
rect 43071 32297 43105 32331
rect 46475 32297 46509 32331
rect 48499 32297 48533 32331
rect 64783 32297 64817 32331
rect 65335 32297 65369 32331
rect 86127 32365 86161 32399
rect 87323 32365 87357 32399
rect 87507 32365 87541 32399
rect 87783 32365 87817 32399
rect 25039 32229 25073 32263
rect 47763 32229 47797 32263
rect 47947 32229 47981 32263
rect 64967 32229 65001 32263
rect 74995 32229 75029 32263
rect 86035 32229 86069 32263
rect 86219 32229 86253 32263
rect 88887 32229 88921 32263
rect 5259 32025 5293 32059
rect 5995 32025 6029 32059
rect 12895 32025 12929 32059
rect 27523 32025 27557 32059
rect 41047 32025 41081 32059
rect 47027 32025 47061 32059
rect 82907 32025 82941 32059
rect 88151 32025 88185 32059
rect 92015 32025 92049 32059
rect 11975 31957 12009 31991
rect 16759 31957 16793 31991
rect 18231 31957 18265 31991
rect 18507 31957 18541 31991
rect 39483 31957 39517 31991
rect 47487 31957 47521 31991
rect 82815 31957 82849 31991
rect 5351 31889 5385 31923
rect 6363 31889 6397 31923
rect 6639 31889 6673 31923
rect 7743 31889 7777 31923
rect 7927 31889 7961 31923
rect 11239 31889 11273 31923
rect 11699 31889 11733 31923
rect 12711 31889 12745 31923
rect 12803 31889 12837 31923
rect 14735 31889 14769 31923
rect 16943 31889 16977 31923
rect 17127 31889 17161 31923
rect 17679 31889 17713 31923
rect 17863 31889 17897 31923
rect 19151 31889 19185 31923
rect 21819 31889 21853 31923
rect 22003 31889 22037 31923
rect 23843 31889 23877 31923
rect 26143 31889 26177 31923
rect 27891 31889 27925 31923
rect 28397 31889 28431 31923
rect 28673 31889 28707 31923
rect 28903 31889 28937 31923
rect 29271 31889 29305 31923
rect 29547 31889 29581 31923
rect 39575 31889 39609 31923
rect 40955 31889 40989 31923
rect 44359 31889 44393 31923
rect 44543 31889 44577 31923
rect 44727 31889 44761 31923
rect 45187 31889 45221 31923
rect 45279 31889 45313 31923
rect 46751 31889 46785 31923
rect 46935 31889 46969 31923
rect 48407 31889 48441 31923
rect 49879 31889 49913 31923
rect 51535 31889 51569 31923
rect 52915 31889 52949 31923
rect 54019 31889 54053 31923
rect 57791 31889 57825 31923
rect 58251 31889 58285 31923
rect 59631 31889 59665 31923
rect 63587 31889 63621 31923
rect 68647 31889 68681 31923
rect 69199 31889 69233 31923
rect 69383 31889 69417 31923
rect 70027 31889 70061 31923
rect 71775 31889 71809 31923
rect 72051 31889 72085 31923
rect 74259 31889 74293 31923
rect 74535 31889 74569 31923
rect 77019 31889 77053 31923
rect 77387 31889 77421 31923
rect 77663 31889 77697 31923
rect 78215 31889 78249 31923
rect 78399 31889 78433 31923
rect 80423 31889 80457 31923
rect 83275 31889 83309 31923
rect 83367 31889 83401 31923
rect 83735 31889 83769 31923
rect 83827 31889 83861 31923
rect 88335 31889 88369 31923
rect 90819 31889 90853 31923
rect 91003 31889 91037 31923
rect 91463 31889 91497 31923
rect 91555 31889 91589 31923
rect 5443 31821 5477 31855
rect 7099 31821 7133 31855
rect 12067 31821 12101 31855
rect 21727 31821 21761 31855
rect 22371 31821 22405 31855
rect 27983 31821 28017 31855
rect 29363 31821 29397 31855
rect 39299 31821 39333 31855
rect 40127 31821 40161 31855
rect 45831 31821 45865 31855
rect 48499 31821 48533 31855
rect 50155 31821 50189 31855
rect 58435 31821 58469 31855
rect 63955 31821 63989 31855
rect 64139 31821 64173 31855
rect 68555 31821 68589 31855
rect 77479 31821 77513 31855
rect 88611 31821 88645 31855
rect 6455 31753 6489 31787
rect 53007 31753 53041 31787
rect 57883 31753 57917 31787
rect 59815 31753 59849 31787
rect 63863 31753 63897 31787
rect 64507 31753 64541 31787
rect 69567 31753 69601 31787
rect 70211 31753 70245 31787
rect 6179 31685 6213 31719
rect 8019 31685 8053 31719
rect 14919 31685 14953 31719
rect 19335 31685 19369 31719
rect 21543 31685 21577 31719
rect 23751 31685 23785 31719
rect 24027 31685 24061 31719
rect 26235 31685 26269 31719
rect 27707 31685 27741 31719
rect 39759 31685 39793 31719
rect 46107 31685 46141 31719
rect 51719 31685 51753 31719
rect 54111 31685 54145 31719
rect 58803 31685 58837 31719
rect 63403 31685 63437 31719
rect 63752 31685 63786 31719
rect 68279 31685 68313 31719
rect 71867 31685 71901 31719
rect 74351 31685 74385 31719
rect 77203 31685 77237 31719
rect 78675 31685 78709 31719
rect 80607 31685 80641 31719
rect 84287 31685 84321 31719
rect 89715 31685 89749 31719
rect 3051 31481 3085 31515
rect 3511 31481 3545 31515
rect 5995 31481 6029 31515
rect 15287 31481 15321 31515
rect 15655 31481 15689 31515
rect 22095 31481 22129 31515
rect 24579 31481 24613 31515
rect 31847 31481 31881 31515
rect 40035 31481 40069 31515
rect 47027 31481 47061 31515
rect 51627 31481 51661 31515
rect 52087 31481 52121 31515
rect 68647 31481 68681 31515
rect 69015 31481 69049 31515
rect 74075 31481 74109 31515
rect 82907 31481 82941 31515
rect 88427 31481 88461 31515
rect 4983 31413 5017 31447
rect 26879 31413 26913 31447
rect 30099 31413 30133 31447
rect 51167 31413 51201 31447
rect 54341 31413 54375 31447
rect 54479 31413 54513 31447
rect 62851 31413 62885 31447
rect 82796 31413 82830 31447
rect 1671 31345 1705 31379
rect 1947 31345 1981 31379
rect 12987 31345 13021 31379
rect 15287 31345 15321 31379
rect 17219 31345 17253 31379
rect 17495 31345 17529 31379
rect 23935 31345 23969 31379
rect 28995 31345 29029 31379
rect 54568 31345 54602 31379
rect 68739 31345 68773 31379
rect 82999 31345 83033 31379
rect 90727 31345 90761 31379
rect 3603 31277 3637 31311
rect 5075 31277 5109 31311
rect 6363 31277 6397 31311
rect 6455 31277 6489 31311
rect 6639 31277 6673 31311
rect 7927 31277 7961 31311
rect 10503 31277 10537 31311
rect 12435 31277 12469 31311
rect 12527 31277 12561 31311
rect 15471 31277 15505 31311
rect 17679 31277 17713 31311
rect 18231 31277 18265 31311
rect 18415 31277 18449 31311
rect 19703 31277 19737 31311
rect 22003 31277 22037 31311
rect 23199 31277 23233 31311
rect 23843 31277 23877 31311
rect 24211 31277 24245 31311
rect 24395 31277 24429 31311
rect 26511 31277 26545 31311
rect 28719 31277 28753 31311
rect 32215 31277 32249 31311
rect 32307 31277 32341 31311
rect 32813 31277 32847 31311
rect 32951 31277 32985 31311
rect 35711 31277 35745 31311
rect 35895 31277 35929 31311
rect 36447 31277 36481 31311
rect 36631 31277 36665 31311
rect 39943 31277 39977 31311
rect 46935 31277 46969 31311
rect 51443 31277 51477 31311
rect 53007 31277 53041 31311
rect 57607 31277 57641 31311
rect 57883 31277 57917 31311
rect 59263 31277 59297 31311
rect 60091 31277 60125 31311
rect 60183 31277 60217 31311
rect 62667 31277 62701 31311
rect 66255 31277 66289 31311
rect 68371 31277 68405 31311
rect 68518 31277 68552 31311
rect 73615 31277 73649 31311
rect 73891 31277 73925 31311
rect 75363 31277 75397 31311
rect 80699 31277 80733 31311
rect 81251 31277 81285 31311
rect 81527 31277 81561 31311
rect 82631 31277 82665 31311
rect 83367 31277 83401 31311
rect 88335 31277 88369 31311
rect 90911 31277 90945 31311
rect 91371 31277 91405 31311
rect 91463 31277 91497 31311
rect 7099 31209 7133 31243
rect 26603 31209 26637 31243
rect 33319 31209 33353 31243
rect 36999 31209 37033 31243
rect 51351 31209 51385 31243
rect 54203 31209 54237 31243
rect 55031 31209 55065 31243
rect 73799 31209 73833 31243
rect 75179 31209 75213 31243
rect 75731 31209 75765 31243
rect 92015 31209 92049 31243
rect 5259 31141 5293 31175
rect 8111 31141 8145 31175
rect 10687 31141 10721 31175
rect 18691 31141 18725 31175
rect 18967 31141 19001 31175
rect 19887 31141 19921 31175
rect 22923 31141 22957 31175
rect 30467 31141 30501 31175
rect 33595 31141 33629 31175
rect 35527 31141 35561 31175
rect 53191 31141 53225 31175
rect 54847 31141 54881 31175
rect 65887 31141 65921 31175
rect 66071 31141 66105 31175
rect 68187 31141 68221 31175
rect 73339 31141 73373 31175
rect 80515 31141 80549 31175
rect 80791 31141 80825 31175
rect 4247 30937 4281 30971
rect 5259 30937 5293 30971
rect 15931 30937 15965 30971
rect 29179 30937 29213 30971
rect 82171 30937 82205 30971
rect 84839 30937 84873 30971
rect 88519 30937 88553 30971
rect 89715 30937 89749 30971
rect 10043 30869 10077 30903
rect 10503 30869 10537 30903
rect 10871 30869 10905 30903
rect 13355 30869 13389 30903
rect 21911 30869 21945 30903
rect 57607 30869 57641 30903
rect 63127 30869 63161 30903
rect 85759 30869 85793 30903
rect 88243 30869 88277 30903
rect 4339 30801 4373 30835
rect 5443 30801 5477 30835
rect 6547 30801 6581 30835
rect 6639 30801 6673 30835
rect 6823 30801 6857 30835
rect 10319 30801 10353 30835
rect 10411 30801 10445 30835
rect 12159 30801 12193 30835
rect 12343 30801 12377 30835
rect 12619 30801 12653 30835
rect 13171 30801 13205 30835
rect 16023 30801 16057 30835
rect 16207 30801 16241 30835
rect 16759 30801 16793 30835
rect 16943 30801 16977 30835
rect 18507 30801 18541 30835
rect 22095 30801 22129 30835
rect 27339 30801 27373 30835
rect 32951 30801 32985 30835
rect 35159 30801 35193 30835
rect 37459 30801 37493 30835
rect 44451 30801 44485 30835
rect 44911 30801 44945 30835
rect 45003 30801 45037 30835
rect 48407 30801 48441 30835
rect 52271 30801 52305 30835
rect 52363 30801 52397 30835
rect 52639 30801 52673 30835
rect 53191 30801 53225 30835
rect 54295 30801 54329 30835
rect 54571 30801 54605 30835
rect 55031 30801 55065 30835
rect 58159 30801 58193 30835
rect 58435 30801 58469 30835
rect 58619 30801 58653 30835
rect 62299 30801 62333 30835
rect 62483 30801 62517 30835
rect 62851 30801 62885 30835
rect 69015 30801 69049 30835
rect 71131 30801 71165 30835
rect 72879 30801 72913 30835
rect 73983 30801 74017 30835
rect 74167 30801 74201 30835
rect 74535 30801 74569 30835
rect 75363 30801 75397 30835
rect 75455 30801 75489 30835
rect 80699 30801 80733 30835
rect 80975 30801 81009 30835
rect 82079 30801 82113 30835
rect 84747 30801 84781 30835
rect 85943 30801 85977 30835
rect 88427 30801 88461 30835
rect 88887 30801 88921 30835
rect 89623 30801 89657 30835
rect 91371 30801 91405 30835
rect 7283 30733 7317 30767
rect 10135 30733 10169 30767
rect 11699 30733 11733 30767
rect 12987 30733 13021 30767
rect 13447 30733 13481 30767
rect 22371 30733 22405 30767
rect 27615 30733 27649 30767
rect 32675 30733 32709 30767
rect 37183 30733 37217 30767
rect 44083 30733 44117 30767
rect 44267 30733 44301 30767
rect 48775 30733 48809 30767
rect 48867 30733 48901 30767
rect 4523 30665 4557 30699
rect 17127 30665 17161 30699
rect 34975 30665 35009 30699
rect 35343 30665 35377 30699
rect 45831 30665 45865 30699
rect 52823 30733 52857 30767
rect 54387 30733 54421 30767
rect 62943 30733 62977 30767
rect 66531 30733 66565 30767
rect 66807 30733 66841 30767
rect 67911 30733 67945 30767
rect 71407 30733 71441 30767
rect 72511 30733 72545 30767
rect 77111 30733 77145 30767
rect 77387 30733 77421 30767
rect 78491 30733 78525 30767
rect 80147 30733 80181 30767
rect 81159 30733 81193 30767
rect 85023 30733 85057 30767
rect 52455 30665 52489 30699
rect 5627 30597 5661 30631
rect 17587 30597 17621 30631
rect 18691 30597 18725 30631
rect 23659 30597 23693 30631
rect 28719 30597 28753 30631
rect 34055 30597 34089 30631
rect 34423 30597 34457 30631
rect 36907 30597 36941 30631
rect 38563 30597 38597 30631
rect 45463 30597 45497 30631
rect 48545 30597 48579 30631
rect 48683 30597 48717 30631
rect 52271 30597 52305 30631
rect 69199 30597 69233 30631
rect 78859 30597 78893 30631
rect 86035 30597 86069 30631
rect 91555 30597 91589 30631
rect 3235 30393 3269 30427
rect 22371 30393 22405 30427
rect 27431 30393 27465 30427
rect 38103 30393 38137 30427
rect 48315 30393 48349 30427
rect 62207 30393 62241 30427
rect 66991 30393 67025 30427
rect 70947 30393 70981 30427
rect 82171 30393 82205 30427
rect 86771 30393 86805 30427
rect 87967 30393 88001 30427
rect 92107 30393 92141 30427
rect 8019 30325 8053 30359
rect 9675 30325 9709 30359
rect 24763 30325 24797 30359
rect 43991 30325 44025 30359
rect 44359 30325 44393 30359
rect 53651 30325 53685 30359
rect 60183 30325 60217 30359
rect 6455 30257 6489 30291
rect 7099 30257 7133 30291
rect 8663 30257 8697 30291
rect 13355 30257 13389 30291
rect 13631 30257 13665 30291
rect 18231 30257 18265 30291
rect 19611 30257 19645 30291
rect 23107 30257 23141 30291
rect 24395 30257 24429 30291
rect 27155 30257 27189 30291
rect 41139 30257 41173 30291
rect 41323 30257 41357 30291
rect 41507 30257 41541 30291
rect 42795 30257 42829 30291
rect 44083 30257 44117 30291
rect 47027 30257 47061 30291
rect 58251 30257 58285 30291
rect 58527 30257 58561 30291
rect 59631 30257 59665 30291
rect 1671 30189 1705 30223
rect 1947 30189 1981 30223
rect 5075 30189 5109 30223
rect 6363 30189 6397 30223
rect 6639 30189 6673 30223
rect 7927 30189 7961 30223
rect 8203 30189 8237 30223
rect 9491 30189 9525 30223
rect 12527 30189 12561 30223
rect 12619 30189 12653 30223
rect 12803 30189 12837 30223
rect 13263 30189 13297 30223
rect 17955 30189 17989 30223
rect 23567 30189 23601 30223
rect 23751 30189 23785 30223
rect 23935 30189 23969 30223
rect 24487 30189 24521 30223
rect 27247 30189 27281 30223
rect 34331 30189 34365 30223
rect 36907 30189 36941 30223
rect 37091 30189 37125 30223
rect 37551 30189 37585 30223
rect 37643 30189 37677 30223
rect 41691 30189 41725 30223
rect 42151 30189 42185 30223
rect 42243 30189 42277 30223
rect 43715 30189 43749 30223
rect 43862 30189 43896 30223
rect 47119 30189 47153 30223
rect 47303 30189 47337 30223
rect 47763 30189 47797 30223
rect 47855 30189 47889 30223
rect 52271 30189 52305 30223
rect 52547 30189 52581 30223
rect 54939 30189 54973 30223
rect 58619 30189 58653 30223
rect 59079 30189 59113 30223
rect 59171 30189 59205 30223
rect 59999 30189 60033 30223
rect 3419 30121 3453 30155
rect 11975 30121 12009 30155
rect 17771 30121 17805 30155
rect 22831 30121 22865 30155
rect 36723 30121 36757 30155
rect 54755 30121 54789 30155
rect 64415 30257 64449 30291
rect 71131 30257 71165 30291
rect 77571 30257 77605 30291
rect 62391 30189 62425 30223
rect 62667 30189 62701 30223
rect 64691 30189 64725 30223
rect 66899 30189 66933 30223
rect 68831 30189 68865 30223
rect 69935 30189 69969 30223
rect 71039 30189 71073 30223
rect 72143 30189 72177 30223
rect 72327 30189 72361 30223
rect 72695 30189 72729 30223
rect 73891 30189 73925 30223
rect 74259 30189 74293 30223
rect 76099 30189 76133 30223
rect 76191 30189 76225 30223
rect 76467 30189 76501 30223
rect 76651 30189 76685 30223
rect 77479 30189 77513 30223
rect 80791 30189 80825 30223
rect 81067 30189 81101 30223
rect 85391 30189 85425 30223
rect 85667 30189 85701 30223
rect 88519 30189 88553 30223
rect 88611 30189 88645 30223
rect 88887 30189 88921 30223
rect 89071 30189 89105 30223
rect 90635 30189 90669 30223
rect 90727 30189 90761 30223
rect 91003 30189 91037 30223
rect 62575 30121 62609 30155
rect 63127 30121 63161 30155
rect 68739 30121 68773 30155
rect 72879 30121 72913 30155
rect 74075 30121 74109 30155
rect 75455 30121 75489 30155
rect 89163 30121 89197 30155
rect 5259 30053 5293 30087
rect 22555 30053 22589 30087
rect 26971 30053 27005 30087
rect 34423 30053 34457 30087
rect 38379 30053 38413 30087
rect 38655 30053 38689 30087
rect 43071 30053 43105 30087
rect 43255 30053 43289 30087
rect 46751 30053 46785 30087
rect 54019 30053 54053 30087
rect 55031 30053 55065 30087
rect 62207 30053 62241 30087
rect 65795 30053 65829 30087
rect 69015 30053 69049 30087
rect 70119 30053 70153 30087
rect 74351 30053 74385 30087
rect 75363 30053 75397 30087
rect 80699 30053 80733 30087
rect 85207 30053 85241 30087
rect 87691 30053 87725 30087
rect 11607 29849 11641 29883
rect 12251 29849 12285 29883
rect 13079 29849 13113 29883
rect 17495 29849 17529 29883
rect 18783 29849 18817 29883
rect 33963 29849 33997 29883
rect 37367 29849 37401 29883
rect 39759 29849 39793 29883
rect 43991 29849 44025 29883
rect 48775 29849 48809 29883
rect 54295 29849 54329 29883
rect 55859 29849 55893 29883
rect 57515 29849 57549 29883
rect 60367 29849 60401 29883
rect 66807 29849 66841 29883
rect 67911 29849 67945 29883
rect 74719 29849 74753 29883
rect 78123 29849 78157 29883
rect 79871 29849 79905 29883
rect 84287 29849 84321 29883
rect 87783 29849 87817 29883
rect 5719 29781 5753 29815
rect 9307 29781 9341 29815
rect 9491 29781 9525 29815
rect 11515 29781 11549 29815
rect 11699 29781 11733 29815
rect 12067 29781 12101 29815
rect 27063 29781 27097 29815
rect 27523 29781 27557 29815
rect 29639 29781 29673 29815
rect 30467 29781 30501 29815
rect 32123 29781 32157 29815
rect 34147 29781 34181 29815
rect 50983 29781 51017 29815
rect 65795 29781 65829 29815
rect 66163 29781 66197 29815
rect 68739 29781 68773 29815
rect 73247 29781 73281 29815
rect 74535 29781 74569 29815
rect 76191 29781 76225 29815
rect 76467 29781 76501 29815
rect 80055 29781 80089 29815
rect 86035 29781 86069 29815
rect 6179 29713 6213 29747
rect 6363 29713 6397 29747
rect 6639 29713 6673 29747
rect 7191 29713 7225 29747
rect 9399 29713 9433 29747
rect 11331 29713 11365 29747
rect 12895 29713 12929 29747
rect 16391 29713 16425 29747
rect 18691 29713 18725 29747
rect 19059 29713 19093 29747
rect 23291 29713 23325 29747
rect 23475 29713 23509 29747
rect 23751 29713 23785 29747
rect 27983 29713 28017 29747
rect 28167 29713 28201 29747
rect 28351 29713 28385 29747
rect 28719 29713 28753 29747
rect 29823 29713 29857 29747
rect 29915 29713 29949 29747
rect 31663 29713 31697 29747
rect 32215 29713 32249 29747
rect 33779 29713 33813 29747
rect 37275 29713 37309 29747
rect 38563 29713 38597 29747
rect 38747 29713 38781 29747
rect 39207 29713 39241 29747
rect 39299 29713 39333 29747
rect 42427 29713 42461 29747
rect 42795 29713 42829 29747
rect 42979 29713 43013 29747
rect 43439 29713 43473 29747
rect 43531 29713 43565 29747
rect 48591 29713 48625 29747
rect 48959 29713 48993 29747
rect 51167 29713 51201 29747
rect 51535 29713 51569 29747
rect 52547 29713 52581 29747
rect 52639 29713 52673 29747
rect 54019 29713 54053 29747
rect 54203 29713 54237 29747
rect 54663 29713 54697 29747
rect 55583 29713 55617 29747
rect 55767 29713 55801 29747
rect 57699 29713 57733 29747
rect 60551 29713 60585 29747
rect 61379 29713 61413 29747
rect 62667 29713 62701 29747
rect 65335 29713 65369 29747
rect 65887 29713 65921 29747
rect 66715 29713 66749 29747
rect 67727 29713 67761 29747
rect 68923 29713 68957 29747
rect 69107 29713 69141 29747
rect 69291 29713 69325 29747
rect 70855 29713 70889 29747
rect 72695 29713 72729 29747
rect 72787 29713 72821 29747
rect 74879 29713 74913 29747
rect 74995 29713 75029 29747
rect 75180 29713 75214 29747
rect 78031 29713 78065 29747
rect 79043 29713 79077 29747
rect 79319 29713 79353 29747
rect 80239 29713 80273 29747
rect 84195 29713 84229 29747
rect 84471 29713 84505 29747
rect 86127 29713 86161 29747
rect 87691 29713 87725 29747
rect 90543 29713 90577 29747
rect 90727 29713 90761 29747
rect 6823 29645 6857 29679
rect 9123 29645 9157 29679
rect 9859 29645 9893 29679
rect 16115 29645 16149 29679
rect 22923 29645 22957 29679
rect 23935 29645 23969 29679
rect 27247 29645 27281 29679
rect 28903 29645 28937 29679
rect 30375 29645 30409 29679
rect 31571 29645 31605 29679
rect 42611 29645 42645 29679
rect 57883 29645 57917 29679
rect 62391 29645 62425 29679
rect 63771 29645 63805 29679
rect 65243 29645 65277 29679
rect 69659 29645 69693 29679
rect 75455 29645 75489 29679
rect 76835 29645 76869 29679
rect 79135 29645 79169 29679
rect 80607 29645 80641 29679
rect 85759 29645 85793 29679
rect 85851 29645 85885 29679
rect 86587 29645 86621 29679
rect 27339 29577 27373 29611
rect 53191 29577 53225 29611
rect 72327 29577 72361 29611
rect 72511 29577 72545 29611
rect 76605 29577 76639 29611
rect 15931 29509 15965 29543
rect 29179 29509 29213 29543
rect 38471 29509 38505 29543
rect 52363 29509 52397 29543
rect 52823 29509 52857 29543
rect 55399 29509 55433 29543
rect 61471 29509 61505 29543
rect 71039 29509 71073 29543
rect 76743 29509 76777 29543
rect 76927 29509 76961 29543
rect 90819 29509 90853 29543
rect 3051 29305 3085 29339
rect 8295 29305 8329 29339
rect 12987 29305 13021 29339
rect 13263 29305 13297 29339
rect 19151 29305 19185 29339
rect 22831 29305 22865 29339
rect 23107 29305 23141 29339
rect 23475 29305 23509 29339
rect 24395 29305 24429 29339
rect 36355 29305 36389 29339
rect 37735 29305 37769 29339
rect 41231 29305 41265 29339
rect 42795 29305 42829 29339
rect 48315 29305 48349 29339
rect 52823 29305 52857 29339
rect 62713 29305 62747 29339
rect 67543 29305 67577 29339
rect 67819 29305 67853 29339
rect 86679 29305 86713 29339
rect 87047 29305 87081 29339
rect 91003 29305 91037 29339
rect 18967 29237 19001 29271
rect 28903 29237 28937 29271
rect 31847 29237 31881 29271
rect 38287 29237 38321 29271
rect 45693 29237 45727 29271
rect 45831 29237 45865 29271
rect 59355 29237 59389 29271
rect 59999 29237 60033 29271
rect 76099 29237 76133 29271
rect 84931 29237 84965 29271
rect 90175 29237 90209 29271
rect 90543 29237 90577 29271
rect 6455 29169 6489 29203
rect 7191 29169 7225 29203
rect 8019 29169 8053 29203
rect 10227 29169 10261 29203
rect 23107 29169 23141 29203
rect 23935 29169 23969 29203
rect 30099 29169 30133 29203
rect 32031 29169 32065 29203
rect 41415 29169 41449 29203
rect 41599 29169 41633 29203
rect 45923 29169 45957 29203
rect 46843 29169 46877 29203
rect 47119 29169 47153 29203
rect 53559 29169 53593 29203
rect 54295 29169 54329 29203
rect 59815 29169 59849 29203
rect 62483 29169 62517 29203
rect 62943 29169 62977 29203
rect 64047 29169 64081 29203
rect 68003 29169 68037 29203
rect 69107 29169 69141 29203
rect 70119 29169 70153 29203
rect 71591 29169 71625 29203
rect 75087 29169 75121 29203
rect 80883 29169 80917 29203
rect 1671 29101 1705 29135
rect 1947 29101 1981 29135
rect 6639 29101 6673 29135
rect 8111 29101 8145 29135
rect 10411 29101 10445 29135
rect 10503 29101 10537 29135
rect 12895 29101 12929 29135
rect 17495 29101 17529 29135
rect 18875 29101 18909 29135
rect 23199 29101 23233 29135
rect 23291 29101 23325 29135
rect 24579 29101 24613 29135
rect 28811 29101 28845 29135
rect 29087 29101 29121 29135
rect 29179 29101 29213 29135
rect 29639 29101 29673 29135
rect 30467 29101 30501 29135
rect 30835 29101 30869 29135
rect 31019 29101 31053 29135
rect 31203 29101 31237 29135
rect 31387 29101 31421 29135
rect 36539 29101 36573 29135
rect 36723 29101 36757 29135
rect 37183 29101 37217 29135
rect 37275 29101 37309 29135
rect 38747 29101 38781 29135
rect 41783 29101 41817 29135
rect 42243 29101 42277 29135
rect 42335 29101 42369 29135
rect 43255 29101 43289 29135
rect 46935 29101 46969 29135
rect 47303 29101 47337 29135
rect 47763 29101 47797 29135
rect 47855 29101 47889 29135
rect 49327 29101 49361 29135
rect 51167 29101 51201 29135
rect 53651 29101 53685 29135
rect 54019 29101 54053 29135
rect 54203 29101 54237 29135
rect 55031 29101 55065 29135
rect 55123 29101 55157 29135
rect 58435 29101 58469 29135
rect 58527 29101 58561 29135
rect 58895 29101 58929 29135
rect 58987 29101 59021 29135
rect 60459 29101 60493 29135
rect 62805 29101 62839 29135
rect 64139 29101 64173 29135
rect 64323 29101 64357 29135
rect 68647 29101 68681 29135
rect 68739 29101 68773 29135
rect 69015 29101 69049 29135
rect 70027 29101 70061 29135
rect 71039 29101 71073 29135
rect 71131 29101 71165 29135
rect 73615 29101 73649 29135
rect 73891 29101 73925 29135
rect 74811 29101 74845 29135
rect 75823 29101 75857 29135
rect 76007 29101 76041 29135
rect 76283 29101 76317 29135
rect 77755 29101 77789 29135
rect 79871 29101 79905 29135
rect 81251 29101 81285 29135
rect 85023 29101 85057 29135
rect 85391 29101 85425 29135
rect 86587 29101 86621 29135
rect 90819 29101 90853 29135
rect 92107 29101 92141 29135
rect 6823 29033 6857 29067
rect 10595 29033 10629 29067
rect 10963 29033 10997 29067
rect 11147 29033 11181 29067
rect 45555 29033 45589 29067
rect 46291 29033 46325 29067
rect 53007 29033 53041 29067
rect 60551 29033 60585 29067
rect 62575 29033 62609 29067
rect 70855 29033 70889 29067
rect 74443 29033 74477 29067
rect 74627 29033 74661 29067
rect 76743 29033 76777 29067
rect 79687 29033 79721 29067
rect 80239 29033 80273 29067
rect 81067 29033 81101 29067
rect 84563 29033 84597 29067
rect 86403 29033 86437 29067
rect 90727 29033 90761 29067
rect 3419 28965 3453 28999
rect 6731 28965 6765 28999
rect 17587 28965 17621 28999
rect 24763 28965 24797 28999
rect 30283 28965 30317 28999
rect 38103 28965 38137 28999
rect 38839 28965 38873 28999
rect 43163 28965 43197 28999
rect 48683 28965 48717 28999
rect 49511 28965 49545 28999
rect 51259 28965 51293 28999
rect 58159 28965 58193 28999
rect 60827 28965 60861 28999
rect 63219 28965 63253 28999
rect 64415 28965 64449 28999
rect 69291 28965 69325 28999
rect 73707 28965 73741 28999
rect 77571 28965 77605 28999
rect 81343 28965 81377 28999
rect 92199 28965 92233 28999
rect 6731 28761 6765 28795
rect 13171 28761 13205 28795
rect 14919 28761 14953 28795
rect 24487 28761 24521 28795
rect 31663 28761 31697 28795
rect 34147 28761 34181 28795
rect 42887 28761 42921 28795
rect 56411 28761 56445 28795
rect 67359 28761 67393 28795
rect 68463 28761 68497 28795
rect 71591 28761 71625 28795
rect 72419 28761 72453 28795
rect 81067 28761 81101 28795
rect 85667 28761 85701 28795
rect 90543 28761 90577 28795
rect 91923 28761 91957 28795
rect 9123 28693 9157 28727
rect 9491 28693 9525 28727
rect 12987 28693 13021 28727
rect 17219 28693 17253 28727
rect 25775 28693 25809 28727
rect 36171 28693 36205 28727
rect 50155 28693 50189 28727
rect 61195 28693 61229 28727
rect 63771 28693 63805 28727
rect 73247 28693 73281 28727
rect 73523 28693 73557 28727
rect 6547 28625 6581 28659
rect 9307 28625 9341 28659
rect 9399 28625 9433 28659
rect 11515 28625 11549 28659
rect 11699 28625 11733 28659
rect 12067 28625 12101 28659
rect 12251 28625 12285 28659
rect 12527 28625 12561 28659
rect 14735 28625 14769 28659
rect 15103 28625 15137 28659
rect 15839 28625 15873 28659
rect 16115 28625 16149 28659
rect 17587 28625 17621 28659
rect 18139 28625 18173 28659
rect 18323 28625 18357 28659
rect 18967 28625 19001 28659
rect 22739 28625 22773 28659
rect 23475 28625 23509 28659
rect 23659 28625 23693 28659
rect 23843 28625 23877 28659
rect 24119 28625 24153 28659
rect 24763 28625 24797 28659
rect 25591 28625 25625 28659
rect 26971 28625 27005 28659
rect 27247 28625 27281 28659
rect 27523 28625 27557 28659
rect 27615 28625 27649 28659
rect 29179 28625 29213 28659
rect 29823 28625 29857 28659
rect 29915 28625 29949 28659
rect 30191 28625 30225 28659
rect 31571 28625 31605 28659
rect 38747 28625 38781 28659
rect 39207 28625 39241 28659
rect 39299 28625 39333 28659
rect 43163 28625 43197 28659
rect 43715 28625 43749 28659
rect 43899 28625 43933 28659
rect 49327 28625 49361 28659
rect 49695 28625 49729 28659
rect 50707 28625 50741 28659
rect 52087 28625 52121 28659
rect 52823 28625 52857 28659
rect 54019 28625 54053 28659
rect 55307 28625 55341 28659
rect 57515 28625 57549 28659
rect 59631 28625 59665 28659
rect 9859 28557 9893 28591
rect 15747 28557 15781 28591
rect 16023 28557 16057 28591
rect 17403 28557 17437 28591
rect 23107 28557 23141 28591
rect 26695 28557 26729 28591
rect 30283 28557 30317 28591
rect 30559 28557 30593 28591
rect 34423 28557 34457 28591
rect 34515 28557 34549 28591
rect 34791 28557 34825 28591
rect 38563 28557 38597 28591
rect 42979 28557 43013 28591
rect 49235 28557 49269 28591
rect 49787 28557 49821 28591
rect 52455 28557 52489 28591
rect 53007 28557 53041 28591
rect 55031 28557 55065 28591
rect 56779 28557 56813 28591
rect 11423 28489 11457 28523
rect 18507 28489 18541 28523
rect 23015 28489 23049 28523
rect 26327 28489 26361 28523
rect 26603 28489 26637 28523
rect 50063 28489 50097 28523
rect 50891 28489 50925 28523
rect 52252 28489 52286 28523
rect 63955 28625 63989 28659
rect 67175 28625 67209 28659
rect 68279 28625 68313 28659
rect 69383 28625 69417 28659
rect 71775 28625 71809 28659
rect 73339 28625 73373 28659
rect 73615 28625 73649 28659
rect 79411 28625 79445 28659
rect 79503 28625 79537 28659
rect 90083 28625 90117 28659
rect 90359 28625 90393 28659
rect 91647 28625 91681 28659
rect 91831 28625 91865 28659
rect 61287 28557 61321 28591
rect 61563 28557 61597 28591
rect 72143 28557 72177 28591
rect 74075 28557 74109 28591
rect 79779 28557 79813 28591
rect 84287 28557 84321 28591
rect 84563 28557 84597 28591
rect 62667 28489 62701 28523
rect 69475 28489 69509 28523
rect 72051 28489 72085 28523
rect 90175 28489 90209 28523
rect 16299 28421 16333 28455
rect 19059 28421 19093 28455
rect 19243 28421 19277 28455
rect 25407 28421 25441 28455
rect 28075 28421 28109 28455
rect 28351 28421 28385 28455
rect 28995 28421 29029 28455
rect 38379 28421 38413 28455
rect 39759 28421 39793 28455
rect 42611 28421 42645 28455
rect 44175 28421 44209 28455
rect 48775 28421 48809 28455
rect 52363 28421 52397 28455
rect 54111 28421 54145 28455
rect 57699 28421 57733 28455
rect 59815 28421 59849 28455
rect 61195 28421 61229 28455
rect 64047 28421 64081 28455
rect 71940 28421 71974 28455
rect 84195 28421 84229 28455
rect 3051 28217 3085 28251
rect 13539 28217 13573 28251
rect 15103 28217 15137 28251
rect 21819 28217 21853 28251
rect 50799 28217 50833 28251
rect 53835 28217 53869 28251
rect 63955 28217 63989 28251
rect 64415 28217 64449 28251
rect 75271 28217 75305 28251
rect 80423 28217 80457 28251
rect 89439 28217 89473 28251
rect 9215 28149 9249 28183
rect 13263 28149 13297 28183
rect 15379 28149 15413 28183
rect 24027 28149 24061 28183
rect 27707 28149 27741 28183
rect 31571 28149 31605 28183
rect 35435 28149 35469 28183
rect 40219 28149 40253 28183
rect 41783 28149 41817 28183
rect 56135 28149 56169 28183
rect 56227 28149 56261 28183
rect 58803 28149 58837 28183
rect 81343 28149 81377 28183
rect 83091 28149 83125 28183
rect 83183 28149 83217 28183
rect 1671 28081 1705 28115
rect 3511 28081 3545 28115
rect 6639 28081 6673 28115
rect 11883 28081 11917 28115
rect 16391 28081 16425 28115
rect 17771 28081 17805 28115
rect 17955 28081 17989 28115
rect 18231 28081 18265 28115
rect 19335 28081 19369 28115
rect 21083 28081 21117 28115
rect 24211 28081 24245 28115
rect 31203 28081 31237 28115
rect 34423 28081 34457 28115
rect 40587 28081 40621 28115
rect 42151 28081 42185 28115
rect 44359 28081 44393 28115
rect 48131 28081 48165 28115
rect 48407 28081 48441 28115
rect 52823 28081 52857 28115
rect 57883 28081 57917 28115
rect 57975 28081 58009 28115
rect 62759 28081 62793 28115
rect 72327 28081 72361 28115
rect 74167 28081 74201 28115
rect 79871 28081 79905 28115
rect 79963 28081 79997 28115
rect 83919 28081 83953 28115
rect 90175 28081 90209 28115
rect 91555 28081 91589 28115
rect 1947 28013 1981 28047
rect 6915 28013 6949 28047
rect 8295 28013 8329 28047
rect 9123 28013 9157 28047
rect 12067 28013 12101 28047
rect 12435 28013 12469 28047
rect 12711 28013 12745 28047
rect 12895 28013 12929 28047
rect 15655 28013 15689 28047
rect 15931 28013 15965 28047
rect 16299 28013 16333 28047
rect 20991 28013 21025 28047
rect 21195 28013 21229 28047
rect 21635 28013 21669 28047
rect 23107 28013 23141 28047
rect 24487 28013 24521 28047
rect 25867 28013 25901 28047
rect 27615 28013 27649 28047
rect 29547 28013 29581 28047
rect 29731 28013 29765 28047
rect 29915 28013 29949 28047
rect 30099 28013 30133 28047
rect 30467 28013 30501 28047
rect 30743 28013 30777 28047
rect 30835 28013 30869 28047
rect 33779 28013 33813 28047
rect 33963 28013 33997 28047
rect 34515 28013 34549 28047
rect 35067 28013 35101 28047
rect 35251 28013 35285 28047
rect 36539 28013 36573 28047
rect 40725 28013 40759 28047
rect 41231 28013 41265 28047
rect 41323 28013 41357 28047
rect 43071 28013 43105 28047
rect 43255 28013 43289 28047
rect 43715 28013 43749 28047
rect 43807 28013 43841 28047
rect 44543 28013 44577 28047
rect 49879 28013 49913 28047
rect 50063 28013 50097 28047
rect 51995 28013 52029 28047
rect 52179 28013 52213 28047
rect 52312 28013 52346 28047
rect 53743 28013 53777 28047
rect 56135 28013 56169 28047
rect 56595 28013 56629 28047
rect 57423 28013 57457 28047
rect 57699 28013 57733 28047
rect 58711 28013 58745 28047
rect 62667 28013 62701 28047
rect 62943 28013 62977 28047
rect 64231 28013 64265 28047
rect 68187 28013 68221 28047
rect 69567 28013 69601 28047
rect 69751 28013 69785 28047
rect 72235 28013 72269 28047
rect 72695 28013 72729 28047
rect 73891 28013 73925 28047
rect 75639 28013 75673 28047
rect 80239 28013 80273 28047
rect 81711 28013 81745 28047
rect 83367 28013 83401 28047
rect 83459 28013 83493 28047
rect 85667 28013 85701 28047
rect 85943 28013 85977 28047
rect 86127 28013 86161 28047
rect 89347 28013 89381 28047
rect 89623 28013 89657 28047
rect 91095 28013 91129 28047
rect 91187 28013 91221 28047
rect 91463 28013 91497 28047
rect 11699 27945 11733 27979
rect 36631 27945 36665 27979
rect 40403 27945 40437 27979
rect 46199 27945 46233 27979
rect 46291 27945 46325 27979
rect 50431 27945 50465 27979
rect 52731 27945 52765 27979
rect 53559 27945 53593 27979
rect 56871 27945 56905 27979
rect 64139 27945 64173 27979
rect 68003 27945 68037 27979
rect 70119 27945 70153 27979
rect 80147 27945 80181 27979
rect 81527 27945 81561 27979
rect 82079 27945 82113 27979
rect 85115 27945 85149 27979
rect 90451 27945 90485 27979
rect 8479 27877 8513 27911
rect 23291 27877 23325 27911
rect 42887 27877 42921 27911
rect 47579 27877 47613 27911
rect 49511 27877 49545 27911
rect 50523 27877 50557 27911
rect 53375 27877 53409 27911
rect 56411 27877 56445 27911
rect 68279 27877 68313 27911
rect 2315 27673 2349 27707
rect 7743 27673 7777 27707
rect 8111 27673 8145 27707
rect 8295 27673 8329 27707
rect 8479 27673 8513 27707
rect 15471 27673 15505 27707
rect 17863 27673 17897 27707
rect 22647 27673 22681 27707
rect 23475 27673 23509 27707
rect 24763 27673 24797 27707
rect 25131 27673 25165 27707
rect 30559 27673 30593 27707
rect 39299 27673 39333 27707
rect 42519 27673 42553 27707
rect 47395 27673 47429 27707
rect 54295 27673 54329 27707
rect 57331 27673 57365 27707
rect 67911 27673 67945 27707
rect 71315 27673 71349 27707
rect 78951 27673 78985 27707
rect 83827 27673 83861 27707
rect 90543 27673 90577 27707
rect 91739 27673 91773 27707
rect 19611 27605 19645 27639
rect 32031 27605 32065 27639
rect 45003 27605 45037 27639
rect 48499 27605 48533 27639
rect 50155 27605 50189 27639
rect 58619 27605 58653 27639
rect 61931 27605 61965 27639
rect 68187 27605 68221 27639
rect 74535 27605 74569 27639
rect 82171 27605 82205 27639
rect 90267 27605 90301 27639
rect 935 27537 969 27571
rect 6731 27537 6765 27571
rect 7283 27537 7317 27571
rect 7467 27537 7501 27571
rect 11515 27537 11549 27571
rect 11883 27537 11917 27571
rect 12067 27537 12101 27571
rect 12711 27537 12745 27571
rect 12895 27537 12929 27571
rect 15655 27537 15689 27571
rect 16023 27537 16057 27571
rect 16115 27537 16149 27571
rect 16483 27537 16517 27571
rect 16575 27537 16609 27571
rect 18231 27537 18265 27571
rect 18783 27537 18817 27571
rect 18967 27537 19001 27571
rect 22555 27537 22589 27571
rect 23751 27537 23785 27571
rect 24211 27537 24245 27571
rect 24303 27537 24337 27571
rect 27339 27537 27373 27571
rect 28903 27537 28937 27571
rect 30467 27537 30501 27571
rect 32675 27537 32709 27571
rect 33043 27537 33077 27571
rect 33227 27537 33261 27571
rect 35987 27537 36021 27571
rect 42795 27537 42829 27571
rect 42979 27537 43013 27571
rect 43439 27537 43473 27571
rect 43531 27537 43565 27571
rect 44543 27537 44577 27571
rect 47303 27537 47337 27571
rect 48407 27537 48441 27571
rect 49971 27537 50005 27571
rect 50247 27537 50281 27571
rect 51535 27537 51569 27571
rect 52087 27537 52121 27571
rect 54019 27537 54053 27571
rect 54203 27537 54237 27571
rect 57423 27537 57457 27571
rect 57791 27537 57825 27571
rect 61839 27537 61873 27571
rect 62207 27537 62241 27571
rect 63679 27537 63713 27571
rect 68095 27537 68129 27571
rect 68279 27537 68313 27571
rect 70947 27537 70981 27571
rect 74719 27537 74753 27571
rect 78123 27537 78157 27571
rect 79779 27537 79813 27571
rect 80147 27537 80181 27571
rect 82079 27537 82113 27571
rect 83183 27537 83217 27571
rect 83330 27537 83364 27571
rect 84563 27537 84597 27571
rect 84747 27537 84781 27571
rect 85299 27537 85333 27571
rect 87691 27537 87725 27571
rect 89255 27537 89289 27571
rect 90451 27537 90485 27571
rect 91647 27537 91681 27571
rect 1211 27469 1245 27503
rect 6639 27469 6673 27503
rect 11055 27469 11089 27503
rect 18047 27469 18081 27503
rect 23659 27469 23693 27503
rect 25223 27469 25257 27503
rect 27063 27469 27097 27503
rect 31939 27469 31973 27503
rect 32767 27469 32801 27503
rect 33411 27469 33445 27503
rect 37919 27469 37953 27503
rect 38195 27469 38229 27503
rect 44083 27469 44117 27503
rect 45150 27469 45184 27503
rect 45371 27469 45405 27503
rect 50707 27469 50741 27503
rect 51903 27469 51937 27503
rect 58067 27469 58101 27503
rect 58435 27469 58469 27503
rect 62851 27469 62885 27503
rect 63403 27469 63437 27503
rect 63863 27469 63897 27503
rect 69843 27469 69877 27503
rect 72051 27469 72085 27503
rect 72327 27469 72361 27503
rect 79871 27469 79905 27503
rect 80239 27469 80273 27503
rect 83551 27469 83585 27503
rect 84103 27469 84137 27503
rect 85759 27469 85793 27503
rect 87783 27469 87817 27503
rect 2775 27401 2809 27435
rect 6455 27401 6489 27435
rect 12251 27401 12285 27435
rect 13079 27401 13113 27435
rect 17311 27401 17345 27435
rect 19243 27401 19277 27435
rect 28627 27401 28661 27435
rect 35803 27401 35837 27435
rect 37735 27401 37769 27435
rect 39759 27401 39793 27435
rect 44359 27401 44393 27435
rect 45279 27401 45313 27435
rect 45647 27401 45681 27435
rect 73615 27401 73649 27435
rect 78215 27401 78249 27435
rect 83459 27401 83493 27435
rect 85023 27401 85057 27435
rect 2959 27333 2993 27367
rect 10871 27333 10905 27367
rect 15379 27333 15413 27367
rect 17035 27333 17069 27367
rect 31755 27333 31789 27367
rect 36171 27333 36205 27367
rect 50799 27333 50833 27367
rect 51351 27333 51385 27367
rect 68463 27333 68497 27367
rect 71131 27333 71165 27367
rect 71499 27333 71533 27367
rect 73799 27333 73833 27367
rect 74811 27333 74845 27367
rect 79227 27333 79261 27367
rect 89347 27333 89381 27367
rect 3879 27129 3913 27163
rect 9307 27129 9341 27163
rect 11699 27129 11733 27163
rect 13171 27129 13205 27163
rect 16483 27129 16517 27163
rect 16759 27129 16793 27163
rect 19611 27129 19645 27163
rect 33963 27129 33997 27163
rect 34055 27129 34089 27163
rect 34331 27129 34365 27163
rect 35711 27129 35745 27163
rect 43439 27129 43473 27163
rect 56503 27129 56537 27163
rect 58343 27129 58377 27163
rect 15011 27061 15045 27095
rect 16115 27061 16149 27095
rect 17863 27061 17897 27095
rect 25591 27061 25625 27095
rect 27983 27061 28017 27095
rect 29179 27061 29213 27095
rect 31571 27061 31605 27095
rect 32951 27061 32985 27095
rect 33043 27061 33077 27095
rect 52915 27061 52949 27095
rect 64967 27061 65001 27095
rect 66163 27061 66197 27095
rect 69383 27061 69417 27095
rect 70763 27061 70797 27095
rect 73707 27061 73741 27095
rect 75639 27061 75673 27095
rect 79043 27061 79077 27095
rect 87691 27061 87725 27095
rect 2315 26993 2349 27027
rect 12803 26993 12837 27027
rect 18323 26993 18357 27027
rect 23199 26993 23233 27027
rect 23935 26993 23969 27027
rect 24119 26993 24153 27027
rect 25315 26993 25349 27027
rect 29455 26993 29489 27027
rect 2591 26925 2625 26959
rect 4799 26925 4833 26959
rect 9399 26925 9433 26959
rect 9583 26925 9617 26959
rect 10135 26925 10169 26959
rect 10319 26925 10353 26959
rect 11975 26925 12009 26959
rect 12435 26925 12469 26959
rect 12711 26925 12745 26959
rect 13263 26925 13297 26959
rect 15195 26925 15229 26959
rect 16299 26925 16333 26959
rect 16391 26925 16425 26959
rect 18047 26925 18081 26959
rect 20531 26925 20565 26959
rect 20899 26925 20933 26959
rect 22923 26925 22957 26959
rect 23843 26925 23877 26959
rect 24211 26925 24245 26959
rect 24579 26925 24613 26959
rect 25223 26925 25257 26959
rect 27615 26925 27649 26959
rect 29915 26925 29949 26959
rect 30099 26925 30133 26959
rect 30467 26925 30501 26959
rect 30651 26925 30685 26959
rect 30743 26925 30777 26959
rect 31479 26925 31513 26959
rect 4155 26857 4189 26891
rect 10687 26857 10721 26891
rect 16943 26857 16977 26891
rect 27707 26857 27741 26891
rect 35895 26993 35929 27027
rect 43807 26993 43841 27027
rect 43991 26993 44025 27027
rect 48867 26993 48901 27027
rect 50155 26993 50189 27027
rect 51443 26993 51477 27027
rect 52547 26993 52581 27027
rect 56779 26993 56813 27027
rect 62391 26993 62425 27027
rect 62667 26993 62701 27027
rect 63771 26993 63805 27027
rect 65703 26993 65737 27027
rect 68003 26993 68037 27027
rect 68279 26993 68313 27027
rect 69751 26993 69785 27027
rect 70119 26993 70153 27027
rect 71683 26993 71717 27027
rect 74443 26993 74477 27027
rect 78215 26993 78249 27027
rect 79503 26993 79537 27027
rect 80607 26993 80641 27027
rect 85391 26993 85425 27027
rect 86587 26993 86621 27027
rect 90727 26993 90761 27027
rect 33227 26925 33261 26959
rect 36355 26925 36389 26959
rect 36539 26925 36573 26959
rect 36907 26925 36941 26959
rect 37091 26925 37125 26959
rect 42427 26925 42461 26959
rect 42519 26925 42553 26959
rect 42887 26925 42921 26959
rect 42979 26925 43013 26959
rect 48499 26925 48533 26959
rect 49879 26925 49913 26959
rect 51167 26925 51201 26959
rect 53651 26925 53685 26959
rect 57055 26925 57089 26959
rect 65059 26925 65093 26959
rect 65427 26925 65461 26959
rect 70671 26925 70705 26959
rect 72235 26925 72269 26959
rect 72511 26925 72545 26959
rect 72695 26925 72729 26959
rect 73063 26925 73097 26959
rect 73339 26925 73373 26959
rect 73799 26925 73833 26959
rect 74167 26925 74201 26959
rect 75547 26925 75581 26959
rect 78123 26925 78157 26959
rect 79227 26925 79261 26959
rect 85023 26925 85057 26959
rect 85483 26925 85517 26959
rect 86219 26925 86253 26959
rect 86311 26925 86345 26959
rect 90267 26925 90301 26959
rect 90451 26925 90485 26959
rect 92107 26925 92141 26959
rect 35619 26857 35653 26891
rect 48315 26857 48349 26891
rect 49695 26857 49729 26891
rect 53743 26857 53777 26891
rect 70303 26857 70337 26891
rect 70579 26857 70613 26891
rect 70947 26857 70981 26891
rect 71223 26857 71257 26891
rect 71315 26857 71349 26891
rect 71499 26857 71533 26891
rect 84839 26857 84873 26891
rect 4983 26789 5017 26823
rect 20715 26789 20749 26823
rect 29271 26789 29305 26823
rect 32951 26789 32985 26823
rect 69935 26789 69969 26823
rect 3971 26585 4005 26619
rect 7283 26585 7317 26619
rect 38103 26585 38137 26619
rect 38287 26585 38321 26619
rect 37183 26517 37217 26551
rect 3695 26449 3729 26483
rect 5535 26449 5569 26483
rect 34423 26449 34457 26483
rect 34607 26449 34641 26483
rect 35159 26449 35193 26483
rect 35343 26449 35377 26483
rect 35895 26449 35929 26483
rect 37091 26449 37125 26483
rect 38839 26449 38873 26483
rect 39299 26449 39333 26483
rect 39391 26449 39425 26483
rect 5811 26381 5845 26415
rect 38563 26381 38597 26415
rect 38655 26381 38689 26415
rect 7099 26313 7133 26347
rect 3787 26245 3821 26279
rect 35619 26245 35653 26279
rect 39851 26245 39885 26279
rect 3879 26041 3913 26075
rect 6639 26041 6673 26075
rect 35987 26041 36021 26075
rect 36723 26041 36757 26075
rect 42059 26041 42093 26075
rect 2591 25905 2625 25939
rect 34699 25905 34733 25939
rect 36631 25905 36665 25939
rect 2867 25837 2901 25871
rect 2959 25837 2993 25871
rect 3419 25837 3453 25871
rect 3603 25837 3637 25871
rect 6271 25837 6305 25871
rect 34423 25837 34457 25871
rect 36907 25837 36941 25871
rect 37367 25837 37401 25871
rect 37551 25837 37585 25871
rect 37919 25837 37953 25871
rect 38011 25837 38045 25871
rect 40955 25837 40989 25871
rect 41967 25837 42001 25871
rect 6363 25769 6397 25803
rect 41047 25701 41081 25735
rect 5811 25429 5845 25463
rect 34423 25429 34457 25463
rect 39943 25429 39977 25463
rect 41783 25429 41817 25463
rect 3511 25361 3545 25395
rect 4707 25361 4741 25395
rect 5259 25361 5293 25395
rect 5443 25361 5477 25395
rect 37459 25361 37493 25395
rect 37643 25361 37677 25395
rect 38103 25361 38137 25395
rect 38655 25361 38689 25395
rect 38839 25361 38873 25395
rect 40127 25361 40161 25395
rect 4431 25293 4465 25327
rect 4615 25293 4649 25327
rect 37735 25293 37769 25327
rect 37919 25293 37953 25327
rect 39207 25293 39241 25327
rect 40403 25293 40437 25327
rect 3603 25225 3637 25259
rect 3879 25157 3913 25191
rect 1855 24953 1889 24987
rect 35159 24953 35193 24987
rect 42243 24953 42277 24987
rect 7283 24885 7317 24919
rect 7559 24885 7593 24919
rect 9031 24885 9065 24919
rect 35987 24885 36021 24919
rect 2775 24817 2809 24851
rect 1671 24749 1705 24783
rect 3051 24749 3085 24783
rect 7099 24749 7133 24783
rect 4431 24681 4465 24715
rect 35619 24817 35653 24851
rect 35803 24817 35837 24851
rect 36171 24817 36205 24851
rect 40955 24817 40989 24851
rect 35343 24749 35377 24783
rect 36355 24749 36389 24783
rect 36907 24749 36941 24783
rect 37091 24749 37125 24783
rect 40679 24749 40713 24783
rect 21543 24681 21577 24715
rect 34975 24681 35009 24715
rect 37459 24681 37493 24715
rect 2131 24613 2165 24647
rect 4615 24613 4649 24647
rect 9031 24613 9065 24647
rect 21451 24613 21485 24647
rect 40495 24613 40529 24647
rect 4707 24409 4741 24443
rect 37183 24409 37217 24443
rect 3327 24341 3361 24375
rect 5075 24341 5109 24375
rect 7559 24341 7593 24375
rect 3695 24273 3729 24307
rect 3787 24273 3821 24307
rect 4155 24273 4189 24307
rect 4247 24273 4281 24307
rect 5995 24273 6029 24307
rect 35343 24273 35377 24307
rect 37091 24273 37125 24307
rect 37367 24273 37401 24307
rect 5719 24205 5753 24239
rect 35159 24137 35193 24171
rect 7283 24069 7317 24103
rect 7559 23865 7593 23899
rect 34515 23865 34549 23899
rect 34699 23865 34733 23899
rect 34883 23865 34917 23899
rect 37091 23865 37125 23899
rect 2039 23729 2073 23763
rect 33963 23729 33997 23763
rect 35067 23729 35101 23763
rect 36355 23729 36389 23763
rect 37551 23729 37585 23763
rect 2315 23661 2349 23695
rect 2407 23661 2441 23695
rect 2867 23661 2901 23695
rect 3051 23661 3085 23695
rect 7191 23661 7225 23695
rect 3327 23525 3361 23559
rect 7283 23525 7317 23559
rect 35251 23661 35285 23695
rect 35711 23661 35745 23695
rect 35803 23661 35837 23695
rect 37275 23661 37309 23695
rect 36539 23593 36573 23627
rect 38839 23525 38873 23559
rect 3603 23321 3637 23355
rect 6547 23321 6581 23355
rect 33963 23321 33997 23355
rect 34791 23321 34825 23355
rect 39483 23321 39517 23355
rect 6455 23253 6489 23287
rect 3511 23185 3545 23219
rect 4799 23185 4833 23219
rect 34423 23185 34457 23219
rect 34975 23185 35009 23219
rect 38195 23185 38229 23219
rect 40495 23185 40529 23219
rect 5075 23117 5109 23151
rect 37919 23117 37953 23151
rect 40863 23117 40897 23151
rect 3787 22981 3821 23015
rect 34607 22981 34641 23015
rect 37735 22981 37769 23015
rect 40587 22981 40621 23015
rect 6639 22777 6673 22811
rect 34607 22777 34641 22811
rect 3235 22709 3269 22743
rect 1947 22641 1981 22675
rect 3419 22641 3453 22675
rect 42335 22641 42369 22675
rect 1671 22573 1705 22607
rect 4247 22573 4281 22607
rect 6271 22573 6305 22607
rect 33963 22573 33997 22607
rect 34423 22573 34457 22607
rect 34975 22573 35009 22607
rect 37367 22573 37401 22607
rect 37551 22573 37585 22607
rect 38655 22573 38689 22607
rect 40679 22573 40713 22607
rect 40955 22573 40989 22607
rect 6363 22505 6397 22539
rect 4431 22437 4465 22471
rect 3695 22233 3729 22267
rect 7191 22233 7225 22267
rect 2315 22097 2349 22131
rect 3971 22097 4005 22131
rect 4523 22097 4557 22131
rect 4707 22097 4741 22131
rect 6179 22097 6213 22131
rect 6271 22097 6305 22131
rect 6639 22097 6673 22131
rect 6731 22097 6765 22131
rect 3879 22029 3913 22063
rect 5903 22029 5937 22063
rect 2499 21893 2533 21927
rect 4983 21893 5017 21927
rect 38747 22505 38781 22539
rect 34791 22437 34825 22471
rect 37735 22437 37769 22471
rect 40495 22437 40529 22471
rect 43071 22437 43105 22471
rect 39575 22233 39609 22267
rect 40955 22233 40989 22267
rect 35343 22097 35377 22131
rect 35619 22097 35653 22131
rect 39943 22097 39977 22131
rect 40495 22097 40529 22131
rect 40679 22097 40713 22131
rect 39759 22029 39793 22063
rect 35435 21893 35469 21927
rect 3695 21689 3729 21723
rect 33963 21689 33997 21723
rect 34975 21689 35009 21723
rect 35527 21689 35561 21723
rect 3879 21553 3913 21587
rect 35619 21553 35653 21587
rect 36999 21553 37033 21587
rect 2683 21485 2717 21519
rect 3971 21485 4005 21519
rect 4523 21485 4557 21519
rect 4707 21485 4741 21519
rect 34423 21485 34457 21519
rect 35895 21485 35929 21519
rect 39851 21485 39885 21519
rect 40127 21485 40161 21519
rect 5075 21417 5109 21451
rect 2867 21349 2901 21383
rect 34607 21349 34641 21383
rect 34791 21349 34825 21383
rect 39943 21349 39977 21383
rect 43071 21349 43105 21383
rect 7099 21145 7133 21179
rect 34423 21145 34457 21179
rect 37551 21145 37585 21179
rect 39759 21145 39793 21179
rect 6179 21077 6213 21111
rect 6915 21077 6949 21111
rect 35895 21077 35929 21111
rect 39023 21077 39057 21111
rect 4523 21009 4557 21043
rect 6363 21009 6397 21043
rect 7007 21009 7041 21043
rect 34607 21009 34641 21043
rect 34791 21009 34825 21043
rect 35251 21009 35285 21043
rect 35343 21009 35377 21043
rect 37919 21009 37953 21043
rect 38471 21009 38505 21043
rect 38655 21009 38689 21043
rect 40219 21009 40253 21043
rect 4799 20941 4833 20975
rect 37735 20941 37769 20975
rect 39943 20941 39977 20975
rect 41507 20805 41541 20839
rect 2407 20601 2441 20635
rect 6363 20601 6397 20635
rect 36079 20601 36113 20635
rect 40403 20601 40437 20635
rect 40495 20601 40529 20635
rect 2591 20465 2625 20499
rect 2775 20397 2809 20431
rect 3327 20397 3361 20431
rect 3511 20397 3545 20431
rect 6271 20397 6305 20431
rect 36263 20397 36297 20431
rect 40403 20397 40437 20431
rect 40679 20397 40713 20431
rect 40955 20397 40989 20431
rect 3879 20329 3913 20363
rect 42335 20329 42369 20363
rect 6639 20261 6673 20295
rect 34423 20261 34457 20295
rect 36447 20261 36481 20295
rect 43071 20261 43105 20295
rect 39115 20057 39149 20091
rect 6823 19989 6857 20023
rect 5443 19921 5477 19955
rect 39391 19921 39425 19955
rect 39851 19921 39885 19955
rect 39943 19921 39977 19955
rect 41599 19921 41633 19955
rect 5167 19853 5201 19887
rect 39207 19853 39241 19887
rect 40495 19853 40529 19887
rect 40679 19785 40713 19819
rect 41691 19785 41725 19819
rect 7007 19717 7041 19751
rect 4247 19513 4281 19547
rect 34607 19513 34641 19547
rect 35527 19513 35561 19547
rect 37367 19513 37401 19547
rect 1947 19377 1981 19411
rect 37459 19377 37493 19411
rect 39023 19377 39057 19411
rect 39943 19377 39977 19411
rect 1671 19309 1705 19343
rect 3327 19309 3361 19343
rect 3971 19309 4005 19343
rect 4155 19309 4189 19343
rect 35435 19309 35469 19343
rect 37643 19309 37677 19343
rect 38195 19309 38229 19343
rect 38379 19309 38413 19343
rect 39851 19309 39885 19343
rect 38747 19241 38781 19275
rect 3511 19173 3545 19207
rect 34423 19173 34457 19207
rect 5903 18969 5937 19003
rect 39023 18969 39057 19003
rect 40679 18969 40713 19003
rect 3327 18901 3361 18935
rect 3695 18833 3729 18867
rect 3787 18833 3821 18867
rect 4247 18833 4281 18867
rect 4431 18833 4465 18867
rect 5995 18833 6029 18867
rect 6179 18833 6213 18867
rect 6731 18833 6765 18867
rect 6915 18833 6949 18867
rect 34423 18833 34457 18867
rect 34592 18833 34626 18867
rect 35067 18833 35101 18867
rect 35159 18833 35193 18867
rect 39115 18833 39149 18867
rect 39391 18833 39425 18867
rect 4615 18697 4649 18731
rect 7099 18697 7133 18731
rect 35527 18697 35561 18731
rect 7283 18425 7317 18459
rect 36631 18425 36665 18459
rect 40311 18425 40345 18459
rect 3971 18289 4005 18323
rect 34791 18289 34825 18323
rect 35067 18289 35101 18323
rect 40495 18289 40529 18323
rect 3695 18221 3729 18255
rect 7191 18221 7225 18255
rect 40771 18221 40805 18255
rect 36447 18153 36481 18187
rect 5075 18085 5109 18119
rect 5535 18085 5569 18119
rect 7467 18085 7501 18119
rect 34423 18085 34457 18119
rect 42059 18085 42093 18119
rect 4799 17881 4833 17915
rect 41047 17881 41081 17915
rect 40771 17813 40805 17847
rect 4707 17745 4741 17779
rect 5995 17745 6029 17779
rect 38655 17745 38689 17779
rect 39207 17745 39241 17779
rect 39391 17745 39425 17779
rect 40679 17745 40713 17779
rect 5719 17677 5753 17711
rect 7467 17677 7501 17711
rect 38471 17677 38505 17711
rect 39759 17677 39793 17711
rect 5075 17541 5109 17575
rect 7283 17541 7317 17575
rect 38287 17541 38321 17575
rect 37275 17201 37309 17235
rect 35987 17133 36021 17167
rect 36171 17133 36205 17167
rect 36631 17133 36665 17167
rect 36723 17133 36757 17167
rect 38747 17133 38781 17167
rect 39023 17133 39057 17167
rect 39851 17133 39885 17167
rect 40035 17133 40069 17167
rect 40587 17133 40621 17167
rect 40771 17133 40805 17167
rect 38839 17065 38873 17099
rect 34423 16997 34457 17031
rect 35895 16997 35929 17031
rect 39575 16997 39609 17031
rect 41047 16997 41081 17031
rect 5075 16793 5109 16827
rect 5259 16793 5293 16827
rect 37643 16793 37677 16827
rect 39851 16793 39885 16827
rect 5811 16657 5845 16691
rect 6363 16657 6397 16691
rect 6547 16657 6581 16691
rect 37551 16657 37585 16691
rect 40311 16657 40345 16691
rect 5535 16589 5569 16623
rect 5719 16589 5753 16623
rect 40035 16589 40069 16623
rect 41691 16589 41725 16623
rect 6731 16521 6765 16555
rect 5443 16249 5477 16283
rect 5627 16249 5661 16283
rect 36355 16249 36389 16283
rect 3879 16181 3913 16215
rect 4063 16113 4097 16147
rect 6547 16113 6581 16147
rect 36539 16113 36573 16147
rect 4155 16045 4189 16079
rect 4707 16045 4741 16079
rect 4891 16045 4925 16079
rect 6455 16045 6489 16079
rect 36723 16045 36757 16079
rect 37183 16045 37217 16079
rect 37275 16045 37309 16079
rect 38747 16045 38781 16079
rect 5259 15977 5293 16011
rect 38839 15977 38873 16011
rect 6823 15909 6857 15943
rect 37735 15909 37769 15943
rect 36815 15705 36849 15739
rect 5719 15569 5753 15603
rect 37091 15569 37125 15603
rect 37367 15569 37401 15603
rect 5443 15501 5477 15535
rect 7191 15501 7225 15535
rect 7007 15365 7041 15399
rect 38655 15365 38689 15399
rect 7191 15161 7225 15195
rect 37091 15161 37125 15195
rect 37275 15025 37309 15059
rect 37551 15025 37585 15059
rect 7099 14957 7133 14991
rect 38931 14889 38965 14923
rect 7375 14821 7409 14855
rect 34423 14821 34457 14855
rect 7467 14617 7501 14651
rect 5719 14481 5753 14515
rect 5995 14481 6029 14515
rect 7375 14481 7409 14515
rect 34423 10469 34457 10503
rect 7559 10197 7593 10231
rect 5719 10129 5753 10163
rect 7651 10129 7685 10163
rect 5995 10061 6029 10095
rect 7099 9925 7133 9959
rect 43071 2649 43105 2683
rect 34423 2309 34457 2343
<< metal1 >>
rect 538 41962 93642 41984
rect 538 41910 6344 41962
rect 6396 41910 6408 41962
rect 6460 41910 6472 41962
rect 6524 41910 6536 41962
rect 6588 41910 11672 41962
rect 11724 41910 11736 41962
rect 11788 41910 11800 41962
rect 11852 41910 11864 41962
rect 11916 41910 17000 41962
rect 17052 41910 17064 41962
rect 17116 41910 17128 41962
rect 17180 41910 17192 41962
rect 17244 41910 22328 41962
rect 22380 41910 22392 41962
rect 22444 41910 22456 41962
rect 22508 41910 22520 41962
rect 22572 41910 27656 41962
rect 27708 41910 27720 41962
rect 27772 41910 27784 41962
rect 27836 41910 27848 41962
rect 27900 41910 32984 41962
rect 33036 41910 33048 41962
rect 33100 41910 33112 41962
rect 33164 41910 33176 41962
rect 33228 41910 38312 41962
rect 38364 41910 38376 41962
rect 38428 41910 38440 41962
rect 38492 41910 38504 41962
rect 38556 41910 43640 41962
rect 43692 41910 43704 41962
rect 43756 41910 43768 41962
rect 43820 41910 43832 41962
rect 43884 41910 48968 41962
rect 49020 41910 49032 41962
rect 49084 41910 49096 41962
rect 49148 41910 49160 41962
rect 49212 41910 54296 41962
rect 54348 41910 54360 41962
rect 54412 41910 54424 41962
rect 54476 41910 54488 41962
rect 54540 41910 59624 41962
rect 59676 41910 59688 41962
rect 59740 41910 59752 41962
rect 59804 41910 59816 41962
rect 59868 41910 64952 41962
rect 65004 41910 65016 41962
rect 65068 41910 65080 41962
rect 65132 41910 65144 41962
rect 65196 41910 70280 41962
rect 70332 41910 70344 41962
rect 70396 41910 70408 41962
rect 70460 41910 70472 41962
rect 70524 41910 75608 41962
rect 75660 41910 75672 41962
rect 75724 41910 75736 41962
rect 75788 41910 75800 41962
rect 75852 41910 80936 41962
rect 80988 41910 81000 41962
rect 81052 41910 81064 41962
rect 81116 41910 81128 41962
rect 81180 41910 86264 41962
rect 86316 41910 86328 41962
rect 86380 41910 86392 41962
rect 86444 41910 86456 41962
rect 86508 41910 91592 41962
rect 91644 41910 91656 41962
rect 91708 41910 91720 41962
rect 91772 41910 91784 41962
rect 91836 41910 93642 41962
rect 538 41888 93642 41910
rect 65320 41604 65326 41656
rect 65378 41644 65384 41656
rect 66059 41647 66117 41653
rect 66059 41644 66071 41647
rect 65378 41616 66071 41644
rect 65378 41604 65384 41616
rect 66059 41613 66071 41616
rect 66105 41644 66117 41647
rect 66243 41647 66301 41653
rect 66243 41644 66255 41647
rect 66105 41616 66255 41644
rect 66105 41613 66117 41616
rect 66059 41607 66117 41613
rect 66243 41613 66255 41616
rect 66289 41613 66301 41647
rect 66243 41607 66301 41613
rect 66519 41647 66577 41653
rect 66519 41613 66531 41647
rect 66565 41644 66577 41647
rect 68540 41644 68546 41656
rect 66565 41616 68546 41644
rect 66565 41613 66577 41616
rect 66519 41607 66577 41613
rect 68540 41604 68546 41616
rect 68598 41604 68604 41656
rect 88136 41604 88142 41656
rect 88194 41644 88200 41656
rect 88875 41647 88933 41653
rect 88875 41644 88887 41647
rect 88194 41616 88887 41644
rect 88194 41604 88200 41616
rect 88875 41613 88887 41616
rect 88921 41644 88933 41647
rect 89059 41647 89117 41653
rect 89059 41644 89071 41647
rect 88921 41616 89071 41644
rect 88921 41613 88933 41616
rect 88875 41607 88933 41613
rect 89059 41613 89071 41616
rect 89105 41613 89117 41647
rect 89332 41644 89338 41656
rect 89293 41616 89338 41644
rect 89059 41607 89117 41613
rect 89332 41604 89338 41616
rect 89390 41604 89396 41656
rect 3496 41468 3502 41520
rect 3554 41508 3560 41520
rect 20608 41508 20614 41520
rect 3554 41480 20614 41508
rect 3554 41468 3560 41480
rect 20608 41468 20614 41480
rect 20666 41468 20672 41520
rect 67436 41468 67442 41520
rect 67494 41508 67500 41520
rect 67623 41511 67681 41517
rect 67623 41508 67635 41511
rect 67494 41480 67635 41508
rect 67494 41468 67500 41480
rect 67623 41477 67635 41480
rect 67669 41477 67681 41511
rect 67623 41471 67681 41477
rect 73232 41468 73238 41520
rect 73290 41508 73296 41520
rect 90439 41511 90497 41517
rect 90439 41508 90451 41511
rect 73290 41480 90451 41508
rect 73290 41468 73296 41480
rect 90439 41477 90451 41480
rect 90485 41477 90497 41511
rect 90439 41471 90497 41477
rect 538 41418 93642 41440
rect 538 41366 3680 41418
rect 3732 41366 3744 41418
rect 3796 41366 3808 41418
rect 3860 41366 3872 41418
rect 3924 41366 9008 41418
rect 9060 41366 9072 41418
rect 9124 41366 9136 41418
rect 9188 41366 9200 41418
rect 9252 41366 14336 41418
rect 14388 41366 14400 41418
rect 14452 41366 14464 41418
rect 14516 41366 14528 41418
rect 14580 41366 19664 41418
rect 19716 41366 19728 41418
rect 19780 41366 19792 41418
rect 19844 41366 19856 41418
rect 19908 41366 24992 41418
rect 25044 41366 25056 41418
rect 25108 41366 25120 41418
rect 25172 41366 25184 41418
rect 25236 41366 30320 41418
rect 30372 41366 30384 41418
rect 30436 41366 30448 41418
rect 30500 41366 30512 41418
rect 30564 41366 35648 41418
rect 35700 41366 35712 41418
rect 35764 41366 35776 41418
rect 35828 41366 35840 41418
rect 35892 41366 40976 41418
rect 41028 41366 41040 41418
rect 41092 41366 41104 41418
rect 41156 41366 41168 41418
rect 41220 41366 46304 41418
rect 46356 41366 46368 41418
rect 46420 41366 46432 41418
rect 46484 41366 46496 41418
rect 46548 41366 51632 41418
rect 51684 41366 51696 41418
rect 51748 41366 51760 41418
rect 51812 41366 51824 41418
rect 51876 41366 56960 41418
rect 57012 41366 57024 41418
rect 57076 41366 57088 41418
rect 57140 41366 57152 41418
rect 57204 41366 62288 41418
rect 62340 41366 62352 41418
rect 62404 41366 62416 41418
rect 62468 41366 62480 41418
rect 62532 41366 67616 41418
rect 67668 41366 67680 41418
rect 67732 41366 67744 41418
rect 67796 41366 67808 41418
rect 67860 41366 72944 41418
rect 72996 41366 73008 41418
rect 73060 41366 73072 41418
rect 73124 41366 73136 41418
rect 73188 41366 78272 41418
rect 78324 41366 78336 41418
rect 78388 41366 78400 41418
rect 78452 41366 78464 41418
rect 78516 41366 83600 41418
rect 83652 41366 83664 41418
rect 83716 41366 83728 41418
rect 83780 41366 83792 41418
rect 83844 41366 88928 41418
rect 88980 41366 88992 41418
rect 89044 41366 89056 41418
rect 89108 41366 89120 41418
rect 89172 41366 93642 41418
rect 538 41344 93642 41366
rect 2392 41264 2398 41316
rect 2450 41304 2456 41316
rect 3039 41307 3097 41313
rect 3039 41304 3051 41307
rect 2450 41276 3051 41304
rect 2450 41264 2456 41276
rect 3039 41273 3051 41276
rect 3085 41273 3097 41307
rect 3496 41304 3502 41316
rect 3457 41276 3502 41304
rect 3039 41267 3097 41273
rect 3496 41264 3502 41276
rect 3554 41264 3560 41316
rect 17388 41264 17394 41316
rect 17446 41304 17452 41316
rect 18863 41307 18921 41313
rect 18863 41304 18875 41307
rect 17446 41276 18875 41304
rect 17446 41264 17452 41276
rect 18863 41273 18875 41276
rect 18909 41273 18921 41307
rect 18863 41267 18921 41273
rect 24380 41264 24386 41316
rect 24438 41304 24444 41316
rect 24475 41307 24533 41313
rect 24475 41304 24487 41307
rect 24438 41276 24487 41304
rect 24438 41264 24444 41276
rect 24475 41273 24487 41276
rect 24521 41273 24533 41307
rect 24475 41267 24533 41273
rect 27048 41264 27054 41316
rect 27106 41304 27112 41316
rect 27143 41307 27201 41313
rect 27143 41304 27155 41307
rect 27106 41276 27155 41304
rect 27106 41264 27112 41276
rect 27143 41273 27155 41276
rect 27189 41273 27201 41307
rect 27143 41267 27201 41273
rect 30271 41307 30329 41313
rect 30271 41273 30283 41307
rect 30317 41304 30329 41307
rect 31740 41304 31746 41316
rect 30317 41276 31746 41304
rect 30317 41273 30329 41276
rect 30271 41267 30329 41273
rect 31740 41264 31746 41276
rect 31798 41264 31804 41316
rect 48671 41307 48729 41313
rect 48671 41273 48683 41307
rect 48717 41304 48729 41307
rect 48852 41304 48858 41316
rect 48717 41276 48858 41304
rect 48717 41273 48729 41276
rect 48671 41267 48729 41273
rect 48852 41264 48858 41276
rect 48910 41264 48916 41316
rect 52719 41307 52777 41313
rect 52719 41273 52731 41307
rect 52765 41304 52777 41307
rect 53728 41304 53734 41316
rect 52765 41276 53734 41304
rect 52765 41273 52777 41276
rect 52719 41267 52777 41273
rect 53728 41264 53734 41276
rect 53786 41264 53792 41316
rect 54482 41276 60122 41304
rect 1935 41171 1993 41177
rect 1935 41137 1947 41171
rect 1981 41168 1993 41171
rect 3514 41168 3542 41264
rect 1981 41140 3542 41168
rect 5247 41171 5305 41177
rect 1981 41137 1993 41140
rect 1935 41131 1993 41137
rect 5247 41137 5259 41171
rect 5293 41168 5305 41171
rect 6535 41171 6593 41177
rect 6535 41168 6547 41171
rect 5293 41140 6547 41168
rect 5293 41137 5305 41140
rect 5247 41131 5305 41137
rect 6535 41137 6547 41140
rect 6581 41137 6593 41171
rect 6535 41131 6593 41137
rect 12055 41171 12113 41177
rect 12055 41137 12067 41171
rect 12101 41168 12113 41171
rect 23371 41171 23429 41177
rect 12101 41140 13110 41168
rect 12101 41137 12113 41140
rect 12055 41131 12113 41137
rect 1659 41103 1717 41109
rect 1659 41069 1671 41103
rect 1705 41100 1717 41103
rect 3496 41100 3502 41112
rect 1705 41072 3502 41100
rect 1705 41069 1717 41072
rect 1659 41063 1717 41069
rect 3496 41060 3502 41072
rect 3554 41100 3560 41112
rect 3591 41103 3649 41109
rect 3591 41100 3603 41103
rect 3554 41072 3603 41100
rect 3554 41060 3560 41072
rect 3591 41069 3603 41072
rect 3637 41069 3649 41103
rect 4600 41100 4606 41112
rect 4561 41072 4606 41100
rect 3591 41063 3649 41069
rect 4600 41060 4606 41072
rect 4658 41060 4664 41112
rect 6164 41060 6170 41112
rect 6222 41100 6228 41112
rect 6259 41103 6317 41109
rect 6259 41100 6271 41103
rect 6222 41072 6271 41100
rect 6222 41060 6228 41072
rect 6259 41069 6271 41072
rect 6305 41069 6317 41103
rect 12328 41100 12334 41112
rect 12289 41072 12334 41100
rect 6259 41063 6317 41069
rect 12328 41060 12334 41072
rect 12386 41060 12392 41112
rect 13082 41044 13110 41140
rect 23371 41137 23383 41171
rect 23417 41168 23429 41171
rect 24935 41171 24993 41177
rect 24935 41168 24947 41171
rect 23417 41140 24947 41168
rect 23417 41137 23429 41140
rect 23371 41131 23429 41137
rect 24935 41137 24947 41140
rect 24981 41168 24993 41171
rect 37076 41168 37082 41180
rect 24981 41140 37082 41168
rect 24981 41137 24993 41140
rect 24935 41131 24993 41137
rect 37076 41128 37082 41140
rect 37134 41128 37140 41180
rect 43059 41171 43117 41177
rect 43059 41168 43071 41171
rect 37738 41140 43071 41168
rect 17483 41103 17541 41109
rect 17483 41100 17495 41103
rect 17406 41072 17495 41100
rect 13064 40992 13070 41044
rect 13122 41032 13128 41044
rect 13122 41004 13938 41032
rect 13122 40992 13128 41004
rect 7820 40964 7826 40976
rect 7781 40936 7826 40964
rect 7820 40924 7826 40936
rect 7878 40924 7884 40976
rect 8004 40964 8010 40976
rect 7965 40936 8010 40964
rect 8004 40924 8010 40936
rect 8062 40924 8068 40976
rect 13432 40964 13438 40976
rect 13393 40936 13438 40964
rect 13432 40924 13438 40936
rect 13490 40924 13496 40976
rect 13910 40973 13938 41004
rect 17406 40976 17434 41072
rect 17483 41069 17495 41072
rect 17529 41069 17541 41103
rect 17756 41100 17762 41112
rect 17717 41072 17762 41100
rect 17483 41063 17541 41069
rect 17756 41060 17762 41072
rect 17814 41060 17820 41112
rect 23095 41103 23153 41109
rect 23095 41100 23107 41103
rect 22926 41072 23107 41100
rect 13895 40967 13953 40973
rect 13895 40933 13907 40967
rect 13941 40964 13953 40967
rect 14904 40964 14910 40976
rect 13941 40936 14910 40964
rect 13941 40933 13953 40936
rect 13895 40927 13953 40933
rect 14904 40924 14910 40936
rect 14962 40924 14968 40976
rect 17299 40967 17357 40973
rect 17299 40933 17311 40967
rect 17345 40964 17357 40967
rect 17388 40964 17394 40976
rect 17345 40936 17394 40964
rect 17345 40933 17357 40936
rect 17299 40927 17357 40933
rect 17388 40924 17394 40936
rect 17446 40924 17452 40976
rect 20884 40924 20890 40976
rect 20942 40964 20948 40976
rect 22926 40973 22954 41072
rect 23095 41069 23107 41072
rect 23141 41069 23153 41103
rect 23095 41063 23153 41069
rect 25579 41103 25637 41109
rect 25579 41069 25591 41103
rect 25625 41100 25637 41103
rect 25668 41100 25674 41112
rect 25625 41072 25674 41100
rect 25625 41069 25637 41072
rect 25579 41063 25637 41069
rect 25668 41060 25674 41072
rect 25726 41060 25732 41112
rect 25855 41103 25913 41109
rect 25855 41069 25867 41103
rect 25901 41100 25913 41103
rect 28428 41100 28434 41112
rect 25901 41072 28434 41100
rect 25901 41069 25913 41072
rect 25855 41063 25913 41069
rect 28428 41060 28434 41072
rect 28486 41060 28492 41112
rect 28707 41103 28765 41109
rect 28707 41100 28719 41103
rect 28538 41072 28719 41100
rect 28538 40976 28566 41072
rect 28707 41069 28719 41072
rect 28753 41069 28765 41103
rect 28707 41063 28765 41069
rect 28796 41060 28802 41112
rect 28854 41100 28860 41112
rect 28983 41103 29041 41109
rect 28983 41100 28995 41103
rect 28854 41072 28995 41100
rect 28854 41060 28860 41072
rect 28983 41069 28995 41072
rect 29029 41069 29041 41103
rect 28983 41063 29041 41069
rect 32019 41103 32077 41109
rect 32019 41069 32031 41103
rect 32065 41069 32077 41103
rect 32019 41063 32077 41069
rect 32034 41032 32062 41063
rect 32752 41060 32758 41112
rect 32810 41100 32816 41112
rect 33123 41103 33181 41109
rect 33123 41100 33135 41103
rect 32810 41072 33135 41100
rect 32810 41060 32816 41072
rect 33123 41069 33135 41072
rect 33169 41069 33181 41103
rect 33123 41063 33181 41069
rect 33215 41103 33273 41109
rect 33215 41069 33227 41103
rect 33261 41100 33273 41103
rect 36340 41100 36346 41112
rect 33261 41072 36346 41100
rect 33261 41069 33273 41072
rect 33215 41063 33273 41069
rect 33230 41032 33258 41063
rect 36340 41060 36346 41072
rect 36398 41060 36404 41112
rect 37738 41109 37766 41140
rect 43059 41137 43071 41140
rect 43105 41168 43117 41171
rect 50784 41168 50790 41180
rect 43105 41140 43286 41168
rect 43105 41137 43117 41140
rect 43059 41131 43117 41137
rect 37355 41103 37413 41109
rect 37355 41069 37367 41103
rect 37401 41100 37413 41103
rect 37723 41103 37781 41109
rect 37723 41100 37735 41103
rect 37401 41072 37735 41100
rect 37401 41069 37413 41072
rect 37355 41063 37413 41069
rect 37723 41069 37735 41072
rect 37769 41069 37781 41103
rect 37723 41063 37781 41069
rect 37999 41103 38057 41109
rect 37999 41069 38011 41103
rect 38045 41100 38057 41103
rect 40848 41100 40854 41112
rect 38045 41072 40854 41100
rect 38045 41069 38057 41072
rect 37999 41063 38057 41069
rect 32034 41004 33258 41032
rect 22911 40967 22969 40973
rect 22911 40964 22923 40967
rect 20942 40936 22923 40964
rect 20942 40924 20948 40936
rect 22911 40933 22923 40936
rect 22957 40933 22969 40967
rect 22911 40927 22969 40933
rect 26772 40924 26778 40976
rect 26830 40964 26836 40976
rect 27327 40967 27385 40973
rect 27327 40964 27339 40967
rect 26830 40936 27339 40964
rect 26830 40924 26836 40936
rect 27327 40933 27339 40936
rect 27373 40964 27385 40967
rect 28520 40964 28526 40976
rect 27373 40936 28526 40964
rect 27373 40933 27385 40936
rect 27327 40927 27385 40933
rect 28520 40924 28526 40936
rect 28578 40964 28584 40976
rect 29348 40964 29354 40976
rect 28578 40936 29354 40964
rect 28578 40924 28584 40936
rect 29348 40924 29354 40936
rect 29406 40964 29412 40976
rect 30452 40964 30458 40976
rect 29406 40936 30458 40964
rect 29406 40924 29412 40936
rect 30452 40924 30458 40936
rect 30510 40924 30516 40976
rect 31556 40924 31562 40976
rect 31614 40964 31620 40976
rect 32203 40967 32261 40973
rect 32203 40964 32215 40967
rect 31614 40936 32215 40964
rect 31614 40924 31620 40936
rect 32203 40933 32215 40936
rect 32249 40933 32261 40967
rect 32203 40927 32261 40933
rect 32752 40924 32758 40976
rect 32810 40964 32816 40976
rect 32939 40967 32997 40973
rect 32939 40964 32951 40967
rect 32810 40936 32951 40964
rect 32810 40924 32816 40936
rect 32939 40933 32951 40936
rect 32985 40933 32997 40967
rect 32939 40927 32997 40933
rect 36527 40967 36585 40973
rect 36527 40933 36539 40967
rect 36573 40964 36585 40967
rect 37370 40964 37398 41063
rect 40848 41060 40854 41072
rect 40906 41060 40912 41112
rect 43258 41109 43286 41140
rect 43810 41140 50790 41168
rect 43810 41109 43838 41140
rect 50784 41128 50790 41140
rect 50842 41128 50848 41180
rect 52532 41128 52538 41180
rect 52590 41168 52596 41180
rect 54482 41177 54510 41276
rect 60094 41177 60122 41276
rect 61088 41264 61094 41316
rect 61146 41304 61152 41316
rect 74983 41307 75041 41313
rect 74983 41304 74995 41307
rect 61146 41276 74995 41304
rect 61146 41264 61152 41276
rect 74983 41273 74995 41276
rect 75029 41273 75041 41307
rect 74983 41267 75041 41273
rect 82619 41307 82677 41313
rect 82619 41273 82631 41307
rect 82665 41304 82677 41307
rect 83076 41304 83082 41316
rect 82665 41276 83082 41304
rect 82665 41273 82677 41276
rect 82619 41267 82677 41273
rect 83076 41264 83082 41276
rect 83134 41264 83140 41316
rect 54467 41171 54525 41177
rect 54467 41168 54479 41171
rect 52590 41140 54479 41168
rect 52590 41128 52596 41140
rect 54467 41137 54479 41140
rect 54513 41137 54525 41171
rect 54467 41131 54525 41137
rect 55755 41171 55813 41177
rect 55755 41137 55767 41171
rect 55801 41168 55813 41171
rect 57043 41171 57101 41177
rect 57043 41168 57055 41171
rect 55801 41140 57055 41168
rect 55801 41137 55813 41140
rect 55755 41131 55813 41137
rect 57043 41137 57055 41140
rect 57089 41137 57101 41171
rect 57043 41131 57101 41137
rect 60079 41171 60137 41177
rect 60079 41137 60091 41171
rect 60125 41137 60137 41171
rect 60079 41131 60137 41137
rect 61367 41171 61425 41177
rect 61367 41137 61379 41171
rect 61413 41168 61425 41171
rect 62655 41171 62713 41177
rect 62655 41168 62667 41171
rect 61413 41140 62667 41168
rect 61413 41137 61425 41140
rect 61367 41131 61425 41137
rect 62655 41137 62667 41140
rect 62701 41137 62713 41171
rect 62655 41131 62713 41137
rect 80963 41171 81021 41177
rect 80963 41137 80975 41171
rect 81009 41168 81021 41171
rect 81009 41140 81374 41168
rect 81009 41137 81021 41140
rect 80963 41131 81021 41137
rect 43243 41103 43301 41109
rect 43243 41069 43255 41103
rect 43289 41069 43301 41103
rect 43243 41063 43301 41069
rect 43795 41103 43853 41109
rect 43795 41069 43807 41103
rect 43841 41069 43853 41103
rect 47104 41100 47110 41112
rect 47065 41072 47110 41100
rect 43795 41063 43853 41069
rect 37536 40964 37542 40976
rect 36573 40936 37398 40964
rect 37497 40936 37542 40964
rect 36573 40933 36585 40936
rect 36527 40927 36585 40933
rect 37536 40924 37542 40936
rect 37594 40924 37600 40976
rect 43258 40964 43286 41063
rect 47104 41060 47110 41072
rect 47162 41060 47168 41112
rect 47380 41100 47386 41112
rect 47341 41072 47386 41100
rect 47380 41060 47386 41072
rect 47438 41060 47444 41112
rect 51060 41060 51066 41112
rect 51118 41100 51124 41112
rect 51155 41103 51213 41109
rect 51155 41100 51167 41103
rect 51118 41072 51167 41100
rect 51118 41060 51124 41072
rect 51155 41069 51167 41072
rect 51201 41069 51213 41103
rect 51428 41100 51434 41112
rect 51389 41072 51434 41100
rect 51155 41063 51213 41069
rect 43979 41035 44037 41041
rect 43979 41001 43991 41035
rect 44025 41032 44037 41035
rect 44068 41032 44074 41044
rect 44025 41004 44074 41032
rect 44025 41001 44037 41004
rect 43979 40995 44037 41001
rect 44068 40992 44074 41004
rect 44126 40992 44132 41044
rect 46736 40964 46742 40976
rect 43258 40936 46742 40964
rect 46736 40924 46742 40936
rect 46794 40924 46800 40976
rect 47104 40924 47110 40976
rect 47162 40964 47168 40976
rect 48855 40967 48913 40973
rect 48855 40964 48867 40967
rect 47162 40936 48867 40964
rect 47162 40924 47168 40936
rect 48855 40933 48867 40936
rect 48901 40964 48913 40967
rect 49496 40964 49502 40976
rect 48901 40936 49502 40964
rect 48901 40933 48913 40936
rect 48855 40927 48913 40933
rect 49496 40924 49502 40936
rect 49554 40924 49560 40976
rect 51170 40964 51198 41063
rect 51428 41060 51434 41072
rect 51486 41060 51492 41112
rect 54648 41100 54654 41112
rect 54609 41072 54654 41100
rect 54648 41060 54654 41072
rect 54706 41060 54712 41112
rect 55203 41103 55261 41109
rect 55203 41069 55215 41103
rect 55249 41069 55261 41103
rect 55203 41063 55261 41069
rect 55387 41103 55445 41109
rect 55387 41069 55399 41103
rect 55433 41069 55445 41103
rect 55387 41063 55445 41069
rect 54666 41032 54694 41060
rect 55218 41032 55246 41063
rect 54666 41004 55246 41032
rect 55402 41032 55430 41063
rect 56028 41060 56034 41112
rect 56086 41100 56092 41112
rect 56764 41100 56770 41112
rect 56086 41072 56770 41100
rect 56086 41060 56092 41072
rect 56764 41060 56770 41072
rect 56822 41060 56828 41112
rect 60260 41100 60266 41112
rect 60221 41072 60266 41100
rect 60260 41060 60266 41072
rect 60318 41060 60324 41112
rect 60815 41103 60873 41109
rect 60815 41069 60827 41103
rect 60861 41069 60873 41103
rect 60815 41063 60873 41069
rect 60999 41103 61057 41109
rect 60999 41069 61011 41103
rect 61045 41100 61057 41103
rect 61045 41072 61686 41100
rect 61045 41069 61057 41072
rect 60999 41063 61057 41069
rect 60278 41032 60306 41060
rect 60830 41032 60858 41063
rect 55402 41004 56074 41032
rect 60278 41004 60858 41032
rect 52903 40967 52961 40973
rect 52903 40964 52915 40967
rect 51170 40936 52915 40964
rect 52903 40933 52915 40936
rect 52949 40964 52961 40967
rect 55568 40964 55574 40976
rect 52949 40936 55574 40964
rect 52949 40933 52961 40936
rect 52903 40927 52961 40933
rect 55568 40924 55574 40936
rect 55626 40964 55632 40976
rect 55844 40964 55850 40976
rect 55626 40936 55850 40964
rect 55626 40924 55632 40936
rect 55844 40924 55850 40936
rect 55902 40924 55908 40976
rect 56046 40973 56074 41004
rect 56031 40967 56089 40973
rect 56031 40933 56043 40967
rect 56077 40964 56089 40967
rect 56672 40964 56678 40976
rect 56077 40936 56678 40964
rect 56077 40933 56089 40936
rect 56031 40927 56089 40933
rect 56672 40924 56678 40936
rect 56730 40924 56736 40976
rect 58052 40924 58058 40976
rect 58110 40964 58116 40976
rect 58147 40967 58205 40973
rect 58147 40964 58159 40967
rect 58110 40936 58159 40964
rect 58110 40924 58116 40936
rect 58147 40933 58159 40936
rect 58193 40933 58205 40967
rect 58147 40927 58205 40933
rect 58607 40967 58665 40973
rect 58607 40933 58619 40967
rect 58653 40964 58665 40967
rect 58696 40964 58702 40976
rect 58653 40936 58702 40964
rect 58653 40933 58665 40936
rect 58607 40927 58665 40933
rect 58696 40924 58702 40936
rect 58754 40924 58760 40976
rect 61658 40973 61686 41072
rect 61732 41060 61738 41112
rect 61790 41100 61796 41112
rect 62195 41103 62253 41109
rect 62195 41100 62207 41103
rect 61790 41072 62207 41100
rect 61790 41060 61796 41072
rect 62195 41069 62207 41072
rect 62241 41100 62253 41103
rect 62379 41103 62437 41109
rect 62379 41100 62391 41103
rect 62241 41072 62391 41100
rect 62241 41069 62253 41072
rect 62195 41063 62253 41069
rect 62379 41069 62391 41072
rect 62425 41100 62437 41103
rect 65320 41100 65326 41112
rect 62425 41072 65326 41100
rect 62425 41069 62437 41072
rect 62379 41063 62437 41069
rect 65320 41060 65326 41072
rect 65378 41060 65384 41112
rect 73603 41103 73661 41109
rect 73603 41069 73615 41103
rect 73649 41100 73661 41103
rect 73692 41100 73698 41112
rect 73649 41072 73698 41100
rect 73649 41069 73661 41072
rect 73603 41063 73661 41069
rect 73692 41060 73698 41072
rect 73750 41060 73756 41112
rect 73876 41100 73882 41112
rect 73837 41072 73882 41100
rect 73876 41060 73882 41072
rect 73934 41060 73940 41112
rect 79488 41060 79494 41112
rect 79546 41100 79552 41112
rect 80779 41103 80837 41109
rect 80779 41100 80791 41103
rect 79546 41072 80791 41100
rect 79546 41060 79552 41072
rect 80779 41069 80791 41072
rect 80825 41100 80837 41103
rect 81055 41103 81113 41109
rect 81055 41100 81067 41103
rect 80825 41072 81067 41100
rect 80825 41069 80837 41072
rect 80779 41063 80837 41069
rect 81055 41069 81067 41072
rect 81101 41100 81113 41103
rect 81144 41100 81150 41112
rect 81101 41072 81150 41100
rect 81101 41069 81113 41072
rect 81055 41063 81113 41069
rect 81144 41060 81150 41072
rect 81202 41060 81208 41112
rect 81346 41109 81374 41140
rect 83628 41128 83634 41180
rect 83686 41168 83692 41180
rect 86759 41171 86817 41177
rect 86759 41168 86771 41171
rect 83686 41140 86771 41168
rect 83686 41128 83692 41140
rect 86759 41137 86771 41140
rect 86805 41137 86817 41171
rect 86759 41131 86817 41137
rect 81331 41103 81389 41109
rect 81331 41069 81343 41103
rect 81377 41100 81389 41103
rect 81420 41100 81426 41112
rect 81377 41072 81426 41100
rect 81377 41069 81389 41072
rect 81331 41063 81389 41069
rect 81420 41060 81426 41072
rect 81478 41060 81484 41112
rect 85379 41103 85437 41109
rect 85379 41069 85391 41103
rect 85425 41069 85437 41103
rect 85652 41100 85658 41112
rect 85613 41072 85658 41100
rect 85379 41063 85437 41069
rect 61643 40967 61701 40973
rect 61643 40933 61655 40967
rect 61689 40964 61701 40967
rect 61732 40964 61738 40976
rect 61689 40936 61738 40964
rect 61689 40933 61701 40936
rect 61643 40927 61701 40933
rect 61732 40924 61738 40936
rect 61790 40924 61796 40976
rect 63572 40924 63578 40976
rect 63630 40964 63636 40976
rect 63759 40967 63817 40973
rect 63759 40964 63771 40967
rect 63630 40936 63771 40964
rect 63630 40924 63636 40936
rect 63759 40933 63771 40936
rect 63805 40933 63817 40967
rect 63759 40927 63817 40933
rect 75443 40967 75501 40973
rect 75443 40933 75455 40967
rect 75489 40964 75501 40967
rect 75992 40964 75998 40976
rect 75489 40936 75998 40964
rect 75489 40933 75501 40936
rect 75443 40927 75501 40933
rect 75992 40924 75998 40936
rect 76050 40924 76056 40976
rect 85008 40924 85014 40976
rect 85066 40964 85072 40976
rect 85287 40967 85345 40973
rect 85287 40964 85299 40967
rect 85066 40936 85299 40964
rect 85066 40924 85072 40936
rect 85287 40933 85299 40936
rect 85333 40964 85345 40967
rect 85394 40964 85422 41063
rect 85652 41060 85658 41072
rect 85710 41060 85716 41112
rect 88136 40964 88142 40976
rect 85333 40936 88142 40964
rect 85333 40933 85345 40936
rect 85287 40927 85345 40933
rect 88136 40924 88142 40936
rect 88194 40924 88200 40976
rect 538 40874 93642 40896
rect 538 40822 6344 40874
rect 6396 40822 6408 40874
rect 6460 40822 6472 40874
rect 6524 40822 6536 40874
rect 6588 40822 11672 40874
rect 11724 40822 11736 40874
rect 11788 40822 11800 40874
rect 11852 40822 11864 40874
rect 11916 40822 17000 40874
rect 17052 40822 17064 40874
rect 17116 40822 17128 40874
rect 17180 40822 17192 40874
rect 17244 40822 22328 40874
rect 22380 40822 22392 40874
rect 22444 40822 22456 40874
rect 22508 40822 22520 40874
rect 22572 40822 27656 40874
rect 27708 40822 27720 40874
rect 27772 40822 27784 40874
rect 27836 40822 27848 40874
rect 27900 40822 32984 40874
rect 33036 40822 33048 40874
rect 33100 40822 33112 40874
rect 33164 40822 33176 40874
rect 33228 40822 38312 40874
rect 38364 40822 38376 40874
rect 38428 40822 38440 40874
rect 38492 40822 38504 40874
rect 38556 40822 43640 40874
rect 43692 40822 43704 40874
rect 43756 40822 43768 40874
rect 43820 40822 43832 40874
rect 43884 40822 48968 40874
rect 49020 40822 49032 40874
rect 49084 40822 49096 40874
rect 49148 40822 49160 40874
rect 49212 40822 54296 40874
rect 54348 40822 54360 40874
rect 54412 40822 54424 40874
rect 54476 40822 54488 40874
rect 54540 40822 59624 40874
rect 59676 40822 59688 40874
rect 59740 40822 59752 40874
rect 59804 40822 59816 40874
rect 59868 40822 64952 40874
rect 65004 40822 65016 40874
rect 65068 40822 65080 40874
rect 65132 40822 65144 40874
rect 65196 40822 70280 40874
rect 70332 40822 70344 40874
rect 70396 40822 70408 40874
rect 70460 40822 70472 40874
rect 70524 40822 75608 40874
rect 75660 40822 75672 40874
rect 75724 40822 75736 40874
rect 75788 40822 75800 40874
rect 75852 40822 80936 40874
rect 80988 40822 81000 40874
rect 81052 40822 81064 40874
rect 81116 40822 81128 40874
rect 81180 40822 86264 40874
rect 86316 40822 86328 40874
rect 86380 40822 86392 40874
rect 86444 40822 86456 40874
rect 86508 40822 91592 40874
rect 91644 40822 91656 40874
rect 91708 40822 91720 40874
rect 91772 40822 91784 40874
rect 91836 40822 93642 40874
rect 538 40800 93642 40822
rect 3496 40720 3502 40772
rect 3554 40760 3560 40772
rect 5431 40763 5489 40769
rect 5431 40760 5443 40763
rect 3554 40732 5443 40760
rect 3554 40720 3560 40732
rect 5431 40729 5443 40732
rect 5477 40760 5489 40763
rect 6164 40760 6170 40772
rect 5477 40732 6170 40760
rect 5477 40729 5489 40732
rect 5431 40723 5489 40729
rect 6164 40720 6170 40732
rect 6222 40720 6228 40772
rect 14904 40720 14910 40772
rect 14962 40760 14968 40772
rect 28339 40763 28397 40769
rect 14962 40732 16790 40760
rect 14962 40720 14968 40732
rect 16762 40701 16790 40732
rect 28339 40729 28351 40763
rect 28385 40760 28397 40763
rect 29256 40760 29262 40772
rect 28385 40732 29262 40760
rect 28385 40729 28397 40732
rect 28339 40723 28397 40729
rect 29256 40720 29262 40732
rect 29314 40720 29320 40772
rect 47104 40760 47110 40772
rect 45466 40732 47110 40760
rect 16747 40695 16805 40701
rect 16747 40661 16759 40695
rect 16793 40692 16805 40695
rect 17388 40692 17394 40704
rect 16793 40664 17394 40692
rect 16793 40661 16805 40664
rect 16747 40655 16805 40661
rect 17388 40652 17394 40664
rect 17446 40652 17452 40704
rect 28520 40692 28526 40704
rect 28481 40664 28526 40692
rect 28520 40652 28526 40664
rect 28578 40652 28584 40704
rect 0 40584 6 40636
rect 58 40624 64 40636
rect 2395 40627 2453 40633
rect 2395 40624 2407 40627
rect 58 40596 2407 40624
rect 58 40584 64 40596
rect 2395 40593 2407 40596
rect 2441 40593 2453 40627
rect 3496 40624 3502 40636
rect 3457 40596 3502 40624
rect 2395 40587 2453 40593
rect 3496 40584 3502 40596
rect 3554 40584 3560 40636
rect 4048 40584 4054 40636
rect 4106 40624 4112 40636
rect 5060 40624 5066 40636
rect 4106 40596 5066 40624
rect 4106 40584 4112 40596
rect 5060 40584 5066 40596
rect 5118 40584 5124 40636
rect 6719 40627 6777 40633
rect 6719 40624 6731 40627
rect 5170 40596 6731 40624
rect 3775 40559 3833 40565
rect 3775 40525 3787 40559
rect 3821 40556 3833 40559
rect 3821 40528 4554 40556
rect 3821 40525 3833 40528
rect 3775 40519 3833 40525
rect 2484 40420 2490 40432
rect 2445 40392 2490 40420
rect 2484 40380 2490 40392
rect 2542 40380 2548 40432
rect 4526 40420 4554 40528
rect 4876 40516 4882 40568
rect 4934 40556 4940 40568
rect 4971 40559 5029 40565
rect 4971 40556 4983 40559
rect 4934 40528 4983 40556
rect 4934 40516 4940 40528
rect 4971 40525 4983 40528
rect 5017 40525 5029 40559
rect 4971 40519 5029 40525
rect 4600 40448 4606 40500
rect 4658 40488 4664 40500
rect 5170 40488 5198 40596
rect 6719 40593 6731 40596
rect 6765 40593 6777 40627
rect 8004 40624 8010 40636
rect 6719 40587 6777 40593
rect 7286 40596 8010 40624
rect 6164 40516 6170 40568
rect 6222 40556 6228 40568
rect 6443 40559 6501 40565
rect 6443 40556 6455 40559
rect 6222 40528 6455 40556
rect 6222 40516 6228 40528
rect 6443 40525 6455 40528
rect 6489 40556 6501 40559
rect 7286 40556 7314 40596
rect 8004 40584 8010 40596
rect 8062 40624 8068 40636
rect 8191 40627 8249 40633
rect 8191 40624 8203 40627
rect 8062 40596 8203 40624
rect 8062 40584 8068 40596
rect 8191 40593 8203 40596
rect 8237 40593 8249 40627
rect 8191 40587 8249 40593
rect 9752 40584 9758 40636
rect 9810 40624 9816 40636
rect 13432 40624 13438 40636
rect 9810 40596 13438 40624
rect 9810 40584 9816 40596
rect 13432 40584 13438 40596
rect 13490 40584 13496 40636
rect 14628 40584 14634 40636
rect 14686 40624 14692 40636
rect 14686 40596 18814 40624
rect 14686 40584 14692 40596
rect 6489 40528 7314 40556
rect 6489 40525 6501 40528
rect 6443 40519 6501 40525
rect 7360 40516 7366 40568
rect 7418 40516 7424 40568
rect 11040 40556 11046 40568
rect 11001 40528 11046 40556
rect 11040 40516 11046 40528
rect 11098 40516 11104 40568
rect 11319 40559 11377 40565
rect 11319 40525 11331 40559
rect 11365 40556 11377 40559
rect 14168 40556 14174 40568
rect 11365 40528 14174 40556
rect 11365 40525 11377 40528
rect 11319 40519 11377 40525
rect 14168 40516 14174 40528
rect 14226 40516 14232 40568
rect 14904 40556 14910 40568
rect 14865 40528 14910 40556
rect 14904 40516 14910 40528
rect 14962 40516 14968 40568
rect 15183 40559 15241 40565
rect 15183 40525 15195 40559
rect 15229 40556 15241 40559
rect 17299 40559 17357 40565
rect 15229 40528 17250 40556
rect 15229 40525 15241 40528
rect 15183 40519 15241 40525
rect 4658 40460 5198 40488
rect 7378 40488 7406 40516
rect 7378 40460 9614 40488
rect 4658 40448 4664 40460
rect 5336 40420 5342 40432
rect 4526 40392 5342 40420
rect 5336 40380 5342 40392
rect 5394 40380 5400 40432
rect 8004 40420 8010 40432
rect 7965 40392 8010 40420
rect 8004 40380 8010 40392
rect 8062 40380 8068 40432
rect 9586 40420 9614 40460
rect 12144 40448 12150 40500
rect 12202 40488 12208 40500
rect 12202 40460 14766 40488
rect 12202 40448 12208 40460
rect 12423 40423 12481 40429
rect 12423 40420 12435 40423
rect 9586 40392 12435 40420
rect 12423 40389 12435 40392
rect 12469 40389 12481 40423
rect 12423 40383 12481 40389
rect 12883 40423 12941 40429
rect 12883 40389 12895 40423
rect 12929 40420 12941 40423
rect 13064 40420 13070 40432
rect 12929 40392 13070 40420
rect 12929 40389 12941 40392
rect 12883 40383 12941 40389
rect 13064 40380 13070 40392
rect 13122 40380 13128 40432
rect 14738 40420 14766 40460
rect 16287 40423 16345 40429
rect 16287 40420 16299 40423
rect 14738 40392 16299 40420
rect 16287 40389 16299 40392
rect 16333 40389 16345 40423
rect 17222 40420 17250 40528
rect 17299 40525 17311 40559
rect 17345 40556 17357 40559
rect 17388 40556 17394 40568
rect 17345 40528 17394 40556
rect 17345 40525 17357 40528
rect 17299 40519 17357 40525
rect 17388 40516 17394 40528
rect 17446 40516 17452 40568
rect 17664 40556 17670 40568
rect 17625 40528 17670 40556
rect 17664 40516 17670 40528
rect 17722 40516 17728 40568
rect 18786 40565 18814 40596
rect 25668 40584 25674 40636
rect 25726 40624 25732 40636
rect 26772 40624 26778 40636
rect 25726 40596 26778 40624
rect 25726 40584 25732 40596
rect 26772 40584 26778 40596
rect 26830 40584 26836 40636
rect 30452 40584 30458 40636
rect 30510 40624 30516 40636
rect 31835 40627 31893 40633
rect 31835 40624 31847 40627
rect 30510 40596 31847 40624
rect 30510 40584 30516 40596
rect 31835 40593 31847 40596
rect 31881 40624 31893 40627
rect 33491 40627 33549 40633
rect 31881 40596 32798 40624
rect 31881 40593 31893 40596
rect 31835 40587 31893 40593
rect 18771 40559 18829 40565
rect 18771 40525 18783 40559
rect 18817 40525 18829 40559
rect 20979 40559 21037 40565
rect 20979 40556 20991 40559
rect 18771 40519 18829 40525
rect 20902 40528 20991 40556
rect 20902 40432 20930 40528
rect 20979 40525 20991 40528
rect 21025 40525 21037 40559
rect 21252 40556 21258 40568
rect 21213 40528 21258 40556
rect 20979 40519 21037 40525
rect 21252 40516 21258 40528
rect 21310 40516 21316 40568
rect 21988 40516 21994 40568
rect 22046 40556 22052 40568
rect 22359 40559 22417 40565
rect 22359 40556 22371 40559
rect 22046 40528 22371 40556
rect 22046 40516 22052 40528
rect 22359 40525 22371 40528
rect 22405 40525 22417 40559
rect 27048 40556 27054 40568
rect 27009 40528 27054 40556
rect 22359 40519 22417 40525
rect 27048 40516 27054 40528
rect 27106 40516 27112 40568
rect 32111 40559 32169 40565
rect 32111 40525 32123 40559
rect 32157 40556 32169 40559
rect 32292 40556 32298 40568
rect 32157 40528 32298 40556
rect 32157 40525 32169 40528
rect 32111 40519 32169 40525
rect 32292 40516 32298 40528
rect 32350 40516 32356 40568
rect 32770 40556 32798 40596
rect 33491 40593 33503 40627
rect 33537 40624 33549 40627
rect 34132 40624 34138 40636
rect 33537 40596 34138 40624
rect 33537 40593 33549 40596
rect 33491 40587 33549 40593
rect 34132 40584 34138 40596
rect 34190 40584 34196 40636
rect 35975 40627 36033 40633
rect 35975 40593 35987 40627
rect 36021 40624 36033 40627
rect 36616 40624 36622 40636
rect 36021 40596 36622 40624
rect 36021 40593 36033 40596
rect 35975 40587 36033 40593
rect 36616 40584 36622 40596
rect 36674 40584 36680 40636
rect 37447 40627 37505 40633
rect 37447 40593 37459 40627
rect 37493 40624 37505 40627
rect 37536 40624 37542 40636
rect 37493 40596 37542 40624
rect 37493 40593 37505 40596
rect 37447 40587 37505 40593
rect 37536 40584 37542 40596
rect 37594 40584 37600 40636
rect 38827 40627 38885 40633
rect 38827 40593 38839 40627
rect 38873 40624 38885 40627
rect 39100 40624 39106 40636
rect 38873 40596 39106 40624
rect 38873 40593 38885 40596
rect 38827 40587 38885 40593
rect 39100 40584 39106 40596
rect 39158 40584 39164 40636
rect 41311 40627 41369 40633
rect 41311 40593 41323 40627
rect 41357 40624 41369 40627
rect 41492 40624 41498 40636
rect 41357 40596 41498 40624
rect 41357 40593 41369 40596
rect 41311 40587 41369 40593
rect 41492 40584 41498 40596
rect 41550 40584 41556 40636
rect 43059 40627 43117 40633
rect 43059 40593 43071 40627
rect 43105 40624 43117 40627
rect 44068 40624 44074 40636
rect 43105 40596 44074 40624
rect 43105 40593 43117 40596
rect 43059 40587 43117 40593
rect 44068 40584 44074 40596
rect 44126 40584 44132 40636
rect 45466 40633 45494 40732
rect 47104 40720 47110 40732
rect 47162 40760 47168 40772
rect 47199 40763 47257 40769
rect 47199 40760 47211 40763
rect 47162 40732 47211 40760
rect 47162 40720 47168 40732
rect 47199 40729 47211 40732
rect 47245 40729 47257 40763
rect 71116 40760 71122 40772
rect 47199 40723 47257 40729
rect 70950 40732 71122 40760
rect 51060 40692 51066 40704
rect 50973 40664 51066 40692
rect 51060 40652 51066 40664
rect 51118 40692 51124 40704
rect 51339 40695 51397 40701
rect 51339 40692 51351 40695
rect 51118 40664 51351 40692
rect 51118 40652 51124 40664
rect 51339 40661 51351 40664
rect 51385 40661 51397 40695
rect 51339 40655 51397 40661
rect 56764 40652 56770 40704
rect 56822 40692 56828 40704
rect 57411 40695 57469 40701
rect 57411 40692 57423 40695
rect 56822 40664 57423 40692
rect 56822 40652 56828 40664
rect 57411 40661 57423 40664
rect 57457 40692 57469 40695
rect 57457 40664 58742 40692
rect 57457 40661 57469 40664
rect 57411 40655 57469 40661
rect 45451 40627 45509 40633
rect 45451 40593 45463 40627
rect 45497 40593 45509 40627
rect 49496 40624 49502 40636
rect 49457 40596 49502 40624
rect 45451 40587 45509 40593
rect 49496 40584 49502 40596
rect 49554 40624 49560 40636
rect 51078 40624 51106 40652
rect 58714 40636 58742 40664
rect 49554 40596 51106 40624
rect 51155 40627 51213 40633
rect 49554 40584 49560 40596
rect 51155 40593 51167 40627
rect 51201 40624 51213 40627
rect 51244 40624 51250 40636
rect 51201 40596 51250 40624
rect 51201 40593 51213 40596
rect 51155 40587 51213 40593
rect 51244 40584 51250 40596
rect 51302 40584 51308 40636
rect 55568 40624 55574 40636
rect 55529 40596 55574 40624
rect 55568 40584 55574 40596
rect 55626 40584 55632 40636
rect 56120 40584 56126 40636
rect 56178 40624 56184 40636
rect 57316 40624 57322 40636
rect 56178 40596 57322 40624
rect 56178 40584 56184 40596
rect 57316 40584 57322 40596
rect 57374 40584 57380 40636
rect 58052 40624 58058 40636
rect 58013 40596 58058 40624
rect 58052 40584 58058 40596
rect 58110 40584 58116 40636
rect 58696 40584 58702 40636
rect 58754 40624 58760 40636
rect 60999 40627 61057 40633
rect 60999 40624 61011 40627
rect 58754 40596 61011 40624
rect 58754 40584 58760 40596
rect 60999 40593 61011 40596
rect 61045 40624 61057 40627
rect 61091 40627 61149 40633
rect 61091 40624 61103 40627
rect 61045 40596 61103 40624
rect 61045 40593 61057 40596
rect 60999 40587 61057 40593
rect 61091 40593 61103 40596
rect 61137 40624 61149 40627
rect 61640 40624 61646 40636
rect 61137 40596 61646 40624
rect 61137 40593 61149 40596
rect 61091 40587 61149 40593
rect 61640 40584 61646 40596
rect 61698 40584 61704 40636
rect 62652 40584 62658 40636
rect 62710 40624 62716 40636
rect 62928 40624 62934 40636
rect 62710 40596 62934 40624
rect 62710 40584 62716 40596
rect 62928 40584 62934 40596
rect 62986 40584 62992 40636
rect 63572 40624 63578 40636
rect 63533 40596 63578 40624
rect 63572 40584 63578 40596
rect 63630 40584 63636 40636
rect 66519 40627 66577 40633
rect 66519 40593 66531 40627
rect 66565 40624 66577 40627
rect 68267 40627 68325 40633
rect 68267 40624 68279 40627
rect 66565 40596 68279 40624
rect 66565 40593 66577 40596
rect 66519 40587 66577 40593
rect 68267 40593 68279 40596
rect 68313 40593 68325 40627
rect 68267 40587 68325 40593
rect 33583 40559 33641 40565
rect 33583 40556 33595 40559
rect 32770 40528 33595 40556
rect 33583 40525 33595 40528
rect 33629 40556 33641 40559
rect 34227 40559 34285 40565
rect 34227 40556 34239 40559
rect 33629 40528 34239 40556
rect 33629 40525 33641 40528
rect 33583 40519 33641 40525
rect 34227 40525 34239 40528
rect 34273 40556 34285 40559
rect 34319 40559 34377 40565
rect 34319 40556 34331 40559
rect 34273 40528 34331 40556
rect 34273 40525 34285 40528
rect 34227 40519 34285 40525
rect 34319 40525 34331 40528
rect 34365 40525 34377 40559
rect 34592 40556 34598 40568
rect 34553 40528 34598 40556
rect 34319 40519 34377 40525
rect 17848 40420 17854 40432
rect 17222 40392 17854 40420
rect 16287 40383 16345 40389
rect 17848 40380 17854 40392
rect 17906 40380 17912 40432
rect 20884 40420 20890 40432
rect 20845 40392 20890 40420
rect 20884 40380 20890 40392
rect 20942 40380 20948 40432
rect 34334 40420 34362 40519
rect 34592 40516 34598 40528
rect 34650 40516 34656 40568
rect 37171 40559 37229 40565
rect 37171 40556 37183 40559
rect 36910 40528 37183 40556
rect 34684 40420 34690 40432
rect 34334 40392 34690 40420
rect 34684 40380 34690 40392
rect 34742 40420 34748 40432
rect 36910 40429 36938 40528
rect 37171 40525 37183 40528
rect 37217 40556 37229 40559
rect 39471 40559 39529 40565
rect 39471 40556 39483 40559
rect 37217 40528 39483 40556
rect 37217 40525 37229 40528
rect 37171 40519 37229 40525
rect 39471 40525 39483 40528
rect 39517 40556 39529 40559
rect 39652 40556 39658 40568
rect 39517 40528 39658 40556
rect 39517 40525 39529 40528
rect 39471 40519 39529 40525
rect 39652 40516 39658 40528
rect 39710 40516 39716 40568
rect 39928 40556 39934 40568
rect 39889 40528 39934 40556
rect 39928 40516 39934 40528
rect 39986 40516 39992 40568
rect 41584 40516 41590 40568
rect 41642 40556 41648 40568
rect 42599 40559 42657 40565
rect 42599 40556 42611 40559
rect 41642 40528 42611 40556
rect 41642 40516 41648 40528
rect 42599 40525 42611 40528
rect 42645 40556 42657 40559
rect 42783 40559 42841 40565
rect 42783 40556 42795 40559
rect 42645 40528 42795 40556
rect 42645 40525 42657 40528
rect 42599 40519 42657 40525
rect 42783 40525 42795 40528
rect 42829 40525 42841 40559
rect 42783 40519 42841 40525
rect 43976 40516 43982 40568
rect 44034 40556 44040 40568
rect 44163 40559 44221 40565
rect 44163 40556 44175 40559
rect 44034 40528 44175 40556
rect 44034 40516 44040 40528
rect 44163 40525 44175 40528
rect 44209 40525 44221 40559
rect 45724 40556 45730 40568
rect 45685 40528 45730 40556
rect 44163 40519 44221 40525
rect 45724 40516 45730 40528
rect 45782 40516 45788 40568
rect 46644 40516 46650 40568
rect 46702 40556 46708 40568
rect 46831 40559 46889 40565
rect 46831 40556 46843 40559
rect 46702 40528 46843 40556
rect 46702 40516 46708 40528
rect 46831 40525 46843 40528
rect 46877 40525 46889 40559
rect 49772 40556 49778 40568
rect 49733 40528 49778 40556
rect 46831 40519 46889 40525
rect 49772 40516 49778 40528
rect 49830 40516 49836 40568
rect 55844 40556 55850 40568
rect 55805 40528 55850 40556
rect 55844 40516 55850 40528
rect 55902 40516 55908 40568
rect 56672 40516 56678 40568
rect 56730 40556 56736 40568
rect 58147 40559 58205 40565
rect 58147 40556 58159 40559
rect 56730 40528 58159 40556
rect 56730 40516 56736 40528
rect 58147 40525 58159 40528
rect 58193 40525 58205 40559
rect 61364 40556 61370 40568
rect 61325 40528 61370 40556
rect 58147 40519 58205 40525
rect 61364 40516 61370 40528
rect 61422 40516 61428 40568
rect 61732 40516 61738 40568
rect 61790 40556 61796 40568
rect 62744 40556 62750 40568
rect 61790 40528 62750 40556
rect 61790 40516 61796 40528
rect 62744 40516 62750 40528
rect 62802 40556 62808 40568
rect 63667 40559 63725 40565
rect 63667 40556 63679 40559
rect 62802 40528 63679 40556
rect 62802 40516 62808 40528
rect 63667 40525 63679 40528
rect 63713 40525 63725 40559
rect 63667 40519 63725 40525
rect 66795 40559 66853 40565
rect 66795 40525 66807 40559
rect 66841 40556 66853 40559
rect 68172 40556 68178 40568
rect 66841 40528 68178 40556
rect 66841 40525 66853 40528
rect 66795 40519 66853 40525
rect 68172 40516 68178 40528
rect 68230 40516 68236 40568
rect 68282 40556 68310 40587
rect 68356 40584 68362 40636
rect 68414 40624 68420 40636
rect 70748 40624 70754 40636
rect 68414 40596 70754 40624
rect 68414 40584 68420 40596
rect 70748 40584 70754 40596
rect 70806 40584 70812 40636
rect 70950 40624 70978 40732
rect 71116 40720 71122 40732
rect 71174 40720 71180 40772
rect 81055 40763 81113 40769
rect 79230 40732 79626 40760
rect 71119 40627 71177 40633
rect 71119 40624 71131 40627
rect 70950 40596 71131 40624
rect 71119 40593 71131 40596
rect 71165 40593 71177 40627
rect 71119 40587 71177 40593
rect 71208 40584 71214 40636
rect 71266 40624 71272 40636
rect 71266 40596 75302 40624
rect 71266 40584 71272 40596
rect 69920 40556 69926 40568
rect 68282 40528 69926 40556
rect 69920 40516 69926 40528
rect 69978 40556 69984 40568
rect 70843 40559 70901 40565
rect 70843 40556 70855 40559
rect 69978 40528 70855 40556
rect 69978 40516 69984 40528
rect 70843 40525 70855 40528
rect 70889 40556 70901 40559
rect 73327 40559 73385 40565
rect 70889 40528 72726 40556
rect 70889 40525 70901 40528
rect 70843 40519 70901 40525
rect 41400 40448 41406 40500
rect 41458 40488 41464 40500
rect 42688 40488 42694 40500
rect 41458 40460 42694 40488
rect 41458 40448 41464 40460
rect 42688 40448 42694 40460
rect 42746 40448 42752 40500
rect 59524 40488 59530 40500
rect 56506 40460 59530 40488
rect 36895 40423 36953 40429
rect 36895 40420 36907 40423
rect 34742 40392 36907 40420
rect 34742 40380 34748 40392
rect 36895 40389 36907 40392
rect 36941 40389 36953 40423
rect 36895 40383 36953 40389
rect 51336 40380 51342 40432
rect 51394 40420 51400 40432
rect 56506 40420 56534 40460
rect 59524 40448 59530 40460
rect 59582 40448 59588 40500
rect 51394 40392 56534 40420
rect 51394 40380 51400 40392
rect 56856 40380 56862 40432
rect 56914 40420 56920 40432
rect 56951 40423 57009 40429
rect 56951 40420 56963 40423
rect 56914 40392 56963 40420
rect 56914 40380 56920 40392
rect 56951 40389 56963 40392
rect 56997 40389 57009 40423
rect 62652 40420 62658 40432
rect 62613 40392 62658 40420
rect 56951 40383 57009 40389
rect 62652 40380 62658 40392
rect 62710 40380 62716 40432
rect 64032 40380 64038 40432
rect 64090 40420 64096 40432
rect 67899 40423 67957 40429
rect 67899 40420 67911 40423
rect 64090 40392 67911 40420
rect 64090 40380 64096 40392
rect 67899 40389 67911 40392
rect 67945 40389 67957 40423
rect 72220 40420 72226 40432
rect 72181 40392 72226 40420
rect 67899 40383 67957 40389
rect 72220 40380 72226 40392
rect 72278 40380 72284 40432
rect 72698 40429 72726 40528
rect 73327 40525 73339 40559
rect 73373 40525 73385 40559
rect 73600 40556 73606 40568
rect 73561 40528 73606 40556
rect 73327 40519 73385 40525
rect 72683 40423 72741 40429
rect 72683 40389 72695 40423
rect 72729 40420 72741 40423
rect 73342 40420 73370 40519
rect 73600 40516 73606 40528
rect 73658 40516 73664 40568
rect 73692 40516 73698 40568
rect 73750 40556 73756 40568
rect 73750 40528 75210 40556
rect 73750 40516 73756 40528
rect 73692 40420 73698 40432
rect 72729 40392 73698 40420
rect 72729 40389 72741 40392
rect 72683 40383 72741 40389
rect 73692 40380 73698 40392
rect 73750 40380 73756 40432
rect 74704 40420 74710 40432
rect 74665 40392 74710 40420
rect 74704 40380 74710 40392
rect 74762 40380 74768 40432
rect 75182 40429 75210 40528
rect 75274 40488 75302 40596
rect 78108 40584 78114 40636
rect 78166 40624 78172 40636
rect 78479 40627 78537 40633
rect 78479 40624 78491 40627
rect 78166 40596 78491 40624
rect 78166 40584 78172 40596
rect 78479 40593 78491 40596
rect 78525 40593 78537 40627
rect 78479 40587 78537 40593
rect 78568 40584 78574 40636
rect 78626 40624 78632 40636
rect 79230 40624 79258 40732
rect 79488 40692 79494 40704
rect 78626 40596 79258 40624
rect 79322 40664 79494 40692
rect 78626 40584 78632 40596
rect 75992 40516 75998 40568
rect 76050 40556 76056 40568
rect 76360 40556 76366 40568
rect 76050 40528 76366 40556
rect 76050 40516 76056 40528
rect 76360 40516 76366 40528
rect 76418 40556 76424 40568
rect 77927 40559 77985 40565
rect 77927 40556 77939 40559
rect 76418 40528 77939 40556
rect 76418 40516 76424 40528
rect 77927 40525 77939 40528
rect 77973 40556 77985 40559
rect 78203 40559 78261 40565
rect 78203 40556 78215 40559
rect 77973 40528 78215 40556
rect 77973 40525 77985 40528
rect 77927 40519 77985 40525
rect 78203 40525 78215 40528
rect 78249 40556 78261 40559
rect 79322 40556 79350 40664
rect 79488 40652 79494 40664
rect 79546 40652 79552 40704
rect 78249 40528 79350 40556
rect 79598 40556 79626 40732
rect 81055 40729 81067 40763
rect 81101 40729 81113 40763
rect 82340 40760 82346 40772
rect 82301 40732 82346 40760
rect 81055 40723 81113 40729
rect 79859 40627 79917 40633
rect 79859 40593 79871 40627
rect 79905 40624 79917 40627
rect 80592 40624 80598 40636
rect 79905 40596 80598 40624
rect 79905 40593 79917 40596
rect 79859 40587 79917 40593
rect 80592 40584 80598 40596
rect 80650 40584 80656 40636
rect 80868 40624 80874 40636
rect 80829 40596 80874 40624
rect 80868 40584 80874 40596
rect 80926 40584 80932 40636
rect 81070 40624 81098 40723
rect 82340 40720 82346 40732
rect 82398 40720 82404 40772
rect 88136 40760 88142 40772
rect 88097 40732 88142 40760
rect 88136 40720 88142 40732
rect 88194 40720 88200 40772
rect 81144 40652 81150 40704
rect 81202 40692 81208 40704
rect 81202 40664 82662 40692
rect 81202 40652 81208 40664
rect 82064 40624 82070 40636
rect 81070 40596 82070 40624
rect 82064 40584 82070 40596
rect 82122 40584 82128 40636
rect 82524 40624 82530 40636
rect 82485 40596 82530 40624
rect 82524 40584 82530 40596
rect 82582 40584 82588 40636
rect 82634 40624 82662 40664
rect 83815 40627 83873 40633
rect 83815 40624 83827 40627
rect 82634 40596 83827 40624
rect 83815 40593 83827 40596
rect 83861 40624 83873 40627
rect 83907 40627 83965 40633
rect 83907 40624 83919 40627
rect 83861 40596 83919 40624
rect 83861 40593 83873 40596
rect 83815 40587 83873 40593
rect 83907 40593 83919 40596
rect 83953 40624 83965 40627
rect 85008 40624 85014 40636
rect 83953 40596 85014 40624
rect 83953 40593 83965 40596
rect 83907 40587 83965 40593
rect 85008 40584 85014 40596
rect 85066 40584 85072 40636
rect 85468 40584 85474 40636
rect 85526 40624 85532 40636
rect 85526 40596 92138 40624
rect 85526 40584 85532 40596
rect 83628 40556 83634 40568
rect 79598 40528 83634 40556
rect 78249 40525 78261 40528
rect 78203 40519 78261 40525
rect 83628 40516 83634 40528
rect 83686 40516 83692 40568
rect 84180 40556 84186 40568
rect 84141 40528 84186 40556
rect 84180 40516 84186 40528
rect 84238 40516 84244 40568
rect 88136 40516 88142 40568
rect 88194 40556 88200 40568
rect 88231 40559 88289 40565
rect 88231 40556 88243 40559
rect 88194 40528 88243 40556
rect 88194 40516 88200 40528
rect 88231 40525 88243 40528
rect 88277 40525 88289 40559
rect 88504 40556 88510 40568
rect 88465 40528 88510 40556
rect 88231 40519 88289 40525
rect 88504 40516 88510 40528
rect 88562 40516 88568 40568
rect 90715 40559 90773 40565
rect 90715 40556 90727 40559
rect 90362 40528 90727 40556
rect 75274 40460 78246 40488
rect 75167 40423 75225 40429
rect 75167 40389 75179 40423
rect 75213 40420 75225 40423
rect 75992 40420 75998 40432
rect 75213 40392 75998 40420
rect 75213 40389 75225 40392
rect 75167 40383 75225 40389
rect 75992 40380 75998 40392
rect 76050 40380 76056 40432
rect 78108 40420 78114 40432
rect 78069 40392 78114 40420
rect 78108 40380 78114 40392
rect 78166 40380 78172 40432
rect 78218 40420 78246 40460
rect 79138 40460 83858 40488
rect 79138 40420 79166 40460
rect 78218 40392 79166 40420
rect 79212 40380 79218 40432
rect 79270 40420 79276 40432
rect 80687 40423 80745 40429
rect 80687 40420 80699 40423
rect 79270 40392 80699 40420
rect 79270 40380 79276 40392
rect 80687 40389 80699 40392
rect 80733 40420 80745 40423
rect 80868 40420 80874 40432
rect 80733 40392 80874 40420
rect 80733 40389 80745 40392
rect 80687 40383 80745 40389
rect 80868 40380 80874 40392
rect 80926 40380 80932 40432
rect 83830 40420 83858 40460
rect 85287 40423 85345 40429
rect 85287 40420 85299 40423
rect 83830 40392 85299 40420
rect 85287 40389 85299 40392
rect 85333 40389 85345 40423
rect 85287 40383 85345 40389
rect 88136 40380 88142 40432
rect 88194 40420 88200 40432
rect 89611 40423 89669 40429
rect 89611 40420 89623 40423
rect 88194 40392 89623 40420
rect 88194 40380 88200 40392
rect 89611 40389 89623 40392
rect 89657 40389 89669 40423
rect 89611 40383 89669 40389
rect 90160 40380 90166 40432
rect 90218 40420 90224 40432
rect 90362 40429 90390 40528
rect 90715 40525 90727 40528
rect 90761 40525 90773 40559
rect 90988 40556 90994 40568
rect 90949 40528 90994 40556
rect 90715 40519 90773 40525
rect 90988 40516 90994 40528
rect 91046 40516 91052 40568
rect 92110 40565 92138 40596
rect 92095 40559 92153 40565
rect 92095 40525 92107 40559
rect 92141 40525 92153 40559
rect 92095 40519 92153 40525
rect 90347 40423 90405 40429
rect 90347 40420 90359 40423
rect 90218 40392 90359 40420
rect 90218 40380 90224 40392
rect 90347 40389 90359 40392
rect 90393 40389 90405 40423
rect 90528 40420 90534 40432
rect 90489 40392 90534 40420
rect 90347 40383 90405 40389
rect 90528 40380 90534 40392
rect 90586 40420 90592 40432
rect 90988 40420 90994 40432
rect 90586 40392 90994 40420
rect 90586 40380 90592 40392
rect 90988 40380 90994 40392
rect 91046 40420 91052 40432
rect 92828 40420 92834 40432
rect 91046 40392 92834 40420
rect 91046 40380 91052 40392
rect 92828 40380 92834 40392
rect 92886 40380 92892 40432
rect 538 40330 93642 40352
rect 538 40278 3680 40330
rect 3732 40278 3744 40330
rect 3796 40278 3808 40330
rect 3860 40278 3872 40330
rect 3924 40278 9008 40330
rect 9060 40278 9072 40330
rect 9124 40278 9136 40330
rect 9188 40278 9200 40330
rect 9252 40278 14336 40330
rect 14388 40278 14400 40330
rect 14452 40278 14464 40330
rect 14516 40278 14528 40330
rect 14580 40278 19664 40330
rect 19716 40278 19728 40330
rect 19780 40278 19792 40330
rect 19844 40278 19856 40330
rect 19908 40278 24992 40330
rect 25044 40278 25056 40330
rect 25108 40278 25120 40330
rect 25172 40278 25184 40330
rect 25236 40278 30320 40330
rect 30372 40278 30384 40330
rect 30436 40278 30448 40330
rect 30500 40278 30512 40330
rect 30564 40278 35648 40330
rect 35700 40278 35712 40330
rect 35764 40278 35776 40330
rect 35828 40278 35840 40330
rect 35892 40278 40976 40330
rect 41028 40278 41040 40330
rect 41092 40278 41104 40330
rect 41156 40278 41168 40330
rect 41220 40278 46304 40330
rect 46356 40278 46368 40330
rect 46420 40278 46432 40330
rect 46484 40278 46496 40330
rect 46548 40278 51632 40330
rect 51684 40278 51696 40330
rect 51748 40278 51760 40330
rect 51812 40278 51824 40330
rect 51876 40278 56960 40330
rect 57012 40278 57024 40330
rect 57076 40278 57088 40330
rect 57140 40278 57152 40330
rect 57204 40278 62288 40330
rect 62340 40278 62352 40330
rect 62404 40278 62416 40330
rect 62468 40278 62480 40330
rect 62532 40278 67616 40330
rect 67668 40278 67680 40330
rect 67732 40278 67744 40330
rect 67796 40278 67808 40330
rect 67860 40278 72944 40330
rect 72996 40278 73008 40330
rect 73060 40278 73072 40330
rect 73124 40278 73136 40330
rect 73188 40278 78272 40330
rect 78324 40278 78336 40330
rect 78388 40278 78400 40330
rect 78452 40278 78464 40330
rect 78516 40278 83600 40330
rect 83652 40278 83664 40330
rect 83716 40278 83728 40330
rect 83780 40278 83792 40330
rect 83844 40278 88928 40330
rect 88980 40278 88992 40330
rect 89044 40278 89056 40330
rect 89108 40278 89120 40330
rect 89172 40278 93642 40330
rect 538 40256 93642 40278
rect 2484 40176 2490 40228
rect 2542 40216 2548 40228
rect 11960 40216 11966 40228
rect 2542 40188 11966 40216
rect 2542 40176 2548 40188
rect 11960 40176 11966 40188
rect 12018 40176 12024 40228
rect 12328 40176 12334 40228
rect 12386 40216 12392 40228
rect 12791 40219 12849 40225
rect 12791 40216 12803 40219
rect 12386 40188 12803 40216
rect 12386 40176 12392 40188
rect 12791 40185 12803 40188
rect 12837 40185 12849 40219
rect 14168 40216 14174 40228
rect 14129 40188 14174 40216
rect 12791 40179 12849 40185
rect 14168 40176 14174 40188
rect 14226 40176 14232 40228
rect 19504 40176 19510 40228
rect 19562 40216 19568 40228
rect 20151 40219 20209 40225
rect 20151 40216 20163 40219
rect 19562 40188 20163 40216
rect 19562 40176 19568 40188
rect 20151 40185 20163 40188
rect 20197 40185 20209 40219
rect 20151 40179 20209 40185
rect 39652 40176 39658 40228
rect 39710 40216 39716 40228
rect 41584 40216 41590 40228
rect 39710 40188 41590 40216
rect 39710 40176 39716 40188
rect 41584 40176 41590 40188
rect 41642 40176 41648 40228
rect 46555 40219 46613 40225
rect 46555 40185 46567 40219
rect 46601 40216 46613 40219
rect 46736 40216 46742 40228
rect 46601 40188 46742 40216
rect 46601 40185 46613 40188
rect 46555 40179 46613 40185
rect 46736 40176 46742 40188
rect 46794 40216 46800 40228
rect 49315 40219 49373 40225
rect 49315 40216 49327 40219
rect 46794 40188 49327 40216
rect 46794 40176 46800 40188
rect 49315 40185 49327 40188
rect 49361 40185 49373 40219
rect 49315 40179 49373 40185
rect 55663 40219 55721 40225
rect 55663 40185 55675 40219
rect 55709 40216 55721 40219
rect 55844 40216 55850 40228
rect 55709 40188 55850 40216
rect 55709 40185 55721 40188
rect 55663 40179 55721 40185
rect 8096 40148 8102 40160
rect 8057 40120 8102 40148
rect 8096 40108 8102 40120
rect 8154 40108 8160 40160
rect 11040 40108 11046 40160
rect 11098 40148 11104 40160
rect 13064 40148 13070 40160
rect 11098 40120 13070 40148
rect 11098 40108 11104 40120
rect 13064 40108 13070 40120
rect 13122 40108 13128 40160
rect 13524 40108 13530 40160
rect 13582 40148 13588 40160
rect 16652 40148 16658 40160
rect 13582 40120 16658 40148
rect 13582 40108 13588 40120
rect 16652 40108 16658 40120
rect 16710 40108 16716 40160
rect 21531 40151 21589 40157
rect 21531 40117 21543 40151
rect 21577 40148 21589 40151
rect 32752 40148 32758 40160
rect 21577 40120 32758 40148
rect 21577 40117 21589 40120
rect 21531 40111 21589 40117
rect 6164 40040 6170 40092
rect 6222 40080 6228 40092
rect 6351 40083 6409 40089
rect 6351 40080 6363 40083
rect 6222 40052 6363 40080
rect 6222 40040 6228 40052
rect 6351 40049 6363 40052
rect 6397 40049 6409 40083
rect 6351 40043 6409 40049
rect 6627 40083 6685 40089
rect 6627 40049 6639 40083
rect 6673 40080 6685 40083
rect 7820 40080 7826 40092
rect 6673 40052 7826 40080
rect 6673 40049 6685 40052
rect 6627 40043 6685 40049
rect 7820 40040 7826 40052
rect 7878 40040 7884 40092
rect 8004 40040 8010 40092
rect 8062 40080 8068 40092
rect 9111 40083 9169 40089
rect 9111 40080 9123 40083
rect 8062 40052 9123 40080
rect 8062 40040 8068 40052
rect 9111 40049 9123 40052
rect 9157 40049 9169 40083
rect 9111 40043 9169 40049
rect 12515 40083 12573 40089
rect 12515 40049 12527 40083
rect 12561 40080 12573 40083
rect 12561 40052 13938 40080
rect 12561 40049 12573 40052
rect 12515 40043 12573 40049
rect 13910 40024 13938 40052
rect 17388 40040 17394 40092
rect 17446 40080 17452 40092
rect 18679 40083 18737 40089
rect 18679 40080 18691 40083
rect 17446 40052 18691 40080
rect 17446 40040 17452 40052
rect 18679 40049 18691 40052
rect 18725 40080 18737 40083
rect 18771 40083 18829 40089
rect 18771 40080 18783 40083
rect 18725 40052 18783 40080
rect 18725 40049 18737 40052
rect 18679 40043 18737 40049
rect 18771 40049 18783 40052
rect 18817 40080 18829 40083
rect 20884 40080 20890 40092
rect 18817 40052 20890 40080
rect 18817 40049 18829 40052
rect 18771 40043 18829 40049
rect 20884 40040 20890 40052
rect 20942 40040 20948 40092
rect 8096 39972 8102 40024
rect 8154 40012 8160 40024
rect 8835 40015 8893 40021
rect 8835 40012 8847 40015
rect 8154 39984 8847 40012
rect 8154 39972 8160 39984
rect 8835 39981 8847 39984
rect 8881 40012 8893 40015
rect 10583 40015 10641 40021
rect 10583 40012 10595 40015
rect 8881 39984 10595 40012
rect 8881 39981 8893 39984
rect 8835 39975 8893 39981
rect 10583 39981 10595 39984
rect 10629 40012 10641 40015
rect 11040 40012 11046 40024
rect 10629 39984 11046 40012
rect 10629 39981 10641 39984
rect 10583 39975 10641 39981
rect 11040 39972 11046 39984
rect 11098 39972 11104 40024
rect 12607 40015 12665 40021
rect 12607 39981 12619 40015
rect 12653 40012 12665 40015
rect 13248 40012 13254 40024
rect 12653 39984 13254 40012
rect 12653 39981 12665 39984
rect 12607 39975 12665 39981
rect 13248 39972 13254 39984
rect 13306 39972 13312 40024
rect 13892 40012 13898 40024
rect 13853 39984 13898 40012
rect 13892 39972 13898 39984
rect 13950 39972 13956 40024
rect 13987 40015 14045 40021
rect 13987 39981 13999 40015
rect 14033 39981 14045 40015
rect 19044 40012 19050 40024
rect 19005 39984 19050 40012
rect 13987 39975 14045 39981
rect 8004 39944 8010 39956
rect 7965 39916 8010 39944
rect 8004 39904 8010 39916
rect 8062 39904 8068 39956
rect 10491 39947 10549 39953
rect 10491 39913 10503 39947
rect 10537 39944 10549 39947
rect 12236 39944 12242 39956
rect 10537 39916 12242 39944
rect 10537 39913 10549 39916
rect 10491 39907 10549 39913
rect 12236 39904 12242 39916
rect 12294 39904 12300 39956
rect 12972 39904 12978 39956
rect 13030 39944 13036 39956
rect 14002 39944 14030 39975
rect 19044 39972 19050 39984
rect 19102 39972 19108 40024
rect 21638 40021 21666 40120
rect 32752 40108 32758 40120
rect 32810 40108 32816 40160
rect 26131 40083 26189 40089
rect 26131 40049 26143 40083
rect 26177 40080 26189 40083
rect 27048 40080 27054 40092
rect 26177 40052 27054 40080
rect 26177 40049 26189 40052
rect 26131 40043 26189 40049
rect 27048 40040 27054 40052
rect 27106 40040 27112 40092
rect 27695 40083 27753 40089
rect 27695 40049 27707 40083
rect 27741 40080 27753 40083
rect 28796 40080 28802 40092
rect 27741 40052 28802 40080
rect 27741 40049 27753 40052
rect 27695 40043 27753 40049
rect 28796 40040 28802 40052
rect 28854 40040 28860 40092
rect 32387 40083 32445 40089
rect 32387 40049 32399 40083
rect 32433 40080 32445 40083
rect 34592 40080 34598 40092
rect 32433 40052 34598 40080
rect 32433 40049 32445 40052
rect 32387 40043 32445 40049
rect 34592 40040 34598 40052
rect 34650 40040 34656 40092
rect 38088 40080 38094 40092
rect 37278 40052 38094 40080
rect 21623 40015 21681 40021
rect 21623 39981 21635 40015
rect 21669 39981 21681 40015
rect 21623 39975 21681 39981
rect 25579 40015 25637 40021
rect 25579 39981 25591 40015
rect 25625 39981 25637 40015
rect 25579 39975 25637 39981
rect 25947 40015 26005 40021
rect 25947 39981 25959 40015
rect 25993 40012 26005 40015
rect 27140 40012 27146 40024
rect 25993 39984 27146 40012
rect 25993 39981 26005 39984
rect 25947 39975 26005 39981
rect 13030 39916 14030 39944
rect 25594 39944 25622 39975
rect 27140 39972 27146 39984
rect 27198 39972 27204 40024
rect 27235 40015 27293 40021
rect 27235 39981 27247 40015
rect 27281 39981 27293 40015
rect 27416 40012 27422 40024
rect 27377 39984 27422 40012
rect 27235 39975 27293 39981
rect 27250 39944 27278 39975
rect 27416 39972 27422 39984
rect 27474 39972 27480 40024
rect 28983 40015 29041 40021
rect 28983 39981 28995 40015
rect 29029 39981 29041 40015
rect 28983 39975 29041 39981
rect 29259 40015 29317 40021
rect 29259 39981 29271 40015
rect 29305 40012 29317 40015
rect 31372 40012 31378 40024
rect 29305 39984 31378 40012
rect 29305 39981 29317 39984
rect 29259 39975 29317 39981
rect 28998 39944 29026 39975
rect 31372 39972 31378 39984
rect 31430 39972 31436 40024
rect 31651 40015 31709 40021
rect 31651 39981 31663 40015
rect 31697 39981 31709 40015
rect 32108 40012 32114 40024
rect 32069 39984 32114 40012
rect 31651 39975 31709 39981
rect 31556 39944 31562 39956
rect 25594 39916 31562 39944
rect 13030 39904 13036 39916
rect 31556 39904 31562 39916
rect 31614 39944 31620 39956
rect 31666 39944 31694 39975
rect 32108 39972 32114 39984
rect 32166 39972 32172 40024
rect 37278 40021 37306 40052
rect 38088 40040 38094 40052
rect 38146 40040 38152 40092
rect 41602 40080 41630 40176
rect 41679 40083 41737 40089
rect 41679 40080 41691 40083
rect 41602 40052 41691 40080
rect 41679 40049 41691 40052
rect 41725 40049 41737 40083
rect 41679 40043 41737 40049
rect 45724 40040 45730 40092
rect 45782 40080 45788 40092
rect 47199 40083 47257 40089
rect 47199 40080 47211 40083
rect 45782 40052 47211 40080
rect 45782 40040 45788 40052
rect 47199 40049 47211 40052
rect 47245 40049 47257 40083
rect 47199 40043 47257 40049
rect 37263 40015 37321 40021
rect 37263 39981 37275 40015
rect 37309 39981 37321 40015
rect 37263 39975 37321 39981
rect 37539 40015 37597 40021
rect 37539 39981 37551 40015
rect 37585 40012 37597 40015
rect 39192 40012 39198 40024
rect 37585 39984 39198 40012
rect 37585 39981 37597 39984
rect 37539 39975 37597 39981
rect 39192 39972 39198 39984
rect 39250 39972 39256 40024
rect 41952 40012 41958 40024
rect 41913 39984 41958 40012
rect 41952 39972 41958 39984
rect 42010 39972 42016 40024
rect 46736 40012 46742 40024
rect 46697 39984 46742 40012
rect 46736 39972 46742 39984
rect 46794 39972 46800 40024
rect 47107 40015 47165 40021
rect 47107 39981 47119 40015
rect 47153 39981 47165 40015
rect 49330 40012 49358 40179
rect 55844 40176 55850 40188
rect 55902 40176 55908 40228
rect 61091 40219 61149 40225
rect 61091 40185 61103 40219
rect 61137 40216 61149 40219
rect 61364 40216 61370 40228
rect 61137 40188 61370 40216
rect 61137 40185 61149 40188
rect 61091 40179 61149 40185
rect 61364 40176 61370 40188
rect 61422 40176 61428 40228
rect 63480 40176 63486 40228
rect 63538 40216 63544 40228
rect 67436 40216 67442 40228
rect 63538 40188 67442 40216
rect 63538 40176 63544 40188
rect 67436 40176 67442 40188
rect 67494 40176 67500 40228
rect 72220 40216 72226 40228
rect 67914 40188 72226 40216
rect 50048 40108 50054 40160
rect 50106 40148 50112 40160
rect 50106 40120 54786 40148
rect 50106 40108 50112 40120
rect 50235 40083 50293 40089
rect 50235 40049 50247 40083
rect 50281 40080 50293 40083
rect 51428 40080 51434 40092
rect 50281 40052 51434 40080
rect 50281 40049 50293 40052
rect 50235 40043 50293 40049
rect 51428 40040 51434 40052
rect 51486 40040 51492 40092
rect 49496 40012 49502 40024
rect 49330 39984 49502 40012
rect 47107 39975 47165 39981
rect 31614 39916 31694 39944
rect 31614 39904 31620 39916
rect 34224 39904 34230 39956
rect 34282 39944 34288 39956
rect 35420 39944 35426 39956
rect 34282 39916 35426 39944
rect 34282 39904 34288 39916
rect 35420 39904 35426 39916
rect 35478 39904 35484 39956
rect 40296 39944 40302 39956
rect 36910 39916 40302 39944
rect 20240 39836 20246 39888
rect 20298 39876 20304 39888
rect 21807 39879 21865 39885
rect 21807 39876 21819 39879
rect 20298 39848 21819 39876
rect 20298 39836 20304 39848
rect 21807 39845 21819 39848
rect 21853 39845 21865 39879
rect 21807 39839 21865 39845
rect 25576 39836 25582 39888
rect 25634 39876 25640 39888
rect 27140 39876 27146 39888
rect 25634 39848 27146 39876
rect 25634 39836 25640 39848
rect 27140 39836 27146 39848
rect 27198 39836 27204 39888
rect 28428 39836 28434 39888
rect 28486 39876 28492 39888
rect 28799 39879 28857 39885
rect 28799 39876 28811 39879
rect 28486 39848 28811 39876
rect 28486 39836 28492 39848
rect 28799 39845 28811 39848
rect 28845 39845 28857 39879
rect 28799 39839 28857 39845
rect 33304 39836 33310 39888
rect 33362 39876 33368 39888
rect 36910 39876 36938 39916
rect 40296 39904 40302 39916
rect 40354 39904 40360 39956
rect 47122 39944 47150 39975
rect 49496 39972 49502 39984
rect 49554 39972 49560 40024
rect 50051 40015 50109 40021
rect 50051 39981 50063 40015
rect 50097 40012 50109 40015
rect 51152 40012 51158 40024
rect 50097 39984 51158 40012
rect 50097 39981 50109 39984
rect 50051 39975 50109 39981
rect 51152 39972 51158 39984
rect 51210 39972 51216 40024
rect 54648 40012 54654 40024
rect 54561 39984 54654 40012
rect 54648 39972 54654 39984
rect 54706 39972 54712 40024
rect 54758 40021 54786 40120
rect 57316 40108 57322 40160
rect 57374 40148 57380 40160
rect 64032 40148 64038 40160
rect 57374 40120 64038 40148
rect 57374 40108 57380 40120
rect 64032 40108 64038 40120
rect 64090 40108 64096 40160
rect 62100 40040 62106 40092
rect 62158 40080 62164 40092
rect 62158 40052 62790 40080
rect 62158 40040 62164 40052
rect 54743 40015 54801 40021
rect 54743 39981 54755 40015
rect 54789 39981 54801 40015
rect 54743 39975 54801 39981
rect 49864 39944 49870 39956
rect 47122 39916 49870 39944
rect 49864 39904 49870 39916
rect 49922 39904 49928 39956
rect 37076 39876 37082 39888
rect 33362 39848 36938 39876
rect 37037 39848 37082 39876
rect 33362 39836 33368 39848
rect 37076 39836 37082 39848
rect 37134 39836 37140 39888
rect 37907 39879 37965 39885
rect 37907 39845 37919 39879
rect 37953 39876 37965 39879
rect 38088 39876 38094 39888
rect 37953 39848 38094 39876
rect 37953 39845 37965 39848
rect 37907 39839 37965 39845
rect 38088 39836 38094 39848
rect 38146 39836 38152 39888
rect 43056 39876 43062 39888
rect 43017 39848 43062 39876
rect 43056 39836 43062 39848
rect 43114 39836 43120 39888
rect 54666 39876 54694 39972
rect 54758 39944 54786 39975
rect 55200 39972 55206 40024
rect 55258 40012 55264 40024
rect 55384 40012 55390 40024
rect 55258 39984 55303 40012
rect 55345 39984 55390 40012
rect 55258 39972 55264 39984
rect 55384 39972 55390 39984
rect 55442 39972 55448 40024
rect 56856 39972 56862 40024
rect 56914 40012 56920 40024
rect 57135 40015 57193 40021
rect 57135 40012 57147 40015
rect 56914 39984 57147 40012
rect 56914 39972 56920 39984
rect 57135 39981 57147 39984
rect 57181 39981 57193 40015
rect 57135 39975 57193 39981
rect 59895 40015 59953 40021
rect 59895 39981 59907 40015
rect 59941 39981 59953 40015
rect 59895 39975 59953 39981
rect 60079 40015 60137 40021
rect 60079 39981 60091 40015
rect 60125 40012 60137 40015
rect 60260 40012 60266 40024
rect 60125 39984 60266 40012
rect 60125 39981 60137 39984
rect 60079 39975 60137 39981
rect 59910 39944 59938 39975
rect 60260 39972 60266 39984
rect 60318 40012 60324 40024
rect 60631 40015 60689 40021
rect 60631 40012 60643 40015
rect 60318 39984 60643 40012
rect 60318 39972 60324 39984
rect 60631 39981 60643 39984
rect 60677 39981 60689 40015
rect 60631 39975 60689 39981
rect 60815 40015 60873 40021
rect 60815 39981 60827 40015
rect 60861 39981 60873 40015
rect 60815 39975 60873 39981
rect 62471 40015 62529 40021
rect 62471 39981 62483 40015
rect 62517 40012 62529 40015
rect 62652 40012 62658 40024
rect 62517 39984 62658 40012
rect 62517 39981 62529 39984
rect 62471 39975 62529 39981
rect 54758 39916 59938 39944
rect 59984 39904 59990 39956
rect 60042 39944 60048 39956
rect 60830 39944 60858 39975
rect 62652 39972 62658 39984
rect 62710 39972 62716 40024
rect 62762 40012 62790 40052
rect 65964 40040 65970 40092
rect 66022 40080 66028 40092
rect 67914 40080 67942 40188
rect 72220 40176 72226 40188
rect 72278 40176 72284 40228
rect 75900 40176 75906 40228
rect 75958 40216 75964 40228
rect 82527 40219 82585 40225
rect 82527 40216 82539 40219
rect 75958 40188 82539 40216
rect 75958 40176 75964 40188
rect 82527 40185 82539 40188
rect 82573 40185 82585 40219
rect 82527 40179 82585 40185
rect 74704 40148 74710 40160
rect 66022 40052 67942 40080
rect 68006 40120 74710 40148
rect 66022 40040 66028 40052
rect 68006 40012 68034 40120
rect 74704 40108 74710 40120
rect 74762 40108 74768 40160
rect 83720 40108 83726 40160
rect 83778 40148 83784 40160
rect 90528 40148 90534 40160
rect 83778 40120 90534 40148
rect 83778 40108 83784 40120
rect 90528 40108 90534 40120
rect 90586 40108 90592 40160
rect 68540 40080 68546 40092
rect 68501 40052 68546 40080
rect 68540 40040 68546 40052
rect 68598 40040 68604 40092
rect 71318 40052 71714 40080
rect 62762 39984 68034 40012
rect 68267 40015 68325 40021
rect 68267 39981 68279 40015
rect 68313 39981 68325 40015
rect 68448 40012 68454 40024
rect 68409 39984 68454 40012
rect 68267 39975 68325 39981
rect 62563 39947 62621 39953
rect 62563 39944 62575 39947
rect 60042 39916 62575 39944
rect 60042 39904 60048 39916
rect 62563 39913 62575 39916
rect 62609 39944 62621 39947
rect 63112 39944 63118 39956
rect 62609 39916 63118 39944
rect 62609 39913 62621 39916
rect 62563 39907 62621 39913
rect 63112 39904 63118 39916
rect 63170 39904 63176 39956
rect 67988 39904 67994 39956
rect 68046 39944 68052 39956
rect 68282 39944 68310 39975
rect 68448 39972 68454 39984
rect 68506 39972 68512 40024
rect 71208 40012 71214 40024
rect 68558 39984 71214 40012
rect 68558 39944 68586 39984
rect 71208 39972 71214 39984
rect 71266 40012 71272 40024
rect 71318 40021 71346 40052
rect 71303 40015 71361 40021
rect 71303 40012 71315 40015
rect 71266 39984 71315 40012
rect 71266 39972 71272 39984
rect 71303 39981 71315 39984
rect 71349 39981 71361 40015
rect 71576 40012 71582 40024
rect 71537 39984 71582 40012
rect 71303 39975 71361 39981
rect 71576 39972 71582 39984
rect 71634 39972 71640 40024
rect 71686 40012 71714 40052
rect 72036 40040 72042 40092
rect 72094 40080 72100 40092
rect 73324 40080 73330 40092
rect 72094 40052 73330 40080
rect 72094 40040 72100 40052
rect 73324 40040 73330 40052
rect 73382 40040 73388 40092
rect 75440 40040 75446 40092
rect 75498 40080 75504 40092
rect 75719 40083 75777 40089
rect 75719 40080 75731 40083
rect 75498 40052 75731 40080
rect 75498 40040 75504 40052
rect 75719 40049 75731 40052
rect 75765 40049 75777 40083
rect 78019 40083 78077 40089
rect 78019 40080 78031 40083
rect 75719 40043 75777 40049
rect 76930 40052 78031 40080
rect 72864 40012 72870 40024
rect 71686 39984 72870 40012
rect 72864 39972 72870 39984
rect 72922 40012 72928 40024
rect 73603 40015 73661 40021
rect 73603 40012 73615 40015
rect 72922 39984 73615 40012
rect 72922 39972 72928 39984
rect 73603 39981 73615 39984
rect 73649 39981 73661 40015
rect 74060 40012 74066 40024
rect 74021 39984 74066 40012
rect 73603 39975 73661 39981
rect 74060 39972 74066 39984
rect 74118 39972 74124 40024
rect 75256 39972 75262 40024
rect 75314 40012 75320 40024
rect 75903 40015 75961 40021
rect 75903 40012 75915 40015
rect 75314 39984 75915 40012
rect 75314 39972 75320 39984
rect 75903 39981 75915 39984
rect 75949 40012 75961 40015
rect 76455 40015 76513 40021
rect 76455 40012 76467 40015
rect 75949 39984 76467 40012
rect 75949 39981 75961 39984
rect 75903 39975 75961 39981
rect 76455 39981 76467 39984
rect 76501 39981 76513 40015
rect 76455 39975 76513 39981
rect 76639 40015 76697 40021
rect 76639 39981 76651 40015
rect 76685 40012 76697 40015
rect 76930 40012 76958 40052
rect 78019 40049 78031 40052
rect 78065 40049 78077 40083
rect 78019 40043 78077 40049
rect 78939 40083 78997 40089
rect 78939 40049 78951 40083
rect 78985 40080 78997 40083
rect 81423 40083 81481 40089
rect 78985 40052 81374 40080
rect 78985 40049 78997 40052
rect 78939 40043 78997 40049
rect 76685 39984 76958 40012
rect 76685 39981 76697 39984
rect 76639 39975 76697 39981
rect 72772 39944 72778 39956
rect 68046 39916 68586 39944
rect 70950 39916 72778 39944
rect 68046 39904 68052 39916
rect 55016 39876 55022 39888
rect 54666 39848 55022 39876
rect 55016 39836 55022 39848
rect 55074 39836 55080 39888
rect 55384 39836 55390 39888
rect 55442 39876 55448 39888
rect 55844 39876 55850 39888
rect 55442 39848 55850 39876
rect 55442 39836 55448 39848
rect 55844 39836 55850 39848
rect 55902 39876 55908 39888
rect 57227 39879 57285 39885
rect 57227 39876 57239 39879
rect 55902 39848 57239 39876
rect 55902 39836 55908 39848
rect 57227 39845 57239 39848
rect 57273 39845 57285 39879
rect 57227 39839 57285 39845
rect 67160 39836 67166 39888
rect 67218 39876 67224 39888
rect 70950 39876 70978 39916
rect 72772 39904 72778 39916
rect 72830 39904 72836 39956
rect 74520 39904 74526 39956
rect 74578 39944 74584 39956
rect 74578 39916 75854 39944
rect 74578 39904 74584 39916
rect 71116 39876 71122 39888
rect 67218 39848 70978 39876
rect 71077 39848 71122 39876
rect 67218 39836 67224 39848
rect 71116 39836 71122 39848
rect 71174 39836 71180 39888
rect 73600 39836 73606 39888
rect 73658 39876 73664 39888
rect 73695 39879 73753 39885
rect 73695 39876 73707 39879
rect 73658 39848 73707 39876
rect 73658 39836 73664 39848
rect 73695 39845 73707 39848
rect 73741 39845 73753 39879
rect 73695 39839 73753 39845
rect 74152 39836 74158 39888
rect 74210 39876 74216 39888
rect 75167 39879 75225 39885
rect 75167 39876 75179 39879
rect 74210 39848 75179 39876
rect 74210 39836 74216 39848
rect 75167 39845 75179 39848
rect 75213 39876 75225 39879
rect 75256 39876 75262 39888
rect 75213 39848 75262 39876
rect 75213 39845 75225 39848
rect 75167 39839 75225 39845
rect 75256 39836 75262 39848
rect 75314 39876 75320 39888
rect 75351 39879 75409 39885
rect 75351 39876 75363 39879
rect 75314 39848 75363 39876
rect 75314 39836 75320 39848
rect 75351 39845 75363 39848
rect 75397 39845 75409 39879
rect 75351 39839 75409 39845
rect 75440 39836 75446 39888
rect 75498 39876 75504 39888
rect 75535 39879 75593 39885
rect 75535 39876 75547 39879
rect 75498 39848 75547 39876
rect 75498 39836 75504 39848
rect 75535 39845 75547 39848
rect 75581 39845 75593 39879
rect 75826 39876 75854 39916
rect 76268 39904 76274 39956
rect 76326 39944 76332 39956
rect 76654 39944 76682 39975
rect 77096 39972 77102 40024
rect 77154 40012 77160 40024
rect 77927 40015 77985 40021
rect 77154 39984 77878 40012
rect 77154 39972 77160 39984
rect 76326 39916 76682 39944
rect 77007 39947 77065 39953
rect 76326 39904 76332 39916
rect 77007 39913 77019 39947
rect 77053 39944 77065 39947
rect 77648 39944 77654 39956
rect 77053 39916 77654 39944
rect 77053 39913 77065 39916
rect 77007 39907 77065 39913
rect 77648 39904 77654 39916
rect 77706 39904 77712 39956
rect 77850 39944 77878 39984
rect 77927 39981 77939 40015
rect 77973 40012 77985 40015
rect 79856 40012 79862 40024
rect 77973 39984 79862 40012
rect 77973 39981 77985 39984
rect 77927 39975 77985 39981
rect 79856 39972 79862 39984
rect 79914 39972 79920 40024
rect 81055 40015 81113 40021
rect 81055 39981 81067 40015
rect 81101 40012 81113 40015
rect 81144 40012 81150 40024
rect 81101 39984 81150 40012
rect 81101 39981 81113 39984
rect 81055 39975 81113 39981
rect 81144 39972 81150 39984
rect 81202 39972 81208 40024
rect 81346 40012 81374 40052
rect 81423 40049 81435 40083
rect 81469 40080 81481 40083
rect 82340 40080 82346 40092
rect 81469 40052 82346 40080
rect 81469 40049 81481 40052
rect 81423 40043 81481 40049
rect 82340 40040 82346 40052
rect 82398 40040 82404 40092
rect 88412 40080 88418 40092
rect 82450 40052 88418 40080
rect 82450 40012 82478 40052
rect 88412 40040 88418 40052
rect 88470 40040 88476 40092
rect 89332 40080 89338 40092
rect 89293 40052 89338 40080
rect 89332 40040 89338 40052
rect 89390 40040 89396 40092
rect 81346 39984 82478 40012
rect 83904 39972 83910 40024
rect 83962 40012 83968 40024
rect 85379 40015 85437 40021
rect 85379 40012 85391 40015
rect 83962 39984 85391 40012
rect 83962 39972 83968 39984
rect 85379 39981 85391 39984
rect 85425 39981 85437 40015
rect 85836 40012 85842 40024
rect 85797 39984 85842 40012
rect 85379 39975 85437 39981
rect 85394 39944 85422 39975
rect 85836 39972 85842 39984
rect 85894 39972 85900 40024
rect 88599 40015 88657 40021
rect 88599 39981 88611 40015
rect 88645 39981 88657 40015
rect 88599 39975 88657 39981
rect 88614 39944 88642 39975
rect 88780 39972 88786 40024
rect 88838 40012 88844 40024
rect 89059 40015 89117 40021
rect 89059 40012 89071 40015
rect 88838 39984 89071 40012
rect 88838 39972 88844 39984
rect 89059 39981 89071 39984
rect 89105 39981 89117 40015
rect 89059 39975 89117 39981
rect 88688 39944 88694 39956
rect 77850 39916 81190 39944
rect 85394 39916 88694 39944
rect 78939 39879 78997 39885
rect 78939 39876 78951 39879
rect 75826 39848 78951 39876
rect 75535 39839 75593 39845
rect 78939 39845 78951 39848
rect 78985 39845 78997 39879
rect 81162 39876 81190 39916
rect 88688 39904 88694 39916
rect 88746 39904 88752 39956
rect 82800 39876 82806 39888
rect 81162 39848 82806 39876
rect 78939 39839 78997 39845
rect 82800 39836 82806 39848
rect 82858 39836 82864 39888
rect 85652 39876 85658 39888
rect 85613 39848 85658 39876
rect 85652 39836 85658 39848
rect 85710 39836 85716 39888
rect 538 39786 93642 39808
rect 538 39734 6344 39786
rect 6396 39734 6408 39786
rect 6460 39734 6472 39786
rect 6524 39734 6536 39786
rect 6588 39734 11672 39786
rect 11724 39734 11736 39786
rect 11788 39734 11800 39786
rect 11852 39734 11864 39786
rect 11916 39734 17000 39786
rect 17052 39734 17064 39786
rect 17116 39734 17128 39786
rect 17180 39734 17192 39786
rect 17244 39734 22328 39786
rect 22380 39734 22392 39786
rect 22444 39734 22456 39786
rect 22508 39734 22520 39786
rect 22572 39734 27656 39786
rect 27708 39734 27720 39786
rect 27772 39734 27784 39786
rect 27836 39734 27848 39786
rect 27900 39734 32984 39786
rect 33036 39734 33048 39786
rect 33100 39734 33112 39786
rect 33164 39734 33176 39786
rect 33228 39734 38312 39786
rect 38364 39734 38376 39786
rect 38428 39734 38440 39786
rect 38492 39734 38504 39786
rect 38556 39734 43640 39786
rect 43692 39734 43704 39786
rect 43756 39734 43768 39786
rect 43820 39734 43832 39786
rect 43884 39734 48968 39786
rect 49020 39734 49032 39786
rect 49084 39734 49096 39786
rect 49148 39734 49160 39786
rect 49212 39734 54296 39786
rect 54348 39734 54360 39786
rect 54412 39734 54424 39786
rect 54476 39734 54488 39786
rect 54540 39734 59624 39786
rect 59676 39734 59688 39786
rect 59740 39734 59752 39786
rect 59804 39734 59816 39786
rect 59868 39734 64952 39786
rect 65004 39734 65016 39786
rect 65068 39734 65080 39786
rect 65132 39734 65144 39786
rect 65196 39734 70280 39786
rect 70332 39734 70344 39786
rect 70396 39734 70408 39786
rect 70460 39734 70472 39786
rect 70524 39734 75608 39786
rect 75660 39734 75672 39786
rect 75724 39734 75736 39786
rect 75788 39734 75800 39786
rect 75852 39734 80936 39786
rect 80988 39734 81000 39786
rect 81052 39734 81064 39786
rect 81116 39734 81128 39786
rect 81180 39734 86264 39786
rect 86316 39734 86328 39786
rect 86380 39734 86392 39786
rect 86444 39734 86456 39786
rect 86508 39734 91592 39786
rect 91644 39734 91656 39786
rect 91708 39734 91720 39786
rect 91772 39734 91784 39786
rect 91836 39734 93642 39786
rect 538 39712 93642 39734
rect 4143 39675 4201 39681
rect 4143 39641 4155 39675
rect 4189 39672 4201 39675
rect 4600 39672 4606 39684
rect 4189 39644 4606 39672
rect 4189 39641 4201 39644
rect 4143 39635 4201 39641
rect 4600 39632 4606 39644
rect 4658 39632 4664 39684
rect 10948 39632 10954 39684
rect 11006 39672 11012 39684
rect 15916 39672 15922 39684
rect 11006 39644 15922 39672
rect 11006 39632 11012 39644
rect 15916 39632 15922 39644
rect 15974 39632 15980 39684
rect 37355 39675 37413 39681
rect 37355 39641 37367 39675
rect 37401 39672 37413 39675
rect 38088 39672 38094 39684
rect 37401 39644 38094 39672
rect 37401 39641 37413 39644
rect 37355 39635 37413 39641
rect 38088 39632 38094 39644
rect 38146 39672 38152 39684
rect 39468 39672 39474 39684
rect 38146 39644 39474 39672
rect 38146 39632 38152 39644
rect 39468 39632 39474 39644
rect 39526 39632 39532 39684
rect 41679 39675 41737 39681
rect 41679 39641 41691 39675
rect 41725 39672 41737 39675
rect 41952 39672 41958 39684
rect 41725 39644 41958 39672
rect 41725 39641 41737 39644
rect 41679 39635 41737 39641
rect 41952 39632 41958 39644
rect 42010 39632 42016 39684
rect 42872 39632 42878 39684
rect 42930 39672 42936 39684
rect 47656 39672 47662 39684
rect 42930 39644 47662 39672
rect 42930 39632 42936 39644
rect 47656 39632 47662 39644
rect 47714 39632 47720 39684
rect 49496 39672 49502 39684
rect 49457 39644 49502 39672
rect 49496 39632 49502 39644
rect 49554 39632 49560 39684
rect 49772 39672 49778 39684
rect 49733 39644 49778 39672
rect 49772 39632 49778 39644
rect 49830 39632 49836 39684
rect 49864 39632 49870 39684
rect 49922 39672 49928 39684
rect 54467 39675 54525 39681
rect 54467 39672 54479 39675
rect 49922 39644 54479 39672
rect 49922 39632 49928 39644
rect 54467 39641 54479 39644
rect 54513 39641 54525 39675
rect 54467 39635 54525 39641
rect 55034 39644 55246 39672
rect 13616 39604 13622 39616
rect 12162 39576 13622 39604
rect 5336 39496 5342 39548
rect 5394 39536 5400 39548
rect 12162 39545 12190 39576
rect 13616 39564 13622 39576
rect 13674 39564 13680 39616
rect 13892 39564 13898 39616
rect 13950 39604 13956 39616
rect 18768 39604 18774 39616
rect 13950 39576 18774 39604
rect 13950 39564 13956 39576
rect 12147 39539 12205 39545
rect 5394 39508 12098 39536
rect 5394 39496 5400 39508
rect 3496 39468 3502 39480
rect 3457 39440 3502 39468
rect 3496 39428 3502 39440
rect 3554 39428 3560 39480
rect 11500 39428 11506 39480
rect 11558 39468 11564 39480
rect 11963 39471 12021 39477
rect 11963 39468 11975 39471
rect 11558 39440 11975 39468
rect 11558 39428 11564 39440
rect 11963 39437 11975 39440
rect 12009 39437 12021 39471
rect 11963 39431 12021 39437
rect 12070 39400 12098 39508
rect 12147 39505 12159 39539
rect 12193 39505 12205 39539
rect 12147 39499 12205 39505
rect 12236 39496 12242 39548
rect 12294 39536 12300 39548
rect 17314 39545 17342 39576
rect 18768 39564 18774 39576
rect 18826 39564 18832 39616
rect 21252 39564 21258 39616
rect 21310 39604 21316 39616
rect 21623 39607 21681 39613
rect 21623 39604 21635 39607
rect 21310 39576 21635 39604
rect 21310 39564 21316 39576
rect 21623 39573 21635 39576
rect 21669 39573 21681 39607
rect 32292 39604 32298 39616
rect 21623 39567 21681 39573
rect 27894 39576 32154 39604
rect 32253 39576 32298 39604
rect 12515 39539 12573 39545
rect 12515 39536 12527 39539
rect 12294 39508 12527 39536
rect 12294 39496 12300 39508
rect 12515 39505 12527 39508
rect 12561 39505 12573 39539
rect 12515 39499 12573 39505
rect 17299 39539 17357 39545
rect 17299 39505 17311 39539
rect 17345 39505 17357 39539
rect 17480 39536 17486 39548
rect 17441 39508 17486 39536
rect 17299 39499 17357 39505
rect 17480 39496 17486 39508
rect 17538 39496 17544 39548
rect 27894 39545 27922 39576
rect 17575 39539 17633 39545
rect 17575 39505 17587 39539
rect 17621 39536 17633 39539
rect 21163 39539 21221 39545
rect 17621 39508 18262 39536
rect 17621 39505 17633 39508
rect 17575 39499 17633 39505
rect 12328 39428 12334 39480
rect 12386 39468 12392 39480
rect 12423 39471 12481 39477
rect 12423 39468 12435 39471
rect 12386 39440 12435 39468
rect 12386 39428 12392 39440
rect 12423 39437 12435 39440
rect 12469 39437 12481 39471
rect 12423 39431 12481 39437
rect 17388 39400 17394 39412
rect 12070 39372 17394 39400
rect 17388 39360 17394 39372
rect 17446 39360 17452 39412
rect 11779 39335 11837 39341
rect 11779 39301 11791 39335
rect 11825 39332 11837 39335
rect 12236 39332 12242 39344
rect 11825 39304 12242 39332
rect 11825 39301 11837 39304
rect 11779 39295 11837 39301
rect 12236 39292 12242 39304
rect 12294 39292 12300 39344
rect 17756 39332 17762 39344
rect 17717 39304 17762 39332
rect 17756 39292 17762 39304
rect 17814 39292 17820 39344
rect 18234 39341 18262 39508
rect 21163 39505 21175 39539
rect 21209 39536 21221 39539
rect 27327 39539 27385 39545
rect 21209 39508 21850 39536
rect 21209 39505 21221 39508
rect 21163 39499 21221 39505
rect 21068 39468 21074 39480
rect 21029 39440 21074 39468
rect 21068 39428 21074 39440
rect 21126 39428 21132 39480
rect 21822 39409 21850 39508
rect 27327 39505 27339 39539
rect 27373 39536 27385 39539
rect 27879 39539 27937 39545
rect 27879 39536 27891 39539
rect 27373 39508 27891 39536
rect 27373 39505 27385 39508
rect 27327 39499 27385 39505
rect 27879 39505 27891 39508
rect 27925 39505 27937 39539
rect 27879 39499 27937 39505
rect 27968 39496 27974 39548
rect 28026 39536 28032 39548
rect 28063 39539 28121 39545
rect 28063 39536 28075 39539
rect 28026 39508 28075 39536
rect 28026 39496 28032 39508
rect 28063 39505 28075 39508
rect 28109 39505 28121 39539
rect 31556 39536 31562 39548
rect 31517 39508 31562 39536
rect 28063 39499 28121 39505
rect 31556 39496 31562 39508
rect 31614 39496 31620 39548
rect 32016 39536 32022 39548
rect 31977 39508 32022 39536
rect 32016 39496 32022 39508
rect 32074 39496 32080 39548
rect 32126 39536 32154 39576
rect 32292 39564 32298 39576
rect 32350 39564 32356 39616
rect 32752 39564 32758 39616
rect 32810 39604 32816 39616
rect 55034 39604 55062 39644
rect 32810 39576 55062 39604
rect 55218 39604 55246 39644
rect 55292 39632 55298 39684
rect 55350 39672 55356 39684
rect 55939 39675 55997 39681
rect 55939 39672 55951 39675
rect 55350 39644 55951 39672
rect 55350 39632 55356 39644
rect 55939 39641 55951 39644
rect 55985 39672 55997 39675
rect 56672 39672 56678 39684
rect 55985 39644 56678 39672
rect 55985 39641 55997 39644
rect 55939 39635 55997 39641
rect 56672 39632 56678 39644
rect 56730 39672 56736 39684
rect 57316 39672 57322 39684
rect 56730 39644 57322 39672
rect 56730 39632 56736 39644
rect 57316 39632 57322 39644
rect 57374 39632 57380 39684
rect 58604 39632 58610 39684
rect 58662 39672 58668 39684
rect 62100 39672 62106 39684
rect 58662 39644 62106 39672
rect 58662 39632 58668 39644
rect 62100 39632 62106 39644
rect 62158 39632 62164 39684
rect 62210 39644 78338 39672
rect 62210 39604 62238 39644
rect 55218 39576 62238 39604
rect 32810 39564 32816 39576
rect 70748 39564 70754 39616
rect 70806 39604 70812 39616
rect 73327 39607 73385 39613
rect 70806 39576 73002 39604
rect 70806 39564 70812 39576
rect 33491 39539 33549 39545
rect 33491 39536 33503 39539
rect 32126 39508 33503 39536
rect 33491 39505 33503 39508
rect 33537 39536 33549 39539
rect 34040 39536 34046 39548
rect 33537 39508 34046 39536
rect 33537 39505 33549 39508
rect 33491 39499 33549 39505
rect 34040 39496 34046 39508
rect 34098 39496 34104 39548
rect 34227 39539 34285 39545
rect 34227 39505 34239 39539
rect 34273 39536 34285 39539
rect 34868 39536 34874 39548
rect 34273 39508 34874 39536
rect 34273 39505 34285 39508
rect 34227 39499 34285 39505
rect 34868 39496 34874 39508
rect 34926 39496 34932 39548
rect 36340 39496 36346 39548
rect 36398 39536 36404 39548
rect 37171 39539 37229 39545
rect 37171 39536 37183 39539
rect 36398 39508 37183 39536
rect 36398 39496 36404 39508
rect 37171 39505 37183 39508
rect 37217 39505 37229 39539
rect 37171 39499 37229 39505
rect 40388 39496 40394 39548
rect 40446 39536 40452 39548
rect 40667 39539 40725 39545
rect 40667 39536 40679 39539
rect 40446 39508 40679 39536
rect 40446 39496 40452 39508
rect 40667 39505 40679 39508
rect 40713 39536 40725 39539
rect 41219 39539 41277 39545
rect 41219 39536 41231 39539
rect 40713 39508 41231 39536
rect 40713 39505 40725 39508
rect 40667 39499 40725 39505
rect 41219 39505 41231 39508
rect 41265 39505 41277 39539
rect 41219 39499 41277 39505
rect 41308 39496 41314 39548
rect 41366 39536 41372 39548
rect 41403 39539 41461 39545
rect 41403 39536 41415 39539
rect 41366 39508 41415 39536
rect 41366 39496 41372 39508
rect 41403 39505 41415 39508
rect 41449 39536 41461 39539
rect 42783 39539 42841 39545
rect 41449 39508 41906 39536
rect 41449 39505 41461 39508
rect 41403 39499 41461 39505
rect 27235 39471 27293 39477
rect 27235 39437 27247 39471
rect 27281 39437 27293 39471
rect 27235 39431 27293 39437
rect 21807 39403 21865 39409
rect 21807 39369 21819 39403
rect 21853 39400 21865 39403
rect 24196 39400 24202 39412
rect 21853 39372 24202 39400
rect 21853 39369 21865 39372
rect 21807 39363 21865 39369
rect 24196 39360 24202 39372
rect 24254 39360 24260 39412
rect 27048 39400 27054 39412
rect 26961 39372 27054 39400
rect 27048 39360 27054 39372
rect 27106 39400 27112 39412
rect 27250 39400 27278 39431
rect 31924 39428 31930 39480
rect 31982 39468 31988 39480
rect 33304 39468 33310 39480
rect 31982 39440 33310 39468
rect 31982 39428 31988 39440
rect 33304 39428 33310 39440
rect 33362 39428 33368 39480
rect 40575 39471 40633 39477
rect 40575 39437 40587 39471
rect 40621 39437 40633 39471
rect 41878 39468 41906 39508
rect 42783 39505 42795 39539
rect 42829 39536 42841 39539
rect 43056 39536 43062 39548
rect 42829 39508 43062 39536
rect 42829 39505 42841 39508
rect 42783 39499 42841 39505
rect 42875 39471 42933 39477
rect 42875 39468 42887 39471
rect 41878 39440 42887 39468
rect 40575 39431 40633 39437
rect 42875 39437 42887 39440
rect 42921 39437 42933 39471
rect 42875 39431 42933 39437
rect 28244 39400 28250 39412
rect 27106 39372 27278 39400
rect 28205 39372 28250 39400
rect 27106 39360 27112 39372
rect 18219 39335 18277 39341
rect 18219 39301 18231 39335
rect 18265 39332 18277 39335
rect 18308 39332 18314 39344
rect 18265 39304 18314 39332
rect 18265 39301 18277 39304
rect 18219 39295 18277 39301
rect 18308 39292 18314 39304
rect 18366 39292 18372 39344
rect 27250 39332 27278 39372
rect 28244 39360 28250 39372
rect 28302 39360 28308 39412
rect 37812 39400 37818 39412
rect 28354 39372 37818 39400
rect 28354 39332 28382 39372
rect 37812 39360 37818 39372
rect 37870 39360 37876 39412
rect 40590 39400 40618 39431
rect 42982 39400 43010 39508
rect 43056 39496 43062 39508
rect 43114 39496 43120 39548
rect 49496 39496 49502 39548
rect 49554 39536 49560 39548
rect 49683 39539 49741 39545
rect 49683 39536 49695 39539
rect 49554 39508 49695 39536
rect 49554 39496 49560 39508
rect 49683 39505 49695 39508
rect 49729 39505 49741 39539
rect 49683 39499 49741 39505
rect 50235 39539 50293 39545
rect 50235 39505 50247 39539
rect 50281 39536 50293 39539
rect 50281 39508 52578 39536
rect 50281 39505 50293 39508
rect 50235 39499 50293 39505
rect 52550 39468 52578 39508
rect 53912 39496 53918 39548
rect 53970 39536 53976 39548
rect 54099 39539 54157 39545
rect 54099 39536 54111 39539
rect 53970 39508 54111 39536
rect 53970 39496 53976 39508
rect 54099 39505 54111 39508
rect 54145 39536 54157 39539
rect 55019 39539 55077 39545
rect 55019 39536 55031 39539
rect 54145 39508 55031 39536
rect 54145 39505 54157 39508
rect 54099 39499 54157 39505
rect 55019 39505 55031 39508
rect 55065 39505 55077 39539
rect 55384 39536 55390 39548
rect 55345 39508 55390 39536
rect 55019 39499 55077 39505
rect 55384 39496 55390 39508
rect 55442 39496 55448 39548
rect 56856 39496 56862 39548
rect 56914 39536 56920 39548
rect 57043 39539 57101 39545
rect 57043 39536 57055 39539
rect 56914 39508 57055 39536
rect 56914 39496 56920 39508
rect 57043 39505 57055 39508
rect 57089 39505 57101 39539
rect 57043 39499 57101 39505
rect 64676 39496 64682 39548
rect 64734 39536 64740 39548
rect 67804 39536 67810 39548
rect 64734 39508 67810 39536
rect 64734 39496 64740 39508
rect 67804 39496 67810 39508
rect 67862 39496 67868 39548
rect 67988 39536 67994 39548
rect 67949 39508 67994 39536
rect 67988 39496 67994 39508
rect 68046 39496 68052 39548
rect 68264 39536 68270 39548
rect 68225 39508 68270 39536
rect 68264 39496 68270 39508
rect 68322 39496 68328 39548
rect 70840 39536 70846 39548
rect 70801 39508 70846 39536
rect 70840 39496 70846 39508
rect 70898 39496 70904 39548
rect 72864 39536 72870 39548
rect 72825 39508 72870 39536
rect 72864 39496 72870 39508
rect 72922 39496 72928 39548
rect 54648 39468 54654 39480
rect 52550 39440 54654 39468
rect 54648 39428 54654 39440
rect 54706 39428 54712 39480
rect 55111 39471 55169 39477
rect 55111 39437 55123 39471
rect 55157 39468 55169 39471
rect 55200 39468 55206 39480
rect 55157 39440 55206 39468
rect 55157 39437 55169 39440
rect 55111 39431 55169 39437
rect 55200 39428 55206 39440
rect 55258 39428 55264 39480
rect 55295 39471 55353 39477
rect 55295 39437 55307 39471
rect 55341 39468 55353 39471
rect 55755 39471 55813 39477
rect 55755 39468 55767 39471
rect 55341 39440 55767 39468
rect 55341 39437 55353 39440
rect 55295 39431 55353 39437
rect 55755 39437 55767 39440
rect 55801 39468 55813 39471
rect 65047 39471 65105 39477
rect 55801 39440 57086 39468
rect 55801 39437 55813 39440
rect 55755 39431 55813 39437
rect 43151 39403 43209 39409
rect 43151 39400 43163 39403
rect 40590 39372 42918 39400
rect 42982 39372 43163 39400
rect 27250 39304 28382 39332
rect 30636 39292 30642 39344
rect 30694 39332 30700 39344
rect 31832 39332 31838 39344
rect 30694 39304 31838 39332
rect 30694 39292 30700 39304
rect 31832 39292 31838 39304
rect 31890 39292 31896 39344
rect 34500 39332 34506 39344
rect 34461 39304 34506 39332
rect 34500 39292 34506 39304
rect 34558 39292 34564 39344
rect 34868 39332 34874 39344
rect 34829 39304 34874 39332
rect 34868 39292 34874 39304
rect 34926 39292 34932 39344
rect 42890 39332 42918 39372
rect 43151 39369 43163 39372
rect 43197 39400 43209 39403
rect 56580 39400 56586 39412
rect 43197 39372 56586 39400
rect 43197 39369 43209 39372
rect 43151 39363 43209 39369
rect 56580 39360 56586 39372
rect 56638 39360 56644 39412
rect 56764 39360 56770 39412
rect 56822 39400 56828 39412
rect 56859 39403 56917 39409
rect 56859 39400 56871 39403
rect 56822 39372 56871 39400
rect 56822 39360 56828 39372
rect 56859 39369 56871 39372
rect 56905 39369 56917 39403
rect 56859 39363 56917 39369
rect 43056 39332 43062 39344
rect 42890 39304 43062 39332
rect 43056 39292 43062 39304
rect 43114 39332 43120 39344
rect 45172 39332 45178 39344
rect 43114 39304 45178 39332
rect 43114 39292 43120 39304
rect 45172 39292 45178 39304
rect 45230 39292 45236 39344
rect 54188 39332 54194 39344
rect 54149 39304 54194 39332
rect 54188 39292 54194 39304
rect 54246 39292 54252 39344
rect 57058 39332 57086 39440
rect 65047 39437 65059 39471
rect 65093 39468 65105 39471
rect 65228 39468 65234 39480
rect 65093 39440 65234 39468
rect 65093 39437 65105 39440
rect 65047 39431 65105 39437
rect 65228 39428 65234 39440
rect 65286 39428 65292 39480
rect 65504 39468 65510 39480
rect 65465 39440 65510 39468
rect 65504 39428 65510 39440
rect 65562 39428 65568 39480
rect 68172 39468 68178 39480
rect 68133 39440 68178 39468
rect 68172 39428 68178 39440
rect 68230 39428 68236 39480
rect 71208 39468 71214 39480
rect 71134 39440 71214 39468
rect 71027 39403 71085 39409
rect 71027 39369 71039 39403
rect 71073 39400 71085 39403
rect 71134 39400 71162 39440
rect 71208 39428 71214 39440
rect 71266 39428 71272 39480
rect 72974 39468 73002 39576
rect 73327 39573 73339 39607
rect 73373 39604 73385 39607
rect 73876 39604 73882 39616
rect 73373 39576 73882 39604
rect 73373 39573 73385 39576
rect 73327 39567 73385 39573
rect 73876 39564 73882 39576
rect 73934 39564 73940 39616
rect 77283 39607 77341 39613
rect 77283 39573 77295 39607
rect 77329 39604 77341 39607
rect 77464 39604 77470 39616
rect 77329 39576 77470 39604
rect 77329 39573 77341 39576
rect 77283 39567 77341 39573
rect 73143 39539 73201 39545
rect 73143 39505 73155 39539
rect 73189 39536 73201 39539
rect 73416 39536 73422 39548
rect 73189 39508 73422 39536
rect 73189 39505 73201 39508
rect 73143 39499 73201 39505
rect 73416 39496 73422 39508
rect 73474 39496 73480 39548
rect 77188 39536 77194 39548
rect 73526 39508 77194 39536
rect 73526 39468 73554 39508
rect 77188 39496 77194 39508
rect 77246 39496 77252 39548
rect 77390 39545 77418 39576
rect 77464 39564 77470 39576
rect 77522 39564 77528 39616
rect 78310 39604 78338 39644
rect 79396 39632 79402 39684
rect 79454 39672 79460 39684
rect 84180 39672 84186 39684
rect 79454 39644 83858 39672
rect 84141 39644 84186 39672
rect 79454 39632 79460 39644
rect 83720 39604 83726 39616
rect 78310 39576 83726 39604
rect 83720 39564 83726 39576
rect 83778 39564 83784 39616
rect 83830 39604 83858 39644
rect 84180 39632 84186 39644
rect 84238 39632 84244 39684
rect 88504 39632 88510 39684
rect 88562 39672 88568 39684
rect 88783 39675 88841 39681
rect 88783 39672 88795 39675
rect 88562 39644 88795 39672
rect 88562 39632 88568 39644
rect 88783 39641 88795 39644
rect 88829 39641 88841 39675
rect 88783 39635 88841 39641
rect 88228 39604 88234 39616
rect 83830 39576 88234 39604
rect 88228 39564 88234 39576
rect 88286 39564 88292 39616
rect 88320 39564 88326 39616
rect 88378 39604 88384 39616
rect 90160 39604 90166 39616
rect 88378 39576 90166 39604
rect 88378 39564 88384 39576
rect 90160 39564 90166 39576
rect 90218 39564 90224 39616
rect 77375 39539 77433 39545
rect 77375 39505 77387 39539
rect 77421 39505 77433 39539
rect 77648 39536 77654 39548
rect 77609 39508 77654 39536
rect 77375 39499 77433 39505
rect 77648 39496 77654 39508
rect 77706 39496 77712 39548
rect 82064 39496 82070 39548
rect 82122 39536 82128 39548
rect 83904 39536 83910 39548
rect 82122 39508 83910 39536
rect 82122 39496 82128 39508
rect 83904 39496 83910 39508
rect 83962 39496 83968 39548
rect 84456 39536 84462 39548
rect 84417 39508 84462 39536
rect 84456 39496 84462 39508
rect 84514 39496 84520 39548
rect 88688 39536 88694 39548
rect 88649 39508 88694 39536
rect 88688 39496 88694 39508
rect 88746 39496 88752 39548
rect 89151 39539 89209 39545
rect 89151 39505 89163 39539
rect 89197 39505 89209 39539
rect 89151 39499 89209 39505
rect 72974 39440 73554 39468
rect 77556 39428 77562 39480
rect 77614 39468 77620 39480
rect 88136 39468 88142 39480
rect 77614 39440 88142 39468
rect 77614 39428 77620 39440
rect 88136 39428 88142 39440
rect 88194 39428 88200 39480
rect 88596 39428 88602 39480
rect 88654 39468 88660 39480
rect 89166 39468 89194 39499
rect 88654 39440 89194 39468
rect 88654 39428 88660 39440
rect 79212 39400 79218 39412
rect 71073 39372 71162 39400
rect 78310 39372 79218 39400
rect 71073 39369 71085 39372
rect 71027 39363 71085 39369
rect 62744 39332 62750 39344
rect 57058 39304 62750 39332
rect 62744 39292 62750 39304
rect 62802 39292 62808 39344
rect 66792 39332 66798 39344
rect 66753 39304 66798 39332
rect 66792 39292 66798 39304
rect 66850 39292 66856 39344
rect 67988 39292 67994 39344
rect 68046 39332 68052 39344
rect 69920 39332 69926 39344
rect 68046 39304 69926 39332
rect 68046 39292 68052 39304
rect 69920 39292 69926 39304
rect 69978 39292 69984 39344
rect 71300 39292 71306 39344
rect 71358 39332 71364 39344
rect 78310 39332 78338 39372
rect 79212 39360 79218 39372
rect 79270 39360 79276 39412
rect 71358 39304 78338 39332
rect 78939 39335 78997 39341
rect 71358 39292 71364 39304
rect 78939 39301 78951 39335
rect 78985 39332 78997 39335
rect 79856 39332 79862 39344
rect 78985 39304 79862 39332
rect 78985 39301 78997 39304
rect 78939 39295 78997 39301
rect 79856 39292 79862 39304
rect 79914 39292 79920 39344
rect 538 39242 93642 39264
rect 538 39190 3680 39242
rect 3732 39190 3744 39242
rect 3796 39190 3808 39242
rect 3860 39190 3872 39242
rect 3924 39190 9008 39242
rect 9060 39190 9072 39242
rect 9124 39190 9136 39242
rect 9188 39190 9200 39242
rect 9252 39190 14336 39242
rect 14388 39190 14400 39242
rect 14452 39190 14464 39242
rect 14516 39190 14528 39242
rect 14580 39190 19664 39242
rect 19716 39190 19728 39242
rect 19780 39190 19792 39242
rect 19844 39190 19856 39242
rect 19908 39190 24992 39242
rect 25044 39190 25056 39242
rect 25108 39190 25120 39242
rect 25172 39190 25184 39242
rect 25236 39190 30320 39242
rect 30372 39190 30384 39242
rect 30436 39190 30448 39242
rect 30500 39190 30512 39242
rect 30564 39190 35648 39242
rect 35700 39190 35712 39242
rect 35764 39190 35776 39242
rect 35828 39190 35840 39242
rect 35892 39190 40976 39242
rect 41028 39190 41040 39242
rect 41092 39190 41104 39242
rect 41156 39190 41168 39242
rect 41220 39190 46304 39242
rect 46356 39190 46368 39242
rect 46420 39190 46432 39242
rect 46484 39190 46496 39242
rect 46548 39190 51632 39242
rect 51684 39190 51696 39242
rect 51748 39190 51760 39242
rect 51812 39190 51824 39242
rect 51876 39190 56960 39242
rect 57012 39190 57024 39242
rect 57076 39190 57088 39242
rect 57140 39190 57152 39242
rect 57204 39190 62288 39242
rect 62340 39190 62352 39242
rect 62404 39190 62416 39242
rect 62468 39190 62480 39242
rect 62532 39190 67616 39242
rect 67668 39190 67680 39242
rect 67732 39190 67744 39242
rect 67796 39190 67808 39242
rect 67860 39190 72944 39242
rect 72996 39190 73008 39242
rect 73060 39190 73072 39242
rect 73124 39190 73136 39242
rect 73188 39190 78272 39242
rect 78324 39190 78336 39242
rect 78388 39190 78400 39242
rect 78452 39190 78464 39242
rect 78516 39190 83600 39242
rect 83652 39190 83664 39242
rect 83716 39190 83728 39242
rect 83780 39190 83792 39242
rect 83844 39190 88928 39242
rect 88980 39190 88992 39242
rect 89044 39190 89056 39242
rect 89108 39190 89120 39242
rect 89172 39190 93642 39242
rect 538 39168 93642 39190
rect 19044 39088 19050 39140
rect 19102 39128 19108 39140
rect 19139 39131 19197 39137
rect 19139 39128 19151 39131
rect 19102 39100 19151 39128
rect 19102 39088 19108 39100
rect 19139 39097 19151 39100
rect 19185 39097 19197 39131
rect 19139 39091 19197 39097
rect 20427 39131 20485 39137
rect 20427 39097 20439 39131
rect 20473 39128 20485 39131
rect 21068 39128 21074 39140
rect 20473 39100 21074 39128
rect 20473 39097 20485 39100
rect 20427 39091 20485 39097
rect 18768 39020 18774 39072
rect 18826 39060 18832 39072
rect 20442 39060 20470 39091
rect 21068 39088 21074 39100
rect 21126 39088 21132 39140
rect 26867 39131 26925 39137
rect 26867 39097 26879 39131
rect 26913 39128 26925 39131
rect 27416 39128 27422 39140
rect 26913 39100 27422 39128
rect 26913 39097 26925 39100
rect 26867 39091 26925 39097
rect 27416 39088 27422 39100
rect 27474 39088 27480 39140
rect 32016 39088 32022 39140
rect 32074 39128 32080 39140
rect 32111 39131 32169 39137
rect 32111 39128 32123 39131
rect 32074 39100 32123 39128
rect 32074 39088 32080 39100
rect 32111 39097 32123 39100
rect 32157 39097 32169 39131
rect 34684 39128 34690 39140
rect 34645 39100 34690 39128
rect 32111 39091 32169 39097
rect 34684 39088 34690 39100
rect 34742 39088 34748 39140
rect 41768 39088 41774 39140
rect 41826 39128 41832 39140
rect 42139 39131 42197 39137
rect 42139 39128 42151 39131
rect 41826 39100 42151 39128
rect 41826 39088 41832 39100
rect 42139 39097 42151 39100
rect 42185 39128 42197 39131
rect 44804 39128 44810 39140
rect 42185 39100 44810 39128
rect 42185 39097 42197 39100
rect 42139 39091 42197 39097
rect 44804 39088 44810 39100
rect 44862 39088 44868 39140
rect 50324 39128 50330 39140
rect 47674 39100 50330 39128
rect 18826 39032 20470 39060
rect 33215 39063 33273 39069
rect 18826 39020 18832 39032
rect 33215 39029 33227 39063
rect 33261 39060 33273 39063
rect 34868 39060 34874 39072
rect 33261 39032 34874 39060
rect 33261 39029 33273 39032
rect 33215 39023 33273 39029
rect 2484 38992 2490 39004
rect 2397 38964 2490 38992
rect 2484 38952 2490 38964
rect 2542 38992 2548 39004
rect 3496 38992 3502 39004
rect 2542 38964 3502 38992
rect 2542 38952 2548 38964
rect 3496 38952 3502 38964
rect 3554 38952 3560 39004
rect 8004 38952 8010 39004
rect 8062 38992 8068 39004
rect 8559 38995 8617 39001
rect 8559 38992 8571 38995
rect 8062 38964 8571 38992
rect 8062 38952 8068 38964
rect 8559 38961 8571 38964
rect 8605 38961 8617 38995
rect 8559 38955 8617 38961
rect 8648 38952 8654 39004
rect 8706 38992 8712 39004
rect 9019 38995 9077 39001
rect 9019 38992 9031 38995
rect 8706 38964 9031 38992
rect 8706 38952 8712 38964
rect 9019 38961 9031 38964
rect 9065 38961 9077 38995
rect 12236 38992 12242 39004
rect 12197 38964 12242 38992
rect 9019 38955 9077 38961
rect 12236 38952 12242 38964
rect 12294 38952 12300 39004
rect 16563 38995 16621 39001
rect 16563 38961 16575 38995
rect 16609 38992 16621 38995
rect 17480 38992 17486 39004
rect 16609 38964 17486 38992
rect 16609 38961 16621 38964
rect 16563 38955 16621 38961
rect 17480 38952 17486 38964
rect 17538 38952 17544 39004
rect 2208 38884 2214 38936
rect 2266 38924 2272 38936
rect 3404 38924 3410 38936
rect 2266 38896 3410 38924
rect 2266 38884 2272 38896
rect 3404 38884 3410 38896
rect 3462 38884 3468 38936
rect 8743 38927 8801 38933
rect 8743 38893 8755 38927
rect 8789 38893 8801 38927
rect 9108 38924 9114 38936
rect 9069 38896 9114 38924
rect 8743 38887 8801 38893
rect 3867 38859 3925 38865
rect 3867 38825 3879 38859
rect 3913 38856 3925 38859
rect 4324 38856 4330 38868
rect 3913 38828 4330 38856
rect 3913 38825 3925 38828
rect 3867 38819 3925 38825
rect 4324 38816 4330 38828
rect 4382 38816 4388 38868
rect 8096 38856 8102 38868
rect 8057 38828 8102 38856
rect 8096 38816 8102 38828
rect 8154 38816 8160 38868
rect 8758 38856 8786 38887
rect 9108 38884 9114 38896
rect 9166 38884 9172 38936
rect 11963 38927 12021 38933
rect 11963 38893 11975 38927
rect 12009 38893 12021 38927
rect 13616 38924 13622 38936
rect 13529 38896 13622 38924
rect 11963 38887 12021 38893
rect 9752 38856 9758 38868
rect 8758 38828 9758 38856
rect 9752 38816 9758 38828
rect 9810 38816 9816 38868
rect 3404 38748 3410 38800
rect 3462 38788 3468 38800
rect 4048 38788 4054 38800
rect 3462 38760 4054 38788
rect 3462 38748 3468 38760
rect 4048 38748 4054 38760
rect 4106 38748 4112 38800
rect 8007 38791 8065 38797
rect 8007 38757 8019 38791
rect 8053 38788 8065 38791
rect 9108 38788 9114 38800
rect 8053 38760 9114 38788
rect 8053 38757 8065 38760
rect 8007 38751 8065 38757
rect 9108 38748 9114 38760
rect 9166 38788 9172 38800
rect 9476 38788 9482 38800
rect 9166 38760 9482 38788
rect 9166 38748 9172 38760
rect 9476 38748 9482 38760
rect 9534 38748 9540 38800
rect 11978 38788 12006 38887
rect 13616 38884 13622 38896
rect 13674 38924 13680 38936
rect 18786 38933 18814 39020
rect 32571 38995 32629 39001
rect 32571 38961 32583 38995
rect 32617 38992 32629 38995
rect 32617 38964 32982 38992
rect 32617 38961 32629 38964
rect 32571 38955 32629 38961
rect 16195 38927 16253 38933
rect 16195 38924 16207 38927
rect 13674 38896 16207 38924
rect 13674 38884 13680 38896
rect 16195 38893 16207 38896
rect 16241 38893 16253 38927
rect 16195 38887 16253 38893
rect 18771 38927 18829 38933
rect 18771 38893 18783 38927
rect 18817 38893 18829 38927
rect 18771 38887 18829 38893
rect 18955 38927 19013 38933
rect 18955 38893 18967 38927
rect 19001 38924 19013 38927
rect 19044 38924 19050 38936
rect 19001 38896 19050 38924
rect 19001 38893 19013 38896
rect 18955 38887 19013 38893
rect 19044 38884 19050 38896
rect 19102 38924 19108 38936
rect 19507 38927 19565 38933
rect 19507 38924 19519 38927
rect 19102 38896 19519 38924
rect 19102 38884 19108 38896
rect 19507 38893 19519 38896
rect 19553 38893 19565 38927
rect 20240 38924 20246 38936
rect 20201 38896 20246 38924
rect 19507 38887 19565 38893
rect 20240 38884 20246 38896
rect 20298 38884 20304 38936
rect 25668 38884 25674 38936
rect 25726 38924 25732 38936
rect 27051 38927 27109 38933
rect 27051 38924 27063 38927
rect 25726 38896 27063 38924
rect 25726 38884 25732 38896
rect 27051 38893 27063 38896
rect 27097 38893 27109 38927
rect 27051 38887 27109 38893
rect 27235 38927 27293 38933
rect 27235 38893 27247 38927
rect 27281 38924 27293 38927
rect 27416 38924 27422 38936
rect 27281 38896 27422 38924
rect 27281 38893 27293 38896
rect 27235 38887 27293 38893
rect 27416 38884 27422 38896
rect 27474 38884 27480 38936
rect 27508 38884 27514 38936
rect 27566 38924 27572 38936
rect 27603 38927 27661 38933
rect 27603 38924 27615 38927
rect 27566 38896 27615 38924
rect 27566 38884 27572 38896
rect 27603 38893 27615 38896
rect 27649 38893 27661 38927
rect 27603 38887 27661 38893
rect 27787 38927 27845 38933
rect 27787 38893 27799 38927
rect 27833 38924 27845 38927
rect 27968 38924 27974 38936
rect 27833 38896 27974 38924
rect 27833 38893 27845 38896
rect 27787 38887 27845 38893
rect 27968 38884 27974 38896
rect 28026 38884 28032 38936
rect 32479 38927 32537 38933
rect 32479 38893 32491 38927
rect 32525 38893 32537 38927
rect 32479 38887 32537 38893
rect 16008 38856 16014 38868
rect 15969 38828 16014 38856
rect 16008 38816 16014 38828
rect 16066 38816 16072 38868
rect 16744 38816 16750 38868
rect 16802 38856 16808 38868
rect 18863 38859 18921 38865
rect 18863 38856 18875 38859
rect 16802 38828 18875 38856
rect 16802 38816 16808 38828
rect 18863 38825 18875 38828
rect 18909 38825 18921 38859
rect 27434 38856 27462 38884
rect 32494 38856 32522 38887
rect 32752 38884 32758 38936
rect 32810 38924 32816 38936
rect 32847 38927 32905 38933
rect 32847 38924 32859 38927
rect 32810 38896 32859 38924
rect 32810 38884 32816 38896
rect 32847 38893 32859 38896
rect 32893 38893 32905 38927
rect 32847 38887 32905 38893
rect 32660 38856 32666 38868
rect 27434 38828 32666 38856
rect 18863 38819 18921 38825
rect 32660 38816 32666 38828
rect 32718 38816 32724 38868
rect 32954 38856 32982 38964
rect 33031 38927 33089 38933
rect 33031 38893 33043 38927
rect 33077 38924 33089 38927
rect 33230 38924 33258 39023
rect 34868 39020 34874 39032
rect 34926 39020 34932 39072
rect 39468 39020 39474 39072
rect 39526 39060 39532 39072
rect 47196 39060 47202 39072
rect 39526 39032 47202 39060
rect 39526 39020 39532 39032
rect 47196 39020 47202 39032
rect 47254 39060 47260 39072
rect 47674 39060 47702 39100
rect 50324 39088 50330 39100
rect 50382 39088 50388 39140
rect 50508 39088 50514 39140
rect 50566 39128 50572 39140
rect 50879 39131 50937 39137
rect 50879 39128 50891 39131
rect 50566 39100 50891 39128
rect 50566 39088 50572 39100
rect 50879 39097 50891 39100
rect 50925 39128 50937 39131
rect 52164 39128 52170 39140
rect 50925 39100 52170 39128
rect 50925 39097 50937 39100
rect 50879 39091 50937 39097
rect 52164 39088 52170 39100
rect 52222 39128 52228 39140
rect 54099 39131 54157 39137
rect 54099 39128 54111 39131
rect 52222 39100 54111 39128
rect 52222 39088 52228 39100
rect 54099 39097 54111 39100
rect 54145 39128 54157 39131
rect 54188 39128 54194 39140
rect 54145 39100 54194 39128
rect 54145 39097 54157 39100
rect 54099 39091 54157 39097
rect 54188 39088 54194 39100
rect 54246 39088 54252 39140
rect 55108 39088 55114 39140
rect 55166 39128 55172 39140
rect 55844 39128 55850 39140
rect 55166 39100 55850 39128
rect 55166 39088 55172 39100
rect 55844 39088 55850 39100
rect 55902 39088 55908 39140
rect 65323 39131 65381 39137
rect 65323 39097 65335 39131
rect 65369 39128 65381 39131
rect 65504 39128 65510 39140
rect 65369 39100 65510 39128
rect 65369 39097 65381 39100
rect 65323 39091 65381 39097
rect 65504 39088 65510 39100
rect 65562 39088 65568 39140
rect 68264 39128 68270 39140
rect 68225 39100 68270 39128
rect 68264 39088 68270 39100
rect 68322 39088 68328 39140
rect 74060 39128 74066 39140
rect 74021 39100 74066 39128
rect 74060 39088 74066 39100
rect 74118 39088 74124 39140
rect 75440 39088 75446 39140
rect 75498 39128 75504 39140
rect 75995 39131 76053 39137
rect 75995 39128 76007 39131
rect 75498 39100 76007 39128
rect 75498 39088 75504 39100
rect 75995 39097 76007 39100
rect 76041 39097 76053 39131
rect 90160 39128 90166 39140
rect 90121 39100 90166 39128
rect 75995 39091 76053 39097
rect 47254 39032 47702 39060
rect 54206 39060 54234 39088
rect 55384 39060 55390 39072
rect 54206 39032 55390 39060
rect 47254 39020 47260 39032
rect 34500 38952 34506 39004
rect 34558 38992 34564 39004
rect 35147 38995 35205 39001
rect 35147 38992 35159 38995
rect 34558 38964 35159 38992
rect 34558 38952 34564 38964
rect 35147 38961 35159 38964
rect 35193 38961 35205 38995
rect 35147 38955 35205 38961
rect 40848 38952 40854 39004
rect 40906 38992 40912 39004
rect 41308 38992 41314 39004
rect 40906 38964 40951 38992
rect 41269 38964 41314 38992
rect 40906 38952 40912 38964
rect 41308 38952 41314 38964
rect 41366 38952 41372 39004
rect 43056 38992 43062 39004
rect 43017 38964 43062 38992
rect 43056 38952 43062 38964
rect 43114 38952 43120 39004
rect 45635 38995 45693 39001
rect 45635 38992 45647 38995
rect 43166 38964 43378 38992
rect 43166 38936 43194 38964
rect 33077 38896 33258 38924
rect 33077 38893 33089 38896
rect 33031 38887 33089 38893
rect 34684 38884 34690 38936
rect 34742 38924 34748 38936
rect 34871 38927 34929 38933
rect 34871 38924 34883 38927
rect 34742 38896 34883 38924
rect 34742 38884 34748 38896
rect 34871 38893 34883 38896
rect 34917 38893 34929 38927
rect 34871 38887 34929 38893
rect 41403 38927 41461 38933
rect 41403 38893 41415 38927
rect 41449 38893 41461 38927
rect 41768 38924 41774 38936
rect 41729 38896 41774 38924
rect 41403 38887 41461 38893
rect 36527 38859 36585 38865
rect 32954 38828 33442 38856
rect 33414 38800 33442 38828
rect 36527 38825 36539 38859
rect 36573 38856 36585 38859
rect 41308 38856 41314 38868
rect 36573 38828 41314 38856
rect 36573 38825 36585 38828
rect 36527 38819 36585 38825
rect 41308 38816 41314 38828
rect 41366 38816 41372 38868
rect 13803 38791 13861 38797
rect 13803 38788 13815 38791
rect 11978 38760 13815 38788
rect 13803 38757 13815 38760
rect 13849 38788 13861 38791
rect 14076 38788 14082 38800
rect 13849 38760 14082 38788
rect 13849 38757 13861 38760
rect 13803 38751 13861 38757
rect 14076 38748 14082 38760
rect 14134 38748 14140 38800
rect 33396 38788 33402 38800
rect 33357 38760 33402 38788
rect 33396 38748 33402 38760
rect 33454 38748 33460 38800
rect 41418 38788 41446 38887
rect 41768 38884 41774 38896
rect 41826 38884 41832 38936
rect 41955 38927 42013 38933
rect 41955 38893 41967 38927
rect 42001 38893 42013 38927
rect 43148 38924 43154 38936
rect 43109 38896 43154 38924
rect 41955 38887 42013 38893
rect 41970 38856 41998 38887
rect 43148 38884 43154 38896
rect 43206 38884 43212 38936
rect 43350 38924 43378 38964
rect 44086 38964 45647 38992
rect 43703 38927 43761 38933
rect 43703 38924 43715 38927
rect 43350 38896 43715 38924
rect 43703 38893 43715 38896
rect 43749 38893 43761 38927
rect 43703 38887 43761 38893
rect 43887 38927 43945 38933
rect 43887 38893 43899 38927
rect 43933 38924 43945 38927
rect 44086 38924 44114 38964
rect 45635 38961 45647 38964
rect 45681 38961 45693 38995
rect 45635 38955 45693 38961
rect 47472 38952 47478 39004
rect 47530 38992 47536 39004
rect 48119 38995 48177 39001
rect 48119 38992 48131 38995
rect 47530 38964 48131 38992
rect 47530 38952 47536 38964
rect 48119 38961 48131 38964
rect 48165 38961 48177 38995
rect 51152 38992 51158 39004
rect 51113 38964 51158 38992
rect 48119 38955 48177 38961
rect 51152 38952 51158 38964
rect 51210 38952 51216 39004
rect 53912 38992 53918 39004
rect 51538 38964 53918 38992
rect 43933 38896 44114 38924
rect 45543 38927 45601 38933
rect 43933 38893 43945 38896
rect 43887 38887 43945 38893
rect 45543 38893 45555 38927
rect 45589 38924 45601 38927
rect 45911 38927 45969 38933
rect 45911 38924 45923 38927
rect 45589 38896 45923 38924
rect 45589 38893 45601 38896
rect 45543 38887 45601 38893
rect 45911 38893 45923 38896
rect 45957 38924 45969 38927
rect 46000 38924 46006 38936
rect 45957 38896 46006 38924
rect 45957 38893 45969 38896
rect 45911 38887 45969 38893
rect 43902 38856 43930 38887
rect 46000 38884 46006 38896
rect 46058 38884 46064 38936
rect 47288 38924 47294 38936
rect 47249 38896 47294 38924
rect 47288 38884 47294 38896
rect 47346 38884 47352 38936
rect 48024 38924 48030 38936
rect 47985 38896 48030 38924
rect 48024 38884 48030 38896
rect 48082 38884 48088 38936
rect 50416 38924 50422 38936
rect 50342 38896 50422 38924
rect 41970 38828 43930 38856
rect 44255 38859 44313 38865
rect 44255 38825 44267 38859
rect 44301 38856 44313 38859
rect 44712 38856 44718 38868
rect 44301 38828 44718 38856
rect 44301 38825 44313 38828
rect 44255 38819 44313 38825
rect 44712 38816 44718 38828
rect 44770 38816 44776 38868
rect 44804 38816 44810 38868
rect 44862 38856 44868 38868
rect 50342 38856 50370 38896
rect 50416 38884 50422 38896
rect 50474 38884 50480 38936
rect 51538 38924 51566 38964
rect 50710 38896 51566 38924
rect 51615 38927 51673 38933
rect 44862 38828 50370 38856
rect 44862 38816 44868 38828
rect 42320 38788 42326 38800
rect 41418 38760 42326 38788
rect 42320 38748 42326 38760
rect 42378 38748 42384 38800
rect 47380 38748 47386 38800
rect 47438 38788 47444 38800
rect 47438 38760 47483 38788
rect 47438 38748 47444 38760
rect 47564 38748 47570 38800
rect 47622 38788 47628 38800
rect 50710 38797 50738 38896
rect 51615 38893 51627 38927
rect 51661 38924 51673 38927
rect 51704 38924 51710 38936
rect 51661 38896 51710 38924
rect 51661 38893 51673 38896
rect 51615 38887 51673 38893
rect 51704 38884 51710 38896
rect 51762 38884 51768 38936
rect 51814 38933 51842 38964
rect 53912 38952 53918 38964
rect 53970 38992 53976 39004
rect 55019 38995 55077 39001
rect 53970 38964 54970 38992
rect 53970 38952 53976 38964
rect 51799 38927 51857 38933
rect 51799 38893 51811 38927
rect 51845 38893 51857 38927
rect 52164 38924 52170 38936
rect 52125 38896 52170 38924
rect 51799 38887 51857 38893
rect 52164 38884 52170 38896
rect 52222 38884 52228 38936
rect 52256 38884 52262 38936
rect 52314 38924 52320 38936
rect 54942 38933 54970 38964
rect 55019 38961 55031 38995
rect 55065 38992 55077 38995
rect 55108 38992 55114 39004
rect 55065 38964 55114 38992
rect 55065 38961 55077 38964
rect 55019 38955 55077 38961
rect 55108 38952 55114 38964
rect 55166 38952 55172 39004
rect 54927 38927 54985 38933
rect 52314 38896 52359 38924
rect 52314 38884 52320 38896
rect 54927 38893 54939 38927
rect 54973 38893 54985 38927
rect 55218 38924 55246 39032
rect 55384 39020 55390 39032
rect 55442 39020 55448 39072
rect 55476 39020 55482 39072
rect 55534 39060 55540 39072
rect 70840 39060 70846 39072
rect 55534 39032 70846 39060
rect 55534 39020 55540 39032
rect 70840 39020 70846 39032
rect 70898 39020 70904 39072
rect 59984 38992 59990 39004
rect 55494 38964 59990 38992
rect 55494 38933 55522 38964
rect 59984 38952 59990 38964
rect 60042 38952 60048 39004
rect 63020 38952 63026 39004
rect 63078 38992 63084 39004
rect 73968 38992 73974 39004
rect 63078 38964 64538 38992
rect 63078 38952 63084 38964
rect 55295 38927 55353 38933
rect 55295 38924 55307 38927
rect 55218 38896 55307 38924
rect 54927 38887 54985 38893
rect 55295 38893 55307 38896
rect 55341 38893 55353 38927
rect 55295 38887 55353 38893
rect 55479 38927 55537 38933
rect 55479 38893 55491 38927
rect 55525 38893 55537 38927
rect 55479 38887 55537 38893
rect 60263 38927 60321 38933
rect 60263 38893 60275 38927
rect 60309 38924 60321 38927
rect 60352 38924 60358 38936
rect 60309 38896 60358 38924
rect 60309 38893 60321 38896
rect 60263 38887 60321 38893
rect 60352 38884 60358 38896
rect 60410 38924 60416 38936
rect 61364 38924 61370 38936
rect 60410 38896 61370 38924
rect 60410 38884 60416 38896
rect 61364 38884 61370 38896
rect 61422 38884 61428 38936
rect 62928 38884 62934 38936
rect 62986 38924 62992 38936
rect 64124 38924 64130 38936
rect 62986 38896 64130 38924
rect 62986 38884 62992 38896
rect 64124 38884 64130 38896
rect 64182 38884 64188 38936
rect 64311 38927 64369 38933
rect 64311 38893 64323 38927
rect 64357 38893 64369 38927
rect 64510 38924 64538 38964
rect 65246 38964 73974 38992
rect 64768 38924 64774 38936
rect 64510 38896 64774 38924
rect 64311 38887 64369 38893
rect 50784 38816 50790 38868
rect 50842 38856 50848 38868
rect 54283 38859 54341 38865
rect 54283 38856 54295 38859
rect 50842 38828 54295 38856
rect 50842 38816 50848 38828
rect 54283 38825 54295 38828
rect 54329 38825 54341 38859
rect 54283 38819 54341 38825
rect 63664 38816 63670 38868
rect 63722 38856 63728 38868
rect 63851 38859 63909 38865
rect 63851 38856 63863 38859
rect 63722 38828 63863 38856
rect 63722 38816 63728 38828
rect 63851 38825 63863 38828
rect 63897 38856 63909 38859
rect 64035 38859 64093 38865
rect 64035 38856 64047 38859
rect 63897 38828 64047 38856
rect 63897 38825 63909 38828
rect 63851 38819 63909 38825
rect 64035 38825 64047 38828
rect 64081 38856 64093 38859
rect 64326 38856 64354 38887
rect 64768 38884 64774 38896
rect 64826 38884 64832 38936
rect 64863 38927 64921 38933
rect 64863 38893 64875 38927
rect 64909 38924 64921 38927
rect 65246 38924 65274 38964
rect 73968 38952 73974 38964
rect 74026 38992 74032 39004
rect 74152 38992 74158 39004
rect 74026 38964 74158 38992
rect 74026 38952 74032 38964
rect 74152 38952 74158 38964
rect 74210 38952 74216 39004
rect 74523 38995 74581 39001
rect 74523 38961 74535 38995
rect 74569 38992 74581 38995
rect 76010 38992 76038 39091
rect 90160 39088 90166 39100
rect 90218 39088 90224 39140
rect 76179 38995 76237 39001
rect 76179 38992 76191 38995
rect 74569 38964 75302 38992
rect 76010 38964 76191 38992
rect 74569 38961 74581 38964
rect 74523 38955 74581 38961
rect 66792 38924 66798 38936
rect 64909 38896 65274 38924
rect 66753 38896 66798 38924
rect 64909 38893 64921 38896
rect 64863 38887 64921 38893
rect 64878 38856 64906 38887
rect 66792 38884 66798 38896
rect 66850 38884 66856 38936
rect 68451 38927 68509 38933
rect 68451 38924 68463 38927
rect 66902 38896 68463 38924
rect 64081 38828 64906 38856
rect 64081 38825 64093 38828
rect 64035 38819 64093 38825
rect 50695 38791 50753 38797
rect 50695 38788 50707 38791
rect 47622 38760 50707 38788
rect 47622 38748 47628 38760
rect 50695 38757 50707 38760
rect 50741 38757 50753 38791
rect 50695 38751 50753 38757
rect 60260 38748 60266 38800
rect 60318 38788 60324 38800
rect 60539 38791 60597 38797
rect 60539 38788 60551 38791
rect 60318 38760 60551 38788
rect 60318 38748 60324 38760
rect 60539 38757 60551 38760
rect 60585 38757 60597 38791
rect 60539 38751 60597 38757
rect 64768 38748 64774 38800
rect 64826 38788 64832 38800
rect 66902 38797 66930 38896
rect 68451 38893 68463 38896
rect 68497 38893 68509 38927
rect 68632 38924 68638 38936
rect 68593 38896 68638 38924
rect 68451 38887 68509 38893
rect 68632 38884 68638 38896
rect 68690 38884 68696 38936
rect 69000 38924 69006 38936
rect 68961 38896 69006 38924
rect 69000 38884 69006 38896
rect 69058 38884 69064 38936
rect 69095 38927 69153 38933
rect 69095 38893 69107 38927
rect 69141 38893 69153 38927
rect 69095 38887 69153 38893
rect 66887 38791 66945 38797
rect 66887 38788 66899 38791
rect 64826 38760 66899 38788
rect 64826 38748 64832 38760
rect 66887 38757 66899 38760
rect 66933 38757 66945 38791
rect 66887 38751 66945 38757
rect 68356 38748 68362 38800
rect 68414 38788 68420 38800
rect 69110 38788 69138 38887
rect 73692 38884 73698 38936
rect 73750 38924 73756 38936
rect 74431 38927 74489 38933
rect 74431 38924 74443 38927
rect 73750 38896 74443 38924
rect 73750 38884 73756 38896
rect 74431 38893 74443 38896
rect 74477 38893 74489 38927
rect 74431 38887 74489 38893
rect 74799 38927 74857 38933
rect 74799 38893 74811 38927
rect 74845 38893 74857 38927
rect 74799 38887 74857 38893
rect 74983 38927 75041 38933
rect 74983 38893 74995 38927
rect 75029 38893 75041 38927
rect 75274 38924 75302 38964
rect 76179 38961 76191 38964
rect 76225 38961 76237 38995
rect 76179 38955 76237 38961
rect 77467 38995 77525 39001
rect 77467 38961 77479 38995
rect 77513 38992 77525 38995
rect 79491 38995 79549 39001
rect 79491 38992 79503 38995
rect 77513 38964 79503 38992
rect 77513 38961 77525 38964
rect 77467 38955 77525 38961
rect 79491 38961 79503 38964
rect 79537 38961 79549 38995
rect 79491 38955 79549 38961
rect 90160 38952 90166 39004
rect 90218 38992 90224 39004
rect 90439 38995 90497 39001
rect 90439 38992 90451 38995
rect 90218 38964 90451 38992
rect 90218 38952 90224 38964
rect 90439 38961 90451 38964
rect 90485 38961 90497 38995
rect 90439 38955 90497 38961
rect 76268 38924 76274 38936
rect 75274 38896 76274 38924
rect 74983 38887 75041 38893
rect 73784 38816 73790 38868
rect 73842 38856 73848 38868
rect 74814 38856 74842 38887
rect 73842 38828 74842 38856
rect 74998 38856 75026 38887
rect 76268 38884 76274 38896
rect 76326 38884 76332 38936
rect 76363 38927 76421 38933
rect 76363 38893 76375 38927
rect 76409 38924 76421 38927
rect 76452 38924 76458 38936
rect 76409 38896 76458 38924
rect 76409 38893 76421 38896
rect 76363 38887 76421 38893
rect 76452 38884 76458 38896
rect 76510 38924 76516 38936
rect 76915 38927 76973 38933
rect 76915 38924 76927 38927
rect 76510 38896 76927 38924
rect 76510 38884 76516 38896
rect 76915 38893 76927 38896
rect 76961 38893 76973 38927
rect 77096 38924 77102 38936
rect 77057 38896 77102 38924
rect 76915 38887 76973 38893
rect 77096 38884 77102 38896
rect 77154 38884 77160 38936
rect 79215 38927 79273 38933
rect 79215 38924 79227 38927
rect 78954 38896 79227 38924
rect 77114 38856 77142 38884
rect 74998 38828 77142 38856
rect 73842 38816 73848 38828
rect 69279 38791 69337 38797
rect 69279 38788 69291 38791
rect 68414 38760 69291 38788
rect 68414 38748 68420 38760
rect 69279 38757 69291 38760
rect 69325 38757 69337 38791
rect 69279 38751 69337 38757
rect 77464 38748 77470 38800
rect 77522 38788 77528 38800
rect 78954 38797 78982 38896
rect 79215 38893 79227 38896
rect 79261 38893 79273 38927
rect 90712 38924 90718 38936
rect 90673 38896 90718 38924
rect 79215 38887 79273 38893
rect 90712 38884 90718 38896
rect 90770 38884 90776 38936
rect 78939 38791 78997 38797
rect 78939 38788 78951 38791
rect 77522 38760 78951 38788
rect 77522 38748 77528 38760
rect 78939 38757 78951 38760
rect 78985 38757 78997 38791
rect 78939 38751 78997 38757
rect 80408 38748 80414 38800
rect 80466 38788 80472 38800
rect 80595 38791 80653 38797
rect 80595 38788 80607 38791
rect 80466 38760 80607 38788
rect 80466 38748 80472 38760
rect 80595 38757 80607 38760
rect 80641 38757 80653 38791
rect 80595 38751 80653 38757
rect 91448 38748 91454 38800
rect 91506 38788 91512 38800
rect 91819 38791 91877 38797
rect 91819 38788 91831 38791
rect 91506 38760 91831 38788
rect 91506 38748 91512 38760
rect 91819 38757 91831 38760
rect 91865 38757 91877 38791
rect 91819 38751 91877 38757
rect 538 38698 93642 38720
rect 538 38646 6344 38698
rect 6396 38646 6408 38698
rect 6460 38646 6472 38698
rect 6524 38646 6536 38698
rect 6588 38646 11672 38698
rect 11724 38646 11736 38698
rect 11788 38646 11800 38698
rect 11852 38646 11864 38698
rect 11916 38646 17000 38698
rect 17052 38646 17064 38698
rect 17116 38646 17128 38698
rect 17180 38646 17192 38698
rect 17244 38646 22328 38698
rect 22380 38646 22392 38698
rect 22444 38646 22456 38698
rect 22508 38646 22520 38698
rect 22572 38646 27656 38698
rect 27708 38646 27720 38698
rect 27772 38646 27784 38698
rect 27836 38646 27848 38698
rect 27900 38646 32984 38698
rect 33036 38646 33048 38698
rect 33100 38646 33112 38698
rect 33164 38646 33176 38698
rect 33228 38646 38312 38698
rect 38364 38646 38376 38698
rect 38428 38646 38440 38698
rect 38492 38646 38504 38698
rect 38556 38646 43640 38698
rect 43692 38646 43704 38698
rect 43756 38646 43768 38698
rect 43820 38646 43832 38698
rect 43884 38646 48968 38698
rect 49020 38646 49032 38698
rect 49084 38646 49096 38698
rect 49148 38646 49160 38698
rect 49212 38646 54296 38698
rect 54348 38646 54360 38698
rect 54412 38646 54424 38698
rect 54476 38646 54488 38698
rect 54540 38646 59624 38698
rect 59676 38646 59688 38698
rect 59740 38646 59752 38698
rect 59804 38646 59816 38698
rect 59868 38646 64952 38698
rect 65004 38646 65016 38698
rect 65068 38646 65080 38698
rect 65132 38646 65144 38698
rect 65196 38646 70280 38698
rect 70332 38646 70344 38698
rect 70396 38646 70408 38698
rect 70460 38646 70472 38698
rect 70524 38646 75608 38698
rect 75660 38646 75672 38698
rect 75724 38646 75736 38698
rect 75788 38646 75800 38698
rect 75852 38646 80936 38698
rect 80988 38646 81000 38698
rect 81052 38646 81064 38698
rect 81116 38646 81128 38698
rect 81180 38646 86264 38698
rect 86316 38646 86328 38698
rect 86380 38646 86392 38698
rect 86444 38646 86456 38698
rect 86508 38646 91592 38698
rect 91644 38646 91656 38698
rect 91708 38646 91720 38698
rect 91772 38646 91784 38698
rect 91836 38646 93642 38698
rect 538 38624 93642 38646
rect 2484 38584 2490 38596
rect 2445 38556 2490 38584
rect 2484 38544 2490 38556
rect 2542 38544 2548 38596
rect 11871 38587 11929 38593
rect 11871 38584 11883 38587
rect 10046 38556 11883 38584
rect 4324 38448 4330 38460
rect 4285 38420 4330 38448
rect 4324 38408 4330 38420
rect 4382 38408 4388 38460
rect 9292 38408 9298 38460
rect 9350 38448 9356 38460
rect 10046 38457 10074 38556
rect 11871 38553 11883 38556
rect 11917 38584 11929 38587
rect 13064 38584 13070 38596
rect 11917 38556 13070 38584
rect 11917 38553 11929 38556
rect 11871 38547 11929 38553
rect 13064 38544 13070 38556
rect 13122 38544 13128 38596
rect 29348 38584 29354 38596
rect 27526 38556 29354 38584
rect 16744 38516 16750 38528
rect 16705 38488 16750 38516
rect 16744 38476 16750 38488
rect 16802 38476 16808 38528
rect 23463 38519 23521 38525
rect 23463 38485 23475 38519
rect 23509 38516 23521 38519
rect 27048 38516 27054 38528
rect 23509 38488 27054 38516
rect 23509 38485 23521 38488
rect 23463 38479 23521 38485
rect 10031 38451 10089 38457
rect 10031 38448 10043 38451
rect 9350 38420 10043 38448
rect 9350 38408 9356 38420
rect 10031 38417 10043 38420
rect 10077 38417 10089 38451
rect 10031 38411 10089 38417
rect 16008 38408 16014 38460
rect 16066 38448 16072 38460
rect 16195 38451 16253 38457
rect 16195 38448 16207 38451
rect 16066 38420 16207 38448
rect 16066 38408 16072 38420
rect 16195 38417 16207 38420
rect 16241 38417 16253 38451
rect 16376 38448 16382 38460
rect 16337 38420 16382 38448
rect 16195 38411 16253 38417
rect 16376 38408 16382 38420
rect 16434 38408 16440 38460
rect 17756 38448 17762 38460
rect 17717 38420 17762 38448
rect 17756 38408 17762 38420
rect 17814 38408 17820 38460
rect 23846 38457 23874 38488
rect 27048 38476 27054 38488
rect 27106 38476 27112 38528
rect 17851 38451 17909 38457
rect 17851 38417 17863 38451
rect 17897 38448 17909 38451
rect 23739 38451 23797 38457
rect 17897 38420 18538 38448
rect 17897 38417 17909 38420
rect 17851 38411 17909 38417
rect 1843 38383 1901 38389
rect 1843 38349 1855 38383
rect 1889 38380 1901 38383
rect 2392 38380 2398 38392
rect 1889 38352 2398 38380
rect 1889 38349 1901 38352
rect 1843 38343 1901 38349
rect 2392 38340 2398 38352
rect 2450 38340 2456 38392
rect 4048 38380 4054 38392
rect 4009 38352 4054 38380
rect 4048 38340 4054 38352
rect 4106 38340 4112 38392
rect 5707 38383 5765 38389
rect 5707 38349 5719 38383
rect 5753 38380 5765 38383
rect 7636 38380 7642 38392
rect 5753 38352 7642 38380
rect 5753 38349 5765 38352
rect 5707 38343 5765 38349
rect 7636 38340 7642 38352
rect 7694 38340 7700 38392
rect 10304 38380 10310 38392
rect 10265 38352 10310 38380
rect 10304 38340 10310 38352
rect 10362 38340 10368 38392
rect 5888 38244 5894 38256
rect 5849 38216 5894 38244
rect 5888 38204 5894 38216
rect 5946 38204 5952 38256
rect 10764 38204 10770 38256
rect 10822 38244 10828 38256
rect 11411 38247 11469 38253
rect 11411 38244 11423 38247
rect 10822 38216 11423 38244
rect 10822 38204 10828 38216
rect 11411 38213 11423 38216
rect 11457 38244 11469 38247
rect 11960 38244 11966 38256
rect 11457 38216 11966 38244
rect 11457 38213 11469 38216
rect 11411 38207 11469 38213
rect 11960 38204 11966 38216
rect 12018 38204 12024 38256
rect 15732 38204 15738 38256
rect 15790 38244 15796 38256
rect 15916 38244 15922 38256
rect 15790 38216 15922 38244
rect 15790 38204 15796 38216
rect 15916 38204 15922 38216
rect 15974 38204 15980 38256
rect 17572 38244 17578 38256
rect 17533 38216 17578 38244
rect 17572 38204 17578 38216
rect 17630 38204 17636 38256
rect 17664 38204 17670 38256
rect 17722 38244 17728 38256
rect 18510 38253 18538 38420
rect 23739 38417 23751 38451
rect 23785 38417 23797 38451
rect 23739 38411 23797 38417
rect 23831 38451 23889 38457
rect 23831 38417 23843 38451
rect 23877 38417 23889 38451
rect 24291 38451 24349 38457
rect 24291 38448 24303 38451
rect 23831 38411 23889 38417
rect 23938 38420 24303 38448
rect 23754 38380 23782 38411
rect 23938 38380 23966 38420
rect 24291 38417 24303 38420
rect 24337 38417 24349 38451
rect 24291 38411 24349 38417
rect 24475 38451 24533 38457
rect 24475 38417 24487 38451
rect 24521 38448 24533 38451
rect 25668 38448 25674 38460
rect 24521 38420 25674 38448
rect 24521 38417 24533 38420
rect 24475 38411 24533 38417
rect 25668 38408 25674 38420
rect 25726 38408 25732 38460
rect 27526 38457 27554 38556
rect 29348 38544 29354 38556
rect 29406 38544 29412 38596
rect 32847 38587 32905 38593
rect 32847 38553 32859 38587
rect 32893 38584 32905 38587
rect 33215 38587 33273 38593
rect 33215 38584 33227 38587
rect 32893 38556 33227 38584
rect 32893 38553 32905 38556
rect 32847 38547 32905 38553
rect 33215 38553 33227 38556
rect 33261 38584 33273 38587
rect 34684 38584 34690 38596
rect 33261 38556 34690 38584
rect 33261 38553 33273 38556
rect 33215 38547 33273 38553
rect 27511 38451 27569 38457
rect 27511 38417 27523 38451
rect 27557 38417 27569 38451
rect 27511 38411 27569 38417
rect 27787 38451 27845 38457
rect 27787 38417 27799 38451
rect 27833 38448 27845 38451
rect 28244 38448 28250 38460
rect 27833 38420 28250 38448
rect 27833 38417 27845 38420
rect 27787 38411 27845 38417
rect 28244 38408 28250 38420
rect 28302 38408 28308 38460
rect 33322 38457 33350 38556
rect 34684 38544 34690 38556
rect 34742 38544 34748 38596
rect 41403 38587 41461 38593
rect 41403 38553 41415 38587
rect 41449 38584 41461 38587
rect 41768 38584 41774 38596
rect 41449 38556 41774 38584
rect 41449 38553 41461 38556
rect 41403 38547 41461 38553
rect 41768 38544 41774 38556
rect 41826 38544 41832 38596
rect 42320 38544 42326 38596
rect 42378 38584 42384 38596
rect 47564 38584 47570 38596
rect 42378 38556 47570 38584
rect 42378 38544 42384 38556
rect 47564 38544 47570 38556
rect 47622 38544 47628 38596
rect 48024 38544 48030 38596
rect 48082 38584 48088 38596
rect 48671 38587 48729 38593
rect 48671 38584 48683 38587
rect 48082 38556 48683 38584
rect 48082 38544 48088 38556
rect 48671 38553 48683 38556
rect 48717 38553 48729 38587
rect 48671 38547 48729 38553
rect 51247 38587 51305 38593
rect 51247 38553 51259 38587
rect 51293 38584 51305 38587
rect 51336 38584 51342 38596
rect 51293 38556 51342 38584
rect 51293 38553 51305 38556
rect 51247 38547 51305 38553
rect 51336 38544 51342 38556
rect 51394 38544 51400 38596
rect 53912 38544 53918 38596
rect 53970 38584 53976 38596
rect 54283 38587 54341 38593
rect 54283 38584 54295 38587
rect 53970 38556 54295 38584
rect 53970 38544 53976 38556
rect 54283 38553 54295 38556
rect 54329 38584 54341 38587
rect 60263 38587 60321 38593
rect 54329 38556 55338 38584
rect 54329 38553 54341 38556
rect 54283 38547 54341 38553
rect 34868 38476 34874 38528
rect 34926 38516 34932 38528
rect 43516 38516 43522 38528
rect 34926 38488 43522 38516
rect 34926 38476 34932 38488
rect 43516 38476 43522 38488
rect 43574 38476 43580 38528
rect 33031 38451 33089 38457
rect 33031 38417 33043 38451
rect 33077 38448 33089 38451
rect 33307 38451 33365 38457
rect 33077 38420 33258 38448
rect 33077 38417 33089 38420
rect 33031 38411 33089 38417
rect 23754 38352 23966 38380
rect 18035 38247 18093 38253
rect 18035 38244 18047 38247
rect 17722 38216 18047 38244
rect 17722 38204 17728 38216
rect 18035 38213 18047 38216
rect 18081 38213 18093 38247
rect 18035 38207 18093 38213
rect 18495 38247 18553 38253
rect 18495 38213 18507 38247
rect 18541 38244 18553 38247
rect 18584 38244 18590 38256
rect 18541 38216 18590 38244
rect 18541 38213 18553 38216
rect 18495 38207 18553 38213
rect 18584 38204 18590 38216
rect 18642 38204 18648 38256
rect 23938 38244 23966 38352
rect 29167 38383 29225 38389
rect 29167 38349 29179 38383
rect 29213 38380 29225 38383
rect 29716 38380 29722 38392
rect 29213 38352 29722 38380
rect 29213 38349 29225 38352
rect 29167 38343 29225 38349
rect 29716 38340 29722 38352
rect 29774 38340 29780 38392
rect 24656 38312 24662 38324
rect 24617 38284 24662 38312
rect 24656 38272 24662 38284
rect 24714 38272 24720 38324
rect 25119 38247 25177 38253
rect 25119 38244 25131 38247
rect 23938 38216 25131 38244
rect 25119 38213 25131 38216
rect 25165 38244 25177 38247
rect 25303 38247 25361 38253
rect 25303 38244 25315 38247
rect 25165 38216 25315 38244
rect 25165 38213 25177 38216
rect 25119 38207 25177 38213
rect 25303 38213 25315 38216
rect 25349 38244 25361 38247
rect 29624 38244 29630 38256
rect 25349 38216 29630 38244
rect 25349 38213 25361 38216
rect 25303 38207 25361 38213
rect 29624 38204 29630 38216
rect 29682 38204 29688 38256
rect 33230 38244 33258 38420
rect 33307 38417 33319 38451
rect 33353 38417 33365 38451
rect 33307 38411 33365 38417
rect 39195 38451 39253 38457
rect 39195 38417 39207 38451
rect 39241 38448 39253 38451
rect 39468 38448 39474 38460
rect 39241 38420 39474 38448
rect 39241 38417 39253 38420
rect 39195 38411 39253 38417
rect 39468 38408 39474 38420
rect 39526 38408 39532 38460
rect 40020 38448 40026 38460
rect 39981 38420 40026 38448
rect 40020 38408 40026 38420
rect 40078 38408 40084 38460
rect 41219 38451 41277 38457
rect 41219 38448 41231 38451
rect 41050 38420 41231 38448
rect 33580 38380 33586 38392
rect 33541 38352 33586 38380
rect 33580 38340 33586 38352
rect 33638 38340 33644 38392
rect 40296 38380 40302 38392
rect 40257 38352 40302 38380
rect 40296 38340 40302 38352
rect 40354 38340 40360 38392
rect 39563 38315 39621 38321
rect 39563 38281 39575 38315
rect 39609 38312 39621 38315
rect 39928 38312 39934 38324
rect 39609 38284 39934 38312
rect 39609 38281 39621 38284
rect 39563 38275 39621 38281
rect 39928 38272 39934 38284
rect 39986 38272 39992 38324
rect 33948 38244 33954 38256
rect 33230 38216 33954 38244
rect 33948 38204 33954 38216
rect 34006 38204 34012 38256
rect 34868 38244 34874 38256
rect 34829 38216 34874 38244
rect 34868 38204 34874 38216
rect 34926 38204 34932 38256
rect 40848 38204 40854 38256
rect 40906 38244 40912 38256
rect 41050 38253 41078 38420
rect 41219 38417 41231 38420
rect 41265 38417 41277 38451
rect 44712 38448 44718 38460
rect 44673 38420 44718 38448
rect 41219 38411 41277 38417
rect 44712 38408 44718 38420
rect 44770 38408 44776 38460
rect 48116 38408 48122 38460
rect 48174 38448 48180 38460
rect 51354 38457 51382 38544
rect 51538 38488 52118 38516
rect 51538 38457 51566 38488
rect 48395 38451 48453 38457
rect 48395 38448 48407 38451
rect 48174 38420 48407 38448
rect 48174 38408 48180 38420
rect 48395 38417 48407 38420
rect 48441 38417 48453 38451
rect 48395 38411 48453 38417
rect 48579 38451 48637 38457
rect 48579 38417 48591 38451
rect 48625 38448 48637 38451
rect 51339 38451 51397 38457
rect 48625 38420 49174 38448
rect 48625 38417 48637 38420
rect 48579 38411 48637 38417
rect 44439 38383 44497 38389
rect 44439 38349 44451 38383
rect 44485 38380 44497 38383
rect 44485 38352 46138 38380
rect 44485 38349 44497 38352
rect 44439 38343 44497 38349
rect 46110 38256 46138 38352
rect 41035 38247 41093 38253
rect 41035 38244 41047 38247
rect 40906 38216 41047 38244
rect 40906 38204 40912 38216
rect 41035 38213 41047 38216
rect 41081 38213 41093 38247
rect 41035 38207 41093 38213
rect 41308 38204 41314 38256
rect 41366 38244 41372 38256
rect 45448 38244 45454 38256
rect 41366 38216 45454 38244
rect 41366 38204 41372 38216
rect 45448 38204 45454 38216
rect 45506 38204 45512 38256
rect 46000 38244 46006 38256
rect 45961 38216 46006 38244
rect 46000 38204 46006 38216
rect 46058 38204 46064 38256
rect 46092 38204 46098 38256
rect 46150 38244 46156 38256
rect 46187 38247 46245 38253
rect 46187 38244 46199 38247
rect 46150 38216 46199 38244
rect 46150 38204 46156 38216
rect 46187 38213 46199 38216
rect 46233 38213 46245 38247
rect 48116 38244 48122 38256
rect 48077 38216 48122 38244
rect 46187 38207 46245 38213
rect 48116 38204 48122 38216
rect 48174 38204 48180 38256
rect 49146 38253 49174 38420
rect 51339 38417 51351 38451
rect 51385 38417 51397 38451
rect 51339 38411 51397 38417
rect 51523 38451 51581 38457
rect 51523 38417 51535 38451
rect 51569 38417 51581 38451
rect 51980 38448 51986 38460
rect 51941 38420 51986 38448
rect 51523 38411 51581 38417
rect 51980 38408 51986 38420
rect 52038 38408 52044 38460
rect 52090 38457 52118 38488
rect 54188 38476 54194 38528
rect 54246 38516 54252 38528
rect 54467 38519 54525 38525
rect 54467 38516 54479 38519
rect 54246 38488 54479 38516
rect 54246 38476 54252 38488
rect 54467 38485 54479 38488
rect 54513 38485 54525 38519
rect 54648 38516 54654 38528
rect 54609 38488 54654 38516
rect 54467 38479 54525 38485
rect 54648 38476 54654 38488
rect 54706 38476 54712 38528
rect 52075 38451 52133 38457
rect 52075 38417 52087 38451
rect 52121 38448 52133 38451
rect 55200 38448 55206 38460
rect 52121 38420 55206 38448
rect 52121 38417 52133 38420
rect 52075 38411 52133 38417
rect 55200 38408 55206 38420
rect 55258 38408 55264 38460
rect 55310 38457 55338 38556
rect 60263 38553 60275 38587
rect 60309 38584 60321 38587
rect 61640 38584 61646 38596
rect 60309 38556 61646 38584
rect 60309 38553 60321 38556
rect 60263 38547 60321 38553
rect 55384 38476 55390 38528
rect 55442 38516 55448 38528
rect 55442 38488 55706 38516
rect 55442 38476 55448 38488
rect 55678 38457 55706 38488
rect 55295 38451 55353 38457
rect 55295 38417 55307 38451
rect 55341 38417 55353 38451
rect 55295 38411 55353 38417
rect 55663 38451 55721 38457
rect 55663 38417 55675 38451
rect 55709 38417 55721 38451
rect 55663 38411 55721 38417
rect 55847 38451 55905 38457
rect 55847 38417 55859 38451
rect 55893 38448 55905 38451
rect 55939 38451 55997 38457
rect 55939 38448 55951 38451
rect 55893 38420 55951 38448
rect 55893 38417 55905 38420
rect 55847 38411 55905 38417
rect 55939 38417 55951 38420
rect 55985 38448 55997 38451
rect 59064 38448 59070 38460
rect 55985 38420 59070 38448
rect 55985 38417 55997 38420
rect 55939 38411 55997 38417
rect 59064 38408 59070 38420
rect 59122 38408 59128 38460
rect 60370 38457 60398 38556
rect 61640 38544 61646 38556
rect 61698 38544 61704 38596
rect 63664 38584 63670 38596
rect 63625 38556 63670 38584
rect 63664 38544 63670 38556
rect 63722 38544 63728 38596
rect 68632 38544 68638 38596
rect 68690 38584 68696 38596
rect 72404 38584 72410 38596
rect 68690 38556 72410 38584
rect 68690 38544 68696 38556
rect 72404 38544 72410 38556
rect 72462 38544 72468 38596
rect 72499 38587 72557 38593
rect 72499 38553 72511 38587
rect 72545 38584 72557 38587
rect 74244 38584 74250 38596
rect 72545 38556 74250 38584
rect 72545 38553 72557 38556
rect 72499 38547 72557 38553
rect 61364 38476 61370 38528
rect 61422 38516 61428 38528
rect 72514 38516 72542 38547
rect 74244 38544 74250 38556
rect 74302 38584 74308 38596
rect 76452 38584 76458 38596
rect 74302 38556 76458 38584
rect 74302 38544 74308 38556
rect 76452 38544 76458 38556
rect 76510 38544 76516 38596
rect 77096 38544 77102 38596
rect 77154 38584 77160 38596
rect 80043 38587 80101 38593
rect 80043 38584 80055 38587
rect 77154 38556 80055 38584
rect 77154 38544 77160 38556
rect 80043 38553 80055 38556
rect 80089 38553 80101 38587
rect 80043 38547 80101 38553
rect 88412 38544 88418 38596
rect 88470 38584 88476 38596
rect 88783 38587 88841 38593
rect 88783 38584 88795 38587
rect 88470 38556 88795 38584
rect 88470 38544 88476 38556
rect 88783 38553 88795 38556
rect 88829 38553 88841 38587
rect 88783 38547 88841 38553
rect 90163 38587 90221 38593
rect 90163 38553 90175 38587
rect 90209 38584 90221 38587
rect 90712 38584 90718 38596
rect 90209 38556 90718 38584
rect 90209 38553 90221 38556
rect 90163 38547 90221 38553
rect 73416 38516 73422 38528
rect 61422 38488 63618 38516
rect 61422 38476 61428 38488
rect 60355 38451 60413 38457
rect 60355 38417 60367 38451
rect 60401 38417 60413 38451
rect 63483 38451 63541 38457
rect 63483 38448 63495 38451
rect 60355 38411 60413 38417
rect 63314 38420 63495 38448
rect 55387 38383 55445 38389
rect 55387 38349 55399 38383
rect 55433 38349 55445 38383
rect 60628 38380 60634 38392
rect 60589 38352 60634 38380
rect 55387 38343 55445 38349
rect 52440 38312 52446 38324
rect 52401 38284 52446 38312
rect 52440 38272 52446 38284
rect 52498 38272 52504 38324
rect 49131 38247 49189 38253
rect 49131 38213 49143 38247
rect 49177 38244 49189 38247
rect 53912 38244 53918 38256
rect 49177 38216 53918 38244
rect 49177 38213 49189 38216
rect 49131 38207 49189 38213
rect 53912 38204 53918 38216
rect 53970 38204 53976 38256
rect 55402 38244 55430 38343
rect 60628 38340 60634 38352
rect 60686 38340 60692 38392
rect 56215 38247 56273 38253
rect 56215 38244 56227 38247
rect 55402 38216 56227 38244
rect 56215 38213 56227 38216
rect 56261 38244 56273 38247
rect 57960 38244 57966 38256
rect 56261 38216 57966 38244
rect 56261 38213 56273 38216
rect 56215 38207 56273 38213
rect 57960 38204 57966 38216
rect 58018 38204 58024 38256
rect 61732 38244 61738 38256
rect 61693 38216 61738 38244
rect 61732 38204 61738 38216
rect 61790 38204 61796 38256
rect 63204 38204 63210 38256
rect 63262 38244 63268 38256
rect 63314 38253 63342 38420
rect 63483 38417 63495 38420
rect 63529 38417 63541 38451
rect 63483 38411 63541 38417
rect 63590 38312 63618 38488
rect 67638 38488 72542 38516
rect 73377 38488 73422 38516
rect 64124 38408 64130 38460
rect 64182 38448 64188 38460
rect 67638 38457 67666 38488
rect 73416 38476 73422 38488
rect 73474 38476 73480 38528
rect 73784 38476 73790 38528
rect 73842 38516 73848 38528
rect 73842 38488 74474 38516
rect 73842 38476 73848 38488
rect 66887 38451 66945 38457
rect 66887 38448 66899 38451
rect 64182 38420 66899 38448
rect 64182 38408 64188 38420
rect 66887 38417 66899 38420
rect 66933 38417 66945 38451
rect 66887 38411 66945 38417
rect 67071 38451 67129 38457
rect 67071 38417 67083 38451
rect 67117 38448 67129 38451
rect 67623 38451 67681 38457
rect 67623 38448 67635 38451
rect 67117 38420 67635 38448
rect 67117 38417 67129 38420
rect 67071 38411 67129 38417
rect 67623 38417 67635 38420
rect 67669 38417 67681 38451
rect 67804 38448 67810 38460
rect 67765 38420 67810 38448
rect 67623 38411 67681 38417
rect 67804 38408 67810 38420
rect 67862 38448 67868 38460
rect 68356 38448 68362 38460
rect 67862 38420 68362 38448
rect 67862 38408 67868 38420
rect 68356 38408 68362 38420
rect 68414 38408 68420 38460
rect 69092 38448 69098 38460
rect 69053 38420 69098 38448
rect 69092 38408 69098 38420
rect 69150 38408 69156 38460
rect 72315 38451 72373 38457
rect 72315 38448 72327 38451
rect 72238 38420 72327 38448
rect 68374 38380 68402 38408
rect 69187 38383 69245 38389
rect 69187 38380 69199 38383
rect 68374 38352 69199 38380
rect 69187 38349 69199 38352
rect 69233 38349 69245 38383
rect 69187 38343 69245 38349
rect 72238 38312 72266 38420
rect 72315 38417 72327 38420
rect 72361 38417 72373 38451
rect 72315 38411 72373 38417
rect 72588 38408 72594 38460
rect 72646 38448 72652 38460
rect 73692 38448 73698 38460
rect 72646 38420 73698 38448
rect 72646 38408 72652 38420
rect 73692 38408 73698 38420
rect 73750 38448 73756 38460
rect 74446 38457 74474 38488
rect 83830 38488 88734 38516
rect 74063 38451 74121 38457
rect 74063 38448 74075 38451
rect 73750 38420 74075 38448
rect 73750 38408 73756 38420
rect 74063 38417 74075 38420
rect 74109 38417 74121 38451
rect 74063 38411 74121 38417
rect 74431 38451 74489 38457
rect 74431 38417 74443 38451
rect 74477 38417 74489 38451
rect 74431 38411 74489 38417
rect 74615 38451 74673 38457
rect 74615 38417 74627 38451
rect 74661 38448 74673 38451
rect 74980 38448 74986 38460
rect 74661 38420 74986 38448
rect 74661 38417 74673 38420
rect 74615 38411 74673 38417
rect 74980 38408 74986 38420
rect 75038 38408 75044 38460
rect 75440 38408 75446 38460
rect 75498 38448 75504 38460
rect 77743 38451 77801 38457
rect 77743 38448 77755 38451
rect 75498 38420 77755 38448
rect 75498 38408 75504 38420
rect 77743 38417 77755 38420
rect 77789 38417 77801 38451
rect 77743 38411 77801 38417
rect 79951 38451 80009 38457
rect 79951 38417 79963 38451
rect 79997 38448 80009 38451
rect 80408 38448 80414 38460
rect 79997 38420 80414 38448
rect 79997 38417 80009 38420
rect 79951 38411 80009 38417
rect 80408 38408 80414 38420
rect 80466 38408 80472 38460
rect 82800 38408 82806 38460
rect 82858 38448 82864 38460
rect 83079 38451 83137 38457
rect 83079 38448 83091 38451
rect 82858 38420 83091 38448
rect 82858 38408 82864 38420
rect 83079 38417 83091 38420
rect 83125 38417 83137 38451
rect 83260 38448 83266 38460
rect 83173 38420 83266 38448
rect 83079 38411 83137 38417
rect 83260 38408 83266 38420
rect 83318 38448 83324 38460
rect 83830 38457 83858 38488
rect 83815 38451 83873 38457
rect 83815 38448 83827 38451
rect 83318 38420 83827 38448
rect 83318 38408 83324 38420
rect 83815 38417 83827 38420
rect 83861 38417 83873 38451
rect 83815 38411 83873 38417
rect 83999 38451 84057 38457
rect 83999 38417 84011 38451
rect 84045 38448 84057 38451
rect 85287 38451 85345 38457
rect 84045 38420 84318 38448
rect 84045 38417 84057 38420
rect 83999 38411 84057 38417
rect 74155 38383 74213 38389
rect 74155 38349 74167 38383
rect 74201 38380 74213 38383
rect 74704 38380 74710 38392
rect 74201 38352 74710 38380
rect 74201 38349 74213 38352
rect 74155 38343 74213 38349
rect 74704 38340 74710 38352
rect 74762 38340 74768 38392
rect 77467 38383 77525 38389
rect 77467 38349 77479 38383
rect 77513 38349 77525 38383
rect 77467 38343 77525 38349
rect 63590 38284 72266 38312
rect 72238 38256 72266 38284
rect 77482 38256 77510 38343
rect 84290 38312 84318 38420
rect 85287 38417 85299 38451
rect 85333 38448 85345 38451
rect 86388 38448 86394 38460
rect 85333 38420 86394 38448
rect 85333 38417 85345 38420
rect 85287 38411 85345 38417
rect 86388 38408 86394 38420
rect 86446 38408 86452 38460
rect 88706 38392 88734 38488
rect 88798 38448 88826 38547
rect 90712 38544 90718 38556
rect 90770 38544 90776 38596
rect 91543 38519 91601 38525
rect 91543 38516 91555 38519
rect 89902 38488 91555 38516
rect 89902 38460 89930 38488
rect 91543 38485 91555 38488
rect 91589 38485 91601 38519
rect 91543 38479 91601 38485
rect 88967 38451 89025 38457
rect 88967 38448 88979 38451
rect 88798 38420 88979 38448
rect 88967 38417 88979 38420
rect 89013 38417 89025 38451
rect 88967 38411 89025 38417
rect 89151 38451 89209 38457
rect 89151 38417 89163 38451
rect 89197 38448 89209 38451
rect 89703 38451 89761 38457
rect 89703 38448 89715 38451
rect 89197 38420 89715 38448
rect 89197 38417 89209 38420
rect 89151 38411 89209 38417
rect 89703 38417 89715 38420
rect 89749 38417 89761 38451
rect 89884 38448 89890 38460
rect 89845 38420 89890 38448
rect 89703 38411 89761 38417
rect 84367 38383 84425 38389
rect 84367 38349 84379 38383
rect 84413 38380 84425 38383
rect 85100 38380 85106 38392
rect 84413 38352 85106 38380
rect 84413 38349 84425 38352
rect 84367 38343 84425 38349
rect 85100 38340 85106 38352
rect 85158 38340 85164 38392
rect 88688 38340 88694 38392
rect 88746 38380 88752 38392
rect 89166 38380 89194 38411
rect 89884 38408 89890 38420
rect 89942 38408 89948 38460
rect 91448 38448 91454 38460
rect 91409 38420 91454 38448
rect 91448 38408 91454 38420
rect 91506 38408 91512 38460
rect 88746 38352 89194 38380
rect 88746 38340 88752 38352
rect 84290 38284 84594 38312
rect 63299 38247 63357 38253
rect 63299 38244 63311 38247
rect 63262 38216 63311 38244
rect 63262 38204 63268 38216
rect 63299 38213 63311 38216
rect 63345 38213 63357 38247
rect 63299 38207 63357 38213
rect 68083 38247 68141 38253
rect 68083 38213 68095 38247
rect 68129 38244 68141 38247
rect 68264 38244 68270 38256
rect 68129 38216 68270 38244
rect 68129 38213 68141 38216
rect 68083 38207 68141 38213
rect 68264 38204 68270 38216
rect 68322 38204 68328 38256
rect 68540 38204 68546 38256
rect 68598 38244 68604 38256
rect 69644 38244 69650 38256
rect 68598 38216 69650 38244
rect 68598 38204 68604 38216
rect 69644 38204 69650 38216
rect 69702 38204 69708 38256
rect 72220 38244 72226 38256
rect 72181 38216 72226 38244
rect 72220 38204 72226 38216
rect 72278 38204 72284 38256
rect 77375 38247 77433 38253
rect 77375 38213 77387 38247
rect 77421 38244 77433 38247
rect 77464 38244 77470 38256
rect 77421 38216 77470 38244
rect 77421 38213 77433 38216
rect 77375 38207 77433 38213
rect 77464 38204 77470 38216
rect 77522 38204 77528 38256
rect 79031 38247 79089 38253
rect 79031 38213 79043 38247
rect 79077 38244 79089 38247
rect 79212 38244 79218 38256
rect 79077 38216 79218 38244
rect 79077 38213 79089 38216
rect 79031 38207 79089 38213
rect 79212 38204 79218 38216
rect 79270 38204 79276 38256
rect 84566 38253 84594 38284
rect 84551 38247 84609 38253
rect 84551 38213 84563 38247
rect 84597 38244 84609 38247
rect 85284 38244 85290 38256
rect 84597 38216 85290 38244
rect 84597 38213 84609 38216
rect 84551 38207 84609 38213
rect 85284 38204 85290 38216
rect 85342 38244 85348 38256
rect 85379 38247 85437 38253
rect 85379 38244 85391 38247
rect 85342 38216 85391 38244
rect 85342 38204 85348 38216
rect 85379 38213 85391 38216
rect 85425 38213 85437 38247
rect 85379 38207 85437 38213
rect 538 38154 93642 38176
rect 538 38102 3680 38154
rect 3732 38102 3744 38154
rect 3796 38102 3808 38154
rect 3860 38102 3872 38154
rect 3924 38102 9008 38154
rect 9060 38102 9072 38154
rect 9124 38102 9136 38154
rect 9188 38102 9200 38154
rect 9252 38102 14336 38154
rect 14388 38102 14400 38154
rect 14452 38102 14464 38154
rect 14516 38102 14528 38154
rect 14580 38102 19664 38154
rect 19716 38102 19728 38154
rect 19780 38102 19792 38154
rect 19844 38102 19856 38154
rect 19908 38102 24992 38154
rect 25044 38102 25056 38154
rect 25108 38102 25120 38154
rect 25172 38102 25184 38154
rect 25236 38102 30320 38154
rect 30372 38102 30384 38154
rect 30436 38102 30448 38154
rect 30500 38102 30512 38154
rect 30564 38102 35648 38154
rect 35700 38102 35712 38154
rect 35764 38102 35776 38154
rect 35828 38102 35840 38154
rect 35892 38102 40976 38154
rect 41028 38102 41040 38154
rect 41092 38102 41104 38154
rect 41156 38102 41168 38154
rect 41220 38102 46304 38154
rect 46356 38102 46368 38154
rect 46420 38102 46432 38154
rect 46484 38102 46496 38154
rect 46548 38102 51632 38154
rect 51684 38102 51696 38154
rect 51748 38102 51760 38154
rect 51812 38102 51824 38154
rect 51876 38102 56960 38154
rect 57012 38102 57024 38154
rect 57076 38102 57088 38154
rect 57140 38102 57152 38154
rect 57204 38102 62288 38154
rect 62340 38102 62352 38154
rect 62404 38102 62416 38154
rect 62468 38102 62480 38154
rect 62532 38102 67616 38154
rect 67668 38102 67680 38154
rect 67732 38102 67744 38154
rect 67796 38102 67808 38154
rect 67860 38102 72944 38154
rect 72996 38102 73008 38154
rect 73060 38102 73072 38154
rect 73124 38102 73136 38154
rect 73188 38102 78272 38154
rect 78324 38102 78336 38154
rect 78388 38102 78400 38154
rect 78452 38102 78464 38154
rect 78516 38102 83600 38154
rect 83652 38102 83664 38154
rect 83716 38102 83728 38154
rect 83780 38102 83792 38154
rect 83844 38102 88928 38154
rect 88980 38102 88992 38154
rect 89044 38102 89056 38154
rect 89108 38102 89120 38154
rect 89172 38102 93642 38154
rect 538 38080 93642 38102
rect 9292 38040 9298 38052
rect 9253 38012 9298 38040
rect 9292 38000 9298 38012
rect 9350 38000 9356 38052
rect 9752 38000 9758 38052
rect 9810 38040 9816 38052
rect 10396 38040 10402 38052
rect 9810 38012 10402 38040
rect 9810 38000 9816 38012
rect 10396 38000 10402 38012
rect 10454 38000 10460 38052
rect 17483 38043 17541 38049
rect 17483 38009 17495 38043
rect 17529 38040 17541 38043
rect 17572 38040 17578 38052
rect 17529 38012 17578 38040
rect 17529 38009 17541 38012
rect 17483 38003 17541 38009
rect 17572 38000 17578 38012
rect 17630 38040 17636 38052
rect 20151 38043 20209 38049
rect 20151 38040 20163 38043
rect 17630 38012 20163 38040
rect 17630 38000 17636 38012
rect 20151 38009 20163 38012
rect 20197 38040 20209 38043
rect 20240 38040 20246 38052
rect 20197 38012 20246 38040
rect 20197 38009 20209 38012
rect 20151 38003 20209 38009
rect 20240 38000 20246 38012
rect 20298 38000 20304 38052
rect 27416 38000 27422 38052
rect 27474 38040 27480 38052
rect 27603 38043 27661 38049
rect 27603 38040 27615 38043
rect 27474 38012 27615 38040
rect 27474 38000 27480 38012
rect 27603 38009 27615 38012
rect 27649 38009 27661 38043
rect 27603 38003 27661 38009
rect 33215 38043 33273 38049
rect 33215 38009 33227 38043
rect 33261 38040 33273 38043
rect 33580 38040 33586 38052
rect 33261 38012 33586 38040
rect 33261 38009 33273 38012
rect 33215 38003 33273 38009
rect 33580 38000 33586 38012
rect 33638 38000 33644 38052
rect 40020 38000 40026 38052
rect 40078 38040 40084 38052
rect 40851 38043 40909 38049
rect 40851 38040 40863 38043
rect 40078 38012 40863 38040
rect 40078 38000 40084 38012
rect 40851 38009 40863 38012
rect 40897 38009 40909 38043
rect 42139 38043 42197 38049
rect 40851 38003 40909 38009
rect 41142 38012 41354 38040
rect 8648 37932 8654 37984
rect 8706 37972 8712 37984
rect 8835 37975 8893 37981
rect 8835 37972 8847 37975
rect 8706 37944 8847 37972
rect 8706 37932 8712 37944
rect 8835 37941 8847 37944
rect 8881 37972 8893 37975
rect 9108 37972 9114 37984
rect 8881 37944 9114 37972
rect 8881 37941 8893 37944
rect 8835 37935 8893 37941
rect 9108 37932 9114 37944
rect 9166 37932 9172 37984
rect 17756 37972 17762 37984
rect 16578 37944 17762 37972
rect 7731 37907 7789 37913
rect 7731 37873 7743 37907
rect 7777 37904 7789 37907
rect 8096 37904 8102 37916
rect 7777 37876 8102 37904
rect 7777 37873 7789 37876
rect 7731 37867 7789 37873
rect 8096 37864 8102 37876
rect 8154 37864 8160 37916
rect 11960 37864 11966 37916
rect 12018 37904 12024 37916
rect 16578 37913 16606 37944
rect 17756 37932 17762 37944
rect 17814 37932 17820 37984
rect 29624 37932 29630 37984
rect 29682 37972 29688 37984
rect 29682 37944 30038 37972
rect 29682 37932 29688 37944
rect 16563 37907 16621 37913
rect 12018 37876 16238 37904
rect 12018 37864 12024 37876
rect 2119 37839 2177 37845
rect 2119 37805 2131 37839
rect 2165 37836 2177 37839
rect 2208 37836 2214 37848
rect 2165 37808 2214 37836
rect 2165 37805 2177 37808
rect 2119 37799 2177 37805
rect 2208 37796 2214 37808
rect 2266 37796 2272 37848
rect 2392 37836 2398 37848
rect 2353 37808 2398 37836
rect 2392 37796 2398 37808
rect 2450 37796 2456 37848
rect 7452 37836 7458 37848
rect 7413 37808 7458 37836
rect 7452 37796 7458 37808
rect 7510 37796 7516 37848
rect 12515 37839 12573 37845
rect 12515 37805 12527 37839
rect 12561 37805 12573 37839
rect 12788 37836 12794 37848
rect 12749 37808 12794 37836
rect 12515 37799 12573 37805
rect 3775 37771 3833 37777
rect 3775 37737 3787 37771
rect 3821 37768 3833 37771
rect 4416 37768 4422 37780
rect 3821 37740 4422 37768
rect 3821 37737 3833 37740
rect 3775 37731 3833 37737
rect 4416 37728 4422 37740
rect 4474 37728 4480 37780
rect 3956 37700 3962 37712
rect 3917 37672 3962 37700
rect 3956 37660 3962 37672
rect 4014 37660 4020 37712
rect 12530 37700 12558 37799
rect 12788 37796 12794 37808
rect 12846 37796 12852 37848
rect 16210 37845 16238 37876
rect 16563 37873 16575 37907
rect 16609 37873 16621 37907
rect 16563 37867 16621 37873
rect 17940 37864 17946 37916
rect 17998 37904 18004 37916
rect 18219 37907 18277 37913
rect 18219 37904 18231 37907
rect 17998 37876 18231 37904
rect 17998 37864 18004 37876
rect 18219 37873 18231 37876
rect 18265 37873 18277 37907
rect 18219 37867 18277 37873
rect 20608 37864 20614 37916
rect 20666 37904 20672 37916
rect 20887 37907 20945 37913
rect 20887 37904 20899 37907
rect 20666 37876 20899 37904
rect 20666 37864 20672 37876
rect 20887 37873 20899 37876
rect 20933 37873 20945 37907
rect 20887 37867 20945 37873
rect 21068 37864 21074 37916
rect 21126 37904 21132 37916
rect 22911 37907 22969 37913
rect 22911 37904 22923 37907
rect 21126 37876 22923 37904
rect 21126 37864 21132 37876
rect 22911 37873 22923 37876
rect 22957 37904 22969 37907
rect 23095 37907 23153 37913
rect 23095 37904 23107 37907
rect 22957 37876 23107 37904
rect 22957 37873 22969 37876
rect 22911 37867 22969 37873
rect 23095 37873 23107 37876
rect 23141 37873 23153 37907
rect 23095 37867 23153 37873
rect 23371 37907 23429 37913
rect 23371 37873 23383 37907
rect 23417 37904 23429 37907
rect 24656 37904 24662 37916
rect 23417 37876 24662 37904
rect 23417 37873 23429 37876
rect 23371 37867 23429 37873
rect 24656 37864 24662 37876
rect 24714 37864 24720 37916
rect 25668 37904 25674 37916
rect 25629 37876 25674 37904
rect 25668 37864 25674 37876
rect 25726 37864 25732 37916
rect 27968 37864 27974 37916
rect 28026 37904 28032 37916
rect 29903 37907 29961 37913
rect 29903 37904 29915 37907
rect 28026 37876 29915 37904
rect 28026 37864 28032 37876
rect 29903 37873 29915 37876
rect 29949 37873 29961 37907
rect 29903 37867 29961 37873
rect 16195 37839 16253 37845
rect 16195 37805 16207 37839
rect 16241 37805 16253 37839
rect 16195 37799 16253 37805
rect 17759 37839 17817 37845
rect 17759 37805 17771 37839
rect 17805 37805 17817 37839
rect 20424 37836 20430 37848
rect 20385 37808 20430 37836
rect 17759 37799 17817 37805
rect 14168 37768 14174 37780
rect 14081 37740 14174 37768
rect 14168 37728 14174 37740
rect 14226 37768 14232 37780
rect 15824 37768 15830 37780
rect 14226 37740 15830 37768
rect 14226 37728 14232 37740
rect 15824 37728 15830 37740
rect 15882 37728 15888 37780
rect 16008 37768 16014 37780
rect 15969 37740 16014 37768
rect 16008 37728 16014 37740
rect 16066 37728 16072 37780
rect 17664 37768 17670 37780
rect 17625 37740 17670 37768
rect 17664 37728 17670 37740
rect 17722 37728 17728 37780
rect 17774 37768 17802 37799
rect 20424 37796 20430 37808
rect 20482 37796 20488 37848
rect 24751 37839 24809 37845
rect 24751 37805 24763 37839
rect 24797 37836 24809 37839
rect 25487 37839 25545 37845
rect 25487 37836 25499 37839
rect 24797 37808 25499 37836
rect 24797 37805 24809 37808
rect 24751 37799 24809 37805
rect 25487 37805 25499 37808
rect 25533 37836 25545 37839
rect 25576 37836 25582 37848
rect 25533 37808 25582 37836
rect 25533 37805 25545 37808
rect 25487 37799 25545 37805
rect 25576 37796 25582 37808
rect 25634 37796 25640 37848
rect 27324 37796 27330 37848
rect 27382 37836 27388 37848
rect 27419 37839 27477 37845
rect 27419 37836 27431 37839
rect 27382 37808 27431 37836
rect 27382 37796 27388 37808
rect 27419 37805 27431 37808
rect 27465 37805 27477 37839
rect 27419 37799 27477 37805
rect 28707 37839 28765 37845
rect 28707 37805 28719 37839
rect 28753 37805 28765 37839
rect 28707 37799 28765 37805
rect 17940 37768 17946 37780
rect 17774 37740 17946 37768
rect 17940 37728 17946 37740
rect 17998 37768 18004 37780
rect 18311 37771 18369 37777
rect 18311 37768 18323 37771
rect 17998 37740 18323 37768
rect 17998 37728 18004 37740
rect 18311 37737 18323 37740
rect 18357 37737 18369 37771
rect 20332 37768 20338 37780
rect 20293 37740 20338 37768
rect 18311 37731 18369 37737
rect 20332 37728 20338 37740
rect 20390 37728 20396 37780
rect 27048 37728 27054 37780
rect 27106 37768 27112 37780
rect 28722 37768 28750 37799
rect 29716 37796 29722 37848
rect 29774 37836 29780 37848
rect 29811 37839 29869 37845
rect 29811 37836 29823 37839
rect 29774 37808 29823 37836
rect 29774 37796 29780 37808
rect 29811 37805 29823 37808
rect 29857 37805 29869 37839
rect 30010 37836 30038 37944
rect 34868 37932 34874 37984
rect 34926 37972 34932 37984
rect 41142 37972 41170 38012
rect 34926 37944 41170 37972
rect 41326 37972 41354 38012
rect 42139 38009 42151 38043
rect 42185 38040 42197 38043
rect 42320 38040 42326 38052
rect 42185 38012 42326 38040
rect 42185 38009 42197 38012
rect 42139 38003 42197 38009
rect 42320 38000 42326 38012
rect 42378 38000 42384 38052
rect 69092 38000 69098 38052
rect 69150 38040 69156 38052
rect 69371 38043 69429 38049
rect 69371 38040 69383 38043
rect 69150 38012 69383 38040
rect 69150 38000 69156 38012
rect 69371 38009 69383 38012
rect 69417 38009 69429 38043
rect 69371 38003 69429 38009
rect 72220 38000 72226 38052
rect 72278 38040 72284 38052
rect 82064 38040 82070 38052
rect 72278 38012 82070 38040
rect 72278 38000 72284 38012
rect 82064 38000 82070 38012
rect 82122 38000 82128 38052
rect 86388 38040 86394 38052
rect 86349 38012 86394 38040
rect 86388 38000 86394 38012
rect 86446 38000 86452 38052
rect 90160 38040 90166 38052
rect 90121 38012 90166 38040
rect 90160 38000 90166 38012
rect 90218 38000 90224 38052
rect 45356 37972 45362 37984
rect 41326 37944 45362 37972
rect 34926 37932 34932 37944
rect 45356 37932 45362 37944
rect 45414 37932 45420 37984
rect 47199 37975 47257 37981
rect 47199 37941 47211 37975
rect 47245 37972 47257 37975
rect 47380 37972 47386 37984
rect 47245 37944 47386 37972
rect 47245 37941 47257 37944
rect 47199 37935 47257 37941
rect 47380 37932 47386 37944
rect 47438 37932 47444 37984
rect 50894 37944 52302 37972
rect 31924 37864 31930 37916
rect 31982 37904 31988 37916
rect 32019 37907 32077 37913
rect 32019 37904 32031 37907
rect 31982 37876 32031 37904
rect 31982 37864 31988 37876
rect 32019 37873 32031 37876
rect 32065 37873 32077 37907
rect 32019 37867 32077 37873
rect 34040 37864 34046 37916
rect 34098 37904 34104 37916
rect 34960 37904 34966 37916
rect 34098 37876 34966 37904
rect 34098 37864 34104 37876
rect 34960 37864 34966 37876
rect 35018 37864 35024 37916
rect 36616 37904 36622 37916
rect 36577 37876 36622 37904
rect 36616 37864 36622 37876
rect 36674 37864 36680 37916
rect 37812 37864 37818 37916
rect 37870 37904 37876 37916
rect 37870 37876 40526 37904
rect 37870 37864 37876 37876
rect 31743 37839 31801 37845
rect 31743 37836 31755 37839
rect 30010 37808 31755 37836
rect 29811 37799 29869 37805
rect 31743 37805 31755 37808
rect 31789 37836 31801 37839
rect 31835 37839 31893 37845
rect 31835 37836 31847 37839
rect 31789 37808 31847 37836
rect 31789 37805 31801 37808
rect 31743 37799 31801 37805
rect 31835 37805 31847 37808
rect 31881 37836 31893 37839
rect 32203 37839 32261 37845
rect 32203 37836 32215 37839
rect 31881 37808 32215 37836
rect 31881 37805 31893 37808
rect 31835 37799 31893 37805
rect 32203 37805 32215 37808
rect 32249 37836 32261 37839
rect 32755 37839 32813 37845
rect 32755 37836 32767 37839
rect 32249 37808 32767 37836
rect 32249 37805 32261 37808
rect 32203 37799 32261 37805
rect 32755 37805 32767 37808
rect 32801 37805 32813 37839
rect 32755 37799 32813 37805
rect 32939 37839 32997 37845
rect 32939 37805 32951 37839
rect 32985 37836 32997 37839
rect 33396 37836 33402 37848
rect 32985 37808 33402 37836
rect 32985 37805 32997 37808
rect 32939 37799 32997 37805
rect 29075 37771 29133 37777
rect 29075 37768 29087 37771
rect 27106 37740 29087 37768
rect 27106 37728 27112 37740
rect 29075 37737 29087 37740
rect 29121 37768 29133 37771
rect 32292 37768 32298 37780
rect 29121 37740 32298 37768
rect 29121 37737 29133 37740
rect 29075 37731 29133 37737
rect 32292 37728 32298 37740
rect 32350 37728 32356 37780
rect 32770 37768 32798 37799
rect 33396 37796 33402 37808
rect 33454 37836 33460 37848
rect 33580 37836 33586 37848
rect 33454 37808 33586 37836
rect 33454 37796 33460 37808
rect 33580 37796 33586 37808
rect 33638 37796 33644 37848
rect 34687 37839 34745 37845
rect 34687 37805 34699 37839
rect 34733 37836 34745 37839
rect 34779 37839 34837 37845
rect 34779 37836 34791 37839
rect 34733 37808 34791 37836
rect 34733 37805 34745 37808
rect 34687 37799 34745 37805
rect 34779 37805 34791 37808
rect 34825 37836 34837 37839
rect 35144 37836 35150 37848
rect 34825 37808 35150 37836
rect 34825 37805 34837 37808
rect 34779 37799 34837 37805
rect 35144 37796 35150 37808
rect 35202 37796 35208 37848
rect 36435 37839 36493 37845
rect 36435 37805 36447 37839
rect 36481 37836 36493 37839
rect 36711 37839 36769 37845
rect 36711 37836 36723 37839
rect 36481 37808 36723 37836
rect 36481 37805 36493 37808
rect 36435 37799 36493 37805
rect 36711 37805 36723 37808
rect 36757 37805 36769 37839
rect 36711 37799 36769 37805
rect 37171 37839 37229 37845
rect 37171 37805 37183 37839
rect 37217 37805 37229 37839
rect 37171 37799 37229 37805
rect 37263 37839 37321 37845
rect 37263 37805 37275 37839
rect 37309 37836 37321 37839
rect 40388 37836 40394 37848
rect 37309 37808 40394 37836
rect 37309 37805 37321 37808
rect 37263 37799 37321 37805
rect 36450 37768 36478 37799
rect 32770 37740 36478 37768
rect 14076 37700 14082 37712
rect 12530 37672 14082 37700
rect 14076 37660 14082 37672
rect 14134 37700 14140 37712
rect 14263 37703 14321 37709
rect 14263 37700 14275 37703
rect 14134 37672 14275 37700
rect 14134 37660 14140 37672
rect 14263 37669 14275 37672
rect 14309 37669 14321 37703
rect 27324 37700 27330 37712
rect 27285 37672 27330 37700
rect 14263 37663 14321 37669
rect 27324 37660 27330 37672
rect 27382 37660 27388 37712
rect 28888 37700 28894 37712
rect 28849 37672 28894 37700
rect 28888 37660 28894 37672
rect 28946 37660 28952 37712
rect 29716 37700 29722 37712
rect 29677 37672 29722 37700
rect 29716 37660 29722 37672
rect 29774 37660 29780 37712
rect 33580 37700 33586 37712
rect 33541 37672 33586 37700
rect 33580 37660 33586 37672
rect 33638 37660 33644 37712
rect 34960 37700 34966 37712
rect 34921 37672 34966 37700
rect 34960 37660 34966 37672
rect 35018 37660 35024 37712
rect 35052 37660 35058 37712
rect 35110 37700 35116 37712
rect 37186 37700 37214 37799
rect 37646 37780 37674 37808
rect 40388 37796 40394 37808
rect 40446 37796 40452 37848
rect 40498 37836 40526 37876
rect 40572 37864 40578 37916
rect 40630 37904 40636 37916
rect 47291 37907 47349 37913
rect 47291 37904 47303 37907
rect 40630 37876 47303 37904
rect 40630 37864 40636 37876
rect 47291 37873 47303 37876
rect 47337 37873 47349 37907
rect 47472 37904 47478 37916
rect 47433 37876 47478 37904
rect 47291 37867 47349 37873
rect 40759 37839 40817 37845
rect 40498 37808 40710 37836
rect 37628 37728 37634 37780
rect 37686 37728 37692 37780
rect 37812 37768 37818 37780
rect 37773 37740 37818 37768
rect 37812 37728 37818 37740
rect 37870 37728 37876 37780
rect 40572 37768 40578 37780
rect 40406 37740 40578 37768
rect 38091 37703 38149 37709
rect 38091 37700 38103 37703
rect 35110 37672 38103 37700
rect 35110 37660 35116 37672
rect 38091 37669 38103 37672
rect 38137 37700 38149 37703
rect 39560 37700 39566 37712
rect 38137 37672 39566 37700
rect 38137 37669 38149 37672
rect 38091 37663 38149 37669
rect 39560 37660 39566 37672
rect 39618 37660 39624 37712
rect 39836 37660 39842 37712
rect 39894 37700 39900 37712
rect 40406 37709 40434 37740
rect 40572 37728 40578 37740
rect 40630 37728 40636 37780
rect 40682 37768 40710 37808
rect 40759 37805 40771 37839
rect 40805 37836 40817 37839
rect 41216 37836 41222 37848
rect 40805 37808 41222 37836
rect 40805 37805 40817 37808
rect 40759 37799 40817 37805
rect 41216 37796 41222 37808
rect 41274 37796 41280 37848
rect 41768 37796 41774 37848
rect 41826 37836 41832 37848
rect 41955 37839 42013 37845
rect 41955 37836 41967 37839
rect 41826 37808 41967 37836
rect 41826 37796 41832 37808
rect 41955 37805 41967 37808
rect 42001 37805 42013 37839
rect 41955 37799 42013 37805
rect 43516 37796 43522 37848
rect 43574 37836 43580 37848
rect 45359 37839 45417 37845
rect 45359 37836 45371 37839
rect 43574 37808 45371 37836
rect 43574 37796 43580 37808
rect 45359 37805 45371 37808
rect 45405 37805 45417 37839
rect 45359 37799 45417 37805
rect 45448 37796 45454 37848
rect 45506 37836 45512 37848
rect 45543 37839 45601 37845
rect 45543 37836 45555 37839
rect 45506 37808 45555 37836
rect 45506 37796 45512 37808
rect 45543 37805 45555 37808
rect 45589 37836 45601 37839
rect 46828 37836 46834 37848
rect 45589 37808 46834 37836
rect 45589 37805 45601 37808
rect 45543 37799 45601 37805
rect 46828 37796 46834 37808
rect 46886 37796 46892 37848
rect 47306 37836 47334 37867
rect 47472 37864 47478 37876
rect 47530 37864 47536 37916
rect 50894 37904 50922 37944
rect 47950 37876 50922 37904
rect 50971 37907 51029 37913
rect 47950 37836 47978 37876
rect 48318 37845 48346 37876
rect 50971 37873 50983 37907
rect 51017 37904 51029 37907
rect 51244 37904 51250 37916
rect 51017 37876 51250 37904
rect 51017 37873 51029 37876
rect 50971 37867 51029 37873
rect 51244 37864 51250 37876
rect 51302 37864 51308 37916
rect 52274 37904 52302 37944
rect 53912 37932 53918 37984
rect 53970 37972 53976 37984
rect 60536 37972 60542 37984
rect 53970 37944 60542 37972
rect 53970 37932 53976 37944
rect 60536 37932 60542 37944
rect 60594 37932 60600 37984
rect 69000 37932 69006 37984
rect 69058 37972 69064 37984
rect 72591 37975 72649 37981
rect 72591 37972 72603 37975
rect 69058 37944 72603 37972
rect 69058 37932 69064 37944
rect 72591 37941 72603 37944
rect 72637 37972 72649 37975
rect 73048 37972 73054 37984
rect 72637 37944 73054 37972
rect 72637 37941 72649 37944
rect 72591 37935 72649 37941
rect 73048 37932 73054 37944
rect 73106 37972 73112 37984
rect 73784 37972 73790 37984
rect 73106 37944 73790 37972
rect 73106 37932 73112 37944
rect 73784 37932 73790 37944
rect 73842 37932 73848 37984
rect 82800 37972 82806 37984
rect 82634 37944 82806 37972
rect 52274 37876 56994 37904
rect 47306 37808 47978 37836
rect 48027 37839 48085 37845
rect 48027 37805 48039 37839
rect 48073 37805 48085 37839
rect 48027 37799 48085 37805
rect 48303 37839 48361 37845
rect 48303 37805 48315 37839
rect 48349 37805 48361 37839
rect 48484 37836 48490 37848
rect 48445 37808 48490 37836
rect 48303 37799 48361 37805
rect 40682 37740 45770 37768
rect 40391 37703 40449 37709
rect 40391 37700 40403 37703
rect 39894 37672 40403 37700
rect 39894 37660 39900 37672
rect 40391 37669 40403 37672
rect 40437 37669 40449 37703
rect 40391 37663 40449 37669
rect 40480 37660 40486 37712
rect 40538 37700 40544 37712
rect 41032 37700 41038 37712
rect 40538 37672 41038 37700
rect 40538 37660 40544 37672
rect 41032 37660 41038 37672
rect 41090 37660 41096 37712
rect 41216 37700 41222 37712
rect 41177 37672 41222 37700
rect 41216 37660 41222 37672
rect 41274 37660 41280 37712
rect 41768 37700 41774 37712
rect 41729 37672 41774 37700
rect 41768 37660 41774 37672
rect 41826 37660 41832 37712
rect 45359 37703 45417 37709
rect 45359 37669 45371 37703
rect 45405 37700 45417 37703
rect 45540 37700 45546 37712
rect 45405 37672 45546 37700
rect 45405 37669 45417 37672
rect 45359 37663 45417 37669
rect 45540 37660 45546 37672
rect 45598 37700 45604 37712
rect 45635 37703 45693 37709
rect 45635 37700 45647 37703
rect 45598 37672 45647 37700
rect 45598 37660 45604 37672
rect 45635 37669 45647 37672
rect 45681 37669 45693 37703
rect 45742 37700 45770 37740
rect 47380 37728 47386 37780
rect 47438 37768 47444 37780
rect 48042 37768 48070 37799
rect 48484 37796 48490 37808
rect 48542 37796 48548 37848
rect 51339 37839 51397 37845
rect 51339 37805 51351 37839
rect 51385 37836 51397 37839
rect 51888 37836 51894 37848
rect 51385 37808 51894 37836
rect 51385 37805 51397 37808
rect 51339 37799 51397 37805
rect 51888 37796 51894 37808
rect 51946 37796 51952 37848
rect 52075 37839 52133 37845
rect 52075 37805 52087 37839
rect 52121 37836 52133 37839
rect 52256 37836 52262 37848
rect 52121 37808 52262 37836
rect 52121 37805 52133 37808
rect 52075 37799 52133 37805
rect 52256 37796 52262 37808
rect 52314 37796 52320 37848
rect 54740 37796 54746 37848
rect 54798 37836 54804 37848
rect 54927 37839 54985 37845
rect 54927 37836 54939 37839
rect 54798 37808 54939 37836
rect 54798 37796 54804 37808
rect 54927 37805 54939 37808
rect 54973 37836 54985 37839
rect 55019 37839 55077 37845
rect 55019 37836 55031 37839
rect 54973 37808 55031 37836
rect 54973 37805 54985 37808
rect 54927 37799 54985 37805
rect 55019 37805 55031 37808
rect 55065 37836 55077 37839
rect 55200 37836 55206 37848
rect 55065 37808 55206 37836
rect 55065 37805 55077 37808
rect 55019 37799 55077 37805
rect 55200 37796 55206 37808
rect 55258 37796 55264 37848
rect 56307 37839 56365 37845
rect 56307 37805 56319 37839
rect 56353 37836 56365 37839
rect 56856 37836 56862 37848
rect 56353 37808 56862 37836
rect 56353 37805 56365 37808
rect 56307 37799 56365 37805
rect 56856 37796 56862 37808
rect 56914 37796 56920 37848
rect 55292 37768 55298 37780
rect 47438 37740 48070 37768
rect 52182 37740 55298 37768
rect 47438 37728 47444 37740
rect 52182 37700 52210 37740
rect 55292 37728 55298 37740
rect 55350 37728 55356 37780
rect 52348 37700 52354 37712
rect 45742 37672 52210 37700
rect 52309 37672 52354 37700
rect 45635 37663 45693 37669
rect 52348 37660 52354 37672
rect 52406 37660 52412 37712
rect 55016 37660 55022 37712
rect 55074 37700 55080 37712
rect 55203 37703 55261 37709
rect 55203 37700 55215 37703
rect 55074 37672 55215 37700
rect 55074 37660 55080 37672
rect 55203 37669 55215 37672
rect 55249 37669 55261 37703
rect 56120 37700 56126 37712
rect 56081 37672 56126 37700
rect 55203 37663 55261 37669
rect 56120 37660 56126 37672
rect 56178 37660 56184 37712
rect 56874 37700 56902 37796
rect 56966 37768 56994 37876
rect 57132 37864 57138 37916
rect 57190 37904 57196 37916
rect 57684 37904 57690 37916
rect 57190 37876 57690 37904
rect 57190 37864 57196 37876
rect 57684 37864 57690 37876
rect 57742 37904 57748 37916
rect 58239 37907 58297 37913
rect 58239 37904 58251 37907
rect 57742 37876 58251 37904
rect 57742 37864 57748 37876
rect 58239 37873 58251 37876
rect 58285 37873 58297 37907
rect 58239 37867 58297 37873
rect 59527 37907 59585 37913
rect 59527 37873 59539 37907
rect 59573 37904 59585 37907
rect 60628 37904 60634 37916
rect 59573 37876 60634 37904
rect 59573 37873 59585 37876
rect 59527 37867 59585 37873
rect 60628 37864 60634 37876
rect 60686 37864 60692 37916
rect 67988 37904 67994 37916
rect 60738 37876 62790 37904
rect 67949 37876 67994 37904
rect 57871 37839 57929 37845
rect 57871 37805 57883 37839
rect 57917 37836 57929 37839
rect 58052 37836 58058 37848
rect 57917 37808 58058 37836
rect 57917 37805 57929 37808
rect 57871 37799 57929 37805
rect 58052 37796 58058 37808
rect 58110 37796 58116 37848
rect 58144 37796 58150 37848
rect 58202 37836 58208 37848
rect 58377 37839 58435 37845
rect 58377 37836 58389 37839
rect 58202 37808 58389 37836
rect 58202 37796 58208 37808
rect 58377 37805 58389 37808
rect 58423 37836 58435 37839
rect 58880 37836 58886 37848
rect 58423 37808 58886 37836
rect 58423 37805 58435 37808
rect 58377 37799 58435 37805
rect 58880 37796 58886 37808
rect 58938 37836 58944 37848
rect 58975 37839 59033 37845
rect 58975 37836 58987 37839
rect 58938 37808 58987 37836
rect 58938 37796 58944 37808
rect 58975 37805 58987 37808
rect 59021 37805 59033 37839
rect 58975 37799 59033 37805
rect 59064 37796 59070 37848
rect 59122 37836 59128 37848
rect 59159 37839 59217 37845
rect 59159 37836 59171 37839
rect 59122 37808 59171 37836
rect 59122 37796 59128 37808
rect 59159 37805 59171 37808
rect 59205 37805 59217 37839
rect 59159 37799 59217 37805
rect 59432 37796 59438 37848
rect 59490 37836 59496 37848
rect 60738 37836 60766 37876
rect 59490 37808 60766 37836
rect 61275 37839 61333 37845
rect 59490 37796 59496 37808
rect 61275 37805 61287 37839
rect 61321 37836 61333 37839
rect 61732 37836 61738 37848
rect 61321 37808 61738 37836
rect 61321 37805 61333 37808
rect 61275 37799 61333 37805
rect 61732 37796 61738 37808
rect 61790 37796 61796 37848
rect 62100 37796 62106 37848
rect 62158 37836 62164 37848
rect 62379 37839 62437 37845
rect 62379 37836 62391 37839
rect 62158 37808 62391 37836
rect 62158 37796 62164 37808
rect 62379 37805 62391 37808
rect 62425 37805 62437 37839
rect 62379 37799 62437 37805
rect 62468 37796 62474 37848
rect 62526 37836 62532 37848
rect 62655 37839 62713 37845
rect 62655 37836 62667 37839
rect 62526 37808 62667 37836
rect 62526 37796 62532 37808
rect 62655 37805 62667 37808
rect 62701 37805 62713 37839
rect 62762 37836 62790 37876
rect 67988 37864 67994 37876
rect 68046 37864 68052 37916
rect 68264 37904 68270 37916
rect 68225 37876 68270 37904
rect 68264 37864 68270 37876
rect 68322 37864 68328 37916
rect 69831 37907 69889 37913
rect 69831 37873 69843 37907
rect 69877 37904 69889 37907
rect 69920 37904 69926 37916
rect 69877 37876 69926 37904
rect 69877 37873 69889 37876
rect 69831 37867 69889 37873
rect 69920 37864 69926 37876
rect 69978 37864 69984 37916
rect 74063 37907 74121 37913
rect 74063 37873 74075 37907
rect 74109 37873 74121 37907
rect 76636 37904 76642 37916
rect 74063 37867 74121 37873
rect 76286 37876 76642 37904
rect 72407 37839 72465 37845
rect 72407 37836 72419 37839
rect 62762 37808 72419 37836
rect 62655 37799 62713 37805
rect 72407 37805 72419 37808
rect 72453 37805 72465 37839
rect 73968 37836 73974 37848
rect 73929 37808 73974 37836
rect 72407 37799 72465 37805
rect 56966 37740 62514 37768
rect 57687 37703 57745 37709
rect 57687 37700 57699 37703
rect 56874 37672 57699 37700
rect 57687 37669 57699 37672
rect 57733 37669 57745 37703
rect 58052 37700 58058 37712
rect 58013 37672 58058 37700
rect 57687 37663 57745 37669
rect 58052 37660 58058 37672
rect 58110 37660 58116 37712
rect 59064 37660 59070 37712
rect 59122 37700 59128 37712
rect 59711 37703 59769 37709
rect 59711 37700 59723 37703
rect 59122 37672 59723 37700
rect 59122 37660 59128 37672
rect 59711 37669 59723 37672
rect 59757 37700 59769 37703
rect 61364 37700 61370 37712
rect 59757 37672 61370 37700
rect 59757 37669 59769 37672
rect 59711 37663 59769 37669
rect 61364 37660 61370 37672
rect 61422 37660 61428 37712
rect 62100 37700 62106 37712
rect 62061 37672 62106 37700
rect 62100 37660 62106 37672
rect 62158 37660 62164 37712
rect 62486 37700 62514 37740
rect 63314 37740 64998 37768
rect 63314 37700 63342 37740
rect 63756 37700 63762 37712
rect 62486 37672 63342 37700
rect 63717 37672 63762 37700
rect 63756 37660 63762 37672
rect 63814 37660 63820 37712
rect 64970 37700 64998 37740
rect 72220 37700 72226 37712
rect 64970 37672 72226 37700
rect 72220 37660 72226 37672
rect 72278 37660 72284 37712
rect 72315 37703 72373 37709
rect 72315 37669 72327 37703
rect 72361 37700 72373 37703
rect 72422 37700 72450 37799
rect 73968 37796 73974 37808
rect 74026 37796 74032 37848
rect 72772 37728 72778 37780
rect 72830 37768 72836 37780
rect 73876 37768 73882 37780
rect 72830 37740 73882 37768
rect 72830 37728 72836 37740
rect 73876 37728 73882 37740
rect 73934 37768 73940 37780
rect 74078 37768 74106 37867
rect 74152 37796 74158 37848
rect 74210 37836 74216 37848
rect 74247 37839 74305 37845
rect 74247 37836 74259 37839
rect 74210 37808 74259 37836
rect 74210 37796 74216 37808
rect 74247 37805 74259 37808
rect 74293 37805 74305 37839
rect 74704 37836 74710 37848
rect 74665 37808 74710 37836
rect 74247 37799 74305 37805
rect 74704 37796 74710 37808
rect 74762 37796 74768 37848
rect 74799 37839 74857 37845
rect 74799 37805 74811 37839
rect 74845 37805 74857 37839
rect 74799 37799 74857 37805
rect 73934 37740 74106 37768
rect 73934 37728 73940 37740
rect 74060 37700 74066 37712
rect 72361 37672 74066 37700
rect 72361 37669 72373 37672
rect 72315 37663 72373 37669
rect 74060 37660 74066 37672
rect 74118 37660 74124 37712
rect 74152 37660 74158 37712
rect 74210 37700 74216 37712
rect 74814 37700 74842 37799
rect 74980 37796 74986 37848
rect 75038 37836 75044 37848
rect 76286 37836 76314 37876
rect 76636 37864 76642 37876
rect 76694 37864 76700 37916
rect 76820 37864 76826 37916
rect 76878 37904 76884 37916
rect 77924 37904 77930 37916
rect 76878 37876 77930 37904
rect 76878 37864 76884 37876
rect 77924 37864 77930 37876
rect 77982 37904 77988 37916
rect 82634 37913 82662 37944
rect 82800 37932 82806 37944
rect 82858 37932 82864 37984
rect 79307 37907 79365 37913
rect 79307 37904 79319 37907
rect 77982 37876 79319 37904
rect 77982 37864 77988 37876
rect 79307 37873 79319 37876
rect 79353 37873 79365 37907
rect 79307 37867 79365 37873
rect 82619 37907 82677 37913
rect 82619 37873 82631 37907
rect 82665 37873 82677 37907
rect 85100 37904 85106 37916
rect 85061 37876 85106 37904
rect 82619 37867 82677 37873
rect 85100 37864 85106 37876
rect 85158 37864 85164 37916
rect 88596 37904 88602 37916
rect 88557 37876 88602 37904
rect 88596 37864 88602 37876
rect 88654 37864 88660 37916
rect 89059 37907 89117 37913
rect 89059 37873 89071 37907
rect 89105 37904 89117 37907
rect 89516 37904 89522 37916
rect 89105 37876 89522 37904
rect 89105 37873 89117 37876
rect 89059 37867 89117 37873
rect 89516 37864 89522 37876
rect 89574 37864 89580 37916
rect 90178 37904 90206 38000
rect 90439 37907 90497 37913
rect 90439 37904 90451 37907
rect 90178 37876 90451 37904
rect 90439 37873 90451 37876
rect 90485 37873 90497 37907
rect 90439 37867 90497 37873
rect 76452 37836 76458 37848
rect 75038 37808 76314 37836
rect 76413 37808 76458 37836
rect 75038 37796 75044 37808
rect 76452 37796 76458 37808
rect 76510 37796 76516 37848
rect 79212 37836 79218 37848
rect 79173 37808 79218 37836
rect 79212 37796 79218 37808
rect 79270 37796 79276 37848
rect 82156 37796 82162 37848
rect 82214 37836 82220 37848
rect 82711 37839 82769 37845
rect 82711 37836 82723 37839
rect 82214 37808 82723 37836
rect 82214 37796 82220 37808
rect 82711 37805 82723 37808
rect 82757 37836 82769 37839
rect 83263 37839 83321 37845
rect 83263 37836 83275 37839
rect 82757 37808 83275 37836
rect 82757 37805 82769 37808
rect 82711 37799 82769 37805
rect 83263 37805 83275 37808
rect 83309 37805 83321 37839
rect 83263 37799 83321 37805
rect 83447 37839 83505 37845
rect 83447 37805 83459 37839
rect 83493 37836 83505 37839
rect 84643 37839 84701 37845
rect 83493 37808 83582 37836
rect 83493 37805 83505 37808
rect 83447 37799 83505 37805
rect 75348 37768 75354 37780
rect 75309 37740 75354 37768
rect 75348 37728 75354 37740
rect 75406 37728 75412 37780
rect 74210 37672 74842 37700
rect 76271 37703 76329 37709
rect 74210 37660 74216 37672
rect 76271 37669 76283 37703
rect 76317 37700 76329 37703
rect 76360 37700 76366 37712
rect 76317 37672 76366 37700
rect 76317 37669 76329 37672
rect 76271 37663 76329 37669
rect 76360 37660 76366 37672
rect 76418 37660 76424 37712
rect 76728 37660 76734 37712
rect 76786 37700 76792 37712
rect 83554 37700 83582 37808
rect 84643 37805 84655 37839
rect 84689 37836 84701 37839
rect 84827 37839 84885 37845
rect 84827 37836 84839 37839
rect 84689 37808 84839 37836
rect 84689 37805 84701 37808
rect 84643 37799 84701 37805
rect 84827 37805 84839 37808
rect 84873 37836 84885 37839
rect 84916 37836 84922 37848
rect 84873 37808 84922 37836
rect 84873 37805 84885 37808
rect 84827 37799 84885 37805
rect 84916 37796 84922 37808
rect 84974 37796 84980 37848
rect 88504 37796 88510 37848
rect 88562 37836 88568 37848
rect 88967 37839 89025 37845
rect 88967 37836 88979 37839
rect 88562 37808 88979 37836
rect 88562 37796 88568 37808
rect 88967 37805 88979 37808
rect 89013 37805 89025 37839
rect 88967 37799 89025 37805
rect 89335 37839 89393 37845
rect 89335 37805 89347 37839
rect 89381 37805 89393 37839
rect 89335 37799 89393 37805
rect 89427 37839 89485 37845
rect 89427 37805 89439 37839
rect 89473 37836 89485 37839
rect 89884 37836 89890 37848
rect 89473 37808 89890 37836
rect 89473 37805 89485 37808
rect 89427 37799 89485 37805
rect 83815 37771 83873 37777
rect 83815 37737 83827 37771
rect 83861 37768 83873 37771
rect 84272 37768 84278 37780
rect 83861 37740 84278 37768
rect 83861 37737 83873 37740
rect 83815 37731 83873 37737
rect 84272 37728 84278 37740
rect 84330 37728 84336 37780
rect 86572 37728 86578 37780
rect 86630 37768 86636 37780
rect 89240 37768 89246 37780
rect 86630 37740 89246 37768
rect 86630 37728 86636 37740
rect 89240 37728 89246 37740
rect 89298 37768 89304 37780
rect 89350 37768 89378 37799
rect 89884 37796 89890 37808
rect 89942 37836 89948 37848
rect 90344 37836 90350 37848
rect 89942 37808 90350 37836
rect 89942 37796 89948 37808
rect 90344 37796 90350 37808
rect 90402 37796 90408 37848
rect 90712 37836 90718 37848
rect 90673 37808 90718 37836
rect 90712 37796 90718 37808
rect 90770 37796 90776 37848
rect 89298 37740 89378 37768
rect 89298 37728 89304 37740
rect 83996 37700 84002 37712
rect 76786 37672 84002 37700
rect 76786 37660 76792 37672
rect 83996 37660 84002 37672
rect 84054 37660 84060 37712
rect 91356 37660 91362 37712
rect 91414 37700 91420 37712
rect 91819 37703 91877 37709
rect 91819 37700 91831 37703
rect 91414 37672 91831 37700
rect 91414 37660 91420 37672
rect 91819 37669 91831 37672
rect 91865 37669 91877 37703
rect 91819 37663 91877 37669
rect 538 37610 93642 37632
rect 538 37558 6344 37610
rect 6396 37558 6408 37610
rect 6460 37558 6472 37610
rect 6524 37558 6536 37610
rect 6588 37558 11672 37610
rect 11724 37558 11736 37610
rect 11788 37558 11800 37610
rect 11852 37558 11864 37610
rect 11916 37558 17000 37610
rect 17052 37558 17064 37610
rect 17116 37558 17128 37610
rect 17180 37558 17192 37610
rect 17244 37558 22328 37610
rect 22380 37558 22392 37610
rect 22444 37558 22456 37610
rect 22508 37558 22520 37610
rect 22572 37558 27656 37610
rect 27708 37558 27720 37610
rect 27772 37558 27784 37610
rect 27836 37558 27848 37610
rect 27900 37558 32984 37610
rect 33036 37558 33048 37610
rect 33100 37558 33112 37610
rect 33164 37558 33176 37610
rect 33228 37558 38312 37610
rect 38364 37558 38376 37610
rect 38428 37558 38440 37610
rect 38492 37558 38504 37610
rect 38556 37558 43640 37610
rect 43692 37558 43704 37610
rect 43756 37558 43768 37610
rect 43820 37558 43832 37610
rect 43884 37558 48968 37610
rect 49020 37558 49032 37610
rect 49084 37558 49096 37610
rect 49148 37558 49160 37610
rect 49212 37558 54296 37610
rect 54348 37558 54360 37610
rect 54412 37558 54424 37610
rect 54476 37558 54488 37610
rect 54540 37558 59624 37610
rect 59676 37558 59688 37610
rect 59740 37558 59752 37610
rect 59804 37558 59816 37610
rect 59868 37558 64952 37610
rect 65004 37558 65016 37610
rect 65068 37558 65080 37610
rect 65132 37558 65144 37610
rect 65196 37558 70280 37610
rect 70332 37558 70344 37610
rect 70396 37558 70408 37610
rect 70460 37558 70472 37610
rect 70524 37558 75608 37610
rect 75660 37558 75672 37610
rect 75724 37558 75736 37610
rect 75788 37558 75800 37610
rect 75852 37558 80936 37610
rect 80988 37558 81000 37610
rect 81052 37558 81064 37610
rect 81116 37558 81128 37610
rect 81180 37558 86264 37610
rect 86316 37558 86328 37610
rect 86380 37558 86392 37610
rect 86444 37558 86456 37610
rect 86508 37558 91592 37610
rect 91644 37558 91656 37610
rect 91708 37558 91720 37610
rect 91772 37558 91784 37610
rect 91836 37558 93642 37610
rect 538 37536 93642 37558
rect 3128 37456 3134 37508
rect 3186 37496 3192 37508
rect 3956 37496 3962 37508
rect 3186 37468 3962 37496
rect 3186 37456 3192 37468
rect 3956 37456 3962 37468
rect 4014 37496 4020 37508
rect 5888 37496 5894 37508
rect 4014 37468 5894 37496
rect 4014 37456 4020 37468
rect 4158 37369 4186 37468
rect 5888 37456 5894 37468
rect 5946 37496 5952 37508
rect 5983 37499 6041 37505
rect 5983 37496 5995 37499
rect 5946 37468 5995 37496
rect 5946 37456 5952 37468
rect 5983 37465 5995 37468
rect 6029 37496 6041 37499
rect 7452 37496 7458 37508
rect 6029 37468 7458 37496
rect 6029 37465 6041 37468
rect 5983 37459 6041 37465
rect 7452 37456 7458 37468
rect 7510 37456 7516 37508
rect 10304 37456 10310 37508
rect 10362 37496 10368 37508
rect 10399 37499 10457 37505
rect 10399 37496 10411 37499
rect 10362 37468 10411 37496
rect 10362 37456 10368 37468
rect 10399 37465 10411 37468
rect 10445 37465 10457 37499
rect 10399 37459 10457 37465
rect 10488 37456 10494 37508
rect 10546 37496 10552 37508
rect 12423 37499 12481 37505
rect 10546 37468 11270 37496
rect 10546 37456 10552 37468
rect 7636 37388 7642 37440
rect 7694 37428 7700 37440
rect 11242 37428 11270 37468
rect 12423 37465 12435 37499
rect 12469 37496 12481 37499
rect 12788 37496 12794 37508
rect 12469 37468 12794 37496
rect 12469 37465 12481 37468
rect 12423 37459 12481 37465
rect 12788 37456 12794 37468
rect 12846 37456 12852 37508
rect 19412 37456 19418 37508
rect 19470 37496 19476 37508
rect 27048 37496 27054 37508
rect 19470 37468 27054 37496
rect 19470 37456 19476 37468
rect 27048 37456 27054 37468
rect 27106 37456 27112 37508
rect 27232 37496 27238 37508
rect 27193 37468 27238 37496
rect 27232 37456 27238 37468
rect 27290 37456 27296 37508
rect 28888 37456 28894 37508
rect 28946 37496 28952 37508
rect 31927 37499 31985 37505
rect 31927 37496 31939 37499
rect 28946 37468 31939 37496
rect 28946 37456 28952 37468
rect 31927 37465 31939 37468
rect 31973 37465 31985 37499
rect 32108 37496 32114 37508
rect 32069 37468 32114 37496
rect 31927 37459 31985 37465
rect 32108 37456 32114 37468
rect 32166 37456 32172 37508
rect 33583 37499 33641 37505
rect 33583 37496 33595 37499
rect 33138 37468 33595 37496
rect 12052 37428 12058 37440
rect 7694 37400 11178 37428
rect 7694 37388 7700 37400
rect 4143 37363 4201 37369
rect 4143 37329 4155 37363
rect 4189 37329 4201 37363
rect 4416 37360 4422 37372
rect 4377 37332 4422 37360
rect 4143 37323 4201 37329
rect 4416 37320 4422 37332
rect 4474 37320 4480 37372
rect 10764 37360 10770 37372
rect 10725 37332 10770 37360
rect 10764 37320 10770 37332
rect 10822 37320 10828 37372
rect 11150 37369 11178 37400
rect 11242 37400 12058 37428
rect 11242 37369 11270 37400
rect 12052 37388 12058 37400
rect 12110 37428 12116 37440
rect 14168 37428 14174 37440
rect 12110 37400 12742 37428
rect 12110 37388 12116 37400
rect 11135 37363 11193 37369
rect 11135 37329 11147 37363
rect 11181 37329 11193 37363
rect 11135 37323 11193 37329
rect 11227 37363 11285 37369
rect 11227 37329 11239 37363
rect 11273 37329 11285 37363
rect 11227 37323 11285 37329
rect 11500 37320 11506 37372
rect 11558 37360 11564 37372
rect 12607 37363 12665 37369
rect 12607 37360 12619 37363
rect 11558 37332 12619 37360
rect 11558 37320 11564 37332
rect 12607 37329 12619 37332
rect 12653 37329 12665 37363
rect 12607 37323 12665 37329
rect 10859 37295 10917 37301
rect 10859 37261 10871 37295
rect 10905 37292 10917 37295
rect 11518 37292 11546 37320
rect 10905 37264 11546 37292
rect 12714 37292 12742 37400
rect 12806 37400 14174 37428
rect 12806 37369 12834 37400
rect 14168 37388 14174 37400
rect 14226 37388 14232 37440
rect 15643 37431 15701 37437
rect 15643 37397 15655 37431
rect 15689 37428 15701 37431
rect 16008 37428 16014 37440
rect 15689 37400 16014 37428
rect 15689 37397 15701 37400
rect 15643 37391 15701 37397
rect 16008 37388 16014 37400
rect 16066 37388 16072 37440
rect 16195 37431 16253 37437
rect 16195 37397 16207 37431
rect 16241 37428 16253 37431
rect 17664 37428 17670 37440
rect 16241 37400 17670 37428
rect 16241 37397 16253 37400
rect 16195 37391 16253 37397
rect 17664 37388 17670 37400
rect 17722 37388 17728 37440
rect 27508 37388 27514 37440
rect 27566 37428 27572 37440
rect 28906 37428 28934 37456
rect 27566 37400 28934 37428
rect 27566 37388 27572 37400
rect 12791 37363 12849 37369
rect 12791 37329 12803 37363
rect 12837 37329 12849 37363
rect 12791 37323 12849 37329
rect 13159 37363 13217 37369
rect 13159 37329 13171 37363
rect 13205 37329 13217 37363
rect 15824 37360 15830 37372
rect 15785 37332 15830 37360
rect 13159 37323 13217 37329
rect 13067 37295 13125 37301
rect 13067 37292 13079 37295
rect 12714 37264 13079 37292
rect 10905 37261 10917 37264
rect 10859 37255 10917 37261
rect 13067 37261 13079 37264
rect 13113 37261 13125 37295
rect 13067 37255 13125 37261
rect 5707 37227 5765 37233
rect 5707 37193 5719 37227
rect 5753 37224 5765 37227
rect 13174 37224 13202 37323
rect 15824 37320 15830 37332
rect 15882 37320 15888 37372
rect 17204 37360 17210 37372
rect 17165 37332 17210 37360
rect 17204 37320 17210 37332
rect 17262 37320 17268 37372
rect 17299 37363 17357 37369
rect 17299 37329 17311 37363
rect 17345 37329 17357 37363
rect 17299 37323 17357 37329
rect 20151 37363 20209 37369
rect 20151 37329 20163 37363
rect 20197 37360 20209 37363
rect 20335 37363 20393 37369
rect 20335 37360 20347 37363
rect 20197 37332 20347 37360
rect 20197 37329 20209 37332
rect 20151 37323 20209 37329
rect 20335 37329 20347 37332
rect 20381 37360 20393 37363
rect 20884 37360 20890 37372
rect 20381 37332 20890 37360
rect 20381 37329 20393 37332
rect 20335 37323 20393 37329
rect 16468 37252 16474 37304
rect 16526 37292 16532 37304
rect 17314 37292 17342 37323
rect 20884 37320 20890 37332
rect 20942 37320 20948 37372
rect 27416 37320 27422 37372
rect 27474 37360 27480 37372
rect 27986 37369 28014 37400
rect 32752 37388 32758 37440
rect 32810 37428 32816 37440
rect 32810 37400 33074 37428
rect 32810 37388 32816 37400
rect 27603 37363 27661 37369
rect 27603 37360 27615 37363
rect 27474 37332 27615 37360
rect 27474 37320 27480 37332
rect 27603 37329 27615 37332
rect 27649 37329 27661 37363
rect 27603 37323 27661 37329
rect 27971 37363 28029 37369
rect 27971 37329 27983 37363
rect 28017 37329 28029 37363
rect 27971 37323 28029 37329
rect 28155 37363 28213 37369
rect 28155 37329 28167 37363
rect 28201 37360 28213 37363
rect 28796 37360 28802 37372
rect 28201 37332 28802 37360
rect 28201 37329 28213 37332
rect 28155 37323 28213 37329
rect 28796 37320 28802 37332
rect 28854 37320 28860 37372
rect 29443 37363 29501 37369
rect 29443 37329 29455 37363
rect 29489 37360 29501 37363
rect 29489 37332 29523 37360
rect 29489 37329 29501 37332
rect 29443 37323 29501 37329
rect 16526 37264 17342 37292
rect 20611 37295 20669 37301
rect 16526 37252 16532 37264
rect 20611 37261 20623 37295
rect 20657 37292 20669 37295
rect 21344 37292 21350 37304
rect 20657 37264 21350 37292
rect 20657 37261 20669 37264
rect 20611 37255 20669 37261
rect 21344 37252 21350 37264
rect 21402 37252 21408 37304
rect 27692 37252 27698 37304
rect 27750 37292 27756 37304
rect 29351 37295 29409 37301
rect 27750 37264 27795 37292
rect 27750 37252 27756 37264
rect 29351 37261 29363 37295
rect 29397 37292 29409 37295
rect 29458 37292 29486 37323
rect 31924 37320 31930 37372
rect 31982 37360 31988 37372
rect 32660 37360 32666 37372
rect 31982 37332 32666 37360
rect 31982 37320 31988 37332
rect 32660 37320 32666 37332
rect 32718 37320 32724 37372
rect 33046 37369 33074 37400
rect 33031 37363 33089 37369
rect 33031 37329 33043 37363
rect 33077 37329 33089 37363
rect 33031 37323 33089 37329
rect 29808 37292 29814 37304
rect 29397 37264 29814 37292
rect 29397 37261 29409 37264
rect 29351 37255 29409 37261
rect 29808 37252 29814 37264
rect 29866 37252 29872 37304
rect 32755 37295 32813 37301
rect 32755 37261 32767 37295
rect 32801 37292 32813 37295
rect 33138 37292 33166 37468
rect 33583 37465 33595 37468
rect 33629 37496 33641 37499
rect 35052 37496 35058 37508
rect 33629 37468 35058 37496
rect 33629 37465 33641 37468
rect 33583 37459 33641 37465
rect 35052 37456 35058 37468
rect 35110 37456 35116 37508
rect 35144 37456 35150 37508
rect 35202 37496 35208 37508
rect 37720 37496 37726 37508
rect 35202 37468 37726 37496
rect 35202 37456 35208 37468
rect 37720 37456 37726 37468
rect 37778 37456 37784 37508
rect 40480 37496 40486 37508
rect 37830 37468 40486 37496
rect 36616 37388 36622 37440
rect 36674 37428 36680 37440
rect 36674 37400 37490 37428
rect 36674 37388 36680 37400
rect 33215 37363 33273 37369
rect 33215 37329 33227 37363
rect 33261 37360 33273 37363
rect 33261 37332 33442 37360
rect 33261 37329 33273 37332
rect 33215 37323 33273 37329
rect 32801 37264 33166 37292
rect 32801 37261 32813 37264
rect 32755 37255 32813 37261
rect 5753 37196 13202 37224
rect 17023 37227 17081 37233
rect 5753 37193 5765 37196
rect 5707 37187 5765 37193
rect 17023 37193 17035 37227
rect 17069 37224 17081 37227
rect 17572 37224 17578 37236
rect 17069 37196 17578 37224
rect 17069 37193 17081 37196
rect 17023 37187 17081 37193
rect 17572 37184 17578 37196
rect 17630 37184 17636 37236
rect 31927 37227 31985 37233
rect 31927 37193 31939 37227
rect 31973 37224 31985 37227
rect 32660 37224 32666 37236
rect 31973 37196 32666 37224
rect 31973 37193 31985 37196
rect 31927 37187 31985 37193
rect 32660 37184 32666 37196
rect 32718 37184 32724 37236
rect 33414 37233 33442 37332
rect 34960 37320 34966 37372
rect 35018 37360 35024 37372
rect 37462 37369 37490 37400
rect 37355 37363 37413 37369
rect 37355 37360 37367 37363
rect 35018 37332 37367 37360
rect 35018 37320 35024 37332
rect 37355 37329 37367 37332
rect 37401 37329 37413 37363
rect 37355 37323 37413 37329
rect 37447 37363 37505 37369
rect 37447 37329 37459 37363
rect 37493 37360 37505 37363
rect 37830 37360 37858 37468
rect 40480 37456 40486 37468
rect 40538 37456 40544 37508
rect 47380 37496 47386 37508
rect 40774 37468 47386 37496
rect 37996 37388 38002 37440
rect 38054 37428 38060 37440
rect 38054 37400 38134 37428
rect 38054 37388 38060 37400
rect 37493 37332 37858 37360
rect 37493 37329 37505 37332
rect 37447 37323 37505 37329
rect 37904 37320 37910 37372
rect 37962 37360 37968 37372
rect 38106 37369 38134 37400
rect 40296 37388 40302 37440
rect 40354 37428 40360 37440
rect 40575 37431 40633 37437
rect 40575 37428 40587 37431
rect 40354 37400 40587 37428
rect 40354 37388 40360 37400
rect 40575 37397 40587 37400
rect 40621 37397 40633 37431
rect 40575 37391 40633 37397
rect 38091 37363 38149 37369
rect 37962 37332 38007 37360
rect 37962 37320 37968 37332
rect 38091 37329 38103 37363
rect 38137 37360 38149 37363
rect 39195 37363 39253 37369
rect 39195 37360 39207 37363
rect 38137 37332 39207 37360
rect 38137 37329 38149 37332
rect 38091 37323 38149 37329
rect 39195 37329 39207 37332
rect 39241 37329 39253 37363
rect 39195 37323 39253 37329
rect 39284 37320 39290 37372
rect 39342 37360 39348 37372
rect 39471 37363 39529 37369
rect 39471 37360 39483 37363
rect 39342 37332 39483 37360
rect 39342 37320 39348 37332
rect 39471 37329 39483 37332
rect 39517 37329 39529 37363
rect 39471 37323 39529 37329
rect 39744 37320 39750 37372
rect 39802 37360 39808 37372
rect 40207 37363 40265 37369
rect 40207 37360 40219 37363
rect 39802 37332 40219 37360
rect 39802 37320 39808 37332
rect 40207 37329 40219 37332
rect 40253 37360 40265 37363
rect 40774 37360 40802 37468
rect 40253 37332 40802 37360
rect 41127 37363 41185 37369
rect 40253 37329 40265 37332
rect 40207 37323 40265 37329
rect 41127 37329 41139 37363
rect 41173 37360 41185 37363
rect 41326 37360 41354 37468
rect 47380 37456 47386 37468
rect 47438 37456 47444 37508
rect 48484 37456 48490 37508
rect 48542 37496 48548 37508
rect 48542 37468 55154 37496
rect 48542 37456 48548 37468
rect 41418 37400 46874 37428
rect 41418 37369 41446 37400
rect 41173 37332 41354 37360
rect 41403 37363 41461 37369
rect 41173 37329 41185 37332
rect 41127 37323 41185 37329
rect 41403 37329 41415 37363
rect 41449 37329 41461 37363
rect 41403 37323 41461 37329
rect 40480 37292 40486 37304
rect 40393 37264 40486 37292
rect 40480 37252 40486 37264
rect 40538 37292 40544 37304
rect 41418 37292 41446 37323
rect 42136 37320 42142 37372
rect 42194 37360 42200 37372
rect 42967 37363 43025 37369
rect 42967 37360 42979 37363
rect 42194 37332 42979 37360
rect 42194 37320 42200 37332
rect 42967 37329 42979 37332
rect 43013 37360 43025 37363
rect 43519 37363 43577 37369
rect 43519 37360 43531 37363
rect 43013 37332 43531 37360
rect 43013 37329 43025 37332
rect 42967 37323 43025 37329
rect 43519 37329 43531 37332
rect 43565 37329 43577 37363
rect 43519 37323 43577 37329
rect 43608 37320 43614 37372
rect 43666 37360 43672 37372
rect 43703 37363 43761 37369
rect 43703 37360 43715 37363
rect 43666 37332 43715 37360
rect 43666 37320 43672 37332
rect 43703 37329 43715 37332
rect 43749 37360 43761 37363
rect 44347 37363 44405 37369
rect 44347 37360 44359 37363
rect 43749 37332 44359 37360
rect 43749 37329 43761 37332
rect 43703 37323 43761 37329
rect 44347 37329 44359 37332
rect 44393 37360 44405 37363
rect 45080 37360 45086 37372
rect 44393 37332 45086 37360
rect 44393 37329 44405 37332
rect 44347 37323 44405 37329
rect 45080 37320 45086 37332
rect 45138 37320 45144 37372
rect 45356 37360 45362 37372
rect 45317 37332 45362 37360
rect 45356 37320 45362 37332
rect 45414 37360 45420 37372
rect 46371 37363 46429 37369
rect 45414 37332 46322 37360
rect 45414 37320 45420 37332
rect 40538 37264 41446 37292
rect 41587 37295 41645 37301
rect 40538 37252 40544 37264
rect 41587 37261 41599 37295
rect 41633 37292 41645 37295
rect 41679 37295 41737 37301
rect 41679 37292 41691 37295
rect 41633 37264 41691 37292
rect 41633 37261 41645 37264
rect 41587 37255 41645 37261
rect 41679 37261 41691 37264
rect 41725 37261 41737 37295
rect 42872 37292 42878 37304
rect 42833 37264 42878 37292
rect 41679 37255 41737 37261
rect 33399 37227 33457 37233
rect 33399 37193 33411 37227
rect 33445 37224 33457 37227
rect 37996 37224 38002 37236
rect 33445 37196 38002 37224
rect 33445 37193 33457 37196
rect 33399 37187 33457 37193
rect 37996 37184 38002 37196
rect 38054 37184 38060 37236
rect 38088 37184 38094 37236
rect 38146 37224 38152 37236
rect 38275 37227 38333 37233
rect 38275 37224 38287 37227
rect 38146 37196 38287 37224
rect 38146 37184 38152 37196
rect 38275 37193 38287 37196
rect 38321 37193 38333 37227
rect 38275 37187 38333 37193
rect 38735 37227 38793 37233
rect 38735 37193 38747 37227
rect 38781 37224 38793 37227
rect 39195 37227 39253 37233
rect 39195 37224 39207 37227
rect 38781 37196 39207 37224
rect 38781 37193 38793 37196
rect 38735 37187 38793 37193
rect 39195 37193 39207 37196
rect 39241 37224 39253 37227
rect 39468 37224 39474 37236
rect 39241 37196 39474 37224
rect 39241 37193 39253 37196
rect 39195 37187 39253 37193
rect 39468 37184 39474 37196
rect 39526 37184 39532 37236
rect 41694 37224 41722 37255
rect 42872 37252 42878 37264
rect 42930 37252 42936 37304
rect 46187 37295 46245 37301
rect 46187 37292 46199 37295
rect 45558 37264 46199 37292
rect 43056 37224 43062 37236
rect 41694 37196 43062 37224
rect 43056 37184 43062 37196
rect 43114 37184 43120 37236
rect 17388 37116 17394 37168
rect 17446 37156 17452 37168
rect 17483 37159 17541 37165
rect 17483 37156 17495 37159
rect 17446 37128 17495 37156
rect 17446 37116 17452 37128
rect 17483 37125 17495 37128
rect 17529 37125 17541 37159
rect 17483 37119 17541 37125
rect 21528 37116 21534 37168
rect 21586 37156 21592 37168
rect 21715 37159 21773 37165
rect 21715 37156 21727 37159
rect 21586 37128 21727 37156
rect 21586 37116 21592 37128
rect 21715 37125 21727 37128
rect 21761 37125 21773 37159
rect 29624 37156 29630 37168
rect 29585 37128 29630 37156
rect 21715 37119 21773 37125
rect 29624 37116 29630 37128
rect 29682 37116 29688 37168
rect 29808 37116 29814 37168
rect 29866 37156 29872 37168
rect 39100 37156 39106 37168
rect 29866 37128 39106 37156
rect 29866 37116 29872 37128
rect 39100 37116 39106 37128
rect 39158 37116 39164 37168
rect 39284 37156 39290 37168
rect 39245 37128 39290 37156
rect 39284 37116 39290 37128
rect 39342 37116 39348 37168
rect 39655 37159 39713 37165
rect 39655 37125 39667 37159
rect 39701 37156 39713 37159
rect 39836 37156 39842 37168
rect 39701 37128 39842 37156
rect 39701 37125 39713 37128
rect 39655 37119 39713 37125
rect 39836 37116 39842 37128
rect 39894 37116 39900 37168
rect 40388 37116 40394 37168
rect 40446 37156 40452 37168
rect 42136 37156 42142 37168
rect 40446 37128 42142 37156
rect 40446 37116 40452 37128
rect 42136 37116 42142 37128
rect 42194 37116 42200 37168
rect 43979 37159 44037 37165
rect 43979 37125 43991 37159
rect 44025 37156 44037 37159
rect 44160 37156 44166 37168
rect 44025 37128 44166 37156
rect 44025 37125 44037 37128
rect 43979 37119 44037 37125
rect 44160 37116 44166 37128
rect 44218 37116 44224 37168
rect 45448 37116 45454 37168
rect 45506 37156 45512 37168
rect 45558 37165 45586 37264
rect 46187 37261 46199 37264
rect 46233 37261 46245 37295
rect 46294 37292 46322 37332
rect 46371 37329 46383 37363
rect 46417 37360 46429 37363
rect 46552 37360 46558 37372
rect 46417 37332 46558 37360
rect 46417 37329 46429 37332
rect 46371 37323 46429 37329
rect 46552 37320 46558 37332
rect 46610 37320 46616 37372
rect 46736 37360 46742 37372
rect 46697 37332 46742 37360
rect 46736 37320 46742 37332
rect 46794 37320 46800 37372
rect 46846 37360 46874 37400
rect 46920 37388 46926 37440
rect 46978 37428 46984 37440
rect 46978 37400 50738 37428
rect 46978 37388 46984 37400
rect 46846 37332 46966 37360
rect 46647 37295 46705 37301
rect 46647 37292 46659 37295
rect 46294 37264 46659 37292
rect 46187 37255 46245 37261
rect 46647 37261 46659 37264
rect 46693 37261 46705 37295
rect 46647 37255 46705 37261
rect 46938 37224 46966 37332
rect 48208 37252 48214 37304
rect 48266 37292 48272 37304
rect 50600 37292 50606 37304
rect 48266 37264 50606 37292
rect 48266 37252 48272 37264
rect 50600 37252 50606 37264
rect 50658 37252 50664 37304
rect 50710 37292 50738 37400
rect 51888 37388 51894 37440
rect 51946 37428 51952 37440
rect 54924 37428 54930 37440
rect 51946 37400 54930 37428
rect 51946 37388 51952 37400
rect 54924 37388 54930 37400
rect 54982 37388 54988 37440
rect 50879 37363 50937 37369
rect 50879 37329 50891 37363
rect 50925 37360 50937 37363
rect 52348 37360 52354 37372
rect 50925 37332 52354 37360
rect 50925 37329 50937 37332
rect 50879 37323 50937 37329
rect 52348 37320 52354 37332
rect 52406 37320 52412 37372
rect 55016 37360 55022 37372
rect 54977 37332 55022 37360
rect 55016 37320 55022 37332
rect 55074 37320 55080 37372
rect 55126 37360 55154 37468
rect 55292 37456 55298 37508
rect 55350 37496 55356 37508
rect 60352 37496 60358 37508
rect 55350 37468 60358 37496
rect 55350 37456 55356 37468
rect 60352 37456 60358 37468
rect 60410 37456 60416 37508
rect 61364 37456 61370 37508
rect 61422 37496 61428 37508
rect 75259 37499 75317 37505
rect 61422 37468 75210 37496
rect 61422 37456 61428 37468
rect 55200 37388 55206 37440
rect 55258 37428 55264 37440
rect 58236 37428 58242 37440
rect 55258 37400 58242 37428
rect 55258 37388 55264 37400
rect 58236 37388 58242 37400
rect 58294 37388 58300 37440
rect 58331 37431 58389 37437
rect 58331 37397 58343 37431
rect 58377 37428 58389 37431
rect 60907 37431 60965 37437
rect 58377 37400 60766 37428
rect 58377 37397 58389 37400
rect 58331 37391 58389 37397
rect 55476 37360 55482 37372
rect 55126 37332 55482 37360
rect 55476 37320 55482 37332
rect 55534 37320 55540 37372
rect 55568 37320 55574 37372
rect 55626 37360 55632 37372
rect 57227 37363 57285 37369
rect 57227 37360 57239 37363
rect 55626 37332 57239 37360
rect 55626 37320 55632 37332
rect 57227 37329 57239 37332
rect 57273 37360 57285 37363
rect 57779 37363 57837 37369
rect 57779 37360 57791 37363
rect 57273 37332 57791 37360
rect 57273 37329 57285 37332
rect 57227 37323 57285 37329
rect 57779 37329 57791 37332
rect 57825 37329 57837 37363
rect 57779 37323 57837 37329
rect 57960 37320 57966 37372
rect 58018 37360 58024 37372
rect 58604 37360 58610 37372
rect 58018 37332 58610 37360
rect 58018 37320 58024 37332
rect 58604 37320 58610 37332
rect 58662 37320 58668 37372
rect 58880 37320 58886 37372
rect 58938 37360 58944 37372
rect 59803 37363 59861 37369
rect 58938 37332 59754 37360
rect 58938 37320 58944 37332
rect 54740 37292 54746 37304
rect 50710 37264 54746 37292
rect 54740 37252 54746 37264
rect 54798 37252 54804 37304
rect 54832 37252 54838 37304
rect 54890 37292 54896 37304
rect 54927 37295 54985 37301
rect 54927 37292 54939 37295
rect 54890 37264 54939 37292
rect 54890 37252 54896 37264
rect 54927 37261 54939 37264
rect 54973 37261 54985 37295
rect 54927 37255 54985 37261
rect 56123 37295 56181 37301
rect 56123 37261 56135 37295
rect 56169 37292 56181 37295
rect 56764 37292 56770 37304
rect 56169 37264 56770 37292
rect 56169 37261 56181 37264
rect 56123 37255 56181 37261
rect 48116 37224 48122 37236
rect 46938 37196 48122 37224
rect 48116 37184 48122 37196
rect 48174 37224 48180 37236
rect 50416 37224 50422 37236
rect 48174 37196 50422 37224
rect 48174 37184 48180 37196
rect 50416 37184 50422 37196
rect 50474 37184 50480 37236
rect 54942 37224 54970 37255
rect 56764 37252 56770 37264
rect 56822 37252 56828 37304
rect 57132 37292 57138 37304
rect 57093 37264 57138 37292
rect 57132 37252 57138 37264
rect 57190 37252 57196 37304
rect 59616 37292 59622 37304
rect 59577 37264 59622 37292
rect 59616 37252 59622 37264
rect 59674 37252 59680 37304
rect 57960 37224 57966 37236
rect 54942 37196 57966 37224
rect 57960 37184 57966 37196
rect 58018 37184 58024 37236
rect 59432 37224 59438 37236
rect 58162 37196 59438 37224
rect 45543 37159 45601 37165
rect 45543 37156 45555 37159
rect 45506 37128 45555 37156
rect 45506 37116 45512 37128
rect 45543 37125 45555 37128
rect 45589 37125 45601 37159
rect 45543 37119 45601 37125
rect 46003 37159 46061 37165
rect 46003 37125 46015 37159
rect 46049 37156 46061 37159
rect 47472 37156 47478 37168
rect 46049 37128 47478 37156
rect 46049 37125 46061 37128
rect 46003 37119 46061 37125
rect 47472 37116 47478 37128
rect 47530 37116 47536 37168
rect 52164 37156 52170 37168
rect 52125 37128 52170 37156
rect 52164 37116 52170 37128
rect 52222 37116 52228 37168
rect 52348 37156 52354 37168
rect 52309 37128 52354 37156
rect 52348 37116 52354 37128
rect 52406 37116 52412 37168
rect 52532 37116 52538 37168
rect 52590 37156 52596 37168
rect 58162 37156 58190 37196
rect 59432 37184 59438 37196
rect 59490 37184 59496 37236
rect 59726 37224 59754 37332
rect 59803 37329 59815 37363
rect 59849 37360 59861 37363
rect 60168 37360 60174 37372
rect 59849 37332 60174 37360
rect 59849 37329 59861 37332
rect 59803 37323 59861 37329
rect 60168 37320 60174 37332
rect 60226 37320 60232 37372
rect 60352 37360 60358 37372
rect 60313 37332 60358 37360
rect 60352 37320 60358 37332
rect 60410 37320 60416 37372
rect 60536 37360 60542 37372
rect 60497 37332 60542 37360
rect 60536 37320 60542 37332
rect 60594 37320 60600 37372
rect 60738 37360 60766 37400
rect 60907 37397 60919 37431
rect 60953 37428 60965 37431
rect 62468 37428 62474 37440
rect 60953 37400 62474 37428
rect 60953 37397 60965 37400
rect 60907 37391 60965 37397
rect 62468 37388 62474 37400
rect 62526 37388 62532 37440
rect 69000 37428 69006 37440
rect 67454 37400 69006 37428
rect 62747 37363 62805 37369
rect 62747 37360 62759 37363
rect 60738 37332 62759 37360
rect 62747 37329 62759 37332
rect 62793 37329 62805 37363
rect 67068 37360 67074 37372
rect 67029 37332 67074 37360
rect 62747 37323 62805 37329
rect 67068 37320 67074 37332
rect 67126 37320 67132 37372
rect 67454 37369 67482 37400
rect 69000 37388 69006 37400
rect 69058 37388 69064 37440
rect 71576 37388 71582 37440
rect 71634 37428 71640 37440
rect 72039 37431 72097 37437
rect 72039 37428 72051 37431
rect 71634 37400 72051 37428
rect 71634 37388 71640 37400
rect 72039 37397 72051 37400
rect 72085 37397 72097 37431
rect 72039 37391 72097 37397
rect 72496 37388 72502 37440
rect 72554 37428 72560 37440
rect 74428 37428 74434 37440
rect 72554 37400 74434 37428
rect 72554 37388 72560 37400
rect 74428 37388 74434 37400
rect 74486 37388 74492 37440
rect 75182 37428 75210 37468
rect 75259 37465 75271 37499
rect 75305 37496 75317 37499
rect 75440 37496 75446 37508
rect 75305 37468 75446 37496
rect 75305 37465 75317 37468
rect 75259 37459 75317 37465
rect 75440 37456 75446 37468
rect 75498 37456 75504 37508
rect 82251 37499 82309 37505
rect 82251 37465 82263 37499
rect 82297 37496 82309 37499
rect 83260 37496 83266 37508
rect 82297 37468 83266 37496
rect 82297 37465 82309 37468
rect 82251 37459 82309 37465
rect 83260 37456 83266 37468
rect 83318 37456 83324 37508
rect 88412 37456 88418 37508
rect 88470 37496 88476 37508
rect 88691 37499 88749 37505
rect 88691 37496 88703 37499
rect 88470 37468 88703 37496
rect 88470 37456 88476 37468
rect 88691 37465 88703 37468
rect 88737 37465 88749 37499
rect 88691 37459 88749 37465
rect 90071 37499 90129 37505
rect 90071 37465 90083 37499
rect 90117 37496 90129 37499
rect 90712 37496 90718 37508
rect 90117 37468 90718 37496
rect 90117 37465 90129 37468
rect 90071 37459 90129 37465
rect 75900 37428 75906 37440
rect 75182 37400 75906 37428
rect 75900 37388 75906 37400
rect 75958 37388 75964 37440
rect 67439 37363 67497 37369
rect 67439 37329 67451 37363
rect 67485 37329 67497 37363
rect 67439 37323 67497 37329
rect 67623 37363 67681 37369
rect 67623 37329 67635 37363
rect 67669 37360 67681 37363
rect 68356 37360 68362 37372
rect 67669 37332 68362 37360
rect 67669 37329 67681 37332
rect 67623 37323 67681 37329
rect 68356 37320 68362 37332
rect 68414 37320 68420 37372
rect 68635 37363 68693 37369
rect 68635 37329 68647 37363
rect 68681 37360 68693 37363
rect 69184 37360 69190 37372
rect 68681 37332 69190 37360
rect 68681 37329 68693 37332
rect 68635 37323 68693 37329
rect 69184 37320 69190 37332
rect 69242 37320 69248 37372
rect 69276 37320 69282 37372
rect 69334 37360 69340 37372
rect 69371 37363 69429 37369
rect 69371 37360 69383 37363
rect 69334 37332 69383 37360
rect 69334 37320 69340 37332
rect 69371 37329 69383 37332
rect 69417 37360 69429 37363
rect 69644 37360 69650 37372
rect 69417 37332 69650 37360
rect 69417 37329 69429 37332
rect 69371 37323 69429 37329
rect 69644 37320 69650 37332
rect 69702 37320 69708 37372
rect 72588 37320 72594 37372
rect 72646 37360 72652 37372
rect 72683 37363 72741 37369
rect 72683 37360 72695 37363
rect 72646 37332 72695 37360
rect 72646 37320 72652 37332
rect 72683 37329 72695 37332
rect 72729 37329 72741 37363
rect 73048 37360 73054 37372
rect 73009 37332 73054 37360
rect 72683 37323 72741 37329
rect 73048 37320 73054 37332
rect 73106 37320 73112 37372
rect 73235 37363 73293 37369
rect 73235 37329 73247 37363
rect 73281 37360 73293 37363
rect 73692 37360 73698 37372
rect 73281 37332 73698 37360
rect 73281 37329 73293 37332
rect 73235 37323 73293 37329
rect 73692 37320 73698 37332
rect 73750 37320 73756 37372
rect 73876 37320 73882 37372
rect 73934 37360 73940 37372
rect 74063 37363 74121 37369
rect 74063 37360 74075 37363
rect 73934 37332 74075 37360
rect 73934 37320 73940 37332
rect 74063 37329 74075 37332
rect 74109 37329 74121 37363
rect 74244 37360 74250 37372
rect 74205 37332 74250 37360
rect 74063 37323 74121 37329
rect 74244 37320 74250 37332
rect 74302 37320 74308 37372
rect 74799 37363 74857 37369
rect 74799 37360 74811 37363
rect 74354 37332 74811 37360
rect 62100 37252 62106 37304
rect 62158 37292 62164 37304
rect 62471 37295 62529 37301
rect 62471 37292 62483 37295
rect 62158 37264 62483 37292
rect 62158 37252 62164 37264
rect 62471 37261 62483 37264
rect 62517 37261 62529 37295
rect 62471 37255 62529 37261
rect 67163 37295 67221 37301
rect 67163 37261 67175 37295
rect 67209 37292 67221 37295
rect 68172 37292 68178 37304
rect 67209 37264 68178 37292
rect 67209 37261 67221 37264
rect 67163 37255 67221 37261
rect 68172 37252 68178 37264
rect 68230 37252 68236 37304
rect 68264 37252 68270 37304
rect 68322 37292 68328 37304
rect 68540 37292 68546 37304
rect 68322 37264 68546 37292
rect 68322 37252 68328 37264
rect 68540 37252 68546 37264
rect 68598 37252 68604 37304
rect 72775 37295 72833 37301
rect 72775 37261 72787 37295
rect 72821 37292 72833 37295
rect 73600 37292 73606 37304
rect 72821 37264 73606 37292
rect 72821 37261 72833 37264
rect 72775 37255 72833 37261
rect 73600 37252 73606 37264
rect 73658 37252 73664 37304
rect 73968 37252 73974 37304
rect 74026 37292 74032 37304
rect 74354 37292 74382 37332
rect 74799 37329 74811 37332
rect 74845 37329 74857 37363
rect 74980 37360 74986 37372
rect 74941 37332 74986 37360
rect 74799 37323 74857 37329
rect 74980 37320 74986 37332
rect 75038 37320 75044 37372
rect 75348 37320 75354 37372
rect 75406 37360 75412 37372
rect 77927 37363 77985 37369
rect 77927 37360 77939 37363
rect 75406 37332 77939 37360
rect 75406 37320 75412 37332
rect 77927 37329 77939 37332
rect 77973 37329 77985 37363
rect 80503 37363 80561 37369
rect 80503 37360 80515 37363
rect 77927 37323 77985 37329
rect 80334 37332 80515 37360
rect 74026 37264 74382 37292
rect 74026 37252 74032 37264
rect 77464 37252 77470 37304
rect 77522 37292 77528 37304
rect 77651 37295 77709 37301
rect 77651 37292 77663 37295
rect 77522 37264 77663 37292
rect 77522 37252 77528 37264
rect 77651 37261 77663 37264
rect 77697 37261 77709 37295
rect 77651 37255 77709 37261
rect 60352 37224 60358 37236
rect 59726 37196 60358 37224
rect 60352 37184 60358 37196
rect 60410 37184 60416 37236
rect 66703 37227 66761 37233
rect 60462 37196 62514 37224
rect 52590 37128 58190 37156
rect 52590 37116 52596 37128
rect 58236 37116 58242 37168
rect 58294 37156 58300 37168
rect 60462 37156 60490 37196
rect 58294 37128 60490 37156
rect 58294 37116 58300 37128
rect 60536 37116 60542 37168
rect 60594 37156 60600 37168
rect 61180 37156 61186 37168
rect 60594 37128 61186 37156
rect 60594 37116 60600 37128
rect 61180 37116 61186 37128
rect 61238 37116 61244 37168
rect 62100 37116 62106 37168
rect 62158 37156 62164 37168
rect 62287 37159 62345 37165
rect 62287 37156 62299 37159
rect 62158 37128 62299 37156
rect 62158 37116 62164 37128
rect 62287 37125 62299 37128
rect 62333 37125 62345 37159
rect 62486 37156 62514 37196
rect 66703 37193 66715 37227
rect 66749 37224 66761 37227
rect 68448 37224 68454 37236
rect 66749 37196 68454 37224
rect 66749 37193 66761 37196
rect 66703 37187 66761 37193
rect 68448 37184 68454 37196
rect 68506 37184 68512 37236
rect 69276 37184 69282 37236
rect 69334 37224 69340 37236
rect 69555 37227 69613 37233
rect 69555 37224 69567 37227
rect 69334 37196 69567 37224
rect 69334 37184 69340 37196
rect 69555 37193 69567 37196
rect 69601 37193 69613 37227
rect 69555 37187 69613 37193
rect 74244 37184 74250 37236
rect 74302 37224 74308 37236
rect 74302 37196 77602 37224
rect 74302 37184 74308 37196
rect 63204 37156 63210 37168
rect 62486 37128 63210 37156
rect 62287 37119 62345 37125
rect 63204 37116 63210 37128
rect 63262 37116 63268 37168
rect 64032 37156 64038 37168
rect 63993 37128 64038 37156
rect 64032 37116 64038 37128
rect 64090 37116 64096 37168
rect 67068 37116 67074 37168
rect 67126 37156 67132 37168
rect 68632 37156 68638 37168
rect 67126 37128 68638 37156
rect 67126 37116 67132 37128
rect 68632 37116 68638 37128
rect 68690 37116 68696 37168
rect 70012 37116 70018 37168
rect 70070 37156 70076 37168
rect 76636 37156 76642 37168
rect 70070 37128 76642 37156
rect 70070 37116 70076 37128
rect 76636 37116 76642 37128
rect 76694 37116 76700 37168
rect 76728 37116 76734 37168
rect 76786 37156 76792 37168
rect 77464 37156 77470 37168
rect 76786 37128 77470 37156
rect 76786 37116 76792 37128
rect 77464 37116 77470 37128
rect 77522 37116 77528 37168
rect 77574 37156 77602 37196
rect 80334 37168 80362 37332
rect 80503 37329 80515 37332
rect 80549 37329 80561 37363
rect 82064 37360 82070 37372
rect 82025 37332 82070 37360
rect 80503 37323 80561 37329
rect 82064 37320 82070 37332
rect 82122 37360 82128 37372
rect 82435 37363 82493 37369
rect 82435 37360 82447 37363
rect 82122 37332 82447 37360
rect 82122 37320 82128 37332
rect 82435 37329 82447 37332
rect 82481 37329 82493 37363
rect 84272 37360 84278 37372
rect 84233 37332 84278 37360
rect 82435 37323 82493 37329
rect 84272 37320 84278 37332
rect 84330 37320 84336 37372
rect 85655 37363 85713 37369
rect 85655 37329 85667 37363
rect 85701 37360 85713 37363
rect 86483 37363 86541 37369
rect 86483 37360 86495 37363
rect 85701 37332 86495 37360
rect 85701 37329 85713 37332
rect 85655 37323 85713 37329
rect 86483 37329 86495 37332
rect 86529 37329 86541 37363
rect 88706 37360 88734 37459
rect 90712 37456 90718 37468
rect 90770 37456 90776 37508
rect 89074 37400 89654 37428
rect 89074 37369 89102 37400
rect 88875 37363 88933 37369
rect 88875 37360 88887 37363
rect 88706 37332 88887 37360
rect 86483 37323 86541 37329
rect 88875 37329 88887 37332
rect 88921 37329 88933 37363
rect 89059 37363 89117 37369
rect 89059 37360 89071 37363
rect 88875 37323 88933 37329
rect 88982 37332 89071 37360
rect 83999 37295 84057 37301
rect 83999 37292 84011 37295
rect 83922 37264 84011 37292
rect 83922 37168 83950 37264
rect 83999 37261 84011 37264
rect 84045 37261 84057 37295
rect 83999 37255 84057 37261
rect 88320 37252 88326 37304
rect 88378 37292 88384 37304
rect 88982 37292 89010 37332
rect 89059 37329 89071 37332
rect 89105 37329 89117 37363
rect 89516 37360 89522 37372
rect 89477 37332 89522 37360
rect 89059 37323 89117 37329
rect 89516 37320 89522 37332
rect 89574 37320 89580 37372
rect 89626 37369 89654 37400
rect 89611 37363 89669 37369
rect 89611 37329 89623 37363
rect 89657 37329 89669 37363
rect 89611 37323 89669 37329
rect 91267 37363 91325 37369
rect 91267 37329 91279 37363
rect 91313 37360 91325 37363
rect 91356 37360 91362 37372
rect 91313 37332 91362 37360
rect 91313 37329 91325 37332
rect 91267 37323 91325 37329
rect 91356 37320 91362 37332
rect 91414 37320 91420 37372
rect 88378 37264 89010 37292
rect 88378 37252 88384 37264
rect 89516 37184 89522 37236
rect 89574 37224 89580 37236
rect 90252 37224 90258 37236
rect 89574 37196 90258 37224
rect 89574 37184 89580 37196
rect 90252 37184 90258 37196
rect 90310 37224 90316 37236
rect 91359 37227 91417 37233
rect 91359 37224 91371 37227
rect 90310 37196 91371 37224
rect 90310 37184 90316 37196
rect 91359 37193 91371 37196
rect 91405 37193 91417 37227
rect 91359 37187 91417 37193
rect 78108 37156 78114 37168
rect 77574 37128 78114 37156
rect 78108 37116 78114 37128
rect 78166 37116 78172 37168
rect 79212 37156 79218 37168
rect 79173 37128 79218 37156
rect 79212 37116 79218 37128
rect 79270 37116 79276 37168
rect 80316 37156 80322 37168
rect 80277 37128 80322 37156
rect 80316 37116 80322 37128
rect 80374 37116 80380 37168
rect 80687 37159 80745 37165
rect 80687 37125 80699 37159
rect 80733 37156 80745 37159
rect 82708 37156 82714 37168
rect 80733 37128 82714 37156
rect 80733 37125 80745 37128
rect 80687 37119 80745 37125
rect 82708 37116 82714 37128
rect 82766 37116 82772 37168
rect 83904 37156 83910 37168
rect 83865 37128 83910 37156
rect 83904 37116 83910 37128
rect 83962 37116 83968 37168
rect 86572 37156 86578 37168
rect 86533 37128 86578 37156
rect 86572 37116 86578 37128
rect 86630 37116 86636 37168
rect 538 37066 93642 37088
rect 538 37014 3680 37066
rect 3732 37014 3744 37066
rect 3796 37014 3808 37066
rect 3860 37014 3872 37066
rect 3924 37014 9008 37066
rect 9060 37014 9072 37066
rect 9124 37014 9136 37066
rect 9188 37014 9200 37066
rect 9252 37014 14336 37066
rect 14388 37014 14400 37066
rect 14452 37014 14464 37066
rect 14516 37014 14528 37066
rect 14580 37014 19664 37066
rect 19716 37014 19728 37066
rect 19780 37014 19792 37066
rect 19844 37014 19856 37066
rect 19908 37014 24992 37066
rect 25044 37014 25056 37066
rect 25108 37014 25120 37066
rect 25172 37014 25184 37066
rect 25236 37014 30320 37066
rect 30372 37014 30384 37066
rect 30436 37014 30448 37066
rect 30500 37014 30512 37066
rect 30564 37014 35648 37066
rect 35700 37014 35712 37066
rect 35764 37014 35776 37066
rect 35828 37014 35840 37066
rect 35892 37014 40976 37066
rect 41028 37014 41040 37066
rect 41092 37014 41104 37066
rect 41156 37014 41168 37066
rect 41220 37014 46304 37066
rect 46356 37014 46368 37066
rect 46420 37014 46432 37066
rect 46484 37014 46496 37066
rect 46548 37014 51632 37066
rect 51684 37014 51696 37066
rect 51748 37014 51760 37066
rect 51812 37014 51824 37066
rect 51876 37014 56960 37066
rect 57012 37014 57024 37066
rect 57076 37014 57088 37066
rect 57140 37014 57152 37066
rect 57204 37014 62288 37066
rect 62340 37014 62352 37066
rect 62404 37014 62416 37066
rect 62468 37014 62480 37066
rect 62532 37014 67616 37066
rect 67668 37014 67680 37066
rect 67732 37014 67744 37066
rect 67796 37014 67808 37066
rect 67860 37014 72944 37066
rect 72996 37014 73008 37066
rect 73060 37014 73072 37066
rect 73124 37014 73136 37066
rect 73188 37014 78272 37066
rect 78324 37014 78336 37066
rect 78388 37014 78400 37066
rect 78452 37014 78464 37066
rect 78516 37014 83600 37066
rect 83652 37014 83664 37066
rect 83716 37014 83728 37066
rect 83780 37014 83792 37066
rect 83844 37014 88928 37066
rect 88980 37014 88992 37066
rect 89044 37014 89056 37066
rect 89108 37014 89120 37066
rect 89172 37014 93642 37066
rect 538 36992 93642 37014
rect 2211 36955 2269 36961
rect 2211 36921 2223 36955
rect 2257 36952 2269 36955
rect 2392 36952 2398 36964
rect 2257 36924 2398 36952
rect 2257 36921 2269 36924
rect 2211 36915 2269 36921
rect 2392 36912 2398 36924
rect 2450 36912 2456 36964
rect 16008 36912 16014 36964
rect 16066 36952 16072 36964
rect 16287 36955 16345 36961
rect 16287 36952 16299 36955
rect 16066 36924 16299 36952
rect 16066 36912 16072 36924
rect 16287 36921 16299 36924
rect 16333 36921 16345 36955
rect 16287 36915 16345 36921
rect 17204 36912 17210 36964
rect 17262 36952 17268 36964
rect 17759 36955 17817 36961
rect 17759 36952 17771 36955
rect 17262 36924 17771 36952
rect 17262 36912 17268 36924
rect 17759 36921 17771 36924
rect 17805 36921 17817 36955
rect 21344 36952 21350 36964
rect 21305 36924 21350 36952
rect 17759 36915 17817 36921
rect 21344 36912 21350 36924
rect 21402 36912 21408 36964
rect 27692 36912 27698 36964
rect 27750 36952 27756 36964
rect 28244 36952 28250 36964
rect 27750 36924 28250 36952
rect 27750 36912 27756 36924
rect 28244 36912 28250 36924
rect 28302 36912 28308 36964
rect 29716 36912 29722 36964
rect 29774 36952 29780 36964
rect 51428 36952 51434 36964
rect 29774 36924 51434 36952
rect 29774 36912 29780 36924
rect 51428 36912 51434 36924
rect 51486 36912 51492 36964
rect 51980 36912 51986 36964
rect 52038 36952 52044 36964
rect 52164 36952 52170 36964
rect 52038 36924 52170 36952
rect 52038 36912 52044 36924
rect 52164 36912 52170 36924
rect 52222 36912 52228 36964
rect 52348 36912 52354 36964
rect 52406 36952 52412 36964
rect 52406 36924 53590 36952
rect 52406 36912 52412 36924
rect 22816 36844 22822 36896
rect 22874 36884 22880 36896
rect 27324 36884 27330 36896
rect 22874 36856 27330 36884
rect 22874 36844 22880 36856
rect 27324 36844 27330 36856
rect 27382 36884 27388 36896
rect 39284 36884 39290 36896
rect 27382 36856 39290 36884
rect 27382 36844 27388 36856
rect 39284 36844 39290 36856
rect 39342 36844 39348 36896
rect 40480 36884 40486 36896
rect 40441 36856 40486 36884
rect 40480 36844 40486 36856
rect 40538 36844 40544 36896
rect 43056 36844 43062 36896
rect 43114 36884 43120 36896
rect 43976 36884 43982 36896
rect 43114 36856 43982 36884
rect 43114 36844 43120 36856
rect 43976 36844 43982 36856
rect 44034 36844 44040 36896
rect 45540 36884 45546 36896
rect 45501 36856 45546 36884
rect 45540 36844 45546 36856
rect 45598 36844 45604 36896
rect 50143 36887 50201 36893
rect 50143 36853 50155 36887
rect 50189 36884 50201 36887
rect 51336 36884 51342 36896
rect 50189 36856 51342 36884
rect 50189 36853 50201 36856
rect 50143 36847 50201 36853
rect 51336 36844 51342 36856
rect 51394 36844 51400 36896
rect 3128 36816 3134 36828
rect 3089 36788 3134 36816
rect 3128 36776 3134 36788
rect 3186 36776 3192 36828
rect 15824 36776 15830 36828
rect 15882 36816 15888 36828
rect 18127 36819 18185 36825
rect 18127 36816 18139 36819
rect 15882 36788 18139 36816
rect 15882 36776 15888 36788
rect 1567 36751 1625 36757
rect 1567 36717 1579 36751
rect 1613 36748 1625 36751
rect 2484 36748 2490 36760
rect 1613 36720 2490 36748
rect 1613 36717 1625 36720
rect 1567 36711 1625 36717
rect 2484 36708 2490 36720
rect 2542 36708 2548 36760
rect 3404 36748 3410 36760
rect 3365 36720 3410 36748
rect 3404 36708 3410 36720
rect 3462 36708 3468 36760
rect 17498 36757 17526 36788
rect 18127 36785 18139 36788
rect 18173 36816 18185 36819
rect 19691 36819 19749 36825
rect 19691 36816 19703 36819
rect 18173 36788 19703 36816
rect 18173 36785 18185 36788
rect 18127 36779 18185 36785
rect 19691 36785 19703 36788
rect 19737 36785 19749 36819
rect 20332 36816 20338 36828
rect 20293 36788 20338 36816
rect 19691 36779 19749 36785
rect 9663 36751 9721 36757
rect 9663 36748 9675 36751
rect 9494 36720 9675 36748
rect 4787 36683 4845 36689
rect 4787 36649 4799 36683
rect 4833 36680 4845 36683
rect 5796 36680 5802 36692
rect 4833 36652 5802 36680
rect 4833 36649 4845 36652
rect 4787 36643 4845 36649
rect 5796 36640 5802 36652
rect 5854 36640 5860 36692
rect 9494 36624 9522 36720
rect 9663 36717 9675 36720
rect 9709 36717 9721 36751
rect 9663 36711 9721 36717
rect 16195 36751 16253 36757
rect 16195 36717 16207 36751
rect 16241 36717 16253 36751
rect 16195 36711 16253 36717
rect 17483 36751 17541 36757
rect 17483 36717 17495 36751
rect 17529 36717 17541 36751
rect 17664 36748 17670 36760
rect 17625 36720 17670 36748
rect 17483 36711 17541 36717
rect 16210 36624 16238 36711
rect 17664 36708 17670 36720
rect 17722 36708 17728 36760
rect 19706 36748 19734 36779
rect 20332 36776 20338 36788
rect 20390 36776 20396 36828
rect 31372 36816 31378 36828
rect 31333 36788 31378 36816
rect 31372 36776 31378 36788
rect 31430 36776 31436 36828
rect 32108 36816 32114 36828
rect 32069 36788 32114 36816
rect 32108 36776 32114 36788
rect 32166 36776 32172 36828
rect 32292 36776 32298 36828
rect 32350 36816 32356 36828
rect 32350 36788 39330 36816
rect 32350 36776 32356 36788
rect 19875 36751 19933 36757
rect 19875 36748 19887 36751
rect 19706 36720 19887 36748
rect 19875 36717 19887 36720
rect 19921 36717 19933 36751
rect 19875 36711 19933 36717
rect 20059 36751 20117 36757
rect 20059 36717 20071 36751
rect 20105 36748 20117 36751
rect 21252 36748 21258 36760
rect 20105 36720 20654 36748
rect 21213 36720 21258 36748
rect 20105 36717 20117 36720
rect 20059 36711 20117 36717
rect 20626 36689 20654 36720
rect 21252 36708 21258 36720
rect 21310 36708 21316 36760
rect 28707 36751 28765 36757
rect 28707 36717 28719 36751
rect 28753 36748 28765 36751
rect 28980 36748 28986 36760
rect 28753 36720 28986 36748
rect 28753 36717 28765 36720
rect 28707 36711 28765 36717
rect 28980 36708 28986 36720
rect 29038 36708 29044 36760
rect 31924 36708 31930 36760
rect 31982 36757 31988 36760
rect 31982 36751 32031 36757
rect 31982 36717 31985 36751
rect 32019 36717 32031 36751
rect 31982 36711 32031 36717
rect 32387 36751 32445 36757
rect 32387 36717 32399 36751
rect 32433 36748 32445 36751
rect 32476 36748 32482 36760
rect 32433 36720 32482 36748
rect 32433 36717 32445 36720
rect 32387 36711 32445 36717
rect 31982 36708 31988 36711
rect 32476 36708 32482 36720
rect 32534 36708 32540 36760
rect 32571 36751 32629 36757
rect 32571 36717 32583 36751
rect 32617 36748 32629 36751
rect 32755 36751 32813 36757
rect 32755 36748 32767 36751
rect 32617 36720 32767 36748
rect 32617 36717 32629 36720
rect 32571 36711 32629 36717
rect 32755 36717 32767 36720
rect 32801 36748 32813 36751
rect 33488 36748 33494 36760
rect 32801 36720 33494 36748
rect 32801 36717 32813 36720
rect 32755 36711 32813 36717
rect 33488 36708 33494 36720
rect 33546 36708 33552 36760
rect 33580 36708 33586 36760
rect 33638 36748 33644 36760
rect 37536 36748 37542 36760
rect 33638 36720 37542 36748
rect 33638 36708 33644 36720
rect 37536 36708 37542 36720
rect 37594 36708 37600 36760
rect 37631 36751 37689 36757
rect 37631 36717 37643 36751
rect 37677 36717 37689 36751
rect 39302 36748 39330 36788
rect 43700 36776 43706 36828
rect 43758 36816 43764 36828
rect 51983 36819 52041 36825
rect 43758 36788 51934 36816
rect 43758 36776 43764 36788
rect 40115 36751 40173 36757
rect 40115 36748 40127 36751
rect 39302 36720 40127 36748
rect 37631 36711 37689 36717
rect 40115 36717 40127 36720
rect 40161 36748 40173 36751
rect 40299 36751 40357 36757
rect 40299 36748 40311 36751
rect 40161 36720 40311 36748
rect 40161 36717 40173 36720
rect 40115 36711 40173 36717
rect 40299 36717 40311 36720
rect 40345 36748 40357 36751
rect 40848 36748 40854 36760
rect 40345 36720 40854 36748
rect 40345 36717 40357 36720
rect 40299 36711 40357 36717
rect 20611 36683 20669 36689
rect 20611 36649 20623 36683
rect 20657 36680 20669 36683
rect 21528 36680 21534 36692
rect 20657 36652 21534 36680
rect 20657 36649 20669 36652
rect 20611 36643 20669 36649
rect 21528 36640 21534 36652
rect 21586 36680 21592 36692
rect 21586 36652 32062 36680
rect 21586 36640 21592 36652
rect 32034 36624 32062 36652
rect 32200 36640 32206 36692
rect 32258 36680 32264 36692
rect 37444 36680 37450 36692
rect 32258 36652 37450 36680
rect 32258 36640 32264 36652
rect 37444 36640 37450 36652
rect 37502 36640 37508 36692
rect 4968 36612 4974 36624
rect 4929 36584 4974 36612
rect 4968 36572 4974 36584
rect 5026 36572 5032 36624
rect 9476 36612 9482 36624
rect 9437 36584 9482 36612
rect 9476 36572 9482 36584
rect 9534 36572 9540 36624
rect 9847 36615 9905 36621
rect 9847 36581 9859 36615
rect 9893 36612 9905 36615
rect 10488 36612 10494 36624
rect 9893 36584 10494 36612
rect 9893 36581 9905 36584
rect 9847 36575 9905 36581
rect 10488 36572 10494 36584
rect 10546 36572 10552 36624
rect 16103 36615 16161 36621
rect 16103 36581 16115 36615
rect 16149 36612 16161 36615
rect 16192 36612 16198 36624
rect 16149 36584 16198 36612
rect 16149 36581 16161 36584
rect 16103 36575 16161 36581
rect 16192 36572 16198 36584
rect 16250 36572 16256 36624
rect 28796 36612 28802 36624
rect 28757 36584 28802 36612
rect 28796 36572 28802 36584
rect 28854 36572 28860 36624
rect 32016 36572 32022 36624
rect 32074 36572 32080 36624
rect 32108 36572 32114 36624
rect 32166 36612 32172 36624
rect 32752 36612 32758 36624
rect 32166 36584 32758 36612
rect 32166 36572 32172 36584
rect 32752 36572 32758 36584
rect 32810 36612 32816 36624
rect 32847 36615 32905 36621
rect 32847 36612 32859 36615
rect 32810 36584 32859 36612
rect 32810 36572 32816 36584
rect 32847 36581 32859 36584
rect 32893 36581 32905 36615
rect 32847 36575 32905 36581
rect 34776 36572 34782 36624
rect 34834 36612 34840 36624
rect 37539 36615 37597 36621
rect 37539 36612 37551 36615
rect 34834 36584 37551 36612
rect 34834 36572 34840 36584
rect 37539 36581 37551 36584
rect 37585 36612 37597 36615
rect 37646 36612 37674 36711
rect 40848 36708 40854 36720
rect 40906 36708 40912 36760
rect 42688 36748 42694 36760
rect 42649 36720 42694 36748
rect 42688 36708 42694 36720
rect 42746 36708 42752 36760
rect 42783 36751 42841 36757
rect 42783 36717 42795 36751
rect 42829 36748 42841 36751
rect 42872 36748 42878 36760
rect 42829 36720 42878 36748
rect 42829 36717 42841 36720
rect 42783 36711 42841 36717
rect 42872 36708 42878 36720
rect 42930 36708 42936 36760
rect 43056 36708 43062 36760
rect 43114 36748 43120 36760
rect 43151 36751 43209 36757
rect 43151 36748 43163 36751
rect 43114 36720 43163 36748
rect 43114 36708 43120 36720
rect 43151 36717 43163 36720
rect 43197 36717 43209 36751
rect 43151 36711 43209 36717
rect 43240 36708 43246 36760
rect 43298 36748 43304 36760
rect 43298 36720 43343 36748
rect 43298 36708 43304 36720
rect 45540 36708 45546 36760
rect 45598 36748 45604 36760
rect 46187 36751 46245 36757
rect 46187 36748 46199 36751
rect 45598 36720 46199 36748
rect 45598 36708 45604 36720
rect 46187 36717 46199 36720
rect 46233 36717 46245 36751
rect 46187 36711 46245 36717
rect 46371 36751 46429 36757
rect 46371 36717 46383 36751
rect 46417 36748 46429 36751
rect 46552 36748 46558 36760
rect 46417 36720 46558 36748
rect 46417 36717 46429 36720
rect 46371 36711 46429 36717
rect 46552 36708 46558 36720
rect 46610 36708 46616 36760
rect 46736 36748 46742 36760
rect 46697 36720 46742 36748
rect 46736 36708 46742 36720
rect 46794 36708 46800 36760
rect 46828 36708 46834 36760
rect 46886 36748 46892 36760
rect 46886 36720 46931 36748
rect 46886 36708 46892 36720
rect 47656 36708 47662 36760
rect 47714 36708 47720 36760
rect 50051 36751 50109 36757
rect 50051 36717 50063 36751
rect 50097 36748 50109 36751
rect 51707 36751 51765 36757
rect 50097 36720 50554 36748
rect 50097 36717 50109 36720
rect 50051 36711 50109 36717
rect 43795 36683 43853 36689
rect 43795 36649 43807 36683
rect 43841 36680 43853 36683
rect 44068 36680 44074 36692
rect 43841 36652 44074 36680
rect 43841 36649 43853 36652
rect 43795 36643 43853 36649
rect 44068 36640 44074 36652
rect 44126 36640 44132 36692
rect 47674 36680 47702 36708
rect 50416 36680 50422 36692
rect 47674 36652 50422 36680
rect 50416 36640 50422 36652
rect 50474 36640 50480 36692
rect 37720 36612 37726 36624
rect 37585 36584 37726 36612
rect 37585 36581 37597 36584
rect 37539 36575 37597 36581
rect 37720 36572 37726 36584
rect 37778 36572 37784 36624
rect 37815 36615 37873 36621
rect 37815 36581 37827 36615
rect 37861 36612 37873 36615
rect 37904 36612 37910 36624
rect 37861 36584 37910 36612
rect 37861 36581 37873 36584
rect 37815 36575 37873 36581
rect 37904 36572 37910 36584
rect 37962 36612 37968 36624
rect 42688 36612 42694 36624
rect 37962 36584 42694 36612
rect 37962 36572 37968 36584
rect 42688 36572 42694 36584
rect 42746 36612 42752 36624
rect 43240 36612 43246 36624
rect 42746 36584 43246 36612
rect 42746 36572 42752 36584
rect 43240 36572 43246 36584
rect 43298 36572 43304 36624
rect 46003 36615 46061 36621
rect 46003 36581 46015 36615
rect 46049 36612 46061 36615
rect 47656 36612 47662 36624
rect 46049 36584 47662 36612
rect 46049 36581 46061 36584
rect 46003 36575 46061 36581
rect 47656 36572 47662 36584
rect 47714 36572 47720 36624
rect 50526 36612 50554 36720
rect 51707 36717 51719 36751
rect 51753 36748 51765 36751
rect 51796 36748 51802 36760
rect 51753 36720 51802 36748
rect 51753 36717 51765 36720
rect 51707 36711 51765 36717
rect 50600 36640 50606 36692
rect 50658 36680 50664 36692
rect 51722 36680 51750 36711
rect 51796 36708 51802 36720
rect 51854 36708 51860 36760
rect 51906 36748 51934 36788
rect 51983 36785 51995 36819
rect 52029 36816 52041 36819
rect 52440 36816 52446 36828
rect 52029 36788 52446 36816
rect 52029 36785 52041 36788
rect 51983 36779 52041 36785
rect 52440 36776 52446 36788
rect 52498 36776 52504 36828
rect 53562 36825 53590 36924
rect 54924 36912 54930 36964
rect 54982 36952 54988 36964
rect 57227 36955 57285 36961
rect 57227 36952 57239 36955
rect 54982 36924 57239 36952
rect 54982 36912 54988 36924
rect 57227 36921 57239 36924
rect 57273 36952 57285 36955
rect 57960 36952 57966 36964
rect 57273 36924 57966 36952
rect 57273 36921 57285 36924
rect 57227 36915 57285 36921
rect 57960 36912 57966 36924
rect 58018 36912 58024 36964
rect 58052 36912 58058 36964
rect 58110 36952 58116 36964
rect 62008 36952 62014 36964
rect 58110 36924 62014 36952
rect 58110 36912 58116 36924
rect 62008 36912 62014 36924
rect 62066 36912 62072 36964
rect 62379 36955 62437 36961
rect 62379 36921 62391 36955
rect 62425 36952 62437 36955
rect 64127 36955 64185 36961
rect 64127 36952 64139 36955
rect 62425 36924 64139 36952
rect 62425 36921 62437 36924
rect 62379 36915 62437 36921
rect 64127 36921 64139 36924
rect 64173 36952 64185 36955
rect 72496 36952 72502 36964
rect 64173 36924 72502 36952
rect 64173 36921 64185 36924
rect 64127 36915 64185 36921
rect 72496 36912 72502 36924
rect 72554 36912 72560 36964
rect 72588 36912 72594 36964
rect 72646 36952 72652 36964
rect 73787 36955 73845 36961
rect 73787 36952 73799 36955
rect 72646 36924 73799 36952
rect 72646 36912 72652 36924
rect 73787 36921 73799 36924
rect 73833 36921 73845 36955
rect 73787 36915 73845 36921
rect 75995 36955 76053 36961
rect 75995 36921 76007 36955
rect 76041 36952 76053 36955
rect 80316 36952 80322 36964
rect 76041 36924 80322 36952
rect 76041 36921 76053 36924
rect 75995 36915 76053 36921
rect 80316 36912 80322 36924
rect 80374 36912 80380 36964
rect 82156 36912 82162 36964
rect 82214 36952 82220 36964
rect 88320 36952 88326 36964
rect 82214 36924 88326 36952
rect 82214 36912 82220 36924
rect 88320 36912 88326 36924
rect 88378 36912 88384 36964
rect 88599 36955 88657 36961
rect 88599 36921 88611 36955
rect 88645 36952 88657 36955
rect 88780 36952 88786 36964
rect 88645 36924 88786 36952
rect 88645 36921 88657 36924
rect 88599 36915 88657 36921
rect 88780 36912 88786 36924
rect 88838 36912 88844 36964
rect 55476 36844 55482 36896
rect 55534 36884 55540 36896
rect 58239 36887 58297 36893
rect 58239 36884 58251 36887
rect 55534 36856 58251 36884
rect 55534 36844 55540 36856
rect 58239 36853 58251 36856
rect 58285 36853 58297 36887
rect 58239 36847 58297 36853
rect 61180 36844 61186 36896
rect 61238 36884 61244 36896
rect 62563 36887 62621 36893
rect 62563 36884 62575 36887
rect 61238 36856 62575 36884
rect 61238 36844 61244 36856
rect 62563 36853 62575 36856
rect 62609 36853 62621 36887
rect 68080 36884 68086 36896
rect 62563 36847 62621 36853
rect 68006 36856 68086 36884
rect 53547 36819 53605 36825
rect 53547 36785 53559 36819
rect 53593 36816 53605 36819
rect 56120 36816 56126 36828
rect 53593 36788 56126 36816
rect 53593 36785 53605 36788
rect 53547 36779 53605 36785
rect 56120 36776 56126 36788
rect 56178 36776 56184 36828
rect 65596 36816 65602 36828
rect 57058 36788 65602 36816
rect 57058 36757 57086 36788
rect 65596 36776 65602 36788
rect 65654 36776 65660 36828
rect 68006 36825 68034 36856
rect 68080 36844 68086 36856
rect 68138 36844 68144 36896
rect 68172 36844 68178 36896
rect 68230 36884 68236 36896
rect 68724 36884 68730 36896
rect 68230 36856 68730 36884
rect 68230 36844 68236 36856
rect 68724 36844 68730 36856
rect 68782 36844 68788 36896
rect 73968 36884 73974 36896
rect 69938 36856 73974 36884
rect 67991 36819 68049 36825
rect 67991 36785 68003 36819
rect 68037 36785 68049 36819
rect 67991 36779 68049 36785
rect 56859 36751 56917 36757
rect 56859 36748 56871 36751
rect 51906 36720 56871 36748
rect 56859 36717 56871 36720
rect 56905 36748 56917 36751
rect 57043 36751 57101 36757
rect 57043 36748 57055 36751
rect 56905 36720 57055 36748
rect 56905 36717 56917 36720
rect 56859 36711 56917 36717
rect 57043 36717 57055 36720
rect 57089 36717 57101 36751
rect 57043 36711 57101 36717
rect 57132 36708 57138 36760
rect 57190 36748 57196 36760
rect 57776 36748 57782 36760
rect 57190 36720 57782 36748
rect 57190 36708 57196 36720
rect 57776 36708 57782 36720
rect 57834 36708 57840 36760
rect 58052 36708 58058 36760
rect 58110 36748 58116 36760
rect 58147 36751 58205 36757
rect 58147 36748 58159 36751
rect 58110 36720 58159 36748
rect 58110 36708 58116 36720
rect 58147 36717 58159 36720
rect 58193 36717 58205 36751
rect 58147 36711 58205 36717
rect 62471 36751 62529 36757
rect 62471 36717 62483 36751
rect 62517 36748 62529 36751
rect 62928 36748 62934 36760
rect 62517 36720 62934 36748
rect 62517 36717 62529 36720
rect 62471 36711 62529 36717
rect 62928 36708 62934 36720
rect 62986 36748 62992 36760
rect 63756 36748 63762 36760
rect 62986 36720 63762 36748
rect 62986 36708 62992 36720
rect 63756 36708 63762 36720
rect 63814 36708 63820 36760
rect 64032 36748 64038 36760
rect 63993 36720 64038 36748
rect 64032 36708 64038 36720
rect 64090 36708 64096 36760
rect 68190 36757 68218 36844
rect 69184 36816 69190 36828
rect 69145 36788 69190 36816
rect 69184 36776 69190 36788
rect 69242 36776 69248 36828
rect 68160 36751 68218 36757
rect 68160 36717 68172 36751
rect 68206 36717 68218 36751
rect 68160 36711 68218 36717
rect 68356 36708 68362 36760
rect 68414 36748 68420 36760
rect 68635 36751 68693 36757
rect 68635 36748 68647 36751
rect 68414 36720 68647 36748
rect 68414 36708 68420 36720
rect 68635 36717 68647 36720
rect 68681 36717 68693 36751
rect 68635 36711 68693 36717
rect 68724 36708 68730 36760
rect 68782 36748 68788 36760
rect 69938 36748 69966 36856
rect 73968 36844 73974 36856
rect 74026 36844 74032 36896
rect 74060 36844 74066 36896
rect 74118 36884 74124 36896
rect 80871 36887 80929 36893
rect 80871 36884 80883 36887
rect 74118 36856 80883 36884
rect 74118 36844 74124 36856
rect 80871 36853 80883 36856
rect 80917 36853 80929 36887
rect 80871 36847 80929 36853
rect 72220 36776 72226 36828
rect 72278 36816 72284 36828
rect 72278 36788 73646 36816
rect 72278 36776 72284 36788
rect 73618 36757 73646 36788
rect 74704 36776 74710 36828
rect 74762 36816 74768 36828
rect 79304 36816 79310 36828
rect 74762 36788 79310 36816
rect 74762 36776 74768 36788
rect 79304 36776 79310 36788
rect 79362 36776 79368 36828
rect 73419 36751 73477 36757
rect 73419 36748 73431 36751
rect 68782 36720 69966 36748
rect 73066 36720 73431 36748
rect 68782 36708 68788 36720
rect 50658 36652 51750 36680
rect 50658 36640 50664 36652
rect 52716 36640 52722 36692
rect 52774 36680 52780 36692
rect 57684 36680 57690 36692
rect 52774 36652 57690 36680
rect 52774 36640 52780 36652
rect 57684 36640 57690 36652
rect 57742 36640 57748 36692
rect 58420 36640 58426 36692
rect 58478 36680 58484 36692
rect 68908 36680 68914 36692
rect 58478 36652 68914 36680
rect 58478 36640 58484 36652
rect 68908 36640 68914 36652
rect 68966 36640 68972 36692
rect 73066 36689 73094 36720
rect 73419 36717 73431 36720
rect 73465 36717 73477 36751
rect 73419 36711 73477 36717
rect 73603 36751 73661 36757
rect 73603 36717 73615 36751
rect 73649 36748 73661 36751
rect 74063 36751 74121 36757
rect 74063 36748 74075 36751
rect 73649 36720 74075 36748
rect 73649 36717 73661 36720
rect 73603 36711 73661 36717
rect 74063 36717 74075 36720
rect 74109 36748 74121 36751
rect 75995 36751 76053 36757
rect 75995 36748 76007 36751
rect 74109 36720 76007 36748
rect 74109 36717 74121 36720
rect 74063 36711 74121 36717
rect 75995 36717 76007 36720
rect 76041 36717 76053 36751
rect 75995 36711 76053 36717
rect 76271 36751 76329 36757
rect 76271 36717 76283 36751
rect 76317 36748 76329 36751
rect 76452 36748 76458 36760
rect 76317 36720 76458 36748
rect 76317 36717 76329 36720
rect 76271 36711 76329 36717
rect 73051 36683 73109 36689
rect 73051 36680 73063 36683
rect 69110 36652 73063 36680
rect 51796 36612 51802 36624
rect 50526 36584 51802 36612
rect 51796 36572 51802 36584
rect 51854 36572 51860 36624
rect 53271 36615 53329 36621
rect 53271 36581 53283 36615
rect 53317 36612 53329 36615
rect 53360 36612 53366 36624
rect 53317 36584 53366 36612
rect 53317 36581 53329 36584
rect 53271 36575 53329 36581
rect 53360 36572 53366 36584
rect 53418 36572 53424 36624
rect 53452 36572 53458 36624
rect 53510 36612 53516 36624
rect 57776 36612 57782 36624
rect 53510 36584 57782 36612
rect 53510 36572 53516 36584
rect 57776 36572 57782 36584
rect 57834 36572 57840 36624
rect 58604 36572 58610 36624
rect 58662 36612 58668 36624
rect 62379 36615 62437 36621
rect 62379 36612 62391 36615
rect 58662 36584 62391 36612
rect 58662 36572 58668 36584
rect 62379 36581 62391 36584
rect 62425 36581 62437 36615
rect 62379 36575 62437 36581
rect 62468 36572 62474 36624
rect 62526 36612 62532 36624
rect 65964 36612 65970 36624
rect 62526 36584 65970 36612
rect 62526 36572 62532 36584
rect 65964 36572 65970 36584
rect 66022 36612 66028 36624
rect 69110 36612 69138 36652
rect 73051 36649 73063 36652
rect 73097 36649 73109 36683
rect 76286 36680 76314 36711
rect 76452 36708 76458 36720
rect 76510 36708 76516 36760
rect 79212 36748 79218 36760
rect 79173 36720 79218 36748
rect 79212 36708 79218 36720
rect 79270 36708 79276 36760
rect 80886 36748 80914 36847
rect 83996 36844 84002 36896
rect 84054 36884 84060 36896
rect 84054 36856 85330 36884
rect 84054 36844 84060 36856
rect 84456 36776 84462 36828
rect 84514 36816 84520 36828
rect 85302 36825 85330 36856
rect 85468 36844 85474 36896
rect 85526 36884 85532 36896
rect 88504 36884 88510 36896
rect 85526 36856 88510 36884
rect 85526 36844 85532 36856
rect 88504 36844 88510 36856
rect 88562 36884 88568 36896
rect 88562 36856 88918 36884
rect 88562 36844 88568 36856
rect 84827 36819 84885 36825
rect 84827 36816 84839 36819
rect 84514 36788 84839 36816
rect 84514 36776 84520 36788
rect 84827 36785 84839 36788
rect 84873 36785 84885 36819
rect 84827 36779 84885 36785
rect 85287 36819 85345 36825
rect 85287 36785 85299 36819
rect 85333 36816 85345 36819
rect 86299 36819 86357 36825
rect 86299 36816 86311 36819
rect 85333 36788 86311 36816
rect 85333 36785 85345 36788
rect 85287 36779 85345 36785
rect 86299 36785 86311 36788
rect 86345 36816 86357 36819
rect 86572 36816 86578 36828
rect 86345 36788 86578 36816
rect 86345 36785 86357 36788
rect 86299 36779 86357 36785
rect 86572 36776 86578 36788
rect 86630 36776 86636 36828
rect 80963 36751 81021 36757
rect 80963 36748 80975 36751
rect 80886 36720 80975 36748
rect 80963 36717 80975 36720
rect 81009 36717 81021 36751
rect 80963 36711 81021 36717
rect 82708 36708 82714 36760
rect 82766 36748 82772 36760
rect 85468 36748 85474 36760
rect 82766 36720 85474 36748
rect 82766 36708 82772 36720
rect 85468 36708 85474 36720
rect 85526 36708 85532 36760
rect 85839 36751 85897 36757
rect 85839 36717 85851 36751
rect 85885 36717 85897 36751
rect 85839 36711 85897 36717
rect 73051 36643 73109 36649
rect 73250 36652 76314 36680
rect 85854 36680 85882 36711
rect 85928 36708 85934 36760
rect 85986 36748 85992 36760
rect 88780 36748 88786 36760
rect 85986 36720 86031 36748
rect 88741 36720 88786 36748
rect 85986 36708 85992 36720
rect 88780 36708 88786 36720
rect 88838 36708 88844 36760
rect 88890 36748 88918 36856
rect 88967 36751 89025 36757
rect 88967 36748 88979 36751
rect 88890 36720 88979 36748
rect 88967 36717 88979 36720
rect 89013 36717 89025 36751
rect 88967 36711 89025 36717
rect 89240 36708 89246 36760
rect 89298 36757 89304 36760
rect 89298 36751 89347 36757
rect 89298 36717 89301 36751
rect 89335 36717 89347 36751
rect 89516 36748 89522 36760
rect 89477 36720 89522 36748
rect 89298 36711 89347 36717
rect 89298 36708 89304 36711
rect 89516 36708 89522 36720
rect 89574 36708 89580 36760
rect 86020 36680 86026 36692
rect 85854 36652 86026 36680
rect 73250 36621 73278 36652
rect 86020 36640 86026 36652
rect 86078 36680 86084 36692
rect 86388 36680 86394 36692
rect 86078 36652 86394 36680
rect 86078 36640 86084 36652
rect 86388 36640 86394 36652
rect 86446 36640 86452 36692
rect 66022 36584 69138 36612
rect 73235 36615 73293 36621
rect 66022 36572 66028 36584
rect 73235 36581 73247 36615
rect 73281 36581 73293 36615
rect 73235 36575 73293 36581
rect 76087 36615 76145 36621
rect 76087 36581 76099 36615
rect 76133 36612 76145 36615
rect 76728 36612 76734 36624
rect 76133 36584 76734 36612
rect 76133 36581 76145 36584
rect 76087 36575 76145 36581
rect 76728 36572 76734 36584
rect 76786 36572 76792 36624
rect 81147 36615 81205 36621
rect 81147 36581 81159 36615
rect 81193 36612 81205 36615
rect 83076 36612 83082 36624
rect 81193 36584 83082 36612
rect 81193 36581 81205 36584
rect 81147 36575 81205 36581
rect 83076 36572 83082 36584
rect 83134 36572 83140 36624
rect 85284 36572 85290 36624
rect 85342 36612 85348 36624
rect 85928 36612 85934 36624
rect 85342 36584 85934 36612
rect 85342 36572 85348 36584
rect 85928 36572 85934 36584
rect 85986 36612 85992 36624
rect 86115 36615 86173 36621
rect 86115 36612 86127 36615
rect 85986 36584 86127 36612
rect 85986 36572 85992 36584
rect 86115 36581 86127 36584
rect 86161 36581 86173 36615
rect 86115 36575 86173 36581
rect 538 36522 93642 36544
rect 538 36470 6344 36522
rect 6396 36470 6408 36522
rect 6460 36470 6472 36522
rect 6524 36470 6536 36522
rect 6588 36470 11672 36522
rect 11724 36470 11736 36522
rect 11788 36470 11800 36522
rect 11852 36470 11864 36522
rect 11916 36470 17000 36522
rect 17052 36470 17064 36522
rect 17116 36470 17128 36522
rect 17180 36470 17192 36522
rect 17244 36470 22328 36522
rect 22380 36470 22392 36522
rect 22444 36470 22456 36522
rect 22508 36470 22520 36522
rect 22572 36470 27656 36522
rect 27708 36470 27720 36522
rect 27772 36470 27784 36522
rect 27836 36470 27848 36522
rect 27900 36470 32984 36522
rect 33036 36470 33048 36522
rect 33100 36470 33112 36522
rect 33164 36470 33176 36522
rect 33228 36470 38312 36522
rect 38364 36470 38376 36522
rect 38428 36470 38440 36522
rect 38492 36470 38504 36522
rect 38556 36470 43640 36522
rect 43692 36470 43704 36522
rect 43756 36470 43768 36522
rect 43820 36470 43832 36522
rect 43884 36470 48968 36522
rect 49020 36470 49032 36522
rect 49084 36470 49096 36522
rect 49148 36470 49160 36522
rect 49212 36470 54296 36522
rect 54348 36470 54360 36522
rect 54412 36470 54424 36522
rect 54476 36470 54488 36522
rect 54540 36470 59624 36522
rect 59676 36470 59688 36522
rect 59740 36470 59752 36522
rect 59804 36470 59816 36522
rect 59868 36470 64952 36522
rect 65004 36470 65016 36522
rect 65068 36470 65080 36522
rect 65132 36470 65144 36522
rect 65196 36470 70280 36522
rect 70332 36470 70344 36522
rect 70396 36470 70408 36522
rect 70460 36470 70472 36522
rect 70524 36470 75608 36522
rect 75660 36470 75672 36522
rect 75724 36470 75736 36522
rect 75788 36470 75800 36522
rect 75852 36470 80936 36522
rect 80988 36470 81000 36522
rect 81052 36470 81064 36522
rect 81116 36470 81128 36522
rect 81180 36470 86264 36522
rect 86316 36470 86328 36522
rect 86380 36470 86392 36522
rect 86444 36470 86456 36522
rect 86508 36470 91592 36522
rect 91644 36470 91656 36522
rect 91708 36470 91720 36522
rect 91772 36470 91784 36522
rect 91836 36470 93642 36522
rect 538 36448 93642 36470
rect 2484 36408 2490 36420
rect 2397 36380 2490 36408
rect 2484 36368 2490 36380
rect 2542 36408 2548 36420
rect 3404 36408 3410 36420
rect 2542 36380 3410 36408
rect 2542 36368 2548 36380
rect 3404 36368 3410 36380
rect 3462 36368 3468 36420
rect 4968 36368 4974 36420
rect 5026 36408 5032 36420
rect 7363 36411 7421 36417
rect 7363 36408 7375 36411
rect 5026 36380 7375 36408
rect 5026 36368 5032 36380
rect 5538 36281 5566 36380
rect 7363 36377 7375 36380
rect 7409 36408 7421 36411
rect 7452 36408 7458 36420
rect 7409 36380 7458 36408
rect 7409 36377 7421 36380
rect 7363 36371 7421 36377
rect 7452 36368 7458 36380
rect 7510 36368 7516 36420
rect 9752 36408 9758 36420
rect 9713 36380 9758 36408
rect 9752 36368 9758 36380
rect 9810 36368 9816 36420
rect 14904 36368 14910 36420
rect 14962 36408 14968 36420
rect 15459 36411 15517 36417
rect 15459 36408 15471 36411
rect 14962 36380 15471 36408
rect 14962 36368 14968 36380
rect 15459 36377 15471 36380
rect 15505 36377 15517 36411
rect 15459 36371 15517 36377
rect 17664 36368 17670 36420
rect 17722 36408 17728 36420
rect 17851 36411 17909 36417
rect 17851 36408 17863 36411
rect 17722 36380 17863 36408
rect 17722 36368 17728 36380
rect 17851 36377 17863 36380
rect 17897 36377 17909 36411
rect 29259 36411 29317 36417
rect 29259 36408 29271 36411
rect 17851 36371 17909 36377
rect 27434 36380 29271 36408
rect 7179 36343 7237 36349
rect 7179 36309 7191 36343
rect 7225 36340 7237 36343
rect 7225 36312 12190 36340
rect 7225 36309 7237 36312
rect 7179 36303 7237 36309
rect 5523 36275 5581 36281
rect 5523 36241 5535 36275
rect 5569 36241 5581 36275
rect 5796 36272 5802 36284
rect 5757 36244 5802 36272
rect 5523 36235 5581 36241
rect 5796 36232 5802 36244
rect 5854 36232 5860 36284
rect 9571 36275 9629 36281
rect 9571 36241 9583 36275
rect 9617 36272 9629 36275
rect 10212 36272 10218 36284
rect 9617 36244 10218 36272
rect 9617 36241 9629 36244
rect 9571 36235 9629 36241
rect 10212 36232 10218 36244
rect 10270 36232 10276 36284
rect 10488 36232 10494 36284
rect 10546 36272 10552 36284
rect 11500 36272 11506 36284
rect 10546 36244 11506 36272
rect 10546 36232 10552 36244
rect 11500 36232 11506 36244
rect 11558 36272 11564 36284
rect 12162 36281 12190 36312
rect 11595 36275 11653 36281
rect 11595 36272 11607 36275
rect 11558 36244 11607 36272
rect 11558 36232 11564 36244
rect 11595 36241 11607 36244
rect 11641 36241 11653 36275
rect 11595 36235 11653 36241
rect 11779 36275 11837 36281
rect 11779 36241 11791 36275
rect 11825 36241 11837 36275
rect 11779 36235 11837 36241
rect 12147 36275 12205 36281
rect 12147 36241 12159 36275
rect 12193 36241 12205 36275
rect 12147 36235 12205 36241
rect 15643 36275 15701 36281
rect 15643 36241 15655 36275
rect 15689 36272 15701 36275
rect 16100 36272 16106 36284
rect 15689 36244 16106 36272
rect 15689 36241 15701 36244
rect 15643 36235 15701 36241
rect 1843 36207 1901 36213
rect 1843 36173 1855 36207
rect 1889 36204 1901 36207
rect 2668 36204 2674 36216
rect 1889 36176 2674 36204
rect 1889 36173 1901 36176
rect 1843 36167 1901 36173
rect 2668 36164 2674 36176
rect 2726 36164 2732 36216
rect 11794 36136 11822 36235
rect 16100 36232 16106 36244
rect 16158 36232 16164 36284
rect 17866 36272 17894 36371
rect 24030 36312 25806 36340
rect 24030 36284 24058 36312
rect 18955 36275 19013 36281
rect 18955 36272 18967 36275
rect 17866 36244 18967 36272
rect 18955 36241 18967 36244
rect 19001 36241 19013 36275
rect 18955 36235 19013 36241
rect 21347 36275 21405 36281
rect 21347 36241 21359 36275
rect 21393 36272 21405 36275
rect 21528 36272 21534 36284
rect 21393 36244 21534 36272
rect 21393 36241 21405 36244
rect 21347 36235 21405 36241
rect 21528 36232 21534 36244
rect 21586 36272 21592 36284
rect 21623 36275 21681 36281
rect 21623 36272 21635 36275
rect 21586 36244 21635 36272
rect 21586 36232 21592 36244
rect 21623 36241 21635 36244
rect 21669 36241 21681 36275
rect 21623 36235 21681 36241
rect 23463 36275 23521 36281
rect 23463 36241 23475 36275
rect 23509 36272 23521 36275
rect 24012 36272 24018 36284
rect 23509 36244 24018 36272
rect 23509 36241 23521 36244
rect 23463 36235 23521 36241
rect 24012 36232 24018 36244
rect 24070 36232 24076 36284
rect 24199 36275 24257 36281
rect 24199 36241 24211 36275
rect 24245 36272 24257 36275
rect 25668 36272 25674 36284
rect 24245 36244 25674 36272
rect 24245 36241 24257 36244
rect 24199 36235 24257 36241
rect 25668 36232 25674 36244
rect 25726 36232 25732 36284
rect 12052 36204 12058 36216
rect 12013 36176 12058 36204
rect 12052 36164 12058 36176
rect 12110 36164 12116 36216
rect 16471 36207 16529 36213
rect 16471 36204 16483 36207
rect 16302 36176 16483 36204
rect 12604 36136 12610 36148
rect 11794 36108 12610 36136
rect 12604 36096 12610 36108
rect 12662 36096 12668 36148
rect 11411 36071 11469 36077
rect 11411 36037 11423 36071
rect 11457 36068 11469 36071
rect 12144 36068 12150 36080
rect 11457 36040 12150 36068
rect 11457 36037 11469 36040
rect 11411 36031 11469 36037
rect 12144 36028 12150 36040
rect 12202 36028 12208 36080
rect 15548 36028 15554 36080
rect 15606 36068 15612 36080
rect 16302 36077 16330 36176
rect 16471 36173 16483 36176
rect 16517 36173 16529 36207
rect 16744 36204 16750 36216
rect 16705 36176 16750 36204
rect 16471 36167 16529 36173
rect 16744 36164 16750 36176
rect 16802 36164 16808 36216
rect 23371 36207 23429 36213
rect 23371 36173 23383 36207
rect 23417 36173 23429 36207
rect 25778 36204 25806 36312
rect 27434 36281 27462 36380
rect 29259 36377 29271 36380
rect 29305 36408 29317 36411
rect 29348 36408 29354 36420
rect 29305 36380 29354 36408
rect 29305 36377 29317 36380
rect 29259 36371 29317 36377
rect 29348 36368 29354 36380
rect 29406 36368 29412 36420
rect 29900 36368 29906 36420
rect 29958 36408 29964 36420
rect 29958 36380 64998 36408
rect 29958 36368 29964 36380
rect 29072 36300 29078 36352
rect 29130 36340 29136 36352
rect 37447 36343 37505 36349
rect 37447 36340 37459 36343
rect 29130 36312 37459 36340
rect 29130 36300 29136 36312
rect 37447 36309 37459 36312
rect 37493 36340 37505 36343
rect 39192 36340 39198 36352
rect 37493 36312 37674 36340
rect 39153 36312 39198 36340
rect 37493 36309 37505 36312
rect 37447 36303 37505 36309
rect 27419 36275 27477 36281
rect 27419 36241 27431 36275
rect 27465 36241 27477 36275
rect 32108 36272 32114 36284
rect 27419 36235 27477 36241
rect 27526 36244 32114 36272
rect 27526 36204 27554 36244
rect 32108 36232 32114 36244
rect 32166 36232 32172 36284
rect 32571 36275 32629 36281
rect 32571 36241 32583 36275
rect 32617 36241 32629 36275
rect 32571 36235 32629 36241
rect 32939 36275 32997 36281
rect 32939 36241 32951 36275
rect 32985 36272 32997 36275
rect 33491 36275 33549 36281
rect 33491 36272 33503 36275
rect 32985 36244 33503 36272
rect 32985 36241 32997 36244
rect 32939 36235 32997 36241
rect 33491 36241 33503 36244
rect 33537 36241 33549 36275
rect 33491 36235 33549 36241
rect 25778 36176 27554 36204
rect 27695 36207 27753 36213
rect 23371 36167 23429 36173
rect 27695 36173 27707 36207
rect 27741 36204 27753 36207
rect 28060 36204 28066 36216
rect 27741 36176 28066 36204
rect 27741 36173 27753 36176
rect 27695 36167 27753 36173
rect 23187 36139 23245 36145
rect 23187 36105 23199 36139
rect 23233 36136 23245 36139
rect 23386 36136 23414 36167
rect 28060 36164 28066 36176
rect 28118 36164 28124 36216
rect 28336 36164 28342 36216
rect 28394 36204 28400 36216
rect 32203 36207 32261 36213
rect 32203 36204 32215 36207
rect 28394 36176 32215 36204
rect 28394 36164 28400 36176
rect 32203 36173 32215 36176
rect 32249 36204 32261 36207
rect 32586 36204 32614 36235
rect 32844 36204 32850 36216
rect 32249 36176 32614 36204
rect 32805 36176 32850 36204
rect 32249 36173 32261 36176
rect 32203 36167 32261 36173
rect 32844 36164 32850 36176
rect 32902 36164 32908 36216
rect 27048 36136 27054 36148
rect 23233 36108 27054 36136
rect 23233 36105 23245 36108
rect 23187 36099 23245 36105
rect 27048 36096 27054 36108
rect 27106 36096 27112 36148
rect 29900 36136 29906 36148
rect 28354 36108 29906 36136
rect 16287 36071 16345 36077
rect 16287 36068 16299 36071
rect 15606 36040 16299 36068
rect 15606 36028 15612 36040
rect 16287 36037 16299 36040
rect 16333 36037 16345 36071
rect 16287 36031 16345 36037
rect 19047 36071 19105 36077
rect 19047 36037 19059 36071
rect 19093 36068 19105 36071
rect 20148 36068 20154 36080
rect 19093 36040 20154 36068
rect 19093 36037 19105 36040
rect 19047 36031 19105 36037
rect 20148 36028 20154 36040
rect 20206 36028 20212 36080
rect 21439 36071 21497 36077
rect 21439 36037 21451 36071
rect 21485 36068 21497 36071
rect 21528 36068 21534 36080
rect 21485 36040 21534 36068
rect 21485 36037 21497 36040
rect 21439 36031 21497 36037
rect 21528 36028 21534 36040
rect 21586 36028 21592 36080
rect 23368 36028 23374 36080
rect 23426 36068 23432 36080
rect 24475 36071 24533 36077
rect 24475 36068 24487 36071
rect 23426 36040 24487 36068
rect 23426 36028 23432 36040
rect 24475 36037 24487 36040
rect 24521 36037 24533 36071
rect 24475 36031 24533 36037
rect 24564 36028 24570 36080
rect 24622 36068 24628 36080
rect 28354 36068 28382 36108
rect 29900 36096 29906 36108
rect 29958 36096 29964 36148
rect 32954 36136 32982 36235
rect 33580 36232 33586 36284
rect 33638 36272 33644 36284
rect 37646 36281 37674 36312
rect 39192 36300 39198 36312
rect 39250 36300 39256 36352
rect 40480 36340 40486 36352
rect 39302 36312 40158 36340
rect 33675 36275 33733 36281
rect 33675 36272 33687 36275
rect 33638 36244 33687 36272
rect 33638 36232 33644 36244
rect 33675 36241 33687 36244
rect 33721 36272 33733 36275
rect 34319 36275 34377 36281
rect 34319 36272 34331 36275
rect 33721 36244 34331 36272
rect 33721 36241 33733 36244
rect 33675 36235 33733 36241
rect 34319 36241 34331 36244
rect 34365 36272 34377 36275
rect 37631 36275 37689 36281
rect 34365 36244 35374 36272
rect 34365 36241 34377 36244
rect 34319 36235 34377 36241
rect 34043 36207 34101 36213
rect 34043 36173 34055 36207
rect 34089 36204 34101 36207
rect 35052 36204 35058 36216
rect 34089 36176 35058 36204
rect 34089 36173 34101 36176
rect 34043 36167 34101 36173
rect 35052 36164 35058 36176
rect 35110 36164 35116 36216
rect 35346 36204 35374 36244
rect 37631 36241 37643 36275
rect 37677 36272 37689 36275
rect 39103 36275 39161 36281
rect 37677 36244 38870 36272
rect 37677 36241 37689 36244
rect 37631 36235 37689 36241
rect 38180 36204 38186 36216
rect 35346 36176 38186 36204
rect 38180 36164 38186 36176
rect 38238 36164 38244 36216
rect 34500 36136 34506 36148
rect 32310 36108 34506 36136
rect 28980 36068 28986 36080
rect 24622 36040 28382 36068
rect 28941 36040 28986 36068
rect 24622 36028 24628 36040
rect 28980 36028 28986 36040
rect 29038 36028 29044 36080
rect 29256 36028 29262 36080
rect 29314 36068 29320 36080
rect 32310 36068 32338 36108
rect 34500 36096 34506 36108
rect 34558 36096 34564 36148
rect 37628 36096 37634 36148
rect 37686 36136 37692 36148
rect 37815 36139 37873 36145
rect 37815 36136 37827 36139
rect 37686 36108 37827 36136
rect 37686 36096 37692 36108
rect 37815 36105 37827 36108
rect 37861 36105 37873 36139
rect 38842 36136 38870 36244
rect 39103 36241 39115 36275
rect 39149 36272 39161 36275
rect 39302 36272 39330 36312
rect 39836 36272 39842 36284
rect 39149 36244 39330 36272
rect 39797 36244 39842 36272
rect 39149 36241 39161 36244
rect 39103 36235 39161 36241
rect 39836 36232 39842 36244
rect 39894 36232 39900 36284
rect 40130 36216 40158 36312
rect 40222 36312 40486 36340
rect 40222 36281 40250 36312
rect 40480 36300 40486 36312
rect 40538 36300 40544 36352
rect 40572 36300 40578 36352
rect 40630 36340 40636 36352
rect 49312 36340 49318 36352
rect 40630 36312 49318 36340
rect 40630 36300 40636 36312
rect 49312 36300 49318 36312
rect 49370 36300 49376 36352
rect 51336 36300 51342 36352
rect 51394 36340 51400 36352
rect 52256 36340 52262 36352
rect 51394 36312 52262 36340
rect 51394 36300 51400 36312
rect 52256 36300 52262 36312
rect 52314 36300 52320 36352
rect 61456 36300 61462 36352
rect 61514 36340 61520 36352
rect 61514 36312 64906 36340
rect 61514 36300 61520 36312
rect 40207 36275 40265 36281
rect 40207 36241 40219 36275
rect 40253 36241 40265 36275
rect 45356 36272 45362 36284
rect 45317 36244 45362 36272
rect 40207 36235 40265 36241
rect 45356 36232 45362 36244
rect 45414 36272 45420 36284
rect 45543 36275 45601 36281
rect 45543 36272 45555 36275
rect 45414 36244 45555 36272
rect 45414 36232 45420 36244
rect 45543 36241 45555 36244
rect 45589 36241 45601 36275
rect 45543 36235 45601 36241
rect 45632 36232 45638 36284
rect 45690 36272 45696 36284
rect 45690 36244 45735 36272
rect 45834 36244 51566 36272
rect 45690 36232 45696 36244
rect 38919 36207 38977 36213
rect 38919 36173 38931 36207
rect 38965 36204 38977 36207
rect 39652 36204 39658 36216
rect 38965 36176 39658 36204
rect 38965 36173 38977 36176
rect 38919 36167 38977 36173
rect 39652 36164 39658 36176
rect 39710 36164 39716 36216
rect 40112 36204 40118 36216
rect 40025 36176 40118 36204
rect 40112 36164 40118 36176
rect 40170 36164 40176 36216
rect 40222 36176 43010 36204
rect 40222 36136 40250 36176
rect 38842 36108 40250 36136
rect 42982 36136 43010 36176
rect 45080 36164 45086 36216
rect 45138 36204 45144 36216
rect 45834 36204 45862 36244
rect 45138 36176 45862 36204
rect 45138 36164 45144 36176
rect 48852 36164 48858 36216
rect 48910 36204 48916 36216
rect 50971 36207 51029 36213
rect 50971 36204 50983 36207
rect 48910 36176 50983 36204
rect 48910 36164 48916 36176
rect 50971 36173 50983 36176
rect 51017 36173 51029 36207
rect 50971 36167 51029 36173
rect 51336 36164 51342 36216
rect 51394 36204 51400 36216
rect 51431 36207 51489 36213
rect 51431 36204 51443 36207
rect 51394 36176 51443 36204
rect 51394 36164 51400 36176
rect 51431 36173 51443 36176
rect 51477 36173 51489 36207
rect 51538 36204 51566 36244
rect 51612 36232 51618 36284
rect 51670 36272 51676 36284
rect 51983 36275 52041 36281
rect 51670 36244 51715 36272
rect 51670 36232 51676 36244
rect 51983 36241 51995 36275
rect 52029 36272 52041 36275
rect 52716 36272 52722 36284
rect 52029 36244 52722 36272
rect 52029 36241 52041 36244
rect 51983 36235 52041 36241
rect 52716 36232 52722 36244
rect 52774 36232 52780 36284
rect 53360 36232 53366 36284
rect 53418 36272 53424 36284
rect 54007 36275 54065 36281
rect 54007 36272 54019 36275
rect 53418 36244 54019 36272
rect 53418 36232 53424 36244
rect 54007 36241 54019 36244
rect 54053 36241 54065 36275
rect 56764 36272 56770 36284
rect 56725 36244 56770 36272
rect 54007 36235 54065 36241
rect 56764 36232 56770 36244
rect 56822 36232 56828 36284
rect 61824 36272 61830 36284
rect 61785 36244 61830 36272
rect 61824 36232 61830 36244
rect 61882 36232 61888 36284
rect 62287 36275 62345 36281
rect 62287 36272 62299 36275
rect 61934 36244 62299 36272
rect 51888 36204 51894 36216
rect 51538 36176 51750 36204
rect 51849 36176 51894 36204
rect 51431 36167 51489 36173
rect 51520 36136 51526 36148
rect 42982 36108 51526 36136
rect 37815 36099 37873 36105
rect 51520 36096 51526 36108
rect 51578 36096 51584 36148
rect 51612 36096 51618 36148
rect 51670 36096 51676 36148
rect 51722 36136 51750 36176
rect 51888 36164 51894 36176
rect 51946 36164 51952 36216
rect 52072 36164 52078 36216
rect 52130 36204 52136 36216
rect 54099 36207 54157 36213
rect 54099 36204 54111 36207
rect 52130 36176 54111 36204
rect 52130 36164 52136 36176
rect 54099 36173 54111 36176
rect 54145 36173 54157 36207
rect 54099 36167 54157 36173
rect 56120 36164 56126 36216
rect 56178 36204 56184 36216
rect 56399 36207 56457 36213
rect 56399 36204 56411 36207
rect 56178 36176 56411 36204
rect 56178 36164 56184 36176
rect 56399 36173 56411 36176
rect 56445 36204 56457 36207
rect 56491 36207 56549 36213
rect 56491 36204 56503 36207
rect 56445 36176 56503 36204
rect 56445 36173 56457 36176
rect 56399 36167 56457 36173
rect 56491 36173 56503 36176
rect 56537 36204 56549 36207
rect 57132 36204 57138 36216
rect 56537 36176 57138 36204
rect 56537 36173 56549 36176
rect 56491 36167 56549 36173
rect 57132 36164 57138 36176
rect 57190 36164 57196 36216
rect 61548 36204 61554 36216
rect 57426 36176 61554 36204
rect 51722 36108 52854 36136
rect 29314 36040 32338 36068
rect 32387 36071 32445 36077
rect 29314 36028 29320 36040
rect 32387 36037 32399 36071
rect 32433 36068 32445 36071
rect 33948 36068 33954 36080
rect 32433 36040 33954 36068
rect 32433 36037 32445 36040
rect 32387 36031 32445 36037
rect 33948 36028 33954 36040
rect 34006 36068 34012 36080
rect 34132 36068 34138 36080
rect 34006 36040 34138 36068
rect 34006 36028 34012 36040
rect 34132 36028 34138 36040
rect 34190 36028 34196 36080
rect 39836 36028 39842 36080
rect 39894 36068 39900 36080
rect 40667 36071 40725 36077
rect 40667 36068 40679 36071
rect 39894 36040 40679 36068
rect 39894 36028 39900 36040
rect 40667 36037 40679 36040
rect 40713 36037 40725 36071
rect 40667 36031 40725 36037
rect 42872 36028 42878 36080
rect 42930 36068 42936 36080
rect 48392 36068 48398 36080
rect 42930 36040 48398 36068
rect 42930 36028 42936 36040
rect 48392 36028 48398 36040
rect 48450 36028 48456 36080
rect 51630 36068 51658 36096
rect 52348 36068 52354 36080
rect 51630 36040 52354 36068
rect 52348 36028 52354 36040
rect 52406 36028 52412 36080
rect 52535 36071 52593 36077
rect 52535 36037 52547 36071
rect 52581 36068 52593 36071
rect 52716 36068 52722 36080
rect 52581 36040 52722 36068
rect 52581 36037 52593 36040
rect 52535 36031 52593 36037
rect 52716 36028 52722 36040
rect 52774 36028 52780 36080
rect 52826 36068 52854 36108
rect 57426 36068 57454 36176
rect 61548 36164 61554 36176
rect 61606 36164 61612 36216
rect 61643 36207 61701 36213
rect 61643 36173 61655 36207
rect 61689 36173 61701 36207
rect 61643 36167 61701 36173
rect 58052 36136 58058 36148
rect 57965 36108 58058 36136
rect 58052 36096 58058 36108
rect 58110 36136 58116 36148
rect 61456 36136 61462 36148
rect 58110 36108 61462 36136
rect 58110 36096 58116 36108
rect 61456 36096 61462 36108
rect 61514 36096 61520 36148
rect 61658 36136 61686 36167
rect 61732 36164 61738 36216
rect 61790 36204 61796 36216
rect 61934 36204 61962 36244
rect 62287 36241 62299 36244
rect 62333 36241 62345 36275
rect 62287 36235 62345 36241
rect 62379 36275 62437 36281
rect 62379 36241 62391 36275
rect 62425 36272 62437 36275
rect 63296 36272 63302 36284
rect 62425 36244 63302 36272
rect 62425 36241 62437 36244
rect 62379 36235 62437 36241
rect 63296 36232 63302 36244
rect 63354 36232 63360 36284
rect 61790 36176 61962 36204
rect 61790 36164 61796 36176
rect 62560 36136 62566 36148
rect 61658 36108 62566 36136
rect 52826 36040 57454 36068
rect 59064 36028 59070 36080
rect 59122 36068 59128 36080
rect 61658 36068 61686 36108
rect 62560 36096 62566 36108
rect 62618 36096 62624 36148
rect 64878 36136 64906 36312
rect 64970 36204 64998 36380
rect 65596 36368 65602 36420
rect 65654 36408 65660 36420
rect 65691 36411 65749 36417
rect 65691 36408 65703 36411
rect 65654 36380 65703 36408
rect 65654 36368 65660 36380
rect 65691 36377 65703 36380
rect 65737 36377 65749 36411
rect 65691 36371 65749 36377
rect 66059 36411 66117 36417
rect 66059 36377 66071 36411
rect 66105 36408 66117 36411
rect 68172 36408 68178 36420
rect 66105 36380 68178 36408
rect 66105 36377 66117 36380
rect 66059 36371 66117 36377
rect 65706 36272 65734 36371
rect 68172 36368 68178 36380
rect 68230 36368 68236 36420
rect 80687 36411 80745 36417
rect 80687 36377 80699 36411
rect 80733 36408 80745 36411
rect 82156 36408 82162 36420
rect 80733 36380 82162 36408
rect 80733 36377 80745 36380
rect 80687 36371 80745 36377
rect 82156 36368 82162 36380
rect 82214 36368 82220 36420
rect 82343 36411 82401 36417
rect 82343 36377 82355 36411
rect 82389 36408 82401 36411
rect 82524 36408 82530 36420
rect 82389 36380 82530 36408
rect 82389 36377 82401 36380
rect 82343 36371 82401 36377
rect 82524 36368 82530 36380
rect 82582 36368 82588 36420
rect 88228 36368 88234 36420
rect 88286 36408 88292 36420
rect 88415 36411 88473 36417
rect 88415 36408 88427 36411
rect 88286 36380 88427 36408
rect 88286 36368 88292 36380
rect 88415 36377 88427 36380
rect 88461 36408 88473 36411
rect 88461 36380 88642 36408
rect 88461 36377 88473 36380
rect 88415 36371 88473 36377
rect 73526 36312 74106 36340
rect 65875 36275 65933 36281
rect 65875 36272 65887 36275
rect 65706 36244 65887 36272
rect 65875 36241 65887 36244
rect 65921 36241 65933 36275
rect 67715 36275 67773 36281
rect 65875 36235 65933 36241
rect 65982 36244 67574 36272
rect 65982 36204 66010 36244
rect 64970 36176 66010 36204
rect 67439 36207 67497 36213
rect 67439 36173 67451 36207
rect 67485 36173 67497 36207
rect 67546 36204 67574 36244
rect 67715 36241 67727 36275
rect 67761 36272 67773 36275
rect 69184 36272 69190 36284
rect 67761 36244 69190 36272
rect 67761 36241 67773 36244
rect 67715 36235 67773 36241
rect 69184 36232 69190 36244
rect 69242 36232 69248 36284
rect 73324 36272 73330 36284
rect 73285 36244 73330 36272
rect 73324 36232 73330 36244
rect 73382 36232 73388 36284
rect 73526 36281 73554 36312
rect 73511 36275 73569 36281
rect 73511 36241 73523 36275
rect 73557 36241 73569 36275
rect 73511 36235 73569 36241
rect 73600 36232 73606 36284
rect 73658 36272 73664 36284
rect 74078 36281 74106 36312
rect 73971 36275 74029 36281
rect 73971 36272 73983 36275
rect 73658 36244 73983 36272
rect 73658 36232 73664 36244
rect 73971 36241 73983 36244
rect 74017 36241 74029 36275
rect 73971 36235 74029 36241
rect 74063 36275 74121 36281
rect 74063 36241 74075 36275
rect 74109 36272 74121 36275
rect 74152 36272 74158 36284
rect 74109 36244 74158 36272
rect 74109 36241 74121 36244
rect 74063 36235 74121 36241
rect 74152 36232 74158 36244
rect 74210 36272 74216 36284
rect 75256 36272 75262 36284
rect 74210 36244 75262 36272
rect 74210 36232 74216 36244
rect 75256 36232 75262 36244
rect 75314 36232 75320 36284
rect 80503 36275 80561 36281
rect 80503 36272 80515 36275
rect 80334 36244 80515 36272
rect 69644 36204 69650 36216
rect 67546 36176 69650 36204
rect 67439 36167 67497 36173
rect 66516 36136 66522 36148
rect 64878 36108 66522 36136
rect 66516 36096 66522 36108
rect 66574 36096 66580 36148
rect 59122 36040 61686 36068
rect 62839 36071 62897 36077
rect 59122 36028 59128 36040
rect 62839 36037 62851 36071
rect 62885 36068 62897 36071
rect 63020 36068 63026 36080
rect 62885 36040 63026 36068
rect 62885 36037 62897 36040
rect 62839 36031 62897 36037
rect 63020 36028 63026 36040
rect 63078 36028 63084 36080
rect 63204 36068 63210 36080
rect 63117 36040 63210 36068
rect 63204 36028 63210 36040
rect 63262 36068 63268 36080
rect 64124 36068 64130 36080
rect 63262 36040 64130 36068
rect 63262 36028 63268 36040
rect 64124 36028 64130 36040
rect 64182 36028 64188 36080
rect 67454 36068 67482 36167
rect 69644 36164 69650 36176
rect 69702 36164 69708 36216
rect 69187 36139 69245 36145
rect 69187 36136 69199 36139
rect 68834 36108 69199 36136
rect 68834 36068 68862 36108
rect 69187 36105 69199 36108
rect 69233 36136 69245 36139
rect 69368 36136 69374 36148
rect 69233 36108 69374 36136
rect 69233 36105 69245 36108
rect 69187 36099 69245 36105
rect 69368 36096 69374 36108
rect 69426 36096 69432 36148
rect 70104 36096 70110 36148
rect 70162 36136 70168 36148
rect 80334 36145 80362 36244
rect 80503 36241 80515 36244
rect 80549 36241 80561 36275
rect 82708 36272 82714 36284
rect 82669 36244 82714 36272
rect 80503 36235 80561 36241
rect 82708 36232 82714 36244
rect 82766 36232 82772 36284
rect 83076 36272 83082 36284
rect 82989 36244 83082 36272
rect 83076 36232 83082 36244
rect 83134 36272 83140 36284
rect 86020 36272 86026 36284
rect 83134 36244 86026 36272
rect 83134 36232 83140 36244
rect 86020 36232 86026 36244
rect 86078 36232 86084 36284
rect 88614 36281 88642 36380
rect 88890 36312 89378 36340
rect 88599 36275 88657 36281
rect 88599 36241 88611 36275
rect 88645 36241 88657 36275
rect 88599 36235 88657 36241
rect 88688 36232 88694 36284
rect 88746 36272 88752 36284
rect 88783 36275 88841 36281
rect 88783 36272 88795 36275
rect 88746 36244 88795 36272
rect 88746 36232 88752 36244
rect 88783 36241 88795 36244
rect 88829 36241 88841 36275
rect 88783 36235 88841 36241
rect 82524 36204 82530 36216
rect 82485 36176 82530 36204
rect 82524 36164 82530 36176
rect 82582 36164 82588 36216
rect 82987 36207 83045 36213
rect 82987 36173 82999 36207
rect 83033 36173 83045 36207
rect 88890 36204 88918 36312
rect 89350 36281 89378 36312
rect 89335 36275 89393 36281
rect 89335 36241 89347 36275
rect 89381 36241 89393 36275
rect 89516 36272 89522 36284
rect 89429 36244 89522 36272
rect 89335 36235 89393 36241
rect 89516 36232 89522 36244
rect 89574 36272 89580 36284
rect 91356 36272 91362 36284
rect 89574 36244 90482 36272
rect 91317 36244 91362 36272
rect 89574 36232 89580 36244
rect 82987 36167 83045 36173
rect 88246 36176 88918 36204
rect 80319 36139 80377 36145
rect 80319 36136 80331 36139
rect 70162 36108 80331 36136
rect 70162 36096 70168 36108
rect 80319 36105 80331 36108
rect 80365 36105 80377 36139
rect 80319 36099 80377 36105
rect 82708 36096 82714 36148
rect 82766 36136 82772 36148
rect 83002 36136 83030 36167
rect 82766 36108 83030 36136
rect 82766 36096 82772 36108
rect 69000 36068 69006 36080
rect 67454 36040 68862 36068
rect 68961 36040 69006 36068
rect 69000 36028 69006 36040
rect 69058 36028 69064 36080
rect 74520 36068 74526 36080
rect 74481 36040 74526 36068
rect 74520 36028 74526 36040
rect 74578 36028 74584 36080
rect 85652 36028 85658 36080
rect 85710 36068 85716 36080
rect 88246 36077 88274 36176
rect 90454 36148 90482 36244
rect 91356 36232 91362 36244
rect 91414 36232 91420 36284
rect 90436 36096 90442 36148
rect 90494 36136 90500 36148
rect 91451 36139 91509 36145
rect 91451 36136 91463 36139
rect 90494 36108 91463 36136
rect 90494 36096 90500 36108
rect 91451 36105 91463 36108
rect 91497 36105 91509 36139
rect 91451 36099 91509 36105
rect 88231 36071 88289 36077
rect 88231 36068 88243 36071
rect 85710 36040 88243 36068
rect 85710 36028 85716 36040
rect 88231 36037 88243 36040
rect 88277 36037 88289 36071
rect 88231 36031 88289 36037
rect 89795 36071 89853 36077
rect 89795 36037 89807 36071
rect 89841 36068 89853 36071
rect 90712 36068 90718 36080
rect 89841 36040 90718 36068
rect 89841 36037 89853 36040
rect 89795 36031 89853 36037
rect 90712 36028 90718 36040
rect 90770 36028 90776 36080
rect 538 35978 93642 36000
rect 538 35926 3680 35978
rect 3732 35926 3744 35978
rect 3796 35926 3808 35978
rect 3860 35926 3872 35978
rect 3924 35926 9008 35978
rect 9060 35926 9072 35978
rect 9124 35926 9136 35978
rect 9188 35926 9200 35978
rect 9252 35926 14336 35978
rect 14388 35926 14400 35978
rect 14452 35926 14464 35978
rect 14516 35926 14528 35978
rect 14580 35926 19664 35978
rect 19716 35926 19728 35978
rect 19780 35926 19792 35978
rect 19844 35926 19856 35978
rect 19908 35926 24992 35978
rect 25044 35926 25056 35978
rect 25108 35926 25120 35978
rect 25172 35926 25184 35978
rect 25236 35926 30320 35978
rect 30372 35926 30384 35978
rect 30436 35926 30448 35978
rect 30500 35926 30512 35978
rect 30564 35926 35648 35978
rect 35700 35926 35712 35978
rect 35764 35926 35776 35978
rect 35828 35926 35840 35978
rect 35892 35926 40976 35978
rect 41028 35926 41040 35978
rect 41092 35926 41104 35978
rect 41156 35926 41168 35978
rect 41220 35926 46304 35978
rect 46356 35926 46368 35978
rect 46420 35926 46432 35978
rect 46484 35926 46496 35978
rect 46548 35926 51632 35978
rect 51684 35926 51696 35978
rect 51748 35926 51760 35978
rect 51812 35926 51824 35978
rect 51876 35926 56960 35978
rect 57012 35926 57024 35978
rect 57076 35926 57088 35978
rect 57140 35926 57152 35978
rect 57204 35926 62288 35978
rect 62340 35926 62352 35978
rect 62404 35926 62416 35978
rect 62468 35926 62480 35978
rect 62532 35926 67616 35978
rect 67668 35926 67680 35978
rect 67732 35926 67744 35978
rect 67796 35926 67808 35978
rect 67860 35926 72944 35978
rect 72996 35926 73008 35978
rect 73060 35926 73072 35978
rect 73124 35926 73136 35978
rect 73188 35926 78272 35978
rect 78324 35926 78336 35978
rect 78388 35926 78400 35978
rect 78452 35926 78464 35978
rect 78516 35926 83600 35978
rect 83652 35926 83664 35978
rect 83716 35926 83728 35978
rect 83780 35926 83792 35978
rect 83844 35926 88928 35978
rect 88980 35926 88992 35978
rect 89044 35926 89056 35978
rect 89108 35926 89120 35978
rect 89172 35926 93642 35978
rect 538 35904 93642 35926
rect 16471 35867 16529 35873
rect 16471 35833 16483 35867
rect 16517 35864 16529 35867
rect 16744 35864 16750 35876
rect 16517 35836 16750 35864
rect 16517 35833 16529 35836
rect 16471 35827 16529 35833
rect 16744 35824 16750 35836
rect 16802 35824 16808 35876
rect 21255 35867 21313 35873
rect 21255 35833 21267 35867
rect 21301 35864 21313 35867
rect 21620 35864 21626 35876
rect 21301 35836 21626 35864
rect 21301 35833 21313 35836
rect 21255 35827 21313 35833
rect 10212 35756 10218 35808
rect 10270 35796 10276 35808
rect 17667 35799 17725 35805
rect 10270 35768 10810 35796
rect 10270 35756 10276 35768
rect 2668 35728 2674 35740
rect 2629 35700 2674 35728
rect 2668 35688 2674 35700
rect 2726 35688 2732 35740
rect 10399 35731 10457 35737
rect 10399 35697 10411 35731
rect 10445 35728 10457 35731
rect 10488 35728 10494 35740
rect 10445 35700 10494 35728
rect 10445 35697 10457 35700
rect 10399 35691 10457 35697
rect 10488 35688 10494 35700
rect 10546 35688 10552 35740
rect 2395 35663 2453 35669
rect 2395 35629 2407 35663
rect 2441 35660 2453 35663
rect 10307 35663 10365 35669
rect 2441 35632 4278 35660
rect 2441 35629 2453 35632
rect 2395 35623 2453 35629
rect 4250 35536 4278 35632
rect 10307 35629 10319 35663
rect 10353 35629 10365 35663
rect 10307 35623 10365 35629
rect 10322 35592 10350 35623
rect 10580 35620 10586 35672
rect 10638 35660 10644 35672
rect 10782 35669 10810 35768
rect 17667 35765 17679 35799
rect 17713 35796 17725 35799
rect 18492 35796 18498 35808
rect 17713 35768 18498 35796
rect 17713 35765 17725 35768
rect 17667 35759 17725 35765
rect 18492 35756 18498 35768
rect 18550 35756 18556 35808
rect 12144 35728 12150 35740
rect 12105 35700 12150 35728
rect 12144 35688 12150 35700
rect 12202 35688 12208 35740
rect 18035 35731 18093 35737
rect 18035 35728 18047 35731
rect 16394 35700 18047 35728
rect 10675 35663 10733 35669
rect 10675 35660 10687 35663
rect 10638 35632 10687 35660
rect 10638 35620 10644 35632
rect 10675 35629 10687 35632
rect 10721 35629 10733 35663
rect 10675 35623 10733 35629
rect 10767 35663 10825 35669
rect 10767 35629 10779 35663
rect 10813 35629 10825 35663
rect 10767 35623 10825 35629
rect 11316 35620 11322 35672
rect 11374 35660 11380 35672
rect 11871 35663 11929 35669
rect 11871 35660 11883 35663
rect 11374 35632 11883 35660
rect 11374 35620 11380 35632
rect 11871 35629 11883 35632
rect 11917 35660 11929 35663
rect 13619 35663 13677 35669
rect 13619 35660 13631 35663
rect 11917 35632 13631 35660
rect 11917 35629 11929 35632
rect 11871 35623 11929 35629
rect 13619 35629 13631 35632
rect 13665 35629 13677 35663
rect 13619 35623 13677 35629
rect 14815 35663 14873 35669
rect 14815 35629 14827 35663
rect 14861 35660 14873 35663
rect 16100 35660 16106 35672
rect 14861 35632 16106 35660
rect 14861 35629 14873 35632
rect 14815 35623 14873 35629
rect 11408 35592 11414 35604
rect 10322 35564 11414 35592
rect 11408 35552 11414 35564
rect 11466 35552 11472 35604
rect 3956 35524 3962 35536
rect 3917 35496 3962 35524
rect 3956 35484 3962 35496
rect 4014 35484 4020 35536
rect 4232 35524 4238 35536
rect 4193 35496 4238 35524
rect 4232 35484 4238 35496
rect 4290 35484 4296 35536
rect 9939 35527 9997 35533
rect 9939 35493 9951 35527
rect 9985 35524 9997 35527
rect 10120 35524 10126 35536
rect 9985 35496 10126 35524
rect 9985 35493 9997 35496
rect 9939 35487 9997 35493
rect 10120 35484 10126 35496
rect 10178 35484 10184 35536
rect 12604 35484 12610 35536
rect 12662 35524 12668 35536
rect 13251 35527 13309 35533
rect 13251 35524 13263 35527
rect 12662 35496 13263 35524
rect 12662 35484 12668 35496
rect 13251 35493 13263 35496
rect 13297 35493 13309 35527
rect 13634 35524 13662 35623
rect 16100 35620 16106 35632
rect 16158 35620 16164 35672
rect 16394 35669 16422 35700
rect 18035 35697 18047 35700
rect 18081 35697 18093 35731
rect 21270 35728 21298 35827
rect 21620 35824 21626 35836
rect 21678 35864 21684 35876
rect 22816 35864 22822 35876
rect 21678 35836 22822 35864
rect 21678 35824 21684 35836
rect 22816 35824 22822 35836
rect 22874 35824 22880 35876
rect 28983 35867 29041 35873
rect 28983 35833 28995 35867
rect 29029 35864 29041 35867
rect 40572 35864 40578 35876
rect 29029 35836 40578 35864
rect 29029 35833 29041 35836
rect 28983 35827 29041 35833
rect 40572 35824 40578 35836
rect 40630 35824 40636 35876
rect 48392 35864 48398 35876
rect 42430 35836 43930 35864
rect 48353 35836 48398 35864
rect 27048 35756 27054 35808
rect 27106 35796 27112 35808
rect 30452 35796 30458 35808
rect 27106 35768 30458 35796
rect 27106 35756 27112 35768
rect 30452 35756 30458 35768
rect 30510 35756 30516 35808
rect 32844 35796 32850 35808
rect 32034 35768 32850 35796
rect 23368 35728 23374 35740
rect 18035 35691 18093 35697
rect 20902 35700 21298 35728
rect 23329 35700 23374 35728
rect 16379 35663 16437 35669
rect 16379 35629 16391 35663
rect 16425 35629 16437 35663
rect 17572 35660 17578 35672
rect 17533 35632 17578 35660
rect 16379 35623 16437 35629
rect 17572 35620 17578 35632
rect 17630 35620 17636 35672
rect 20902 35669 20930 35700
rect 23368 35688 23374 35700
rect 23426 35688 23432 35740
rect 32034 35737 32062 35768
rect 32844 35756 32850 35768
rect 32902 35756 32908 35808
rect 34040 35756 34046 35808
rect 34098 35796 34104 35808
rect 34500 35796 34506 35808
rect 34098 35768 34506 35796
rect 34098 35756 34104 35768
rect 34500 35756 34506 35768
rect 34558 35756 34564 35808
rect 34776 35796 34782 35808
rect 34737 35768 34782 35796
rect 34776 35756 34782 35768
rect 34834 35756 34840 35808
rect 39560 35756 39566 35808
rect 39618 35796 39624 35808
rect 40023 35799 40081 35805
rect 40023 35796 40035 35799
rect 39618 35768 40035 35796
rect 39618 35756 39624 35768
rect 40023 35765 40035 35768
rect 40069 35796 40081 35799
rect 42430 35796 42458 35836
rect 40069 35768 42458 35796
rect 43902 35796 43930 35836
rect 48392 35824 48398 35836
rect 48450 35824 48456 35876
rect 54188 35864 54194 35876
rect 49330 35836 54194 35864
rect 43902 35768 49266 35796
rect 40069 35765 40081 35768
rect 40023 35759 40081 35765
rect 29627 35731 29685 35737
rect 29627 35728 29639 35731
rect 25594 35700 29639 35728
rect 17851 35663 17909 35669
rect 17851 35629 17863 35663
rect 17897 35629 17909 35663
rect 17851 35623 17909 35629
rect 20611 35663 20669 35669
rect 20611 35629 20623 35663
rect 20657 35629 20669 35663
rect 20611 35623 20669 35629
rect 20887 35663 20945 35669
rect 20887 35629 20899 35663
rect 20933 35629 20945 35663
rect 21068 35660 21074 35672
rect 21029 35632 21074 35660
rect 20887 35623 20945 35629
rect 17866 35592 17894 35623
rect 17222 35564 17894 35592
rect 20059 35595 20117 35601
rect 14076 35524 14082 35536
rect 13634 35496 14082 35524
rect 13251 35487 13309 35493
rect 14076 35484 14082 35496
rect 14134 35524 14140 35536
rect 14631 35527 14689 35533
rect 14631 35524 14643 35527
rect 14134 35496 14643 35524
rect 14134 35484 14140 35496
rect 14631 35493 14643 35496
rect 14677 35524 14689 35527
rect 15548 35524 15554 35536
rect 14677 35496 15554 35524
rect 14677 35493 14689 35496
rect 14631 35487 14689 35493
rect 15548 35484 15554 35496
rect 15606 35484 15612 35536
rect 16836 35484 16842 35536
rect 16894 35524 16900 35536
rect 17222 35533 17250 35564
rect 20059 35561 20071 35595
rect 20105 35592 20117 35595
rect 20516 35592 20522 35604
rect 20105 35564 20522 35592
rect 20105 35561 20117 35564
rect 20059 35555 20117 35561
rect 20516 35552 20522 35564
rect 20574 35552 20580 35604
rect 20626 35592 20654 35623
rect 21068 35620 21074 35632
rect 21126 35620 21132 35672
rect 25594 35669 25622 35700
rect 29627 35697 29639 35700
rect 29673 35697 29685 35731
rect 29627 35691 29685 35697
rect 32019 35731 32077 35737
rect 32019 35697 32031 35731
rect 32065 35697 32077 35731
rect 32019 35691 32077 35697
rect 37631 35731 37689 35737
rect 37631 35697 37643 35731
rect 37677 35728 37689 35731
rect 38088 35728 38094 35740
rect 37677 35700 38094 35728
rect 37677 35697 37689 35700
rect 37631 35691 37689 35697
rect 38088 35688 38094 35700
rect 38146 35688 38152 35740
rect 42872 35728 42878 35740
rect 39854 35700 42878 35728
rect 23095 35663 23153 35669
rect 23095 35629 23107 35663
rect 23141 35660 23153 35663
rect 24751 35663 24809 35669
rect 23141 35632 24702 35660
rect 23141 35629 23153 35632
rect 23095 35623 23153 35629
rect 21528 35592 21534 35604
rect 20626 35564 21534 35592
rect 21528 35552 21534 35564
rect 21586 35592 21592 35604
rect 22816 35592 22822 35604
rect 21586 35564 22822 35592
rect 21586 35552 21592 35564
rect 22816 35552 22822 35564
rect 22874 35552 22880 35604
rect 24674 35592 24702 35632
rect 24751 35629 24763 35663
rect 24797 35660 24809 35663
rect 25579 35663 25637 35669
rect 25579 35660 25591 35663
rect 24797 35632 25591 35660
rect 24797 35629 24809 35632
rect 24751 35623 24809 35629
rect 25579 35629 25591 35632
rect 25625 35629 25637 35663
rect 25579 35623 25637 35629
rect 25668 35620 25674 35672
rect 25726 35660 25732 35672
rect 28244 35660 28250 35672
rect 25726 35632 28250 35660
rect 25726 35620 25732 35632
rect 28244 35620 28250 35632
rect 28302 35660 28308 35672
rect 29167 35663 29225 35669
rect 29167 35660 29179 35663
rect 28302 35632 29179 35660
rect 28302 35620 28308 35632
rect 29167 35629 29179 35632
rect 29213 35629 29225 35663
rect 29167 35623 29225 35629
rect 29348 35620 29354 35672
rect 29406 35660 29412 35672
rect 29719 35663 29777 35669
rect 29406 35632 29451 35660
rect 29406 35620 29412 35632
rect 29719 35629 29731 35663
rect 29765 35660 29777 35663
rect 30268 35660 30274 35672
rect 29765 35632 30274 35660
rect 29765 35629 29777 35632
rect 29719 35623 29777 35629
rect 30268 35620 30274 35632
rect 30326 35620 30332 35672
rect 32108 35660 32114 35672
rect 32069 35632 32114 35660
rect 32108 35620 32114 35632
rect 32166 35620 32172 35672
rect 32663 35663 32721 35669
rect 32663 35629 32675 35663
rect 32709 35629 32721 35663
rect 32663 35623 32721 35629
rect 24935 35595 24993 35601
rect 24935 35592 24947 35595
rect 24674 35564 24947 35592
rect 24935 35561 24947 35564
rect 24981 35592 24993 35595
rect 32016 35592 32022 35604
rect 24981 35564 32022 35592
rect 24981 35561 24993 35564
rect 24935 35555 24993 35561
rect 32016 35552 32022 35564
rect 32074 35552 32080 35604
rect 32126 35592 32154 35620
rect 32678 35592 32706 35623
rect 32752 35620 32758 35672
rect 32810 35660 32816 35672
rect 32847 35663 32905 35669
rect 32847 35660 32859 35663
rect 32810 35632 32859 35660
rect 32810 35620 32816 35632
rect 32847 35629 32859 35632
rect 32893 35660 32905 35663
rect 34319 35663 34377 35669
rect 32893 35632 33534 35660
rect 32893 35629 32905 35632
rect 32847 35623 32905 35629
rect 32126 35564 32706 35592
rect 33215 35595 33273 35601
rect 33215 35561 33227 35595
rect 33261 35592 33273 35595
rect 33304 35592 33310 35604
rect 33261 35564 33310 35592
rect 33261 35561 33273 35564
rect 33215 35555 33273 35561
rect 33304 35552 33310 35564
rect 33362 35552 33368 35604
rect 17207 35527 17265 35533
rect 17207 35524 17219 35527
rect 16894 35496 17219 35524
rect 16894 35484 16900 35496
rect 17207 35493 17219 35496
rect 17253 35493 17265 35527
rect 18492 35524 18498 35536
rect 18453 35496 18498 35524
rect 17207 35487 17265 35493
rect 18492 35484 18498 35496
rect 18550 35484 18556 35536
rect 23828 35484 23834 35536
rect 23886 35524 23892 35536
rect 29072 35524 29078 35536
rect 23886 35496 29078 35524
rect 23886 35484 23892 35496
rect 29072 35484 29078 35496
rect 29130 35484 29136 35536
rect 29348 35484 29354 35536
rect 29406 35524 29412 35536
rect 30084 35524 30090 35536
rect 29406 35496 30090 35524
rect 29406 35484 29412 35496
rect 30084 35484 30090 35496
rect 30142 35484 30148 35536
rect 33506 35533 33534 35632
rect 34319 35629 34331 35663
rect 34365 35660 34377 35663
rect 34776 35660 34782 35672
rect 34365 35632 34782 35660
rect 34365 35629 34377 35632
rect 34319 35623 34377 35629
rect 34776 35620 34782 35632
rect 34834 35620 34840 35672
rect 37168 35620 37174 35672
rect 37226 35660 37232 35672
rect 37355 35663 37413 35669
rect 37355 35660 37367 35663
rect 37226 35632 37367 35660
rect 37226 35620 37232 35632
rect 37355 35629 37367 35632
rect 37401 35629 37413 35663
rect 39854 35660 39882 35700
rect 42872 35688 42878 35700
rect 42930 35688 42936 35740
rect 43243 35731 43301 35737
rect 43243 35697 43255 35731
rect 43289 35728 43301 35731
rect 44068 35728 44074 35740
rect 43289 35700 44074 35728
rect 43289 35697 43301 35700
rect 43243 35691 43301 35697
rect 44068 35688 44074 35700
rect 44126 35688 44132 35740
rect 47656 35688 47662 35740
rect 47714 35728 47720 35740
rect 48671 35731 48729 35737
rect 48671 35728 48683 35731
rect 47714 35700 48683 35728
rect 47714 35688 47720 35700
rect 48671 35697 48683 35700
rect 48717 35697 48729 35731
rect 48671 35691 48729 35697
rect 37355 35623 37413 35629
rect 37462 35632 39882 35660
rect 39931 35663 39989 35669
rect 35512 35552 35518 35604
rect 35570 35592 35576 35604
rect 37462 35592 37490 35632
rect 39931 35629 39943 35663
rect 39977 35660 39989 35663
rect 40020 35660 40026 35672
rect 39977 35632 40026 35660
rect 39977 35629 39989 35632
rect 39931 35623 39989 35629
rect 40020 35620 40026 35632
rect 40078 35620 40084 35672
rect 42967 35663 43025 35669
rect 42967 35660 42979 35663
rect 42798 35632 42979 35660
rect 35570 35564 37490 35592
rect 39011 35595 39069 35601
rect 35570 35552 35576 35564
rect 39011 35561 39023 35595
rect 39057 35592 39069 35595
rect 39836 35592 39842 35604
rect 39057 35564 39842 35592
rect 39057 35561 39069 35564
rect 39011 35555 39069 35561
rect 39836 35552 39842 35564
rect 39894 35552 39900 35604
rect 33491 35527 33549 35533
rect 33491 35493 33503 35527
rect 33537 35524 33549 35527
rect 36064 35524 36070 35536
rect 33537 35496 36070 35524
rect 33537 35493 33549 35496
rect 33491 35487 33549 35493
rect 36064 35484 36070 35496
rect 36122 35484 36128 35536
rect 37168 35524 37174 35536
rect 37129 35496 37174 35524
rect 37168 35484 37174 35496
rect 37226 35524 37232 35536
rect 40756 35524 40762 35536
rect 37226 35496 40762 35524
rect 37226 35484 37232 35496
rect 40756 35484 40762 35496
rect 40814 35524 40820 35536
rect 42798 35533 42826 35632
rect 42967 35629 42979 35632
rect 43013 35629 43025 35663
rect 42967 35623 43025 35629
rect 45543 35663 45601 35669
rect 45543 35629 45555 35663
rect 45589 35629 45601 35663
rect 45543 35623 45601 35629
rect 44620 35592 44626 35604
rect 44581 35564 44626 35592
rect 44620 35552 44626 35564
rect 44678 35592 44684 35604
rect 45558 35592 45586 35623
rect 46736 35620 46742 35672
rect 46794 35660 46800 35672
rect 46923 35663 46981 35669
rect 46923 35660 46935 35663
rect 46794 35632 46935 35660
rect 46794 35620 46800 35632
rect 46923 35629 46935 35632
rect 46969 35629 46981 35663
rect 46923 35623 46981 35629
rect 48392 35620 48398 35672
rect 48450 35660 48456 35672
rect 48579 35663 48637 35669
rect 48579 35660 48591 35663
rect 48450 35632 48591 35660
rect 48450 35620 48456 35632
rect 48579 35629 48591 35632
rect 48625 35629 48637 35663
rect 48852 35660 48858 35672
rect 48813 35632 48858 35660
rect 48579 35623 48637 35629
rect 48852 35620 48858 35632
rect 48910 35620 48916 35672
rect 49238 35660 49266 35768
rect 49330 35737 49358 35836
rect 54188 35824 54194 35836
rect 54246 35824 54252 35876
rect 54375 35867 54433 35873
rect 54375 35833 54387 35867
rect 54421 35864 54433 35867
rect 80684 35864 80690 35876
rect 54421 35836 80690 35864
rect 54421 35833 54433 35836
rect 54375 35827 54433 35833
rect 49315 35731 49373 35737
rect 49315 35697 49327 35731
rect 49361 35697 49373 35731
rect 49315 35691 49373 35697
rect 52443 35663 52501 35669
rect 52443 35660 52455 35663
rect 49238 35632 52455 35660
rect 52443 35629 52455 35632
rect 52489 35660 52501 35663
rect 52627 35663 52685 35669
rect 52627 35660 52639 35663
rect 52489 35632 52639 35660
rect 52489 35629 52501 35632
rect 52443 35623 52501 35629
rect 52627 35629 52639 35632
rect 52673 35629 52685 35663
rect 52627 35623 52685 35629
rect 52811 35663 52869 35669
rect 52811 35629 52823 35663
rect 52857 35660 52869 35663
rect 53176 35660 53182 35672
rect 52857 35632 53182 35660
rect 52857 35629 52869 35632
rect 52811 35623 52869 35629
rect 53176 35620 53182 35632
rect 53234 35620 53240 35672
rect 53363 35663 53421 35669
rect 53363 35629 53375 35663
rect 53409 35660 53421 35663
rect 53452 35660 53458 35672
rect 53409 35632 53458 35660
rect 53409 35629 53421 35632
rect 53363 35623 53421 35629
rect 53452 35620 53458 35632
rect 53510 35620 53516 35672
rect 53547 35663 53605 35669
rect 53547 35629 53559 35663
rect 53593 35660 53605 35663
rect 54390 35660 54418 35827
rect 80684 35824 80690 35836
rect 80742 35824 80748 35876
rect 85563 35867 85621 35873
rect 85563 35833 85575 35867
rect 85609 35864 85621 35867
rect 85836 35864 85842 35876
rect 85609 35836 85842 35864
rect 85609 35833 85621 35836
rect 85563 35827 85621 35833
rect 85836 35824 85842 35836
rect 85894 35824 85900 35876
rect 91356 35824 91362 35876
rect 91414 35864 91420 35876
rect 91819 35867 91877 35873
rect 91819 35864 91831 35867
rect 91414 35836 91831 35864
rect 91414 35824 91420 35836
rect 91819 35833 91831 35836
rect 91865 35833 91877 35867
rect 91819 35827 91877 35833
rect 55568 35756 55574 35808
rect 55626 35796 55632 35808
rect 56951 35799 57009 35805
rect 56951 35796 56963 35799
rect 55626 35768 56963 35796
rect 55626 35756 55632 35768
rect 56951 35765 56963 35768
rect 56997 35765 57009 35799
rect 56951 35759 57009 35765
rect 57150 35768 63526 35796
rect 53593 35632 54418 35660
rect 53593 35629 53605 35632
rect 53547 35623 53605 35629
rect 56672 35620 56678 35672
rect 56730 35660 56736 35672
rect 57150 35669 57178 35768
rect 57868 35688 57874 35740
rect 57926 35728 57932 35740
rect 57963 35731 58021 35737
rect 57963 35728 57975 35731
rect 57926 35700 57975 35728
rect 57926 35688 57932 35700
rect 57963 35697 57975 35700
rect 58009 35728 58021 35731
rect 58147 35731 58205 35737
rect 58147 35728 58159 35731
rect 58009 35700 58159 35728
rect 58009 35697 58021 35700
rect 57963 35691 58021 35697
rect 58147 35697 58159 35700
rect 58193 35697 58205 35731
rect 58147 35691 58205 35697
rect 59711 35731 59769 35737
rect 59711 35697 59723 35731
rect 59757 35728 59769 35731
rect 59984 35728 59990 35740
rect 59757 35700 59990 35728
rect 59757 35697 59769 35700
rect 59711 35691 59769 35697
rect 56767 35663 56825 35669
rect 56767 35660 56779 35663
rect 56730 35632 56779 35660
rect 56730 35620 56736 35632
rect 56767 35629 56779 35632
rect 56813 35660 56825 35663
rect 57135 35663 57193 35669
rect 57135 35660 57147 35663
rect 56813 35632 57147 35660
rect 56813 35629 56825 35632
rect 56767 35623 56825 35629
rect 57135 35629 57147 35632
rect 57181 35629 57193 35663
rect 58328 35660 58334 35672
rect 58289 35632 58334 35660
rect 57135 35623 57193 35629
rect 58328 35620 58334 35632
rect 58386 35620 58392 35672
rect 58880 35660 58886 35672
rect 58793 35632 58886 35660
rect 44678 35564 45586 35592
rect 45635 35595 45693 35601
rect 44678 35552 44684 35564
rect 45635 35561 45647 35595
rect 45681 35592 45693 35595
rect 49404 35592 49410 35604
rect 45681 35564 49410 35592
rect 45681 35561 45693 35564
rect 45635 35555 45693 35561
rect 42783 35527 42841 35533
rect 42783 35524 42795 35527
rect 40814 35496 42795 35524
rect 40814 35484 40820 35496
rect 42783 35493 42795 35496
rect 42829 35524 42841 35527
rect 43056 35524 43062 35536
rect 42829 35496 43062 35524
rect 42829 35493 42841 35496
rect 42783 35487 42841 35493
rect 43056 35484 43062 35496
rect 43114 35484 43120 35536
rect 43976 35484 43982 35536
rect 44034 35524 44040 35536
rect 45650 35524 45678 35555
rect 49404 35552 49410 35564
rect 49462 35552 49468 35604
rect 51980 35552 51986 35604
rect 52038 35592 52044 35604
rect 54648 35592 54654 35604
rect 52038 35564 54654 35592
rect 52038 35552 52044 35564
rect 54648 35552 54654 35564
rect 54706 35552 54712 35604
rect 58806 35592 58834 35632
rect 58880 35620 58886 35632
rect 58938 35620 58944 35672
rect 59064 35660 59070 35672
rect 59025 35632 59070 35660
rect 59064 35620 59070 35632
rect 59122 35620 59128 35672
rect 59726 35660 59754 35691
rect 59984 35688 59990 35700
rect 60042 35728 60048 35740
rect 61824 35728 61830 35740
rect 60042 35700 61830 35728
rect 60042 35688 60048 35700
rect 61824 35688 61830 35700
rect 61882 35728 61888 35740
rect 61882 35700 62606 35728
rect 61882 35688 61888 35700
rect 62578 35672 62606 35700
rect 59174 35632 59754 35660
rect 59174 35592 59202 35632
rect 60168 35620 60174 35672
rect 60226 35660 60232 35672
rect 62376 35660 62382 35672
rect 60226 35632 62382 35660
rect 60226 35620 60232 35632
rect 62376 35620 62382 35632
rect 62434 35620 62440 35672
rect 62560 35660 62566 35672
rect 62521 35632 62566 35660
rect 62560 35620 62566 35632
rect 62618 35620 62624 35672
rect 63023 35663 63081 35669
rect 63023 35629 63035 35663
rect 63069 35629 63081 35663
rect 63023 35623 63081 35629
rect 63203 35663 63261 35669
rect 63203 35629 63215 35663
rect 63249 35660 63261 35663
rect 63296 35660 63302 35672
rect 63249 35632 63302 35660
rect 63249 35629 63261 35632
rect 63203 35623 63261 35629
rect 54758 35564 57086 35592
rect 58806 35564 59202 35592
rect 59435 35595 59493 35601
rect 44034 35496 45678 35524
rect 44034 35484 44040 35496
rect 46644 35484 46650 35536
rect 46702 35524 46708 35536
rect 47015 35527 47073 35533
rect 47015 35524 47027 35527
rect 46702 35496 47027 35524
rect 46702 35484 46708 35496
rect 47015 35493 47027 35496
rect 47061 35524 47073 35527
rect 47104 35524 47110 35536
rect 47061 35496 47110 35524
rect 47061 35493 47073 35496
rect 47015 35487 47073 35493
rect 47104 35484 47110 35496
rect 47162 35484 47168 35536
rect 51888 35484 51894 35536
rect 51946 35524 51952 35536
rect 52348 35524 52354 35536
rect 51946 35496 52354 35524
rect 51946 35484 51952 35496
rect 52348 35484 52354 35496
rect 52406 35524 52412 35536
rect 52624 35524 52630 35536
rect 52406 35496 52630 35524
rect 52406 35484 52412 35496
rect 52624 35484 52630 35496
rect 52682 35484 52688 35536
rect 53268 35484 53274 35536
rect 53326 35524 53332 35536
rect 53823 35527 53881 35533
rect 53823 35524 53835 35527
rect 53326 35496 53835 35524
rect 53326 35484 53332 35496
rect 53823 35493 53835 35496
rect 53869 35493 53881 35527
rect 53823 35487 53881 35493
rect 54004 35484 54010 35536
rect 54062 35524 54068 35536
rect 54099 35527 54157 35533
rect 54099 35524 54111 35527
rect 54062 35496 54111 35524
rect 54062 35484 54068 35496
rect 54099 35493 54111 35496
rect 54145 35493 54157 35527
rect 54099 35487 54157 35493
rect 54188 35484 54194 35536
rect 54246 35524 54252 35536
rect 54758 35524 54786 35564
rect 54246 35496 54786 35524
rect 57058 35524 57086 35564
rect 59435 35561 59447 35595
rect 59481 35592 59493 35595
rect 60260 35592 60266 35604
rect 59481 35564 60266 35592
rect 59481 35561 59493 35564
rect 59435 35555 59493 35561
rect 60260 35552 60266 35564
rect 60318 35552 60324 35604
rect 63038 35592 63066 35623
rect 63296 35620 63302 35632
rect 63354 35620 63360 35672
rect 63498 35660 63526 35768
rect 67436 35756 67442 35808
rect 67494 35796 67500 35808
rect 68083 35799 68141 35805
rect 68083 35796 68095 35799
rect 67494 35768 68095 35796
rect 67494 35756 67500 35768
rect 68083 35765 68095 35768
rect 68129 35796 68141 35799
rect 68356 35796 68362 35808
rect 68129 35768 68362 35796
rect 68129 35765 68141 35768
rect 68083 35759 68141 35765
rect 68356 35756 68362 35768
rect 68414 35756 68420 35808
rect 75256 35756 75262 35808
rect 75314 35796 75320 35808
rect 75995 35799 76053 35805
rect 75995 35796 76007 35799
rect 75314 35768 76007 35796
rect 75314 35756 75320 35768
rect 75995 35765 76007 35768
rect 76041 35765 76053 35799
rect 75995 35759 76053 35765
rect 63940 35728 63946 35740
rect 63853 35700 63946 35728
rect 63940 35688 63946 35700
rect 63998 35728 64004 35740
rect 67896 35728 67902 35740
rect 63998 35700 67902 35728
rect 63998 35688 64004 35700
rect 67896 35688 67902 35700
rect 67954 35688 67960 35740
rect 69276 35728 69282 35740
rect 69237 35700 69282 35728
rect 69276 35688 69282 35700
rect 69334 35688 69340 35740
rect 70751 35731 70809 35737
rect 70751 35728 70763 35731
rect 69386 35700 70763 35728
rect 67991 35663 68049 35669
rect 63498 35632 67022 35660
rect 62118 35564 63066 35592
rect 63314 35592 63342 35620
rect 66884 35592 66890 35604
rect 63314 35564 66890 35592
rect 62118 35536 62146 35564
rect 66884 35552 66890 35564
rect 66942 35552 66948 35604
rect 61916 35524 61922 35536
rect 57058 35496 61922 35524
rect 54246 35484 54252 35496
rect 61916 35484 61922 35496
rect 61974 35484 61980 35536
rect 62100 35524 62106 35536
rect 62061 35496 62106 35524
rect 62100 35484 62106 35496
rect 62158 35484 62164 35536
rect 62560 35484 62566 35536
rect 62618 35524 62624 35536
rect 63204 35524 63210 35536
rect 62618 35496 63210 35524
rect 62618 35484 62624 35496
rect 63204 35484 63210 35496
rect 63262 35484 63268 35536
rect 63572 35524 63578 35536
rect 63533 35496 63578 35524
rect 63572 35484 63578 35496
rect 63630 35484 63636 35536
rect 64124 35524 64130 35536
rect 64085 35496 64130 35524
rect 64124 35484 64130 35496
rect 64182 35484 64188 35536
rect 66994 35524 67022 35632
rect 67991 35629 68003 35663
rect 68037 35660 68049 35663
rect 68908 35660 68914 35672
rect 68037 35632 68914 35660
rect 68037 35629 68049 35632
rect 67991 35623 68049 35629
rect 68908 35620 68914 35632
rect 68966 35620 68972 35672
rect 69003 35663 69061 35669
rect 69003 35629 69015 35663
rect 69049 35660 69061 35663
rect 69386 35660 69414 35700
rect 70751 35697 70763 35700
rect 70797 35728 70809 35731
rect 73232 35728 73238 35740
rect 70797 35700 73238 35728
rect 70797 35697 70809 35700
rect 70751 35691 70809 35697
rect 73232 35688 73238 35700
rect 73290 35688 73296 35740
rect 73324 35688 73330 35740
rect 73382 35728 73388 35740
rect 73603 35731 73661 35737
rect 73603 35728 73615 35731
rect 73382 35700 73615 35728
rect 73382 35688 73388 35700
rect 73603 35697 73615 35700
rect 73649 35697 73661 35731
rect 73603 35691 73661 35697
rect 73692 35688 73698 35740
rect 73750 35728 73756 35740
rect 73750 35700 74014 35728
rect 73750 35688 73756 35700
rect 69049 35632 69414 35660
rect 69049 35629 69061 35632
rect 69003 35623 69061 35629
rect 69552 35620 69558 35672
rect 69610 35660 69616 35672
rect 73784 35660 73790 35672
rect 69610 35632 73646 35660
rect 73745 35632 73790 35660
rect 69610 35620 69616 35632
rect 70656 35592 70662 35604
rect 70617 35564 70662 35592
rect 70656 35552 70662 35564
rect 70714 35552 70720 35604
rect 70104 35524 70110 35536
rect 66994 35496 70110 35524
rect 70104 35484 70110 35496
rect 70162 35484 70168 35536
rect 73618 35524 73646 35632
rect 73784 35620 73790 35632
rect 73842 35620 73848 35672
rect 73986 35660 74014 35700
rect 85468 35688 85474 35740
rect 85526 35728 85532 35740
rect 85526 35700 85974 35728
rect 85526 35688 85532 35700
rect 74247 35663 74305 35669
rect 74247 35660 74259 35663
rect 73986 35632 74259 35660
rect 74247 35629 74259 35632
rect 74293 35629 74305 35663
rect 74247 35623 74305 35629
rect 74336 35620 74342 35672
rect 74394 35660 74400 35672
rect 75811 35663 75869 35669
rect 75811 35660 75823 35663
rect 74394 35632 74439 35660
rect 75642 35632 75823 35660
rect 74394 35620 74400 35632
rect 74060 35524 74066 35536
rect 73618 35496 74066 35524
rect 74060 35484 74066 35496
rect 74118 35484 74124 35536
rect 74152 35484 74158 35536
rect 74210 35524 74216 35536
rect 74799 35527 74857 35533
rect 74799 35524 74811 35527
rect 74210 35496 74811 35524
rect 74210 35484 74216 35496
rect 74799 35493 74811 35496
rect 74845 35493 74857 35527
rect 74799 35487 74857 35493
rect 75440 35484 75446 35536
rect 75498 35524 75504 35536
rect 75642 35533 75670 35632
rect 75811 35629 75823 35632
rect 75857 35660 75869 35663
rect 79215 35663 79273 35669
rect 79215 35660 79227 35663
rect 75857 35632 79227 35660
rect 75857 35629 75869 35632
rect 75811 35623 75869 35629
rect 79215 35629 79227 35632
rect 79261 35660 79273 35663
rect 79583 35663 79641 35669
rect 79583 35660 79595 35663
rect 79261 35632 79595 35660
rect 79261 35629 79273 35632
rect 79215 35623 79273 35629
rect 79583 35629 79595 35632
rect 79629 35629 79641 35663
rect 79583 35623 79641 35629
rect 81788 35620 81794 35672
rect 81846 35660 81852 35672
rect 82064 35660 82070 35672
rect 81846 35632 82070 35660
rect 81846 35620 81852 35632
rect 82064 35620 82070 35632
rect 82122 35620 82128 35672
rect 82251 35663 82309 35669
rect 82251 35629 82263 35663
rect 82297 35629 82309 35663
rect 82708 35660 82714 35672
rect 82669 35632 82714 35660
rect 82251 35623 82309 35629
rect 82266 35592 82294 35623
rect 82708 35620 82714 35632
rect 82766 35620 82772 35672
rect 82803 35663 82861 35669
rect 82803 35629 82815 35663
rect 82849 35660 82861 35663
rect 85652 35660 85658 35672
rect 82849 35632 85658 35660
rect 82849 35629 82861 35632
rect 82803 35623 82861 35629
rect 82818 35592 82846 35623
rect 85652 35620 85658 35632
rect 85710 35620 85716 35672
rect 85946 35669 85974 35700
rect 86572 35688 86578 35740
rect 86630 35728 86636 35740
rect 86759 35731 86817 35737
rect 86759 35728 86771 35731
rect 86630 35700 86771 35728
rect 86630 35688 86636 35700
rect 86759 35697 86771 35700
rect 86805 35697 86817 35731
rect 86759 35691 86817 35697
rect 88047 35731 88105 35737
rect 88047 35697 88059 35731
rect 88093 35728 88105 35731
rect 88228 35728 88234 35740
rect 88093 35700 88234 35728
rect 88093 35697 88105 35700
rect 88047 35691 88105 35697
rect 88228 35688 88234 35700
rect 88286 35688 88292 35740
rect 90712 35728 90718 35740
rect 90673 35700 90718 35728
rect 90712 35688 90718 35700
rect 90770 35688 90776 35740
rect 85747 35663 85805 35669
rect 85747 35629 85759 35663
rect 85793 35629 85805 35663
rect 85747 35623 85805 35629
rect 85931 35663 85989 35669
rect 85931 35629 85943 35663
rect 85977 35629 85989 35663
rect 85931 35623 85989 35629
rect 82266 35564 82846 35592
rect 83355 35595 83413 35601
rect 75627 35527 75685 35533
rect 75627 35524 75639 35527
rect 75498 35496 75639 35524
rect 75498 35484 75504 35496
rect 75627 35493 75639 35496
rect 75673 35493 75685 35527
rect 75627 35487 75685 35493
rect 79399 35527 79457 35533
rect 79399 35493 79411 35527
rect 79445 35524 79457 35527
rect 80224 35524 80230 35536
rect 79445 35496 80230 35524
rect 79445 35493 79457 35496
rect 79399 35487 79457 35493
rect 80224 35484 80230 35496
rect 80282 35484 80288 35536
rect 81696 35524 81702 35536
rect 81657 35496 81702 35524
rect 81696 35484 81702 35496
rect 81754 35524 81760 35536
rect 81883 35527 81941 35533
rect 81883 35524 81895 35527
rect 81754 35496 81895 35524
rect 81754 35484 81760 35496
rect 81883 35493 81895 35496
rect 81929 35524 81941 35527
rect 82266 35524 82294 35564
rect 83355 35561 83367 35595
rect 83401 35592 83413 35595
rect 83536 35592 83542 35604
rect 83401 35564 83542 35592
rect 83401 35561 83413 35564
rect 83355 35555 83413 35561
rect 83536 35552 83542 35564
rect 83594 35552 83600 35604
rect 85762 35592 85790 35623
rect 86020 35620 86026 35672
rect 86078 35660 86084 35672
rect 86299 35663 86357 35669
rect 86299 35660 86311 35663
rect 86078 35632 86311 35660
rect 86078 35620 86084 35632
rect 86299 35629 86311 35632
rect 86345 35629 86357 35663
rect 86299 35623 86357 35629
rect 86483 35663 86541 35669
rect 86483 35629 86495 35663
rect 86529 35660 86541 35663
rect 88320 35660 88326 35672
rect 86529 35632 86710 35660
rect 88281 35632 88326 35660
rect 86529 35629 86541 35632
rect 86483 35623 86541 35629
rect 86572 35592 86578 35604
rect 85762 35564 86578 35592
rect 86572 35552 86578 35564
rect 86630 35552 86636 35604
rect 86682 35536 86710 35632
rect 88320 35620 88326 35632
rect 88378 35620 88384 35672
rect 88780 35660 88786 35672
rect 88741 35632 88786 35660
rect 88780 35620 88786 35632
rect 88838 35620 88844 35672
rect 88875 35663 88933 35669
rect 88875 35629 88887 35663
rect 88921 35629 88933 35663
rect 90439 35663 90497 35669
rect 90439 35660 90451 35663
rect 88875 35623 88933 35629
rect 90178 35632 90451 35660
rect 87768 35552 87774 35604
rect 87826 35592 87832 35604
rect 88890 35592 88918 35623
rect 87826 35564 88918 35592
rect 89427 35595 89485 35601
rect 87826 35552 87832 35564
rect 89427 35561 89439 35595
rect 89473 35592 89485 35595
rect 89976 35592 89982 35604
rect 89473 35564 89982 35592
rect 89473 35561 89485 35564
rect 89427 35555 89485 35561
rect 89976 35552 89982 35564
rect 90034 35552 90040 35604
rect 86664 35524 86670 35536
rect 81929 35496 82294 35524
rect 86625 35496 86670 35524
rect 81929 35493 81941 35496
rect 81883 35487 81941 35493
rect 86664 35484 86670 35496
rect 86722 35484 86728 35536
rect 89516 35484 89522 35536
rect 89574 35524 89580 35536
rect 90178 35533 90206 35632
rect 90439 35629 90451 35632
rect 90485 35629 90497 35663
rect 90439 35623 90497 35629
rect 90163 35527 90221 35533
rect 90163 35524 90175 35527
rect 89574 35496 90175 35524
rect 89574 35484 89580 35496
rect 90163 35493 90175 35496
rect 90209 35493 90221 35527
rect 90163 35487 90221 35493
rect 538 35434 93642 35456
rect 538 35382 6344 35434
rect 6396 35382 6408 35434
rect 6460 35382 6472 35434
rect 6524 35382 6536 35434
rect 6588 35382 11672 35434
rect 11724 35382 11736 35434
rect 11788 35382 11800 35434
rect 11852 35382 11864 35434
rect 11916 35382 17000 35434
rect 17052 35382 17064 35434
rect 17116 35382 17128 35434
rect 17180 35382 17192 35434
rect 17244 35382 22328 35434
rect 22380 35382 22392 35434
rect 22444 35382 22456 35434
rect 22508 35382 22520 35434
rect 22572 35382 27656 35434
rect 27708 35382 27720 35434
rect 27772 35382 27784 35434
rect 27836 35382 27848 35434
rect 27900 35382 32984 35434
rect 33036 35382 33048 35434
rect 33100 35382 33112 35434
rect 33164 35382 33176 35434
rect 33228 35382 38312 35434
rect 38364 35382 38376 35434
rect 38428 35382 38440 35434
rect 38492 35382 38504 35434
rect 38556 35382 43640 35434
rect 43692 35382 43704 35434
rect 43756 35382 43768 35434
rect 43820 35382 43832 35434
rect 43884 35382 48968 35434
rect 49020 35382 49032 35434
rect 49084 35382 49096 35434
rect 49148 35382 49160 35434
rect 49212 35382 54296 35434
rect 54348 35382 54360 35434
rect 54412 35382 54424 35434
rect 54476 35382 54488 35434
rect 54540 35382 59624 35434
rect 59676 35382 59688 35434
rect 59740 35382 59752 35434
rect 59804 35382 59816 35434
rect 59868 35382 64952 35434
rect 65004 35382 65016 35434
rect 65068 35382 65080 35434
rect 65132 35382 65144 35434
rect 65196 35382 70280 35434
rect 70332 35382 70344 35434
rect 70396 35382 70408 35434
rect 70460 35382 70472 35434
rect 70524 35382 75608 35434
rect 75660 35382 75672 35434
rect 75724 35382 75736 35434
rect 75788 35382 75800 35434
rect 75852 35382 80936 35434
rect 80988 35382 81000 35434
rect 81052 35382 81064 35434
rect 81116 35382 81128 35434
rect 81180 35382 86264 35434
rect 86316 35382 86328 35434
rect 86380 35382 86392 35434
rect 86444 35382 86456 35434
rect 86508 35382 91592 35434
rect 91644 35382 91656 35434
rect 91708 35382 91720 35434
rect 91772 35382 91784 35434
rect 91836 35382 93642 35434
rect 538 35360 93642 35382
rect 2487 35323 2545 35329
rect 2487 35289 2499 35323
rect 2533 35320 2545 35323
rect 2668 35320 2674 35332
rect 2533 35292 2674 35320
rect 2533 35289 2545 35292
rect 2487 35283 2545 35289
rect 2668 35280 2674 35292
rect 2726 35280 2732 35332
rect 6811 35323 6869 35329
rect 6811 35289 6823 35323
rect 6857 35320 6869 35323
rect 10580 35320 10586 35332
rect 6857 35292 10586 35320
rect 6857 35289 6869 35292
rect 6811 35283 6869 35289
rect 10580 35280 10586 35292
rect 10638 35280 10644 35332
rect 11960 35280 11966 35332
rect 12018 35320 12024 35332
rect 12788 35320 12794 35332
rect 12018 35292 12794 35320
rect 12018 35280 12024 35292
rect 12788 35280 12794 35292
rect 12846 35320 12852 35332
rect 13067 35323 13125 35329
rect 13067 35320 13079 35323
rect 12846 35292 13079 35320
rect 12846 35280 12852 35292
rect 13067 35289 13079 35292
rect 13113 35289 13125 35323
rect 15548 35320 15554 35332
rect 15509 35292 15554 35320
rect 13067 35283 13125 35289
rect 13082 35252 13110 35283
rect 15548 35280 15554 35292
rect 15606 35280 15612 35332
rect 18952 35280 18958 35332
rect 19010 35320 19016 35332
rect 19412 35320 19418 35332
rect 19010 35292 19418 35320
rect 19010 35280 19016 35292
rect 19412 35280 19418 35292
rect 19470 35280 19476 35332
rect 21160 35280 21166 35332
rect 21218 35320 21224 35332
rect 23828 35320 23834 35332
rect 21218 35292 23834 35320
rect 21218 35280 21224 35292
rect 23828 35280 23834 35292
rect 23886 35280 23892 35332
rect 24012 35320 24018 35332
rect 23973 35292 24018 35320
rect 24012 35280 24018 35292
rect 24070 35280 24076 35332
rect 28060 35280 28066 35332
rect 28118 35320 28124 35332
rect 28247 35323 28305 35329
rect 28247 35320 28259 35323
rect 28118 35292 28259 35320
rect 28118 35280 28124 35292
rect 28247 35289 28259 35292
rect 28293 35289 28305 35323
rect 29256 35320 29262 35332
rect 28247 35283 28305 35289
rect 28354 35292 29262 35320
rect 15088 35252 15094 35264
rect 13082 35224 13478 35252
rect 15049 35224 15094 35252
rect 1843 35187 1901 35193
rect 1843 35153 1855 35187
rect 1889 35184 1901 35187
rect 2576 35184 2582 35196
rect 1889 35156 2582 35184
rect 1889 35153 1901 35156
rect 1843 35147 1901 35153
rect 2576 35144 2582 35156
rect 2634 35144 2640 35196
rect 3956 35144 3962 35196
rect 4014 35184 4020 35196
rect 5523 35187 5581 35193
rect 5523 35184 5535 35187
rect 4014 35156 5535 35184
rect 4014 35144 4020 35156
rect 5523 35153 5535 35156
rect 5569 35153 5581 35187
rect 10120 35184 10126 35196
rect 10081 35156 10126 35184
rect 5523 35147 5581 35153
rect 10120 35144 10126 35156
rect 10178 35144 10184 35196
rect 11408 35144 11414 35196
rect 11466 35184 11472 35196
rect 13450 35193 13478 35224
rect 15088 35212 15094 35224
rect 15146 35212 15152 35264
rect 17572 35212 17578 35264
rect 17630 35252 17636 35264
rect 18219 35255 18277 35261
rect 18219 35252 18231 35255
rect 17630 35224 18231 35252
rect 17630 35212 17636 35224
rect 18219 35221 18231 35224
rect 18265 35221 18277 35255
rect 20148 35252 20154 35264
rect 18219 35215 18277 35221
rect 18786 35224 20154 35252
rect 11503 35187 11561 35193
rect 11503 35184 11515 35187
rect 11466 35156 11515 35184
rect 11466 35144 11472 35156
rect 11503 35153 11515 35156
rect 11549 35153 11561 35187
rect 11503 35147 11561 35153
rect 13251 35187 13309 35193
rect 13251 35153 13263 35187
rect 13297 35153 13309 35187
rect 13251 35147 13309 35153
rect 13435 35187 13493 35193
rect 13435 35153 13447 35187
rect 13481 35153 13493 35187
rect 14720 35184 14726 35196
rect 14681 35156 14726 35184
rect 13435 35147 13493 35153
rect 4232 35076 4238 35128
rect 4290 35116 4296 35128
rect 5247 35119 5305 35125
rect 5247 35116 5259 35119
rect 4290 35088 5259 35116
rect 4290 35076 4296 35088
rect 5247 35085 5259 35088
rect 5293 35085 5305 35119
rect 5247 35079 5305 35085
rect 9847 35119 9905 35125
rect 9847 35085 9859 35119
rect 9893 35116 9905 35119
rect 11316 35116 11322 35128
rect 9893 35088 11322 35116
rect 9893 35085 9905 35088
rect 9847 35079 9905 35085
rect 5262 34980 5290 35079
rect 11316 35076 11322 35088
rect 11374 35076 11380 35128
rect 13266 35116 13294 35147
rect 14720 35144 14726 35156
rect 14778 35144 14784 35196
rect 18786 35193 18814 35224
rect 20148 35212 20154 35224
rect 20206 35212 20212 35264
rect 23187 35255 23245 35261
rect 23187 35252 23199 35255
rect 22374 35224 23199 35252
rect 14815 35187 14873 35193
rect 14815 35153 14827 35187
rect 14861 35184 14873 35187
rect 18771 35187 18829 35193
rect 14861 35156 16146 35184
rect 14861 35153 14873 35156
rect 14815 35147 14873 35153
rect 14830 35116 14858 35147
rect 13266 35088 14858 35116
rect 15548 35076 15554 35128
rect 15606 35116 15612 35128
rect 15735 35119 15793 35125
rect 15735 35116 15747 35119
rect 15606 35088 15747 35116
rect 15606 35076 15612 35088
rect 15735 35085 15747 35088
rect 15781 35085 15793 35119
rect 16008 35116 16014 35128
rect 15969 35088 16014 35116
rect 15735 35079 15793 35085
rect 16008 35076 16014 35088
rect 16066 35076 16072 35128
rect 16118 35116 16146 35156
rect 18771 35153 18783 35187
rect 18817 35153 18829 35187
rect 18771 35147 18829 35153
rect 18952 35144 18958 35196
rect 19010 35184 19016 35196
rect 19047 35187 19105 35193
rect 19047 35184 19059 35187
rect 19010 35156 19059 35184
rect 19010 35144 19016 35156
rect 19047 35153 19059 35156
rect 19093 35153 19105 35187
rect 19231 35187 19289 35193
rect 19231 35184 19243 35187
rect 19047 35147 19105 35153
rect 19154 35156 19243 35184
rect 19154 35116 19182 35156
rect 19231 35153 19243 35156
rect 19277 35184 19289 35187
rect 21068 35184 21074 35196
rect 19277 35156 21074 35184
rect 19277 35153 19289 35156
rect 19231 35147 19289 35153
rect 21068 35144 21074 35156
rect 21126 35144 21132 35196
rect 21712 35144 21718 35196
rect 21770 35184 21776 35196
rect 22374 35193 22402 35224
rect 23187 35221 23199 35224
rect 23233 35252 23245 35255
rect 23371 35255 23429 35261
rect 23371 35252 23383 35255
rect 23233 35224 23383 35252
rect 23233 35221 23245 35224
rect 23187 35215 23245 35221
rect 23371 35221 23383 35224
rect 23417 35252 23429 35255
rect 24564 35252 24570 35264
rect 23417 35224 24570 35252
rect 23417 35221 23429 35224
rect 23371 35215 23429 35221
rect 24564 35212 24570 35224
rect 24622 35212 24628 35264
rect 28354 35252 28382 35292
rect 29256 35280 29262 35292
rect 29314 35280 29320 35332
rect 29535 35323 29593 35329
rect 29535 35289 29547 35323
rect 29581 35320 29593 35323
rect 35512 35320 35518 35332
rect 29581 35292 35518 35320
rect 29581 35289 29593 35292
rect 29535 35283 29593 35289
rect 35512 35280 35518 35292
rect 35570 35280 35576 35332
rect 39103 35323 39161 35329
rect 35622 35292 38502 35320
rect 27802 35224 28382 35252
rect 21807 35187 21865 35193
rect 21807 35184 21819 35187
rect 21770 35156 21819 35184
rect 21770 35144 21776 35156
rect 21807 35153 21819 35156
rect 21853 35184 21865 35187
rect 22359 35187 22417 35193
rect 22359 35184 22371 35187
rect 21853 35156 22371 35184
rect 21853 35153 21865 35156
rect 21807 35147 21865 35153
rect 22359 35153 22371 35156
rect 22405 35153 22417 35187
rect 22359 35147 22417 35153
rect 22543 35187 22601 35193
rect 22543 35153 22555 35187
rect 22589 35184 22601 35187
rect 23276 35184 23282 35196
rect 22589 35156 23282 35184
rect 22589 35153 22601 35156
rect 22543 35147 22601 35153
rect 23276 35144 23282 35156
rect 23334 35144 23340 35196
rect 23828 35184 23834 35196
rect 23789 35156 23834 35184
rect 23828 35144 23834 35156
rect 23886 35184 23892 35196
rect 24199 35187 24257 35193
rect 24199 35184 24211 35187
rect 23886 35156 24211 35184
rect 23886 35144 23892 35156
rect 24199 35153 24211 35156
rect 24245 35153 24257 35187
rect 24199 35147 24257 35153
rect 26959 35187 27017 35193
rect 26959 35153 26971 35187
rect 27005 35184 27017 35187
rect 27048 35184 27054 35196
rect 27005 35156 27054 35184
rect 27005 35153 27017 35156
rect 26959 35147 27017 35153
rect 27048 35144 27054 35156
rect 27106 35144 27112 35196
rect 27802 35193 27830 35224
rect 28980 35212 28986 35264
rect 29038 35252 29044 35264
rect 29038 35224 30406 35252
rect 29038 35212 29044 35224
rect 27235 35187 27293 35193
rect 27235 35153 27247 35187
rect 27281 35184 27293 35187
rect 27787 35187 27845 35193
rect 27787 35184 27799 35187
rect 27281 35156 27799 35184
rect 27281 35153 27293 35156
rect 27235 35147 27293 35153
rect 27787 35153 27799 35156
rect 27833 35153 27845 35187
rect 27787 35147 27845 35153
rect 27971 35187 28029 35193
rect 27971 35153 27983 35187
rect 28017 35184 28029 35187
rect 28796 35184 28802 35196
rect 28017 35156 28802 35184
rect 28017 35153 28029 35156
rect 27971 35147 28029 35153
rect 28796 35144 28802 35156
rect 28854 35184 28860 35196
rect 29719 35187 29777 35193
rect 29719 35184 29731 35187
rect 28854 35156 29731 35184
rect 28854 35144 28860 35156
rect 29719 35153 29731 35156
rect 29765 35153 29777 35187
rect 29719 35147 29777 35153
rect 29903 35187 29961 35193
rect 29903 35153 29915 35187
rect 29949 35153 29961 35187
rect 30268 35184 30274 35196
rect 30229 35156 30274 35184
rect 29903 35147 29961 35153
rect 16118 35088 19182 35116
rect 21623 35119 21681 35125
rect 21623 35085 21635 35119
rect 21669 35085 21681 35119
rect 29918 35116 29946 35147
rect 30268 35144 30274 35156
rect 30326 35144 30332 35196
rect 30378 35193 30406 35224
rect 30452 35212 30458 35264
rect 30510 35252 30516 35264
rect 30510 35224 33258 35252
rect 30510 35212 30516 35224
rect 30363 35187 30421 35193
rect 30363 35153 30375 35187
rect 30409 35153 30421 35187
rect 30363 35147 30421 35153
rect 32016 35144 32022 35196
rect 32074 35184 32080 35196
rect 33120 35184 33126 35196
rect 32074 35156 33126 35184
rect 32074 35144 32080 35156
rect 33120 35144 33126 35156
rect 33178 35144 33184 35196
rect 30084 35116 30090 35128
rect 29918 35088 30090 35116
rect 21623 35079 21681 35085
rect 21638 35048 21666 35079
rect 30084 35076 30090 35088
rect 30142 35116 30148 35128
rect 30639 35119 30697 35125
rect 30639 35116 30651 35119
rect 30142 35088 30651 35116
rect 30142 35076 30148 35088
rect 30639 35085 30651 35088
rect 30685 35116 30697 35119
rect 30728 35116 30734 35128
rect 30685 35088 30734 35116
rect 30685 35085 30697 35088
rect 30639 35079 30697 35085
rect 30728 35076 30734 35088
rect 30786 35076 30792 35128
rect 33230 35116 33258 35224
rect 33396 35184 33402 35196
rect 33357 35156 33402 35184
rect 33396 35144 33402 35156
rect 33454 35144 33460 35196
rect 34224 35184 34230 35196
rect 33506 35156 34230 35184
rect 33506 35116 33534 35156
rect 34224 35144 34230 35156
rect 34282 35144 34288 35196
rect 35622 35193 35650 35292
rect 38474 35252 38502 35292
rect 39103 35289 39115 35323
rect 39149 35320 39161 35323
rect 40020 35320 40026 35332
rect 39149 35292 40026 35320
rect 39149 35289 39161 35292
rect 39103 35283 39161 35289
rect 40020 35280 40026 35292
rect 40078 35280 40084 35332
rect 43056 35320 43062 35332
rect 43017 35292 43062 35320
rect 43056 35280 43062 35292
rect 43114 35280 43120 35332
rect 46092 35280 46098 35332
rect 46150 35320 46156 35332
rect 47567 35323 47625 35329
rect 47567 35320 47579 35323
rect 46150 35292 47579 35320
rect 46150 35280 46156 35292
rect 47567 35289 47579 35292
rect 47613 35320 47625 35323
rect 48208 35320 48214 35332
rect 47613 35292 48214 35320
rect 47613 35289 47625 35292
rect 47567 35283 47625 35289
rect 48208 35280 48214 35292
rect 48266 35280 48272 35332
rect 49312 35320 49318 35332
rect 49273 35292 49318 35320
rect 49312 35280 49318 35292
rect 49370 35280 49376 35332
rect 49404 35280 49410 35332
rect 49462 35320 49468 35332
rect 62100 35320 62106 35332
rect 49462 35292 62106 35320
rect 49462 35280 49468 35292
rect 62100 35280 62106 35292
rect 62158 35280 62164 35332
rect 62379 35323 62437 35329
rect 62379 35289 62391 35323
rect 62425 35320 62437 35323
rect 64032 35320 64038 35332
rect 62425 35292 64038 35320
rect 62425 35289 62437 35292
rect 62379 35283 62437 35289
rect 64032 35280 64038 35292
rect 64090 35280 64096 35332
rect 64124 35280 64130 35332
rect 64182 35320 64188 35332
rect 69552 35320 69558 35332
rect 64182 35292 69558 35320
rect 64182 35280 64188 35292
rect 69552 35280 69558 35292
rect 69610 35280 69616 35332
rect 69644 35280 69650 35332
rect 69702 35320 69708 35332
rect 75440 35320 75446 35332
rect 69702 35292 75446 35320
rect 69702 35280 69708 35292
rect 75440 35280 75446 35292
rect 75498 35280 75504 35332
rect 80684 35280 80690 35332
rect 80742 35320 80748 35332
rect 80963 35323 81021 35329
rect 80963 35320 80975 35323
rect 80742 35292 80975 35320
rect 80742 35280 80748 35292
rect 80963 35289 80975 35292
rect 81009 35289 81021 35323
rect 83904 35320 83910 35332
rect 80963 35283 81021 35289
rect 83278 35292 83910 35320
rect 40572 35252 40578 35264
rect 38474 35224 40578 35252
rect 40572 35212 40578 35224
rect 40630 35212 40636 35264
rect 34779 35187 34837 35193
rect 34779 35153 34791 35187
rect 34825 35184 34837 35187
rect 35607 35187 35665 35193
rect 35607 35184 35619 35187
rect 34825 35156 35619 35184
rect 34825 35153 34837 35156
rect 34779 35147 34837 35153
rect 35607 35153 35619 35156
rect 35653 35153 35665 35187
rect 35607 35147 35665 35153
rect 35699 35187 35757 35193
rect 35699 35153 35711 35187
rect 35745 35184 35757 35187
rect 36064 35184 36070 35196
rect 35745 35156 36070 35184
rect 35745 35153 35757 35156
rect 35699 35147 35757 35153
rect 36064 35144 36070 35156
rect 36122 35144 36128 35196
rect 37812 35184 37818 35196
rect 37773 35156 37818 35184
rect 37812 35144 37818 35156
rect 37870 35144 37876 35196
rect 39836 35144 39842 35196
rect 39894 35184 39900 35196
rect 40023 35187 40081 35193
rect 40023 35184 40035 35187
rect 39894 35156 40035 35184
rect 39894 35144 39900 35156
rect 40023 35153 40035 35156
rect 40069 35153 40081 35187
rect 43074 35184 43102 35280
rect 47472 35212 47478 35264
rect 47530 35252 47536 35264
rect 50235 35255 50293 35261
rect 47530 35224 49634 35252
rect 47530 35212 47536 35224
rect 43243 35187 43301 35193
rect 43243 35184 43255 35187
rect 43074 35156 43255 35184
rect 40023 35147 40081 35153
rect 43243 35153 43255 35156
rect 43289 35153 43301 35187
rect 43243 35147 43301 35153
rect 43519 35187 43577 35193
rect 43519 35153 43531 35187
rect 43565 35184 43577 35187
rect 44160 35184 44166 35196
rect 43565 35156 44166 35184
rect 43565 35153 43577 35156
rect 43519 35147 43577 35153
rect 44160 35144 44166 35156
rect 44218 35144 44224 35196
rect 44899 35187 44957 35193
rect 44899 35153 44911 35187
rect 44945 35184 44957 35187
rect 45172 35184 45178 35196
rect 44945 35156 45178 35184
rect 44945 35153 44957 35156
rect 44899 35147 44957 35153
rect 45172 35144 45178 35156
rect 45230 35144 45236 35196
rect 46003 35187 46061 35193
rect 46003 35153 46015 35187
rect 46049 35184 46061 35187
rect 47564 35184 47570 35196
rect 46049 35156 47570 35184
rect 46049 35153 46061 35156
rect 46003 35147 46061 35153
rect 47564 35144 47570 35156
rect 47622 35144 47628 35196
rect 49312 35144 49318 35196
rect 49370 35184 49376 35196
rect 49606 35193 49634 35224
rect 50235 35221 50247 35255
rect 50281 35252 50293 35255
rect 50281 35224 53958 35252
rect 50281 35221 50293 35224
rect 50235 35215 50293 35221
rect 49499 35187 49557 35193
rect 49499 35184 49511 35187
rect 49370 35156 49511 35184
rect 49370 35144 49376 35156
rect 49499 35153 49511 35156
rect 49545 35153 49557 35187
rect 49499 35147 49557 35153
rect 49591 35187 49649 35193
rect 49591 35153 49603 35187
rect 49637 35153 49649 35187
rect 49591 35147 49649 35153
rect 49775 35187 49833 35193
rect 49775 35153 49787 35187
rect 49821 35184 49833 35187
rect 51247 35187 51305 35193
rect 51247 35184 51259 35187
rect 49821 35156 51259 35184
rect 49821 35153 49833 35156
rect 49775 35147 49833 35153
rect 51247 35153 51259 35156
rect 51293 35153 51305 35187
rect 51888 35184 51894 35196
rect 51849 35156 51894 35184
rect 51247 35147 51305 35153
rect 51888 35144 51894 35156
rect 51946 35144 51952 35196
rect 52072 35184 52078 35196
rect 51998 35156 52078 35184
rect 33230 35088 33534 35116
rect 37539 35119 37597 35125
rect 37539 35085 37551 35119
rect 37585 35085 37597 35119
rect 37539 35079 37597 35085
rect 22724 35048 22730 35060
rect 10782 35020 15778 35048
rect 7084 34980 7090 34992
rect 5262 34952 7090 34980
rect 7084 34940 7090 34952
rect 7142 34940 7148 34992
rect 8372 34940 8378 34992
rect 8430 34980 8436 34992
rect 10782 34980 10810 35020
rect 8430 34952 10810 34980
rect 8430 34940 8436 34952
rect 11316 34940 11322 34992
rect 11374 34980 11380 34992
rect 11595 34983 11653 34989
rect 11595 34980 11607 34983
rect 11374 34952 11607 34980
rect 11374 34940 11380 34952
rect 11595 34949 11607 34952
rect 11641 34949 11653 34983
rect 13524 34980 13530 34992
rect 13485 34952 13530 34980
rect 11595 34943 11653 34949
rect 13524 34940 13530 34952
rect 13582 34940 13588 34992
rect 15750 34980 15778 35020
rect 17130 35020 21666 35048
rect 22685 35020 22730 35048
rect 17130 34980 17158 35020
rect 17296 34980 17302 34992
rect 15750 34952 17158 34980
rect 17257 34952 17302 34980
rect 17296 34940 17302 34952
rect 17354 34940 17360 34992
rect 21531 34983 21589 34989
rect 21531 34949 21543 34983
rect 21577 34980 21589 34983
rect 21638 34980 21666 35020
rect 22724 35008 22730 35020
rect 22782 35008 22788 35060
rect 34592 35008 34598 35060
rect 34650 35048 34656 35060
rect 34871 35051 34929 35057
rect 34871 35048 34883 35051
rect 34650 35020 34883 35048
rect 34650 35008 34656 35020
rect 34871 35017 34883 35020
rect 34917 35048 34929 35051
rect 37168 35048 37174 35060
rect 34917 35020 37174 35048
rect 34917 35017 34929 35020
rect 34871 35011 34929 35017
rect 37168 35008 37174 35020
rect 37226 35048 37232 35060
rect 37355 35051 37413 35057
rect 37355 35048 37367 35051
rect 37226 35020 37367 35048
rect 37226 35008 37232 35020
rect 37355 35017 37367 35020
rect 37401 35048 37413 35051
rect 37554 35048 37582 35079
rect 40112 35076 40118 35128
rect 40170 35116 40176 35128
rect 43424 35116 43430 35128
rect 40170 35088 43430 35116
rect 40170 35076 40176 35088
rect 43424 35076 43430 35088
rect 43482 35076 43488 35128
rect 45727 35119 45785 35125
rect 45727 35085 45739 35119
rect 45773 35116 45785 35119
rect 46092 35116 46098 35128
rect 45773 35088 46098 35116
rect 45773 35085 45785 35088
rect 45727 35079 45785 35085
rect 46092 35076 46098 35088
rect 46150 35076 46156 35128
rect 51998 35125 52026 35156
rect 52072 35144 52078 35156
rect 52130 35144 52136 35196
rect 52259 35187 52317 35193
rect 52259 35153 52271 35187
rect 52305 35184 52317 35187
rect 52443 35187 52501 35193
rect 52305 35156 52394 35184
rect 52305 35153 52317 35156
rect 52259 35147 52317 35153
rect 51983 35119 52041 35125
rect 46662 35088 49726 35116
rect 37401 35020 37582 35048
rect 38474 35020 43286 35048
rect 37401 35017 37413 35020
rect 37355 35011 37413 35017
rect 24288 34980 24294 34992
rect 21577 34952 24294 34980
rect 21577 34949 21589 34952
rect 21531 34943 21589 34949
rect 24288 34940 24294 34952
rect 24346 34940 24352 34992
rect 30636 34940 30642 34992
rect 30694 34980 30700 34992
rect 38474 34980 38502 35020
rect 30694 34952 38502 34980
rect 30694 34940 30700 34952
rect 39468 34940 39474 34992
rect 39526 34980 39532 34992
rect 40115 34983 40173 34989
rect 40115 34980 40127 34983
rect 39526 34952 40127 34980
rect 39526 34940 39532 34952
rect 40115 34949 40127 34952
rect 40161 34980 40173 34983
rect 41308 34980 41314 34992
rect 40161 34952 41314 34980
rect 40161 34949 40173 34952
rect 40115 34943 40173 34949
rect 41308 34940 41314 34952
rect 41366 34940 41372 34992
rect 43258 34980 43286 35020
rect 44178 35020 45586 35048
rect 44178 34980 44206 35020
rect 43258 34952 44206 34980
rect 45558 34980 45586 35020
rect 46662 34980 46690 35088
rect 49698 35048 49726 35088
rect 51983 35085 51995 35119
rect 52029 35085 52041 35119
rect 52366 35116 52394 35156
rect 52443 35153 52455 35187
rect 52489 35184 52501 35187
rect 53360 35184 53366 35196
rect 52489 35156 53366 35184
rect 52489 35153 52501 35156
rect 52443 35147 52501 35153
rect 53360 35144 53366 35156
rect 53418 35144 53424 35196
rect 52716 35116 52722 35128
rect 52366 35088 52722 35116
rect 51983 35079 52041 35085
rect 52716 35076 52722 35088
rect 52774 35076 52780 35128
rect 53930 35116 53958 35224
rect 54096 35212 54102 35264
rect 54154 35252 54160 35264
rect 54927 35255 54985 35261
rect 54927 35252 54939 35255
rect 54154 35224 54939 35252
rect 54154 35212 54160 35224
rect 54927 35221 54939 35224
rect 54973 35252 54985 35255
rect 60812 35252 60818 35264
rect 54973 35224 60818 35252
rect 54973 35221 54985 35224
rect 54927 35215 54985 35221
rect 60812 35212 60818 35224
rect 60870 35212 60876 35264
rect 63296 35212 63302 35264
rect 63354 35252 63360 35264
rect 68543 35255 68601 35261
rect 68543 35252 68555 35255
rect 63354 35224 68555 35252
rect 63354 35212 63360 35224
rect 68543 35221 68555 35224
rect 68589 35221 68601 35255
rect 68543 35215 68601 35221
rect 80868 35212 80874 35264
rect 80926 35252 80932 35264
rect 82064 35252 82070 35264
rect 80926 35224 82070 35252
rect 80926 35212 80932 35224
rect 82064 35212 82070 35224
rect 82122 35212 82128 35264
rect 54007 35187 54065 35193
rect 54007 35153 54019 35187
rect 54053 35184 54065 35187
rect 62379 35187 62437 35193
rect 62379 35184 62391 35187
rect 54053 35156 62391 35184
rect 54053 35153 54065 35156
rect 54007 35147 54065 35153
rect 62379 35153 62391 35156
rect 62425 35153 62437 35187
rect 62379 35147 62437 35153
rect 62560 35144 62566 35196
rect 62618 35193 62624 35196
rect 62618 35187 62667 35193
rect 62618 35153 62621 35187
rect 62655 35153 62667 35187
rect 62618 35147 62667 35153
rect 62747 35187 62805 35193
rect 62747 35153 62759 35187
rect 62793 35184 62805 35187
rect 63112 35184 63118 35196
rect 62793 35156 63118 35184
rect 62793 35153 62805 35156
rect 62747 35147 62805 35153
rect 62618 35144 62624 35147
rect 63112 35144 63118 35156
rect 63170 35144 63176 35196
rect 63204 35144 63210 35196
rect 63262 35184 63268 35196
rect 65872 35184 65878 35196
rect 63262 35156 63783 35184
rect 65833 35156 65878 35184
rect 63262 35144 63268 35156
rect 54375 35119 54433 35125
rect 54375 35116 54387 35119
rect 53930 35088 54387 35116
rect 54375 35085 54387 35088
rect 54421 35085 54433 35119
rect 54648 35116 54654 35128
rect 54609 35088 54654 35116
rect 54375 35079 54433 35085
rect 54648 35076 54654 35088
rect 54706 35076 54712 35128
rect 55844 35076 55850 35128
rect 55902 35116 55908 35128
rect 62100 35116 62106 35128
rect 55902 35088 62106 35116
rect 55902 35076 55908 35088
rect 62100 35076 62106 35088
rect 62158 35076 62164 35128
rect 63755 35116 63783 35156
rect 65872 35144 65878 35156
rect 65930 35184 65936 35196
rect 66151 35187 66209 35193
rect 66151 35184 66163 35187
rect 65930 35156 66163 35184
rect 65930 35144 65936 35156
rect 66151 35153 66163 35156
rect 66197 35153 66209 35187
rect 66151 35147 66209 35153
rect 68356 35144 68362 35196
rect 68414 35184 68420 35196
rect 69187 35187 69245 35193
rect 69187 35184 69199 35187
rect 68414 35156 69199 35184
rect 68414 35144 68420 35156
rect 69187 35153 69199 35156
rect 69233 35153 69245 35187
rect 69187 35147 69245 35153
rect 69555 35187 69613 35193
rect 69555 35153 69567 35187
rect 69601 35184 69613 35187
rect 70656 35184 70662 35196
rect 69601 35156 70662 35184
rect 69601 35153 69613 35156
rect 69555 35147 69613 35153
rect 70656 35144 70662 35156
rect 70714 35184 70720 35196
rect 70843 35187 70901 35193
rect 70843 35184 70855 35187
rect 70714 35156 70855 35184
rect 70714 35144 70720 35156
rect 70843 35153 70855 35156
rect 70889 35153 70901 35187
rect 70843 35147 70901 35153
rect 73232 35144 73238 35196
rect 73290 35184 73296 35196
rect 73879 35187 73937 35193
rect 73879 35184 73891 35187
rect 73290 35156 73891 35184
rect 73290 35144 73296 35156
rect 73879 35153 73891 35156
rect 73925 35184 73937 35187
rect 73968 35184 73974 35196
rect 73925 35156 73974 35184
rect 73925 35153 73937 35156
rect 73879 35147 73937 35153
rect 73968 35144 73974 35156
rect 74026 35144 74032 35196
rect 74152 35184 74158 35196
rect 74113 35156 74158 35184
rect 74152 35144 74158 35156
rect 74210 35144 74216 35196
rect 79215 35187 79273 35193
rect 79215 35184 79227 35187
rect 76746 35156 79227 35184
rect 67896 35116 67902 35128
rect 63755 35088 67902 35116
rect 67896 35076 67902 35088
rect 67954 35076 67960 35128
rect 68172 35076 68178 35128
rect 68230 35116 68236 35128
rect 69276 35116 69282 35128
rect 68230 35088 69138 35116
rect 69237 35088 69282 35116
rect 68230 35076 68236 35088
rect 63388 35048 63394 35060
rect 49698 35020 63394 35048
rect 63388 35008 63394 35020
rect 63446 35008 63452 35060
rect 69110 35048 69138 35088
rect 69276 35076 69282 35088
rect 69334 35076 69340 35128
rect 69647 35119 69705 35125
rect 69647 35085 69659 35119
rect 69693 35116 69705 35119
rect 69920 35116 69926 35128
rect 69693 35088 69926 35116
rect 69693 35085 69705 35088
rect 69647 35079 69705 35085
rect 69920 35076 69926 35088
rect 69978 35076 69984 35128
rect 73986 35116 74014 35144
rect 76746 35128 76774 35156
rect 79215 35153 79227 35156
rect 79261 35184 79273 35187
rect 79399 35187 79457 35193
rect 79399 35184 79411 35187
rect 79261 35156 79411 35184
rect 79261 35153 79273 35156
rect 79215 35147 79273 35153
rect 79399 35153 79411 35156
rect 79445 35184 79457 35187
rect 79675 35187 79733 35193
rect 79445 35156 79626 35184
rect 79445 35153 79457 35156
rect 79399 35147 79457 35153
rect 75627 35119 75685 35125
rect 75627 35116 75639 35119
rect 73986 35088 75639 35116
rect 75627 35085 75639 35088
rect 75673 35116 75685 35119
rect 76728 35116 76734 35128
rect 75673 35088 76734 35116
rect 75673 35085 75685 35088
rect 75627 35079 75685 35085
rect 76728 35076 76734 35088
rect 76786 35076 76792 35128
rect 79598 35116 79626 35156
rect 79675 35153 79687 35187
rect 79721 35184 79733 35187
rect 81144 35184 81150 35196
rect 79721 35156 81150 35184
rect 79721 35153 79733 35156
rect 79675 35147 79733 35153
rect 81144 35144 81150 35156
rect 81202 35144 81208 35196
rect 83278 35193 83306 35292
rect 83904 35280 83910 35292
rect 83962 35320 83968 35332
rect 89516 35320 89522 35332
rect 83962 35292 89522 35320
rect 83962 35280 83968 35292
rect 89516 35280 89522 35292
rect 89574 35280 89580 35332
rect 83079 35187 83137 35193
rect 83079 35184 83091 35187
rect 81254 35156 83091 35184
rect 81254 35116 81282 35156
rect 83079 35153 83091 35156
rect 83125 35184 83137 35187
rect 83263 35187 83321 35193
rect 83263 35184 83275 35187
rect 83125 35156 83275 35184
rect 83125 35153 83137 35156
rect 83079 35147 83137 35153
rect 83263 35153 83275 35156
rect 83309 35153 83321 35187
rect 83536 35184 83542 35196
rect 83497 35156 83542 35184
rect 83263 35147 83321 35153
rect 83536 35144 83542 35156
rect 83594 35144 83600 35196
rect 89534 35184 89562 35280
rect 89703 35187 89761 35193
rect 89703 35184 89715 35187
rect 89534 35156 89715 35184
rect 89703 35153 89715 35156
rect 89749 35153 89761 35187
rect 89976 35184 89982 35196
rect 89937 35156 89982 35184
rect 89703 35147 89761 35153
rect 89976 35144 89982 35156
rect 90034 35144 90040 35196
rect 79598 35088 81282 35116
rect 69736 35048 69742 35060
rect 63590 35020 68770 35048
rect 69110 35020 69742 35048
rect 45558 34952 46690 34980
rect 46920 34940 46926 34992
rect 46978 34980 46984 34992
rect 47107 34983 47165 34989
rect 47107 34980 47119 34983
rect 46978 34952 47119 34980
rect 46978 34940 46984 34952
rect 47107 34949 47119 34952
rect 47153 34949 47165 34983
rect 52624 34980 52630 34992
rect 52585 34952 52630 34980
rect 47107 34943 47165 34949
rect 52624 34940 52630 34952
rect 52682 34940 52688 34992
rect 52716 34940 52722 34992
rect 52774 34980 52780 34992
rect 52774 34952 52819 34980
rect 52774 34940 52780 34952
rect 54096 34940 54102 34992
rect 54154 34989 54160 34992
rect 54154 34983 54203 34989
rect 54154 34949 54157 34983
rect 54191 34949 54203 34983
rect 54280 34980 54286 34992
rect 54241 34952 54286 34980
rect 54154 34943 54203 34949
rect 54154 34940 54160 34943
rect 54280 34940 54286 34952
rect 54338 34940 54344 34992
rect 55292 34940 55298 34992
rect 55350 34980 55356 34992
rect 63590 34980 63618 35020
rect 55350 34952 63618 34980
rect 63667 34983 63725 34989
rect 55350 34940 55356 34952
rect 63667 34949 63679 34983
rect 63713 34980 63725 34983
rect 63848 34980 63854 34992
rect 63713 34952 63854 34980
rect 63713 34949 63725 34952
rect 63667 34943 63725 34949
rect 63848 34940 63854 34952
rect 63906 34940 63912 34992
rect 65964 34980 65970 34992
rect 65925 34952 65970 34980
rect 65964 34940 65970 34952
rect 66022 34940 66028 34992
rect 68356 34980 68362 34992
rect 68317 34952 68362 34980
rect 68356 34940 68362 34952
rect 68414 34940 68420 34992
rect 68742 34980 68770 35020
rect 69736 35008 69742 35020
rect 69794 35048 69800 35060
rect 70935 35051 70993 35057
rect 70935 35048 70947 35051
rect 69794 35020 70947 35048
rect 69794 35008 69800 35020
rect 70935 35017 70947 35020
rect 70981 35017 70993 35051
rect 70935 35011 70993 35017
rect 74814 35020 75578 35048
rect 74814 34980 74842 35020
rect 68742 34952 74842 34980
rect 75259 34983 75317 34989
rect 75259 34949 75271 34983
rect 75305 34980 75317 34983
rect 75440 34980 75446 34992
rect 75305 34952 75446 34980
rect 75305 34949 75317 34952
rect 75259 34943 75317 34949
rect 75440 34940 75446 34952
rect 75498 34940 75504 34992
rect 75550 34980 75578 35020
rect 84272 35008 84278 35060
rect 84330 35048 84336 35060
rect 84330 35020 89654 35048
rect 84330 35008 84336 35020
rect 82892 34980 82898 34992
rect 75550 34952 82898 34980
rect 82892 34940 82898 34952
rect 82950 34940 82956 34992
rect 84640 34980 84646 34992
rect 84601 34952 84646 34980
rect 84640 34940 84646 34952
rect 84698 34940 84704 34992
rect 89626 34980 89654 35020
rect 90620 34980 90626 34992
rect 89626 34952 90626 34980
rect 90620 34940 90626 34952
rect 90678 34940 90684 34992
rect 91080 34980 91086 34992
rect 91041 34952 91086 34980
rect 91080 34940 91086 34952
rect 91138 34940 91144 34992
rect 538 34890 93642 34912
rect 538 34838 3680 34890
rect 3732 34838 3744 34890
rect 3796 34838 3808 34890
rect 3860 34838 3872 34890
rect 3924 34838 9008 34890
rect 9060 34838 9072 34890
rect 9124 34838 9136 34890
rect 9188 34838 9200 34890
rect 9252 34838 14336 34890
rect 14388 34838 14400 34890
rect 14452 34838 14464 34890
rect 14516 34838 14528 34890
rect 14580 34838 19664 34890
rect 19716 34838 19728 34890
rect 19780 34838 19792 34890
rect 19844 34838 19856 34890
rect 19908 34838 24992 34890
rect 25044 34838 25056 34890
rect 25108 34838 25120 34890
rect 25172 34838 25184 34890
rect 25236 34838 30320 34890
rect 30372 34838 30384 34890
rect 30436 34838 30448 34890
rect 30500 34838 30512 34890
rect 30564 34838 35648 34890
rect 35700 34838 35712 34890
rect 35764 34838 35776 34890
rect 35828 34838 35840 34890
rect 35892 34838 40976 34890
rect 41028 34838 41040 34890
rect 41092 34838 41104 34890
rect 41156 34838 41168 34890
rect 41220 34838 46304 34890
rect 46356 34838 46368 34890
rect 46420 34838 46432 34890
rect 46484 34838 46496 34890
rect 46548 34838 51632 34890
rect 51684 34838 51696 34890
rect 51748 34838 51760 34890
rect 51812 34838 51824 34890
rect 51876 34838 56960 34890
rect 57012 34838 57024 34890
rect 57076 34838 57088 34890
rect 57140 34838 57152 34890
rect 57204 34838 62288 34890
rect 62340 34838 62352 34890
rect 62404 34838 62416 34890
rect 62468 34838 62480 34890
rect 62532 34838 67616 34890
rect 67668 34838 67680 34890
rect 67732 34838 67744 34890
rect 67796 34838 67808 34890
rect 67860 34838 72944 34890
rect 72996 34838 73008 34890
rect 73060 34838 73072 34890
rect 73124 34838 73136 34890
rect 73188 34838 78272 34890
rect 78324 34838 78336 34890
rect 78388 34838 78400 34890
rect 78452 34838 78464 34890
rect 78516 34838 83600 34890
rect 83652 34838 83664 34890
rect 83716 34838 83728 34890
rect 83780 34838 83792 34890
rect 83844 34838 88928 34890
rect 88980 34838 88992 34890
rect 89044 34838 89056 34890
rect 89108 34838 89120 34890
rect 89172 34838 93642 34890
rect 538 34816 93642 34838
rect 4143 34779 4201 34785
rect 4143 34776 4155 34779
rect 2318 34748 4155 34776
rect 2318 34649 2346 34748
rect 4143 34745 4155 34748
rect 4189 34776 4201 34779
rect 4232 34776 4238 34788
rect 4189 34748 4238 34776
rect 4189 34745 4201 34748
rect 4143 34739 4201 34745
rect 4232 34736 4238 34748
rect 4290 34736 4296 34788
rect 12788 34776 12794 34788
rect 12749 34748 12794 34776
rect 12788 34736 12794 34748
rect 12846 34736 12852 34788
rect 16100 34736 16106 34788
rect 16158 34776 16164 34788
rect 17023 34779 17081 34785
rect 17023 34776 17035 34779
rect 16158 34748 17035 34776
rect 16158 34736 16164 34748
rect 17023 34745 17035 34748
rect 17069 34745 17081 34779
rect 17023 34739 17081 34745
rect 18679 34779 18737 34785
rect 18679 34745 18691 34779
rect 18725 34776 18737 34779
rect 21160 34776 21166 34788
rect 18725 34748 21166 34776
rect 18725 34745 18737 34748
rect 18679 34739 18737 34745
rect 2303 34643 2361 34649
rect 2303 34609 2315 34643
rect 2349 34609 2361 34643
rect 2303 34603 2361 34609
rect 16836 34600 16842 34652
rect 16894 34640 16900 34652
rect 16894 34612 17710 34640
rect 16894 34600 16900 34612
rect 2576 34572 2582 34584
rect 2537 34544 2582 34572
rect 2576 34532 2582 34544
rect 2634 34532 2640 34584
rect 3220 34532 3226 34584
rect 3278 34572 3284 34584
rect 6351 34575 6409 34581
rect 6351 34572 6363 34575
rect 3278 34544 6363 34572
rect 3278 34532 3284 34544
rect 6351 34541 6363 34544
rect 6397 34572 6409 34575
rect 6443 34575 6501 34581
rect 6443 34572 6455 34575
rect 6397 34544 6455 34572
rect 6397 34541 6409 34544
rect 6351 34535 6409 34541
rect 6443 34541 6455 34544
rect 6489 34572 6501 34575
rect 9108 34572 9114 34584
rect 6489 34544 9114 34572
rect 6489 34541 6501 34544
rect 6443 34535 6501 34541
rect 9108 34532 9114 34544
rect 9166 34572 9172 34584
rect 9476 34572 9482 34584
rect 9166 34544 9482 34572
rect 9166 34532 9172 34544
rect 9476 34532 9482 34544
rect 9534 34532 9540 34584
rect 12788 34532 12794 34584
rect 12846 34572 12852 34584
rect 12883 34575 12941 34581
rect 12883 34572 12895 34575
rect 12846 34544 12895 34572
rect 12846 34532 12852 34544
rect 12883 34541 12895 34544
rect 12929 34541 12941 34575
rect 12883 34535 12941 34541
rect 17207 34575 17265 34581
rect 17207 34541 17219 34575
rect 17253 34572 17265 34575
rect 17253 34544 17618 34572
rect 17253 34541 17265 34544
rect 17207 34535 17265 34541
rect 6535 34507 6593 34513
rect 6535 34473 6547 34507
rect 6581 34504 6593 34507
rect 6624 34504 6630 34516
rect 6581 34476 6630 34504
rect 6581 34473 6593 34476
rect 6535 34467 6593 34473
rect 6624 34464 6630 34476
rect 6682 34464 6688 34516
rect 3864 34436 3870 34448
rect 3825 34408 3870 34436
rect 3864 34396 3870 34408
rect 3922 34396 3928 34448
rect 13064 34436 13070 34448
rect 13025 34408 13070 34436
rect 13064 34396 13070 34408
rect 13122 34436 13128 34448
rect 16836 34436 16842 34448
rect 13122 34408 16842 34436
rect 13122 34396 13128 34408
rect 16836 34396 16842 34408
rect 16894 34396 16900 34448
rect 17590 34445 17618 34544
rect 17682 34504 17710 34612
rect 18219 34575 18277 34581
rect 18219 34541 18231 34575
rect 18265 34572 18277 34575
rect 18694 34572 18722 34739
rect 21160 34736 21166 34748
rect 21218 34736 21224 34788
rect 22816 34736 22822 34788
rect 22874 34776 22880 34788
rect 26039 34779 26097 34785
rect 26039 34776 26051 34779
rect 22874 34748 26051 34776
rect 22874 34736 22880 34748
rect 26039 34745 26051 34748
rect 26085 34745 26097 34779
rect 26039 34739 26097 34745
rect 26572 34779 26630 34785
rect 26572 34745 26584 34779
rect 26618 34776 26630 34779
rect 27327 34779 27385 34785
rect 27327 34776 27339 34779
rect 26618 34748 27339 34776
rect 26618 34745 26630 34748
rect 26572 34739 26630 34745
rect 27327 34745 27339 34748
rect 27373 34776 27385 34779
rect 30636 34776 30642 34788
rect 27373 34748 30642 34776
rect 27373 34745 27385 34748
rect 27327 34739 27385 34745
rect 30636 34736 30642 34748
rect 30694 34736 30700 34788
rect 33120 34736 33126 34788
rect 33178 34776 33184 34788
rect 33396 34776 33402 34788
rect 33178 34748 33402 34776
rect 33178 34736 33184 34748
rect 33396 34736 33402 34748
rect 33454 34776 33460 34788
rect 33951 34779 34009 34785
rect 33951 34776 33963 34779
rect 33454 34748 33963 34776
rect 33454 34736 33460 34748
rect 33951 34745 33963 34748
rect 33997 34776 34009 34779
rect 34592 34776 34598 34788
rect 33997 34748 34598 34776
rect 33997 34745 34009 34748
rect 33951 34739 34009 34745
rect 34592 34736 34598 34748
rect 34650 34736 34656 34788
rect 35512 34736 35518 34788
rect 35570 34776 35576 34788
rect 40112 34776 40118 34788
rect 35570 34748 40118 34776
rect 35570 34736 35576 34748
rect 40112 34736 40118 34748
rect 40170 34736 40176 34788
rect 40204 34736 40210 34788
rect 40262 34776 40268 34788
rect 55292 34776 55298 34788
rect 40262 34748 55298 34776
rect 40262 34736 40268 34748
rect 55292 34736 55298 34748
rect 55350 34736 55356 34788
rect 55384 34736 55390 34788
rect 55442 34776 55448 34788
rect 60996 34776 61002 34788
rect 55442 34748 61002 34776
rect 55442 34736 55448 34748
rect 60996 34736 61002 34748
rect 61054 34736 61060 34788
rect 63388 34736 63394 34788
rect 63446 34776 63452 34788
rect 63446 34748 69414 34776
rect 63446 34736 63452 34748
rect 26683 34711 26741 34717
rect 26683 34677 26695 34711
rect 26729 34677 26741 34711
rect 26683 34671 26741 34677
rect 29627 34711 29685 34717
rect 29627 34677 29639 34711
rect 29673 34708 29685 34711
rect 29808 34708 29814 34720
rect 29673 34680 29814 34708
rect 29673 34677 29685 34680
rect 29627 34671 29685 34677
rect 21252 34640 21258 34652
rect 21213 34612 21258 34640
rect 21252 34600 21258 34612
rect 21310 34600 21316 34652
rect 24659 34643 24717 34649
rect 24659 34609 24671 34643
rect 24705 34640 24717 34643
rect 25852 34640 25858 34652
rect 24705 34612 25346 34640
rect 24705 34609 24717 34612
rect 24659 34603 24717 34609
rect 20516 34572 20522 34584
rect 18265 34544 18722 34572
rect 20477 34544 20522 34572
rect 18265 34541 18277 34544
rect 18219 34535 18277 34541
rect 20516 34532 20522 34544
rect 20574 34532 20580 34584
rect 20608 34532 20614 34584
rect 20666 34572 20672 34584
rect 20795 34575 20853 34581
rect 20666 34544 20711 34572
rect 20666 34532 20672 34544
rect 20795 34541 20807 34575
rect 20841 34541 20853 34575
rect 20795 34535 20853 34541
rect 20335 34507 20393 34513
rect 20335 34504 20347 34507
rect 17682 34476 20347 34504
rect 20335 34473 20347 34476
rect 20381 34504 20393 34507
rect 20810 34504 20838 34535
rect 23276 34532 23282 34584
rect 23334 34572 23340 34584
rect 24843 34575 24901 34581
rect 24843 34572 24855 34575
rect 23334 34544 24855 34572
rect 23334 34532 23340 34544
rect 24843 34541 24855 34544
rect 24889 34541 24901 34575
rect 24843 34535 24901 34541
rect 25027 34575 25085 34581
rect 25027 34541 25039 34575
rect 25073 34541 25085 34575
rect 25027 34535 25085 34541
rect 24932 34504 24938 34516
rect 20381 34476 24938 34504
rect 20381 34473 20393 34476
rect 20335 34467 20393 34473
rect 24932 34464 24938 34476
rect 24990 34464 24996 34516
rect 17575 34439 17633 34445
rect 17575 34405 17587 34439
rect 17621 34436 17633 34439
rect 17664 34436 17670 34448
rect 17621 34408 17670 34436
rect 17621 34405 17633 34408
rect 17575 34399 17633 34405
rect 17664 34396 17670 34408
rect 17722 34396 17728 34448
rect 18400 34436 18406 34448
rect 18361 34408 18406 34436
rect 18400 34396 18406 34408
rect 18458 34396 18464 34448
rect 20608 34396 20614 34448
rect 20666 34436 20672 34448
rect 21439 34439 21497 34445
rect 21439 34436 21451 34439
rect 20666 34408 21451 34436
rect 20666 34396 20672 34408
rect 21439 34405 21451 34408
rect 21485 34436 21497 34439
rect 23000 34436 23006 34448
rect 21485 34408 23006 34436
rect 21485 34405 21497 34408
rect 21439 34399 21497 34405
rect 23000 34396 23006 34408
rect 23058 34396 23064 34448
rect 25042 34436 25070 34535
rect 25318 34504 25346 34612
rect 25410 34612 25858 34640
rect 25410 34581 25438 34612
rect 25852 34600 25858 34612
rect 25910 34600 25916 34652
rect 26220 34640 26226 34652
rect 26181 34612 26226 34640
rect 26220 34600 26226 34612
rect 26278 34640 26284 34652
rect 26698 34640 26726 34671
rect 29808 34668 29814 34680
rect 29866 34668 29872 34720
rect 29900 34668 29906 34720
rect 29958 34708 29964 34720
rect 39376 34708 39382 34720
rect 29958 34680 30003 34708
rect 35990 34680 39382 34708
rect 29958 34668 29964 34680
rect 26278 34612 26726 34640
rect 26775 34643 26833 34649
rect 26278 34600 26284 34612
rect 26775 34609 26787 34643
rect 26821 34609 26833 34643
rect 26775 34603 26833 34609
rect 25395 34575 25453 34581
rect 25395 34541 25407 34575
rect 25441 34541 25453 34575
rect 25395 34535 25453 34541
rect 25484 34532 25490 34584
rect 25542 34572 25548 34584
rect 26039 34575 26097 34581
rect 25542 34544 25587 34572
rect 25542 34532 25548 34544
rect 26039 34541 26051 34575
rect 26085 34572 26097 34575
rect 26790 34572 26818 34603
rect 26864 34600 26870 34652
rect 26922 34640 26928 34652
rect 35990 34640 36018 34680
rect 39376 34668 39382 34680
rect 39434 34668 39440 34720
rect 48119 34711 48177 34717
rect 48119 34677 48131 34711
rect 48165 34708 48177 34711
rect 48208 34708 48214 34720
rect 48165 34680 48214 34708
rect 48165 34677 48177 34680
rect 48119 34671 48177 34677
rect 48208 34668 48214 34680
rect 48266 34668 48272 34720
rect 51888 34708 51894 34720
rect 48778 34680 51894 34708
rect 40020 34640 40026 34652
rect 26922 34612 36018 34640
rect 39981 34612 40026 34640
rect 26922 34600 26928 34612
rect 40020 34600 40026 34612
rect 40078 34600 40084 34652
rect 41308 34600 41314 34652
rect 41366 34640 41372 34652
rect 47656 34640 47662 34652
rect 41366 34612 47242 34640
rect 47617 34612 47662 34640
rect 41366 34600 41372 34612
rect 26085 34544 26818 34572
rect 29719 34575 29777 34581
rect 26085 34541 26097 34544
rect 26039 34535 26097 34541
rect 29719 34541 29731 34575
rect 29765 34572 29777 34575
rect 29808 34572 29814 34584
rect 29765 34544 29814 34572
rect 29765 34541 29777 34544
rect 29719 34535 29777 34541
rect 29808 34532 29814 34544
rect 29866 34532 29872 34584
rect 34132 34572 34138 34584
rect 34093 34544 34138 34572
rect 34132 34532 34138 34544
rect 34190 34532 34196 34584
rect 34592 34532 34598 34584
rect 34650 34572 34656 34584
rect 34779 34575 34837 34581
rect 34779 34572 34791 34575
rect 34650 34544 34791 34572
rect 34650 34532 34656 34544
rect 34779 34541 34791 34544
rect 34825 34541 34837 34575
rect 35052 34572 35058 34584
rect 35013 34544 35058 34572
rect 34779 34535 34837 34541
rect 35052 34532 35058 34544
rect 35110 34532 35116 34584
rect 36435 34575 36493 34581
rect 36435 34541 36447 34575
rect 36481 34572 36493 34575
rect 38183 34575 38241 34581
rect 38183 34572 38195 34575
rect 36481 34544 38195 34572
rect 36481 34541 36493 34544
rect 36435 34535 36493 34541
rect 38183 34541 38195 34544
rect 38229 34541 38241 34575
rect 40112 34572 40118 34584
rect 40073 34544 40118 34572
rect 38183 34535 38241 34541
rect 26407 34507 26465 34513
rect 26407 34504 26419 34507
rect 25318 34476 26419 34504
rect 26407 34473 26419 34476
rect 26453 34473 26465 34507
rect 38198 34504 38226 34535
rect 40112 34532 40118 34544
rect 40170 34532 40176 34584
rect 40572 34572 40578 34584
rect 40533 34544 40578 34572
rect 40572 34532 40578 34544
rect 40630 34532 40636 34584
rect 40664 34532 40670 34584
rect 40722 34572 40728 34584
rect 40722 34544 40767 34572
rect 40722 34532 40728 34544
rect 46092 34532 46098 34584
rect 46150 34572 46156 34584
rect 46279 34575 46337 34581
rect 46279 34572 46291 34575
rect 46150 34544 46291 34572
rect 46150 34532 46156 34544
rect 46279 34541 46291 34544
rect 46325 34541 46337 34575
rect 46279 34535 46337 34541
rect 46555 34575 46613 34581
rect 46555 34541 46567 34575
rect 46601 34572 46613 34575
rect 46828 34572 46834 34584
rect 46601 34544 46834 34572
rect 46601 34541 46613 34544
rect 46555 34535 46613 34541
rect 46828 34532 46834 34544
rect 46886 34532 46892 34584
rect 40296 34504 40302 34516
rect 38198 34476 40302 34504
rect 26407 34467 26465 34473
rect 40296 34464 40302 34476
rect 40354 34464 40360 34516
rect 41219 34507 41277 34513
rect 41219 34473 41231 34507
rect 41265 34504 41277 34507
rect 44436 34504 44442 34516
rect 41265 34476 44442 34504
rect 41265 34473 41277 34476
rect 41219 34467 41277 34473
rect 44436 34464 44442 34476
rect 44494 34464 44500 34516
rect 25760 34436 25766 34448
rect 25042 34408 25766 34436
rect 25760 34396 25766 34408
rect 25818 34396 25824 34448
rect 25852 34396 25858 34448
rect 25910 34436 25916 34448
rect 25947 34439 26005 34445
rect 25947 34436 25959 34439
rect 25910 34408 25959 34436
rect 25910 34396 25916 34408
rect 25947 34405 25959 34408
rect 25993 34436 26005 34439
rect 26772 34436 26778 34448
rect 25993 34408 26778 34436
rect 25993 34405 26005 34408
rect 25947 34399 26005 34405
rect 26772 34396 26778 34408
rect 26830 34396 26836 34448
rect 27048 34436 27054 34448
rect 27009 34408 27054 34436
rect 27048 34396 27054 34408
rect 27106 34396 27112 34448
rect 31832 34396 31838 34448
rect 31890 34436 31896 34448
rect 32476 34436 32482 34448
rect 31890 34408 32482 34436
rect 31890 34396 31896 34408
rect 32476 34396 32482 34408
rect 32534 34396 32540 34448
rect 38180 34396 38186 34448
rect 38238 34436 38244 34448
rect 38275 34439 38333 34445
rect 38275 34436 38287 34439
rect 38238 34408 38287 34436
rect 38238 34396 38244 34408
rect 38275 34405 38287 34408
rect 38321 34436 38333 34439
rect 40204 34436 40210 34448
rect 38321 34408 40210 34436
rect 38321 34405 38333 34408
rect 38275 34399 38333 34405
rect 40204 34396 40210 34408
rect 40262 34396 40268 34448
rect 43516 34396 43522 34448
rect 43574 34436 43580 34448
rect 46920 34436 46926 34448
rect 43574 34408 46926 34436
rect 43574 34396 43580 34408
rect 46920 34396 46926 34408
rect 46978 34396 46984 34448
rect 47214 34436 47242 34612
rect 47656 34600 47662 34612
rect 47714 34600 47720 34652
rect 48778 34581 48806 34680
rect 51888 34668 51894 34680
rect 51946 34668 51952 34720
rect 51983 34711 52041 34717
rect 51983 34677 51995 34711
rect 52029 34708 52041 34711
rect 52808 34708 52814 34720
rect 52029 34680 52814 34708
rect 52029 34677 52041 34680
rect 51983 34671 52041 34677
rect 52808 34668 52814 34680
rect 52866 34668 52872 34720
rect 53176 34668 53182 34720
rect 53234 34708 53240 34720
rect 53234 34680 53498 34708
rect 53234 34668 53240 34680
rect 52075 34643 52133 34649
rect 51354 34612 52026 34640
rect 48763 34575 48821 34581
rect 48763 34541 48775 34575
rect 48809 34541 48821 34575
rect 48763 34535 48821 34541
rect 47564 34464 47570 34516
rect 47622 34504 47628 34516
rect 48855 34507 48913 34513
rect 48855 34504 48867 34507
rect 47622 34476 48867 34504
rect 47622 34464 47628 34476
rect 48855 34473 48867 34476
rect 48901 34473 48913 34507
rect 48855 34467 48913 34473
rect 51354 34436 51382 34612
rect 51854 34575 51912 34581
rect 51854 34572 51866 34575
rect 51538 34544 51866 34572
rect 51538 34448 51566 34544
rect 51854 34541 51866 34544
rect 51900 34541 51912 34575
rect 51998 34572 52026 34612
rect 52075 34609 52087 34643
rect 52121 34640 52133 34643
rect 53268 34640 53274 34652
rect 52121 34612 53274 34640
rect 52121 34609 52133 34612
rect 52075 34603 52133 34609
rect 53268 34600 53274 34612
rect 53326 34600 53332 34652
rect 53363 34643 53421 34649
rect 53363 34609 53375 34643
rect 53409 34609 53421 34643
rect 53363 34603 53421 34609
rect 53087 34575 53145 34581
rect 53087 34572 53099 34575
rect 51998 34544 53099 34572
rect 51854 34535 51912 34541
rect 53087 34541 53099 34544
rect 53133 34572 53145 34575
rect 53378 34572 53406 34603
rect 53470 34581 53498 34680
rect 54004 34668 54010 34720
rect 54062 34708 54068 34720
rect 54835 34711 54893 34717
rect 54835 34708 54847 34711
rect 54062 34680 54847 34708
rect 54062 34668 54068 34680
rect 54835 34677 54847 34680
rect 54881 34708 54893 34711
rect 64768 34708 64774 34720
rect 54881 34680 64774 34708
rect 54881 34677 54893 34680
rect 54835 34671 54893 34677
rect 64768 34668 64774 34680
rect 64826 34668 64832 34720
rect 67988 34708 67994 34720
rect 67949 34680 67994 34708
rect 67988 34668 67994 34680
rect 68046 34668 68052 34720
rect 69276 34708 69282 34720
rect 69237 34680 69282 34708
rect 69276 34668 69282 34680
rect 69334 34668 69340 34720
rect 69386 34708 69414 34748
rect 69460 34736 69466 34788
rect 69518 34776 69524 34788
rect 84272 34776 84278 34788
rect 69518 34748 84278 34776
rect 69518 34736 69524 34748
rect 84272 34736 84278 34748
rect 84330 34736 84336 34788
rect 88780 34736 88786 34788
rect 88838 34776 88844 34788
rect 90712 34776 90718 34788
rect 88838 34748 90718 34776
rect 88838 34736 88844 34748
rect 90712 34736 90718 34748
rect 90770 34776 90776 34788
rect 91175 34779 91233 34785
rect 91175 34776 91187 34779
rect 90770 34748 91187 34776
rect 90770 34736 90776 34748
rect 91175 34745 91187 34748
rect 91221 34745 91233 34779
rect 91175 34739 91233 34745
rect 74152 34708 74158 34720
rect 69386 34680 74158 34708
rect 74152 34668 74158 34680
rect 74210 34668 74216 34720
rect 80868 34708 80874 34720
rect 80150 34680 80874 34708
rect 57776 34600 57782 34652
rect 57834 34640 57840 34652
rect 58055 34643 58113 34649
rect 58055 34640 58067 34643
rect 57834 34612 58067 34640
rect 57834 34600 57840 34612
rect 58055 34609 58067 34612
rect 58101 34640 58113 34643
rect 59432 34640 59438 34652
rect 58101 34612 58466 34640
rect 59393 34612 59438 34640
rect 58101 34609 58113 34612
rect 58055 34603 58113 34609
rect 58438 34584 58466 34612
rect 59432 34600 59438 34612
rect 59490 34600 59496 34652
rect 59895 34643 59953 34649
rect 59895 34609 59907 34643
rect 59941 34640 59953 34643
rect 59984 34640 59990 34652
rect 59941 34612 59990 34640
rect 59941 34609 59953 34612
rect 59895 34603 59953 34609
rect 59984 34600 59990 34612
rect 60042 34600 60048 34652
rect 62100 34600 62106 34652
rect 62158 34640 62164 34652
rect 62379 34643 62437 34649
rect 62379 34640 62391 34643
rect 62158 34612 62391 34640
rect 62158 34600 62164 34612
rect 62379 34609 62391 34612
rect 62425 34640 62437 34643
rect 68006 34640 68034 34668
rect 62425 34612 62698 34640
rect 68006 34612 68494 34640
rect 62425 34609 62437 34612
rect 62379 34603 62437 34609
rect 53133 34544 53406 34572
rect 53455 34575 53513 34581
rect 53133 34541 53145 34544
rect 53087 34535 53145 34541
rect 53455 34541 53467 34575
rect 53501 34541 53513 34575
rect 54004 34572 54010 34584
rect 53965 34544 54010 34572
rect 53455 34535 53513 34541
rect 54004 34532 54010 34544
rect 54062 34532 54068 34584
rect 54191 34575 54249 34581
rect 54191 34541 54203 34575
rect 54237 34572 54249 34575
rect 54237 34544 55062 34572
rect 54237 34541 54249 34544
rect 54191 34535 54249 34541
rect 51707 34507 51765 34513
rect 51707 34473 51719 34507
rect 51753 34473 51765 34507
rect 51707 34467 51765 34473
rect 52443 34507 52501 34513
rect 52443 34473 52455 34507
rect 52489 34504 52501 34507
rect 54280 34504 54286 34516
rect 52489 34476 54286 34504
rect 52489 34473 52501 34476
rect 52443 34467 52501 34473
rect 51520 34436 51526 34448
rect 47214 34408 51382 34436
rect 51481 34408 51526 34436
rect 51520 34396 51526 34408
rect 51578 34396 51584 34448
rect 51722 34436 51750 34467
rect 54280 34464 54286 34476
rect 54338 34464 54344 34516
rect 54188 34436 54194 34448
rect 51722 34408 54194 34436
rect 54188 34396 54194 34408
rect 54246 34396 54252 34448
rect 54467 34439 54525 34445
rect 54467 34405 54479 34439
rect 54513 34436 54525 34439
rect 54648 34436 54654 34448
rect 54513 34408 54654 34436
rect 54513 34405 54525 34408
rect 54467 34399 54525 34405
rect 54648 34396 54654 34408
rect 54706 34396 54712 34448
rect 55034 34445 55062 34544
rect 57408 34532 57414 34584
rect 57466 34572 57472 34584
rect 58328 34572 58334 34584
rect 57466 34544 58334 34572
rect 57466 34532 57472 34544
rect 58328 34532 58334 34544
rect 58386 34532 58392 34584
rect 58420 34532 58426 34584
rect 58478 34572 58484 34584
rect 58880 34572 58886 34584
rect 58478 34544 58523 34572
rect 58841 34544 58886 34572
rect 58478 34532 58484 34544
rect 58880 34532 58886 34544
rect 58938 34532 58944 34584
rect 59067 34575 59125 34581
rect 59067 34541 59079 34575
rect 59113 34572 59125 34575
rect 59711 34575 59769 34581
rect 59711 34572 59723 34575
rect 59113 34544 59723 34572
rect 59113 34541 59125 34544
rect 59067 34535 59125 34541
rect 59711 34541 59723 34544
rect 59757 34572 59769 34575
rect 60168 34572 60174 34584
rect 59757 34544 60174 34572
rect 59757 34541 59769 34544
rect 59711 34535 59769 34541
rect 60168 34532 60174 34544
rect 60226 34532 60232 34584
rect 62560 34572 62566 34584
rect 62521 34544 62566 34572
rect 62560 34532 62566 34544
rect 62618 34532 62624 34584
rect 62670 34572 62698 34612
rect 63204 34581 63210 34584
rect 63023 34575 63081 34581
rect 63023 34572 63035 34575
rect 62670 34544 63035 34572
rect 63023 34541 63035 34544
rect 63069 34541 63081 34575
rect 63203 34572 63210 34581
rect 63165 34544 63210 34572
rect 63023 34535 63081 34541
rect 63203 34535 63210 34544
rect 63204 34532 63210 34535
rect 63262 34532 63268 34584
rect 67804 34572 67810 34584
rect 67765 34544 67810 34572
rect 67804 34532 67810 34544
rect 67862 34532 67868 34584
rect 68172 34572 68178 34584
rect 68133 34544 68178 34572
rect 68172 34532 68178 34544
rect 68230 34532 68236 34584
rect 68264 34532 68270 34584
rect 68322 34572 68328 34584
rect 68359 34575 68417 34581
rect 68359 34572 68371 34575
rect 68322 34544 68371 34572
rect 68322 34532 68328 34544
rect 68359 34541 68371 34544
rect 68405 34541 68417 34575
rect 68466 34572 68494 34612
rect 73968 34600 73974 34652
rect 74026 34640 74032 34652
rect 74247 34643 74305 34649
rect 74247 34640 74259 34643
rect 74026 34612 74259 34640
rect 74026 34600 74032 34612
rect 74247 34609 74259 34612
rect 74293 34609 74305 34643
rect 74520 34640 74526 34652
rect 74481 34612 74526 34640
rect 74247 34603 74305 34609
rect 68819 34575 68877 34581
rect 68819 34572 68831 34575
rect 68466 34544 68831 34572
rect 68359 34535 68417 34541
rect 68819 34541 68831 34544
rect 68865 34541 68877 34575
rect 68819 34535 68877 34541
rect 68908 34532 68914 34584
rect 68966 34572 68972 34584
rect 68966 34544 69011 34572
rect 68966 34532 68972 34544
rect 69644 34532 69650 34584
rect 69702 34572 69708 34584
rect 74262 34572 74290 34603
rect 74520 34600 74526 34612
rect 74578 34600 74584 34652
rect 80150 34649 80178 34680
rect 80868 34668 80874 34680
rect 80926 34668 80932 34720
rect 81144 34708 81150 34720
rect 81105 34680 81150 34708
rect 81144 34668 81150 34680
rect 81202 34668 81208 34720
rect 80135 34643 80193 34649
rect 80135 34609 80147 34643
rect 80181 34609 80193 34643
rect 80135 34603 80193 34609
rect 81328 34600 81334 34652
rect 81386 34640 81392 34652
rect 81386 34612 86158 34640
rect 81386 34600 81392 34612
rect 75995 34575 76053 34581
rect 75995 34572 76007 34575
rect 69702 34544 74198 34572
rect 74262 34544 76007 34572
rect 69702 34532 69708 34544
rect 74170 34504 74198 34544
rect 75995 34541 76007 34544
rect 76041 34541 76053 34575
rect 80224 34572 80230 34584
rect 80137 34544 80230 34572
rect 75995 34535 76053 34541
rect 80224 34532 80230 34544
rect 80282 34572 80288 34584
rect 80776 34572 80782 34584
rect 80282 34544 80782 34572
rect 80282 34532 80288 34544
rect 80776 34532 80782 34544
rect 80834 34532 80840 34584
rect 80963 34575 81021 34581
rect 80963 34541 80975 34575
rect 81009 34572 81021 34575
rect 81236 34572 81242 34584
rect 81009 34544 81242 34572
rect 81009 34541 81021 34544
rect 80963 34535 81021 34541
rect 81236 34532 81242 34544
rect 81294 34572 81300 34584
rect 82524 34572 82530 34584
rect 81294 34544 82530 34572
rect 81294 34532 81300 34544
rect 82524 34532 82530 34544
rect 82582 34532 82588 34584
rect 82711 34575 82769 34581
rect 82711 34541 82723 34575
rect 82757 34572 82769 34575
rect 82987 34575 83045 34581
rect 82987 34572 82999 34575
rect 82757 34544 82999 34572
rect 82757 34541 82769 34544
rect 82711 34535 82769 34541
rect 82987 34541 82999 34544
rect 83033 34572 83045 34575
rect 84640 34572 84646 34584
rect 83033 34544 84646 34572
rect 83033 34541 83045 34544
rect 82987 34535 83045 34541
rect 74336 34504 74342 34516
rect 62302 34476 71898 34504
rect 74170 34476 74342 34504
rect 55019 34439 55077 34445
rect 55019 34405 55031 34439
rect 55065 34436 55077 34439
rect 62302 34436 62330 34476
rect 55065 34408 62330 34436
rect 55065 34405 55077 34408
rect 55019 34399 55077 34405
rect 62560 34396 62566 34448
rect 62618 34436 62624 34448
rect 63204 34436 63210 34448
rect 62618 34408 63210 34436
rect 62618 34396 62624 34408
rect 63204 34396 63210 34408
rect 63262 34396 63268 34448
rect 63480 34396 63486 34448
rect 63538 34436 63544 34448
rect 63575 34439 63633 34445
rect 63575 34436 63587 34439
rect 63538 34408 63587 34436
rect 63538 34396 63544 34408
rect 63575 34405 63587 34408
rect 63621 34405 63633 34439
rect 63575 34399 63633 34405
rect 63664 34396 63670 34448
rect 63722 34436 63728 34448
rect 69460 34436 69466 34448
rect 63722 34408 69466 34436
rect 63722 34396 63728 34408
rect 69460 34396 69466 34408
rect 69518 34396 69524 34448
rect 69644 34436 69650 34448
rect 69605 34408 69650 34436
rect 69644 34396 69650 34408
rect 69702 34396 69708 34448
rect 71870 34436 71898 34476
rect 74336 34464 74342 34476
rect 74394 34464 74400 34516
rect 82726 34504 82754 34535
rect 84640 34532 84646 34544
rect 84698 34532 84704 34584
rect 86130 34581 86158 34612
rect 85931 34575 85989 34581
rect 85931 34541 85943 34575
rect 85977 34541 85989 34575
rect 85931 34535 85989 34541
rect 86115 34575 86173 34581
rect 86115 34541 86127 34575
rect 86161 34541 86173 34575
rect 86572 34572 86578 34584
rect 86533 34544 86578 34572
rect 86115 34535 86173 34541
rect 75182 34476 82754 34504
rect 75182 34436 75210 34476
rect 71870 34408 75210 34436
rect 75348 34396 75354 34448
rect 75406 34436 75412 34448
rect 75627 34439 75685 34445
rect 75627 34436 75639 34439
rect 75406 34408 75639 34436
rect 75406 34396 75412 34408
rect 75627 34405 75639 34408
rect 75673 34405 75685 34439
rect 75627 34399 75685 34405
rect 80776 34396 80782 34448
rect 80834 34436 80840 34448
rect 81328 34436 81334 34448
rect 80834 34408 81334 34436
rect 80834 34396 80840 34408
rect 81328 34396 81334 34408
rect 81386 34396 81392 34448
rect 82340 34396 82346 34448
rect 82398 34436 82404 34448
rect 82708 34436 82714 34448
rect 82398 34408 82714 34436
rect 82398 34396 82404 34408
rect 82708 34396 82714 34408
rect 82766 34436 82772 34448
rect 82803 34439 82861 34445
rect 82803 34436 82815 34439
rect 82766 34408 82815 34436
rect 82766 34396 82772 34408
rect 82803 34405 82815 34408
rect 82849 34405 82861 34439
rect 82803 34399 82861 34405
rect 85839 34439 85897 34445
rect 85839 34405 85851 34439
rect 85885 34436 85897 34439
rect 85946 34436 85974 34535
rect 86130 34504 86158 34535
rect 86572 34532 86578 34544
rect 86630 34532 86636 34584
rect 86667 34575 86725 34581
rect 86667 34541 86679 34575
rect 86713 34572 86725 34575
rect 87768 34572 87774 34584
rect 86713 34544 87774 34572
rect 86713 34541 86725 34544
rect 86667 34535 86725 34541
rect 86682 34504 86710 34535
rect 87768 34532 87774 34544
rect 87826 34532 87832 34584
rect 91080 34572 91086 34584
rect 91041 34544 91086 34572
rect 91080 34532 91086 34544
rect 91138 34532 91144 34584
rect 86130 34476 86710 34504
rect 87219 34507 87277 34513
rect 87219 34473 87231 34507
rect 87265 34504 87277 34507
rect 87952 34504 87958 34516
rect 87265 34476 87958 34504
rect 87265 34473 87277 34476
rect 87219 34467 87277 34473
rect 87952 34464 87958 34476
rect 88010 34464 88016 34516
rect 86020 34436 86026 34448
rect 85885 34408 86026 34436
rect 85885 34405 85897 34408
rect 85839 34399 85897 34405
rect 86020 34396 86026 34408
rect 86078 34396 86084 34448
rect 86572 34396 86578 34448
rect 86630 34436 86636 34448
rect 87403 34439 87461 34445
rect 87403 34436 87415 34439
rect 86630 34408 87415 34436
rect 86630 34396 86636 34408
rect 87403 34405 87415 34408
rect 87449 34405 87461 34439
rect 87403 34399 87461 34405
rect 538 34346 93642 34368
rect 538 34294 6344 34346
rect 6396 34294 6408 34346
rect 6460 34294 6472 34346
rect 6524 34294 6536 34346
rect 6588 34294 11672 34346
rect 11724 34294 11736 34346
rect 11788 34294 11800 34346
rect 11852 34294 11864 34346
rect 11916 34294 17000 34346
rect 17052 34294 17064 34346
rect 17116 34294 17128 34346
rect 17180 34294 17192 34346
rect 17244 34294 22328 34346
rect 22380 34294 22392 34346
rect 22444 34294 22456 34346
rect 22508 34294 22520 34346
rect 22572 34294 27656 34346
rect 27708 34294 27720 34346
rect 27772 34294 27784 34346
rect 27836 34294 27848 34346
rect 27900 34294 32984 34346
rect 33036 34294 33048 34346
rect 33100 34294 33112 34346
rect 33164 34294 33176 34346
rect 33228 34294 38312 34346
rect 38364 34294 38376 34346
rect 38428 34294 38440 34346
rect 38492 34294 38504 34346
rect 38556 34294 43640 34346
rect 43692 34294 43704 34346
rect 43756 34294 43768 34346
rect 43820 34294 43832 34346
rect 43884 34294 48968 34346
rect 49020 34294 49032 34346
rect 49084 34294 49096 34346
rect 49148 34294 49160 34346
rect 49212 34294 54296 34346
rect 54348 34294 54360 34346
rect 54412 34294 54424 34346
rect 54476 34294 54488 34346
rect 54540 34294 59624 34346
rect 59676 34294 59688 34346
rect 59740 34294 59752 34346
rect 59804 34294 59816 34346
rect 59868 34294 64952 34346
rect 65004 34294 65016 34346
rect 65068 34294 65080 34346
rect 65132 34294 65144 34346
rect 65196 34294 70280 34346
rect 70332 34294 70344 34346
rect 70396 34294 70408 34346
rect 70460 34294 70472 34346
rect 70524 34294 75608 34346
rect 75660 34294 75672 34346
rect 75724 34294 75736 34346
rect 75788 34294 75800 34346
rect 75852 34294 80936 34346
rect 80988 34294 81000 34346
rect 81052 34294 81064 34346
rect 81116 34294 81128 34346
rect 81180 34294 86264 34346
rect 86316 34294 86328 34346
rect 86380 34294 86392 34346
rect 86444 34294 86456 34346
rect 86508 34294 91592 34346
rect 91644 34294 91656 34346
rect 91708 34294 91720 34346
rect 91772 34294 91784 34346
rect 91836 34294 93642 34346
rect 538 34272 93642 34294
rect 10212 34232 10218 34244
rect 6642 34204 10218 34232
rect 6642 34176 6670 34204
rect 10212 34192 10218 34204
rect 10270 34192 10276 34244
rect 15732 34192 15738 34244
rect 15790 34232 15796 34244
rect 15919 34235 15977 34241
rect 15919 34232 15931 34235
rect 15790 34204 15931 34232
rect 15790 34192 15796 34204
rect 15919 34201 15931 34204
rect 15965 34201 15977 34235
rect 15919 34195 15977 34201
rect 6624 34124 6630 34176
rect 6682 34124 6688 34176
rect 6719 34167 6777 34173
rect 6719 34133 6731 34167
rect 6765 34164 6777 34167
rect 6765 34136 10166 34164
rect 6765 34133 6777 34136
rect 6719 34127 6777 34133
rect 3864 34056 3870 34108
rect 3922 34096 3928 34108
rect 5339 34099 5397 34105
rect 5339 34096 5351 34099
rect 3922 34068 5351 34096
rect 3922 34056 3928 34068
rect 5339 34065 5351 34068
rect 5385 34065 5397 34099
rect 5339 34059 5397 34065
rect 8927 34099 8985 34105
rect 8927 34065 8939 34099
rect 8973 34096 8985 34099
rect 9108 34096 9114 34108
rect 8973 34068 9114 34096
rect 8973 34065 8985 34068
rect 8927 34059 8985 34065
rect 9108 34056 9114 34068
rect 9166 34096 9172 34108
rect 10138 34105 10166 34136
rect 10230 34105 10258 34192
rect 9571 34099 9629 34105
rect 9571 34096 9583 34099
rect 9166 34068 9583 34096
rect 9166 34056 9172 34068
rect 9571 34065 9583 34068
rect 9617 34065 9629 34099
rect 9571 34059 9629 34065
rect 9755 34099 9813 34105
rect 9755 34065 9767 34099
rect 9801 34065 9813 34099
rect 9755 34059 9813 34065
rect 10123 34099 10181 34105
rect 10123 34065 10135 34099
rect 10169 34065 10181 34099
rect 10123 34059 10181 34065
rect 10215 34099 10273 34105
rect 10215 34065 10227 34099
rect 10261 34065 10273 34099
rect 15934 34096 15962 34195
rect 16008 34192 16014 34244
rect 16066 34232 16072 34244
rect 17299 34235 17357 34241
rect 17299 34232 17311 34235
rect 16066 34204 17311 34232
rect 16066 34192 16072 34204
rect 17299 34201 17311 34204
rect 17345 34201 17357 34235
rect 17299 34195 17357 34201
rect 17572 34192 17578 34244
rect 17630 34232 17636 34244
rect 17667 34235 17725 34241
rect 17667 34232 17679 34235
rect 17630 34204 17679 34232
rect 17630 34192 17636 34204
rect 17667 34201 17679 34204
rect 17713 34232 17725 34235
rect 26864 34232 26870 34244
rect 17713 34204 26870 34232
rect 17713 34201 17725 34204
rect 17667 34195 17725 34201
rect 26864 34192 26870 34204
rect 26922 34192 26928 34244
rect 27048 34192 27054 34244
rect 27106 34232 27112 34244
rect 51520 34232 51526 34244
rect 27106 34204 51526 34232
rect 27106 34192 27112 34204
rect 51520 34192 51526 34204
rect 51578 34192 51584 34244
rect 52808 34232 52814 34244
rect 52769 34204 52814 34232
rect 52808 34192 52814 34204
rect 52866 34192 52872 34244
rect 54188 34192 54194 34244
rect 54246 34232 54252 34244
rect 60444 34232 60450 34244
rect 54246 34204 60450 34232
rect 54246 34192 54252 34204
rect 60444 34192 60450 34204
rect 60502 34192 60508 34244
rect 60996 34192 61002 34244
rect 61054 34232 61060 34244
rect 63756 34232 63762 34244
rect 61054 34204 63762 34232
rect 61054 34192 61060 34204
rect 63756 34192 63762 34204
rect 63814 34192 63820 34244
rect 64768 34192 64774 34244
rect 64826 34232 64832 34244
rect 64826 34204 80638 34232
rect 64826 34192 64832 34204
rect 17756 34164 17762 34176
rect 16854 34136 17762 34164
rect 16008 34096 16014 34108
rect 15921 34068 16014 34096
rect 10215 34059 10273 34065
rect 4692 33988 4698 34040
rect 4750 34028 4756 34040
rect 5063 34031 5121 34037
rect 5063 34028 5075 34031
rect 4750 34000 5075 34028
rect 4750 33988 4756 34000
rect 5063 33997 5075 34000
rect 5109 34028 5121 34031
rect 5109 34000 6946 34028
rect 5109 33997 5121 34000
rect 5063 33991 5121 33997
rect 6918 33969 6946 34000
rect 6903 33963 6961 33969
rect 6903 33929 6915 33963
rect 6949 33960 6961 33963
rect 7084 33960 7090 33972
rect 6949 33932 7090 33960
rect 6949 33929 6961 33932
rect 6903 33923 6961 33929
rect 7084 33920 7090 33932
rect 7142 33920 7148 33972
rect 9770 33960 9798 34059
rect 16008 34056 16014 34068
rect 16066 34096 16072 34108
rect 16854 34105 16882 34136
rect 17756 34124 17762 34136
rect 17814 34164 17820 34176
rect 18400 34164 18406 34176
rect 17814 34136 18406 34164
rect 17814 34124 17820 34136
rect 18400 34124 18406 34136
rect 18458 34124 18464 34176
rect 23000 34124 23006 34176
rect 23058 34164 23064 34176
rect 36987 34167 37045 34173
rect 36987 34164 36999 34167
rect 23058 34136 36999 34164
rect 23058 34124 23064 34136
rect 36987 34133 36999 34136
rect 37033 34133 37045 34167
rect 40112 34164 40118 34176
rect 36987 34127 37045 34133
rect 39808 34136 40118 34164
rect 16103 34099 16161 34105
rect 16103 34096 16115 34099
rect 16066 34068 16115 34096
rect 16066 34056 16072 34068
rect 16103 34065 16115 34068
rect 16149 34065 16161 34099
rect 16103 34059 16161 34065
rect 16287 34099 16345 34105
rect 16287 34065 16299 34099
rect 16333 34096 16345 34099
rect 16839 34099 16897 34105
rect 16333 34068 16514 34096
rect 16333 34065 16345 34068
rect 16287 34059 16345 34065
rect 10396 33960 10402 33972
rect 9770 33932 10402 33960
rect 10396 33920 10402 33932
rect 10454 33920 10460 33972
rect 16486 33960 16514 34068
rect 16839 34065 16851 34099
rect 16885 34065 16897 34099
rect 16839 34059 16897 34065
rect 17023 34099 17081 34105
rect 17023 34065 17035 34099
rect 17069 34096 17081 34099
rect 17572 34096 17578 34108
rect 17069 34068 17578 34096
rect 17069 34065 17081 34068
rect 17023 34059 17081 34065
rect 17572 34056 17578 34068
rect 17630 34056 17636 34108
rect 20148 34056 20154 34108
rect 20206 34096 20212 34108
rect 22267 34099 22325 34105
rect 20206 34068 22218 34096
rect 20206 34056 20212 34068
rect 17480 33988 17486 34040
rect 17538 34028 17544 34040
rect 21807 34031 21865 34037
rect 21807 34028 21819 34031
rect 17538 34000 21819 34028
rect 17538 33988 17544 34000
rect 21807 33997 21819 34000
rect 21853 34028 21865 34031
rect 21991 34031 22049 34037
rect 21991 34028 22003 34031
rect 21853 34000 22003 34028
rect 21853 33997 21865 34000
rect 21807 33991 21865 33997
rect 21991 33997 22003 34000
rect 22037 33997 22049 34031
rect 22190 34028 22218 34068
rect 22267 34065 22279 34099
rect 22313 34096 22325 34099
rect 22724 34096 22730 34108
rect 22313 34068 22730 34096
rect 22313 34065 22325 34068
rect 22267 34059 22325 34065
rect 22724 34056 22730 34068
rect 22782 34056 22788 34108
rect 23368 34056 23374 34108
rect 23426 34096 23432 34108
rect 23647 34099 23705 34105
rect 23647 34096 23659 34099
rect 23426 34068 23659 34096
rect 23426 34056 23432 34068
rect 23647 34065 23659 34068
rect 23693 34096 23705 34099
rect 25484 34096 25490 34108
rect 23693 34068 25490 34096
rect 23693 34065 23705 34068
rect 23647 34059 23705 34065
rect 25484 34056 25490 34068
rect 25542 34056 25548 34108
rect 25944 34096 25950 34108
rect 25905 34068 25950 34096
rect 25944 34056 25950 34068
rect 26002 34056 26008 34108
rect 28888 34096 28894 34108
rect 28849 34068 28894 34096
rect 28888 34056 28894 34068
rect 28946 34056 28952 34108
rect 29808 34056 29814 34108
rect 29866 34096 29872 34108
rect 31651 34099 31709 34105
rect 31651 34096 31663 34099
rect 29866 34068 31663 34096
rect 29866 34056 29872 34068
rect 31651 34065 31663 34068
rect 31697 34096 31709 34099
rect 32019 34099 32077 34105
rect 32019 34096 32031 34099
rect 31697 34068 32031 34096
rect 31697 34065 31709 34068
rect 31651 34059 31709 34065
rect 32019 34065 32031 34068
rect 32065 34065 32077 34099
rect 32019 34059 32077 34065
rect 32476 34056 32482 34108
rect 32534 34096 32540 34108
rect 33307 34099 33365 34105
rect 33307 34096 33319 34099
rect 32534 34068 33319 34096
rect 32534 34056 32540 34068
rect 33307 34065 33319 34068
rect 33353 34065 33365 34099
rect 33307 34059 33365 34065
rect 33491 34099 33549 34105
rect 33491 34065 33503 34099
rect 33537 34065 33549 34099
rect 34040 34096 34046 34108
rect 34001 34068 34046 34096
rect 33491 34059 33549 34065
rect 26315 34031 26373 34037
rect 26315 34028 26327 34031
rect 22190 34000 26327 34028
rect 21991 33991 22049 33997
rect 26315 33997 26327 34000
rect 26361 33997 26373 34031
rect 26315 33991 26373 33997
rect 26683 34031 26741 34037
rect 26683 33997 26695 34031
rect 26729 34028 26741 34031
rect 26729 34000 33258 34028
rect 26729 33997 26741 34000
rect 26683 33991 26741 33997
rect 17851 33963 17909 33969
rect 17851 33960 17863 33963
rect 16486 33932 17863 33960
rect 17851 33929 17863 33932
rect 17897 33960 17909 33963
rect 21712 33960 21718 33972
rect 17897 33932 21718 33960
rect 17897 33929 17909 33932
rect 17851 33923 17909 33929
rect 21712 33920 21718 33932
rect 21770 33920 21776 33972
rect 24932 33920 24938 33972
rect 24990 33960 24996 33972
rect 25671 33963 25729 33969
rect 25671 33960 25683 33963
rect 24990 33932 25683 33960
rect 24990 33920 24996 33932
rect 25671 33929 25683 33932
rect 25717 33929 25729 33963
rect 25671 33923 25729 33929
rect 26112 33963 26170 33969
rect 26112 33929 26124 33963
rect 26158 33960 26170 33963
rect 26864 33960 26870 33972
rect 26158 33932 26870 33960
rect 26158 33929 26170 33932
rect 26112 33923 26170 33929
rect 9384 33892 9390 33904
rect 9345 33864 9390 33892
rect 9384 33852 9390 33864
rect 9442 33852 9448 33904
rect 17664 33852 17670 33904
rect 17722 33892 17728 33904
rect 25392 33892 25398 33904
rect 17722 33864 25398 33892
rect 17722 33852 17728 33864
rect 25392 33852 25398 33864
rect 25450 33852 25456 33904
rect 25686 33892 25714 33923
rect 26864 33920 26870 33932
rect 26922 33920 26928 33972
rect 29072 33960 29078 33972
rect 29033 33932 29078 33960
rect 29072 33920 29078 33932
rect 29130 33920 29136 33972
rect 26220 33892 26226 33904
rect 25686 33864 26226 33892
rect 26220 33852 26226 33864
rect 26278 33852 26284 33904
rect 31464 33852 31470 33904
rect 31522 33892 31528 33904
rect 31835 33895 31893 33901
rect 31835 33892 31847 33895
rect 31522 33864 31847 33892
rect 31522 33852 31528 33864
rect 31835 33861 31847 33864
rect 31881 33861 31893 33895
rect 33230 33892 33258 34000
rect 33506 33960 33534 34059
rect 34040 34056 34046 34068
rect 34098 34056 34104 34108
rect 34227 34099 34285 34105
rect 34227 34065 34239 34099
rect 34273 34096 34285 34099
rect 34871 34099 34929 34105
rect 34871 34096 34883 34099
rect 34273 34068 34883 34096
rect 34273 34065 34285 34068
rect 34227 34059 34285 34065
rect 34871 34065 34883 34068
rect 34917 34096 34929 34099
rect 35512 34096 35518 34108
rect 34917 34068 35518 34096
rect 34917 34065 34929 34068
rect 34871 34059 34929 34065
rect 35512 34056 35518 34068
rect 35570 34056 35576 34108
rect 39808 34105 39836 34136
rect 40112 34124 40118 34136
rect 40170 34124 40176 34176
rect 40664 34164 40670 34176
rect 40406 34136 40670 34164
rect 40406 34108 40434 34136
rect 40664 34124 40670 34136
rect 40722 34124 40728 34176
rect 45080 34164 45086 34176
rect 45041 34136 45086 34164
rect 45080 34124 45086 34136
rect 45138 34124 45144 34176
rect 46644 34124 46650 34176
rect 46702 34164 46708 34176
rect 46739 34167 46797 34173
rect 46739 34164 46751 34167
rect 46702 34136 46751 34164
rect 46702 34124 46708 34136
rect 46739 34133 46751 34136
rect 46785 34133 46797 34167
rect 47656 34164 47662 34176
rect 46739 34127 46797 34133
rect 46938 34136 47662 34164
rect 39793 34099 39851 34105
rect 39793 34065 39805 34099
rect 39839 34065 39851 34099
rect 39928 34096 39934 34108
rect 39889 34068 39934 34096
rect 39793 34059 39851 34065
rect 39928 34056 39934 34068
rect 39986 34056 39992 34108
rect 40296 34096 40302 34108
rect 40257 34068 40302 34096
rect 40296 34056 40302 34068
rect 40354 34056 40360 34108
rect 40388 34056 40394 34108
rect 40446 34096 40452 34108
rect 44991 34099 45049 34105
rect 40446 34068 40491 34096
rect 40866 34068 41078 34096
rect 40446 34056 40452 34068
rect 33948 33960 33954 33972
rect 33506 33932 33954 33960
rect 33948 33920 33954 33932
rect 34006 33920 34012 33972
rect 34408 33960 34414 33972
rect 34369 33932 34414 33960
rect 34408 33920 34414 33932
rect 34466 33920 34472 33972
rect 40866 33960 40894 34068
rect 40943 34031 41001 34037
rect 40943 33997 40955 34031
rect 40989 33997 41001 34031
rect 41050 34028 41078 34068
rect 44991 34065 45003 34099
rect 45037 34096 45049 34099
rect 45172 34096 45178 34108
rect 45037 34068 45178 34096
rect 45037 34065 45049 34068
rect 44991 34059 45049 34065
rect 45172 34056 45178 34068
rect 45230 34056 45236 34108
rect 46552 34056 46558 34108
rect 46610 34096 46616 34108
rect 46938 34105 46966 34136
rect 47656 34124 47662 34136
rect 47714 34124 47720 34176
rect 54375 34167 54433 34173
rect 51630 34136 52578 34164
rect 46923 34099 46981 34105
rect 46923 34096 46935 34099
rect 46610 34068 46935 34096
rect 46610 34056 46616 34068
rect 46923 34065 46935 34068
rect 46969 34065 46981 34099
rect 46923 34059 46981 34065
rect 47012 34056 47018 34108
rect 47070 34096 47076 34108
rect 51630 34105 51658 34136
rect 51247 34099 51305 34105
rect 51247 34096 51259 34099
rect 47070 34068 51259 34096
rect 47070 34056 47076 34068
rect 51247 34065 51259 34068
rect 51293 34096 51305 34099
rect 51431 34099 51489 34105
rect 51431 34096 51443 34099
rect 51293 34068 51443 34096
rect 51293 34065 51305 34068
rect 51247 34059 51305 34065
rect 51431 34065 51443 34068
rect 51477 34096 51489 34099
rect 51615 34099 51673 34105
rect 51615 34096 51627 34099
rect 51477 34068 51627 34096
rect 51477 34065 51489 34068
rect 51431 34059 51489 34065
rect 51615 34065 51627 34068
rect 51661 34065 51673 34099
rect 51615 34059 51673 34065
rect 51799 34099 51857 34105
rect 51799 34065 51811 34099
rect 51845 34096 51857 34099
rect 52351 34099 52409 34105
rect 52351 34096 52363 34099
rect 51845 34068 52363 34096
rect 51845 34065 51857 34068
rect 51799 34059 51857 34065
rect 52351 34065 52363 34068
rect 52397 34096 52409 34099
rect 52440 34096 52446 34108
rect 52397 34068 52446 34096
rect 52397 34065 52409 34068
rect 52351 34059 52409 34065
rect 52440 34056 52446 34068
rect 52498 34056 52504 34108
rect 52550 34105 52578 34136
rect 54375 34133 54387 34167
rect 54421 34164 54433 34167
rect 60355 34167 60413 34173
rect 60355 34164 60367 34167
rect 54421 34136 60367 34164
rect 54421 34133 54433 34136
rect 54375 34127 54433 34133
rect 60355 34133 60367 34136
rect 60401 34133 60413 34167
rect 63572 34164 63578 34176
rect 63533 34136 63578 34164
rect 60355 34127 60413 34133
rect 63572 34124 63578 34136
rect 63630 34124 63636 34176
rect 64124 34124 64130 34176
rect 64182 34164 64188 34176
rect 67531 34167 67589 34173
rect 67531 34164 67543 34167
rect 64182 34136 67543 34164
rect 64182 34124 64188 34136
rect 67531 34133 67543 34136
rect 67577 34133 67589 34167
rect 68264 34164 68270 34176
rect 67531 34127 67589 34133
rect 68098 34136 68270 34164
rect 52535 34099 52593 34105
rect 52535 34065 52547 34099
rect 52581 34065 52593 34099
rect 52535 34059 52593 34065
rect 52808 34056 52814 34108
rect 52866 34096 52872 34108
rect 55111 34099 55169 34105
rect 52866 34068 54878 34096
rect 52866 34056 52872 34068
rect 54191 34031 54249 34037
rect 54191 34028 54203 34031
rect 41050 34000 52026 34028
rect 40943 33991 41001 33997
rect 34518 33932 40894 33960
rect 40958 33960 40986 33991
rect 51998 33960 52026 34000
rect 52734 34000 54203 34028
rect 52734 33960 52762 34000
rect 54191 33997 54203 34000
rect 54237 34028 54249 34031
rect 54522 34031 54580 34037
rect 54522 34028 54534 34031
rect 54237 34000 54534 34028
rect 54237 33997 54249 34000
rect 54191 33991 54249 33997
rect 54522 33997 54534 34000
rect 54568 33997 54580 34031
rect 54522 33991 54580 33997
rect 54648 33988 54654 34040
rect 54706 34028 54712 34040
rect 54743 34031 54801 34037
rect 54743 34028 54755 34031
rect 54706 34000 54755 34028
rect 54706 33988 54712 34000
rect 54743 33997 54755 34000
rect 54789 33997 54801 34031
rect 54850 34028 54878 34068
rect 55111 34065 55123 34099
rect 55157 34096 55169 34099
rect 55384 34096 55390 34108
rect 55157 34068 55390 34096
rect 55157 34065 55169 34068
rect 55111 34059 55169 34065
rect 55384 34056 55390 34068
rect 55442 34056 55448 34108
rect 59619 34099 59677 34105
rect 59619 34065 59631 34099
rect 59665 34096 59677 34099
rect 60539 34099 60597 34105
rect 60539 34096 60551 34099
rect 59665 34068 60551 34096
rect 59665 34065 59677 34068
rect 59619 34059 59677 34065
rect 60539 34065 60551 34068
rect 60585 34096 60597 34099
rect 63664 34096 63670 34108
rect 60585 34068 63670 34096
rect 60585 34065 60597 34068
rect 60539 34059 60597 34065
rect 63664 34056 63670 34068
rect 63722 34056 63728 34108
rect 63848 34105 63854 34108
rect 63805 34099 63854 34105
rect 63805 34065 63817 34099
rect 63851 34065 63854 34099
rect 63805 34059 63854 34065
rect 63848 34056 63854 34059
rect 63906 34056 63912 34108
rect 59800 34028 59806 34040
rect 54850 34000 59806 34028
rect 54743 33991 54801 33997
rect 59800 33988 59806 34000
rect 59858 33988 59864 34040
rect 59987 34031 60045 34037
rect 59987 33997 59999 34031
rect 60033 33997 60045 34031
rect 63943 34031 64001 34037
rect 63943 34028 63955 34031
rect 59987 33991 60045 33997
rect 63774 34000 63955 34028
rect 40958 33932 51934 33960
rect 51998 33932 52762 33960
rect 34518 33892 34546 33932
rect 35052 33892 35058 33904
rect 33230 33864 34546 33892
rect 35013 33864 35058 33892
rect 31835 33855 31893 33861
rect 35052 33852 35058 33864
rect 35110 33852 35116 33904
rect 36987 33895 37045 33901
rect 36987 33861 36999 33895
rect 37033 33892 37045 33895
rect 43332 33892 43338 33904
rect 37033 33864 43338 33892
rect 37033 33861 37045 33864
rect 36987 33855 37045 33861
rect 43332 33852 43338 33864
rect 43390 33892 43396 33904
rect 43516 33892 43522 33904
rect 43390 33864 43522 33892
rect 43390 33852 43396 33864
rect 43516 33852 43522 33864
rect 43574 33852 43580 33904
rect 47015 33895 47073 33901
rect 47015 33861 47027 33895
rect 47061 33892 47073 33895
rect 47196 33892 47202 33904
rect 47061 33864 47202 33892
rect 47061 33861 47073 33864
rect 47015 33855 47073 33861
rect 47196 33852 47202 33864
rect 47254 33852 47260 33904
rect 51906 33892 51934 33932
rect 59432 33920 59438 33972
rect 59490 33960 59496 33972
rect 59895 33963 59953 33969
rect 59895 33960 59907 33963
rect 59490 33932 59907 33960
rect 59490 33920 59496 33932
rect 59895 33929 59907 33932
rect 59941 33929 59953 33963
rect 59895 33923 59953 33929
rect 60002 33904 60030 33991
rect 60076 33920 60082 33972
rect 60134 33960 60140 33972
rect 63391 33963 63449 33969
rect 63391 33960 63403 33963
rect 60134 33932 63403 33960
rect 60134 33920 60140 33932
rect 63391 33929 63403 33932
rect 63437 33960 63449 33963
rect 63774 33960 63802 34000
rect 63943 33997 63955 34000
rect 63989 33997 64001 34031
rect 63943 33991 64001 33997
rect 64311 34031 64369 34037
rect 64311 33997 64323 34031
rect 64357 34028 64369 34031
rect 65596 34028 65602 34040
rect 64357 34000 65602 34028
rect 64357 33997 64369 34000
rect 64311 33991 64369 33997
rect 65596 33988 65602 34000
rect 65654 33988 65660 34040
rect 67546 34028 67574 34127
rect 67620 34056 67626 34108
rect 67678 34096 67684 34108
rect 68098 34105 68126 34136
rect 68264 34124 68270 34136
rect 68322 34164 68328 34176
rect 69371 34167 69429 34173
rect 69371 34164 69383 34167
rect 68322 34136 69383 34164
rect 68322 34124 68328 34136
rect 69371 34133 69383 34136
rect 69417 34164 69429 34167
rect 69644 34164 69650 34176
rect 69417 34136 69650 34164
rect 69417 34133 69429 34136
rect 69371 34127 69429 34133
rect 69644 34124 69650 34136
rect 69702 34124 69708 34176
rect 73692 34124 73698 34176
rect 73750 34164 73756 34176
rect 74983 34167 75041 34173
rect 74983 34164 74995 34167
rect 73750 34136 74995 34164
rect 73750 34124 73756 34136
rect 74983 34133 74995 34136
rect 75029 34133 75041 34167
rect 79948 34164 79954 34176
rect 74983 34127 75041 34133
rect 78678 34136 79954 34164
rect 67899 34099 67957 34105
rect 67899 34096 67911 34099
rect 67678 34068 67911 34096
rect 67678 34056 67684 34068
rect 67899 34065 67911 34068
rect 67945 34065 67957 34099
rect 67899 34059 67957 34065
rect 68083 34099 68141 34105
rect 68083 34065 68095 34099
rect 68129 34065 68141 34099
rect 68543 34099 68601 34105
rect 68543 34096 68555 34099
rect 68083 34059 68141 34065
rect 68190 34068 68555 34096
rect 68190 34028 68218 34068
rect 68543 34065 68555 34068
rect 68589 34065 68601 34099
rect 68543 34059 68601 34065
rect 68632 34056 68638 34108
rect 68690 34096 68696 34108
rect 73603 34099 73661 34105
rect 68690 34068 68735 34096
rect 68690 34056 68696 34068
rect 73603 34065 73615 34099
rect 73649 34096 73661 34099
rect 73876 34096 73882 34108
rect 73649 34068 73882 34096
rect 73649 34065 73661 34068
rect 73603 34059 73661 34065
rect 73876 34056 73882 34068
rect 73934 34056 73940 34108
rect 74891 34099 74949 34105
rect 74891 34065 74903 34099
rect 74937 34096 74949 34099
rect 75440 34096 75446 34108
rect 74937 34068 75446 34096
rect 74937 34065 74949 34068
rect 74891 34059 74949 34065
rect 75440 34056 75446 34068
rect 75498 34096 75504 34108
rect 76084 34096 76090 34108
rect 75498 34068 76090 34096
rect 75498 34056 75504 34068
rect 76084 34056 76090 34068
rect 76142 34056 76148 34108
rect 77924 34096 77930 34108
rect 77885 34068 77930 34096
rect 77924 34056 77930 34068
rect 77982 34056 77988 34108
rect 78111 34099 78169 34105
rect 78111 34065 78123 34099
rect 78157 34096 78169 34099
rect 78568 34096 78574 34108
rect 78157 34068 78574 34096
rect 78157 34065 78169 34068
rect 78111 34059 78169 34065
rect 78568 34056 78574 34068
rect 78626 34056 78632 34108
rect 78678 34105 78706 34136
rect 79948 34124 79954 34136
rect 80006 34124 80012 34176
rect 78663 34099 78721 34105
rect 78663 34065 78675 34099
rect 78709 34065 78721 34099
rect 78663 34059 78721 34065
rect 78847 34099 78905 34105
rect 78847 34065 78859 34099
rect 78893 34096 78905 34099
rect 80408 34096 80414 34108
rect 78893 34068 80414 34096
rect 78893 34065 78905 34068
rect 78847 34059 78905 34065
rect 80408 34056 80414 34068
rect 80466 34056 80472 34108
rect 67546 34000 68218 34028
rect 73511 34031 73569 34037
rect 73511 33997 73523 34031
rect 73557 34028 73569 34031
rect 73692 34028 73698 34040
rect 73557 34000 73698 34028
rect 73557 33997 73569 34000
rect 73511 33991 73569 33997
rect 73692 33988 73698 34000
rect 73750 33988 73756 34040
rect 74060 34028 74066 34040
rect 74021 34000 74066 34028
rect 74060 33988 74066 34000
rect 74118 33988 74124 34040
rect 80610 34028 80638 34204
rect 80684 34192 80690 34244
rect 80742 34232 80748 34244
rect 81055 34235 81113 34241
rect 81055 34232 81067 34235
rect 80742 34204 81067 34232
rect 80742 34192 80748 34204
rect 80794 34105 80822 34204
rect 81055 34201 81067 34204
rect 81101 34201 81113 34235
rect 81055 34195 81113 34201
rect 80871 34167 80929 34173
rect 80871 34133 80883 34167
rect 80917 34164 80929 34167
rect 81236 34164 81242 34176
rect 80917 34136 81242 34164
rect 80917 34133 80929 34136
rect 80871 34127 80929 34133
rect 81236 34124 81242 34136
rect 81294 34124 81300 34176
rect 90252 34124 90258 34176
rect 90310 34164 90316 34176
rect 90310 34136 91218 34164
rect 90310 34124 90316 34136
rect 80779 34099 80837 34105
rect 80779 34065 80791 34099
rect 80825 34065 80837 34099
rect 80779 34059 80837 34065
rect 89792 34056 89798 34108
rect 89850 34096 89856 34108
rect 91190 34105 91218 34136
rect 90439 34099 90497 34105
rect 90439 34096 90451 34099
rect 89850 34068 90451 34096
rect 89850 34056 89856 34068
rect 90439 34065 90451 34068
rect 90485 34096 90497 34099
rect 90991 34099 91049 34105
rect 90991 34096 91003 34099
rect 90485 34068 91003 34096
rect 90485 34065 90497 34068
rect 90439 34059 90497 34065
rect 90991 34065 91003 34068
rect 91037 34065 91049 34099
rect 90991 34059 91049 34065
rect 91175 34099 91233 34105
rect 91175 34065 91187 34099
rect 91221 34065 91233 34099
rect 91175 34059 91233 34065
rect 88412 34028 88418 34040
rect 80610 34000 88418 34028
rect 88412 33988 88418 34000
rect 88470 33988 88476 34040
rect 90252 34028 90258 34040
rect 90213 34000 90258 34028
rect 90252 33988 90258 34000
rect 90310 33988 90316 34040
rect 63437 33932 63802 33960
rect 63437 33929 63449 33932
rect 63391 33923 63449 33929
rect 64124 33920 64130 33972
rect 64182 33960 64188 33972
rect 66056 33960 66062 33972
rect 64182 33932 66062 33960
rect 64182 33920 64188 33932
rect 66056 33920 66062 33932
rect 66114 33920 66120 33972
rect 67807 33963 67865 33969
rect 67807 33929 67819 33963
rect 67853 33960 67865 33963
rect 67896 33960 67902 33972
rect 67853 33932 67902 33960
rect 67853 33929 67865 33932
rect 67807 33923 67865 33929
rect 67896 33920 67902 33932
rect 67954 33960 67960 33972
rect 68632 33960 68638 33972
rect 67954 33932 68638 33960
rect 67954 33920 67960 33932
rect 68632 33920 68638 33932
rect 68690 33920 68696 33972
rect 68724 33920 68730 33972
rect 68782 33960 68788 33972
rect 69003 33963 69061 33969
rect 69003 33960 69015 33963
rect 68782 33932 69015 33960
rect 68782 33920 68788 33932
rect 69003 33929 69015 33932
rect 69049 33929 69061 33963
rect 79031 33963 79089 33969
rect 79031 33960 79043 33963
rect 69003 33923 69061 33929
rect 69938 33932 79043 33960
rect 52808 33892 52814 33904
rect 51906 33864 52814 33892
rect 52808 33852 52814 33864
rect 52866 33852 52872 33904
rect 52900 33852 52906 33904
rect 52958 33892 52964 33904
rect 53179 33895 53237 33901
rect 53179 33892 53191 33895
rect 52958 33864 53191 33892
rect 52958 33852 52964 33864
rect 53179 33861 53191 33864
rect 53225 33892 53237 33895
rect 53363 33895 53421 33901
rect 53363 33892 53375 33895
rect 53225 33864 53375 33892
rect 53225 33861 53237 33864
rect 53179 33855 53237 33861
rect 53363 33861 53375 33864
rect 53409 33892 53421 33895
rect 53452 33892 53458 33904
rect 53409 33864 53458 33892
rect 53409 33861 53421 33864
rect 53363 33855 53421 33861
rect 53452 33852 53458 33864
rect 53510 33852 53516 33904
rect 54648 33892 54654 33904
rect 54609 33864 54654 33892
rect 54648 33852 54654 33864
rect 54706 33852 54712 33904
rect 59524 33852 59530 33904
rect 59582 33892 59588 33904
rect 59757 33895 59815 33901
rect 59757 33892 59769 33895
rect 59582 33864 59769 33892
rect 59582 33852 59588 33864
rect 59757 33861 59769 33864
rect 59803 33861 59815 33895
rect 59757 33855 59815 33861
rect 59984 33852 59990 33904
rect 60042 33852 60048 33904
rect 63740 33895 63798 33901
rect 63740 33861 63752 33895
rect 63786 33892 63798 33895
rect 64495 33895 64553 33901
rect 64495 33892 64507 33895
rect 63786 33864 64507 33892
rect 63786 33861 63798 33864
rect 63740 33855 63798 33861
rect 64495 33861 64507 33864
rect 64541 33892 64553 33895
rect 69938 33892 69966 33932
rect 79031 33929 79043 33932
rect 79077 33929 79089 33963
rect 91356 33960 91362 33972
rect 91317 33932 91362 33960
rect 79031 33923 79089 33929
rect 91356 33920 91362 33932
rect 91414 33920 91420 33972
rect 64541 33864 69966 33892
rect 64541 33861 64553 33864
rect 64495 33855 64553 33861
rect 73876 33852 73882 33904
rect 73934 33892 73940 33904
rect 74155 33895 74213 33901
rect 74155 33892 74167 33895
rect 73934 33864 74167 33892
rect 73934 33852 73940 33864
rect 74155 33861 74167 33864
rect 74201 33861 74213 33895
rect 74155 33855 74213 33861
rect 74336 33852 74342 33904
rect 74394 33892 74400 33904
rect 78936 33892 78942 33904
rect 74394 33864 78942 33892
rect 74394 33852 74400 33864
rect 78936 33852 78942 33864
rect 78994 33852 79000 33904
rect 538 33802 93642 33824
rect 538 33750 3680 33802
rect 3732 33750 3744 33802
rect 3796 33750 3808 33802
rect 3860 33750 3872 33802
rect 3924 33750 9008 33802
rect 9060 33750 9072 33802
rect 9124 33750 9136 33802
rect 9188 33750 9200 33802
rect 9252 33750 14336 33802
rect 14388 33750 14400 33802
rect 14452 33750 14464 33802
rect 14516 33750 14528 33802
rect 14580 33750 19664 33802
rect 19716 33750 19728 33802
rect 19780 33750 19792 33802
rect 19844 33750 19856 33802
rect 19908 33750 24992 33802
rect 25044 33750 25056 33802
rect 25108 33750 25120 33802
rect 25172 33750 25184 33802
rect 25236 33750 30320 33802
rect 30372 33750 30384 33802
rect 30436 33750 30448 33802
rect 30500 33750 30512 33802
rect 30564 33750 35648 33802
rect 35700 33750 35712 33802
rect 35764 33750 35776 33802
rect 35828 33750 35840 33802
rect 35892 33750 40976 33802
rect 41028 33750 41040 33802
rect 41092 33750 41104 33802
rect 41156 33750 41168 33802
rect 41220 33750 46304 33802
rect 46356 33750 46368 33802
rect 46420 33750 46432 33802
rect 46484 33750 46496 33802
rect 46548 33750 51632 33802
rect 51684 33750 51696 33802
rect 51748 33750 51760 33802
rect 51812 33750 51824 33802
rect 51876 33750 56960 33802
rect 57012 33750 57024 33802
rect 57076 33750 57088 33802
rect 57140 33750 57152 33802
rect 57204 33750 62288 33802
rect 62340 33750 62352 33802
rect 62404 33750 62416 33802
rect 62468 33750 62480 33802
rect 62532 33750 67616 33802
rect 67668 33750 67680 33802
rect 67732 33750 67744 33802
rect 67796 33750 67808 33802
rect 67860 33750 72944 33802
rect 72996 33750 73008 33802
rect 73060 33750 73072 33802
rect 73124 33750 73136 33802
rect 73188 33750 78272 33802
rect 78324 33750 78336 33802
rect 78388 33750 78400 33802
rect 78452 33750 78464 33802
rect 78516 33750 83600 33802
rect 83652 33750 83664 33802
rect 83716 33750 83728 33802
rect 83780 33750 83792 33802
rect 83844 33750 88928 33802
rect 88980 33750 88992 33802
rect 89044 33750 89056 33802
rect 89108 33750 89120 33802
rect 89172 33750 93642 33802
rect 538 33728 93642 33750
rect 2576 33648 2582 33700
rect 2634 33688 2640 33700
rect 2763 33691 2821 33697
rect 2763 33688 2775 33691
rect 2634 33660 2775 33688
rect 2634 33648 2640 33660
rect 2763 33657 2775 33660
rect 2809 33657 2821 33691
rect 17572 33688 17578 33700
rect 17533 33660 17578 33688
rect 2763 33651 2821 33657
rect 17572 33648 17578 33660
rect 17630 33648 17636 33700
rect 23276 33688 23282 33700
rect 23237 33660 23282 33688
rect 23276 33648 23282 33660
rect 23334 33648 23340 33700
rect 25392 33648 25398 33700
rect 25450 33688 25456 33700
rect 28336 33688 28342 33700
rect 25450 33660 28342 33688
rect 25450 33648 25456 33660
rect 28336 33648 28342 33660
rect 28394 33648 28400 33700
rect 29351 33691 29409 33697
rect 29351 33657 29363 33691
rect 29397 33688 29409 33691
rect 29716 33688 29722 33700
rect 29397 33660 29722 33688
rect 29397 33657 29409 33660
rect 29351 33651 29409 33657
rect 29716 33648 29722 33660
rect 29774 33648 29780 33700
rect 30176 33648 30182 33700
rect 30234 33688 30240 33700
rect 39284 33688 39290 33700
rect 30234 33660 39290 33688
rect 30234 33648 30240 33660
rect 39284 33648 39290 33660
rect 39342 33648 39348 33700
rect 39652 33648 39658 33700
rect 39710 33688 39716 33700
rect 40664 33688 40670 33700
rect 39710 33660 40670 33688
rect 39710 33648 39716 33660
rect 40664 33648 40670 33660
rect 40722 33648 40728 33700
rect 46000 33648 46006 33700
rect 46058 33688 46064 33700
rect 49312 33688 49318 33700
rect 46058 33660 49318 33688
rect 46058 33648 46064 33660
rect 49312 33648 49318 33660
rect 49370 33648 49376 33700
rect 53915 33691 53973 33697
rect 52366 33660 53866 33688
rect 13064 33620 13070 33632
rect 12622 33592 13070 33620
rect 2119 33555 2177 33561
rect 2119 33521 2131 33555
rect 2165 33552 2177 33555
rect 9019 33555 9077 33561
rect 2165 33524 3082 33552
rect 2165 33521 2177 33524
rect 2119 33515 2177 33521
rect 3054 33493 3082 33524
rect 9019 33521 9031 33555
rect 9065 33552 9077 33555
rect 9384 33552 9390 33564
rect 9065 33524 9390 33552
rect 9065 33521 9077 33524
rect 9019 33515 9077 33521
rect 9384 33512 9390 33524
rect 9442 33512 9448 33564
rect 12622 33561 12650 33592
rect 13064 33580 13070 33592
rect 13122 33620 13128 33632
rect 13159 33623 13217 33629
rect 13159 33620 13171 33623
rect 13122 33592 13171 33620
rect 13122 33580 13128 33592
rect 13159 33589 13171 33592
rect 13205 33589 13217 33623
rect 26775 33623 26833 33629
rect 13159 33583 13217 33589
rect 24582 33592 26634 33620
rect 12607 33555 12665 33561
rect 12607 33521 12619 33555
rect 12653 33521 12665 33555
rect 12975 33555 13033 33561
rect 12975 33552 12987 33555
rect 12607 33515 12665 33521
rect 12714 33524 12987 33552
rect 3039 33487 3097 33493
rect 3039 33453 3051 33487
rect 3085 33484 3097 33487
rect 3496 33484 3502 33496
rect 3085 33456 3502 33484
rect 3085 33453 3097 33456
rect 3039 33447 3097 33453
rect 3496 33444 3502 33456
rect 3554 33444 3560 33496
rect 4603 33487 4661 33493
rect 4603 33453 4615 33487
rect 4649 33453 4661 33487
rect 4603 33447 4661 33453
rect 4787 33487 4845 33493
rect 4787 33453 4799 33487
rect 4833 33453 4845 33487
rect 5152 33484 5158 33496
rect 5113 33456 5158 33484
rect 4787 33447 4845 33453
rect 3220 33376 3226 33428
rect 3278 33416 3284 33428
rect 3959 33419 4017 33425
rect 3959 33416 3971 33419
rect 3278 33388 3971 33416
rect 3278 33376 3284 33388
rect 3959 33385 3971 33388
rect 4005 33416 4017 33419
rect 4618 33416 4646 33447
rect 4005 33388 4646 33416
rect 4802 33416 4830 33447
rect 5152 33444 5158 33456
rect 5210 33444 5216 33496
rect 5339 33487 5397 33493
rect 5339 33453 5351 33487
rect 5385 33484 5397 33487
rect 6624 33484 6630 33496
rect 5385 33456 6630 33484
rect 5385 33453 5397 33456
rect 5339 33447 5397 33453
rect 6624 33444 6630 33456
rect 6682 33444 6688 33496
rect 7084 33444 7090 33496
rect 7142 33484 7148 33496
rect 8743 33487 8801 33493
rect 8743 33484 8755 33487
rect 7142 33456 8755 33484
rect 7142 33444 7148 33456
rect 8743 33453 8755 33456
rect 8789 33484 8801 33487
rect 10028 33484 10034 33496
rect 8789 33456 10034 33484
rect 8789 33453 8801 33456
rect 8743 33447 8801 33453
rect 10028 33444 10034 33456
rect 10086 33484 10092 33496
rect 10491 33487 10549 33493
rect 10491 33484 10503 33487
rect 10086 33456 10503 33484
rect 10086 33444 10092 33456
rect 10491 33453 10503 33456
rect 10537 33453 10549 33487
rect 12512 33484 12518 33496
rect 12473 33456 12518 33484
rect 10491 33447 10549 33453
rect 12512 33444 12518 33456
rect 12570 33444 12576 33496
rect 6164 33416 6170 33428
rect 4802 33388 6170 33416
rect 4005 33385 4017 33388
rect 3959 33379 4017 33385
rect 6164 33376 6170 33388
rect 6222 33376 6228 33428
rect 10396 33416 10402 33428
rect 10357 33388 10402 33416
rect 10396 33376 10402 33388
rect 10454 33376 10460 33428
rect 11871 33419 11929 33425
rect 11871 33385 11883 33419
rect 11917 33416 11929 33419
rect 12420 33416 12426 33428
rect 11917 33388 12426 33416
rect 11917 33385 11929 33388
rect 11871 33379 11929 33385
rect 12420 33376 12426 33388
rect 12478 33376 12484 33428
rect 4419 33351 4477 33357
rect 4419 33317 4431 33351
rect 4465 33348 4477 33351
rect 4968 33348 4974 33360
rect 4465 33320 4974 33348
rect 4465 33317 4477 33320
rect 4419 33311 4477 33317
rect 4968 33308 4974 33320
rect 5026 33308 5032 33360
rect 11500 33308 11506 33360
rect 11558 33348 11564 33360
rect 12714 33348 12742 33524
rect 12975 33521 12987 33524
rect 13021 33521 13033 33555
rect 12975 33515 13033 33521
rect 24107 33555 24165 33561
rect 24107 33521 24119 33555
rect 24153 33552 24165 33555
rect 24288 33552 24294 33564
rect 24153 33524 24294 33552
rect 24153 33521 24165 33524
rect 24107 33515 24165 33521
rect 24288 33512 24294 33524
rect 24346 33512 24352 33564
rect 12883 33487 12941 33493
rect 12883 33453 12895 33487
rect 12929 33453 12941 33487
rect 12883 33447 12941 33453
rect 13803 33487 13861 33493
rect 13803 33453 13815 33487
rect 13849 33484 13861 33487
rect 13892 33484 13898 33496
rect 13849 33456 13898 33484
rect 13849 33453 13861 33456
rect 13803 33447 13861 33453
rect 12898 33416 12926 33447
rect 13892 33444 13898 33456
rect 13950 33444 13956 33496
rect 17296 33444 17302 33496
rect 17354 33484 17360 33496
rect 17483 33487 17541 33493
rect 17483 33484 17495 33487
rect 17354 33456 17495 33484
rect 17354 33444 17360 33456
rect 17483 33453 17495 33456
rect 17529 33453 17541 33487
rect 18768 33484 18774 33496
rect 18729 33456 18774 33484
rect 17483 33447 17541 33453
rect 18768 33444 18774 33456
rect 18826 33444 18832 33496
rect 20792 33444 20798 33496
rect 20850 33484 20856 33496
rect 20979 33487 21037 33493
rect 20979 33484 20991 33487
rect 20850 33456 20991 33484
rect 20850 33444 20856 33456
rect 20979 33453 20991 33456
rect 21025 33453 21037 33487
rect 20979 33447 21037 33453
rect 23187 33487 23245 33493
rect 23187 33453 23199 33487
rect 23233 33484 23245 33487
rect 23368 33484 23374 33496
rect 23233 33456 23374 33484
rect 23233 33453 23245 33456
rect 23187 33447 23245 33453
rect 23368 33444 23374 33456
rect 23426 33444 23432 33496
rect 24012 33444 24018 33496
rect 24070 33484 24076 33496
rect 24383 33487 24441 33493
rect 24383 33484 24395 33487
rect 24070 33456 24395 33484
rect 24070 33444 24076 33456
rect 24383 33453 24395 33456
rect 24429 33484 24441 33487
rect 24582 33484 24610 33592
rect 24935 33487 24993 33493
rect 24935 33484 24947 33487
rect 24429 33456 24947 33484
rect 24429 33453 24441 33456
rect 24383 33447 24441 33453
rect 24935 33453 24947 33456
rect 24981 33453 24993 33487
rect 24935 33447 24993 33453
rect 25119 33487 25177 33493
rect 25119 33453 25131 33487
rect 25165 33484 25177 33487
rect 26128 33484 26134 33496
rect 25165 33456 26134 33484
rect 25165 33453 25177 33456
rect 25119 33447 25177 33453
rect 26128 33444 26134 33456
rect 26186 33444 26192 33496
rect 26606 33493 26634 33592
rect 26775 33589 26787 33623
rect 26821 33620 26833 33623
rect 26821 33592 41998 33620
rect 26821 33589 26833 33592
rect 26775 33583 26833 33589
rect 30360 33552 30366 33564
rect 30321 33524 30366 33552
rect 30360 33512 30366 33524
rect 30418 33512 30424 33564
rect 33948 33512 33954 33564
rect 34006 33552 34012 33564
rect 35052 33552 35058 33564
rect 34006 33524 35058 33552
rect 34006 33512 34012 33524
rect 35052 33512 35058 33524
rect 35110 33512 35116 33564
rect 35236 33512 35242 33564
rect 35294 33552 35300 33564
rect 41970 33552 41998 33592
rect 44436 33580 44442 33632
rect 44494 33620 44500 33632
rect 52366 33620 52394 33660
rect 53636 33620 53642 33632
rect 44494 33592 52394 33620
rect 52458 33592 53642 33620
rect 44494 33580 44500 33592
rect 52458 33552 52486 33592
rect 53636 33580 53642 33592
rect 53694 33580 53700 33632
rect 35294 33524 40158 33552
rect 41970 33524 52486 33552
rect 35294 33512 35300 33524
rect 26591 33487 26649 33493
rect 26591 33453 26603 33487
rect 26637 33453 26649 33487
rect 26591 33447 26649 33453
rect 28888 33444 28894 33496
rect 28946 33484 28952 33496
rect 29167 33487 29225 33493
rect 29167 33484 29179 33487
rect 28946 33456 29179 33484
rect 28946 33444 28952 33456
rect 29167 33453 29179 33456
rect 29213 33453 29225 33487
rect 29167 33447 29225 33453
rect 30176 33444 30182 33496
rect 30234 33484 30240 33496
rect 30271 33487 30329 33493
rect 30271 33484 30283 33487
rect 30234 33456 30283 33484
rect 30234 33444 30240 33456
rect 30271 33453 30283 33456
rect 30317 33453 30329 33487
rect 31464 33484 31470 33496
rect 31425 33456 31470 33484
rect 30271 33447 30329 33453
rect 31464 33444 31470 33456
rect 31522 33444 31528 33496
rect 31559 33487 31617 33493
rect 31559 33453 31571 33487
rect 31605 33484 31617 33487
rect 31832 33484 31838 33496
rect 31605 33456 31838 33484
rect 31605 33453 31617 33456
rect 31559 33447 31617 33453
rect 31832 33444 31838 33456
rect 31890 33444 31896 33496
rect 32019 33487 32077 33493
rect 32019 33453 32031 33487
rect 32065 33484 32077 33487
rect 32108 33484 32114 33496
rect 32065 33456 32114 33484
rect 32065 33453 32077 33456
rect 32019 33447 32077 33453
rect 32108 33444 32114 33456
rect 32166 33444 32172 33496
rect 32203 33487 32261 33493
rect 32203 33453 32215 33487
rect 32249 33484 32261 33487
rect 32568 33484 32574 33496
rect 32249 33456 32574 33484
rect 32249 33453 32261 33456
rect 32203 33447 32261 33453
rect 32568 33444 32574 33456
rect 32626 33444 32632 33496
rect 35420 33484 35426 33496
rect 35381 33456 35426 33484
rect 35420 33444 35426 33456
rect 35478 33444 35484 33496
rect 35512 33444 35518 33496
rect 35570 33484 35576 33496
rect 40130 33493 40158 33524
rect 52532 33512 52538 33564
rect 52590 33552 52596 33564
rect 53838 33552 53866 33660
rect 53915 33657 53927 33691
rect 53961 33688 53973 33691
rect 54648 33688 54654 33700
rect 53961 33660 54654 33688
rect 53961 33657 53973 33660
rect 53915 33651 53973 33657
rect 54648 33648 54654 33660
rect 54706 33648 54712 33700
rect 57503 33691 57561 33697
rect 57503 33657 57515 33691
rect 57549 33688 57561 33691
rect 58880 33688 58886 33700
rect 57549 33660 58886 33688
rect 57549 33657 57561 33660
rect 57503 33651 57561 33657
rect 58880 33648 58886 33660
rect 58938 33648 58944 33700
rect 58975 33691 59033 33697
rect 58975 33657 58987 33691
rect 59021 33688 59033 33691
rect 59984 33688 59990 33700
rect 59021 33660 59990 33688
rect 59021 33657 59033 33660
rect 58975 33651 59033 33657
rect 59984 33648 59990 33660
rect 60042 33648 60048 33700
rect 60076 33648 60082 33700
rect 60134 33697 60140 33700
rect 60134 33691 60183 33697
rect 60134 33657 60137 33691
rect 60171 33688 60183 33691
rect 60171 33660 60227 33688
rect 60171 33657 60183 33660
rect 60134 33651 60183 33657
rect 60134 33648 60140 33651
rect 60260 33648 60266 33700
rect 60318 33688 60324 33700
rect 60444 33688 60450 33700
rect 60318 33660 60363 33688
rect 60405 33660 60450 33688
rect 60318 33648 60324 33660
rect 60444 33648 60450 33660
rect 60502 33648 60508 33700
rect 63480 33688 63486 33700
rect 63441 33660 63486 33688
rect 63480 33648 63486 33660
rect 63538 33648 63544 33700
rect 64124 33688 64130 33700
rect 63682 33660 64130 33688
rect 54004 33580 54010 33632
rect 54062 33620 54068 33632
rect 62652 33620 62658 33632
rect 54062 33592 62658 33620
rect 54062 33580 54068 33592
rect 62652 33580 62658 33592
rect 62710 33580 62716 33632
rect 63372 33623 63430 33629
rect 63372 33589 63384 33623
rect 63418 33620 63430 33623
rect 63682 33620 63710 33660
rect 64124 33648 64130 33660
rect 64182 33648 64188 33700
rect 65761 33660 65918 33688
rect 63418 33592 63710 33620
rect 63418 33589 63430 33592
rect 63372 33583 63430 33589
rect 63756 33580 63762 33632
rect 63814 33620 63820 33632
rect 65761 33620 65789 33660
rect 65890 33629 65918 33660
rect 65964 33648 65970 33700
rect 66022 33688 66028 33700
rect 66022 33660 70150 33688
rect 66022 33648 66028 33660
rect 63814 33592 65789 33620
rect 65875 33623 65933 33629
rect 63814 33580 63820 33592
rect 65875 33589 65887 33623
rect 65921 33589 65933 33623
rect 65875 33583 65933 33589
rect 66056 33580 66062 33632
rect 66114 33620 66120 33632
rect 70122 33620 70150 33660
rect 73600 33648 73606 33700
rect 73658 33688 73664 33700
rect 75075 33691 75133 33697
rect 75075 33688 75087 33691
rect 73658 33660 75087 33688
rect 73658 33648 73664 33660
rect 75075 33657 75087 33660
rect 75121 33657 75133 33691
rect 75075 33651 75133 33657
rect 81512 33648 81518 33700
rect 81570 33688 81576 33700
rect 85284 33688 85290 33700
rect 81570 33660 85290 33688
rect 81570 33648 81576 33660
rect 85284 33648 85290 33660
rect 85342 33648 85348 33700
rect 85652 33688 85658 33700
rect 85613 33660 85658 33688
rect 85652 33648 85658 33660
rect 85710 33688 85716 33700
rect 85839 33691 85897 33697
rect 85839 33688 85851 33691
rect 85710 33660 85851 33688
rect 85710 33648 85716 33660
rect 85839 33657 85851 33660
rect 85885 33688 85897 33691
rect 85885 33660 86434 33688
rect 85885 33657 85897 33660
rect 85839 33651 85897 33657
rect 81696 33620 81702 33632
rect 66114 33592 69690 33620
rect 70122 33592 81702 33620
rect 66114 33580 66120 33592
rect 57503 33555 57561 33561
rect 57503 33552 57515 33555
rect 52590 33524 52946 33552
rect 53838 33524 57515 33552
rect 52590 33512 52596 33524
rect 52918 33496 52946 33524
rect 57503 33521 57515 33524
rect 57549 33521 57561 33555
rect 59251 33555 59309 33561
rect 59251 33552 59263 33555
rect 57503 33515 57561 33521
rect 59082 33524 59263 33552
rect 40115 33487 40173 33493
rect 35570 33456 35615 33484
rect 35714 33456 40066 33484
rect 35570 33444 35576 33456
rect 13987 33419 14045 33425
rect 13987 33416 13999 33419
rect 12898 33388 13999 33416
rect 13987 33385 13999 33388
rect 14033 33385 14045 33419
rect 13987 33379 14045 33385
rect 18676 33376 18682 33428
rect 18734 33416 18740 33428
rect 18863 33419 18921 33425
rect 18863 33416 18875 33419
rect 18734 33388 18875 33416
rect 18734 33376 18740 33388
rect 18863 33385 18875 33388
rect 18909 33416 18921 33419
rect 35714 33416 35742 33456
rect 39652 33416 39658 33428
rect 18909 33388 35742 33416
rect 35806 33388 39658 33416
rect 18909 33385 18921 33388
rect 18863 33379 18921 33385
rect 20792 33348 20798 33360
rect 11558 33320 12742 33348
rect 20753 33320 20798 33348
rect 11558 33308 11564 33320
rect 20792 33308 20798 33320
rect 20850 33308 20856 33360
rect 21163 33351 21221 33357
rect 21163 33317 21175 33351
rect 21209 33348 21221 33351
rect 21620 33348 21626 33360
rect 21209 33320 21626 33348
rect 21209 33317 21221 33320
rect 21163 33311 21221 33317
rect 21620 33308 21626 33320
rect 21678 33308 21684 33360
rect 25395 33351 25453 33357
rect 25395 33317 25407 33351
rect 25441 33348 25453 33351
rect 25484 33348 25490 33360
rect 25441 33320 25490 33348
rect 25441 33317 25453 33320
rect 25395 33311 25453 33317
rect 25484 33308 25490 33320
rect 25542 33308 25548 33360
rect 31832 33308 31838 33360
rect 31890 33348 31896 33360
rect 32479 33351 32537 33357
rect 32479 33348 32491 33351
rect 31890 33320 32491 33348
rect 31890 33308 31896 33320
rect 32479 33317 32491 33320
rect 32525 33317 32537 33351
rect 32479 33311 32537 33317
rect 32568 33308 32574 33360
rect 32626 33348 32632 33360
rect 32847 33351 32905 33357
rect 32847 33348 32859 33351
rect 32626 33320 32859 33348
rect 32626 33308 32632 33320
rect 32847 33317 32859 33320
rect 32893 33348 32905 33351
rect 35806 33348 35834 33388
rect 39652 33376 39658 33388
rect 39710 33376 39716 33428
rect 39928 33416 39934 33428
rect 39889 33388 39934 33416
rect 39928 33376 39934 33388
rect 39986 33376 39992 33428
rect 40038 33416 40066 33456
rect 40115 33453 40127 33487
rect 40161 33484 40173 33487
rect 40572 33484 40578 33496
rect 40161 33456 40578 33484
rect 40161 33453 40173 33456
rect 40115 33447 40173 33453
rect 40572 33444 40578 33456
rect 40630 33444 40636 33496
rect 40664 33444 40670 33496
rect 40722 33484 40728 33496
rect 43516 33484 43522 33496
rect 40722 33456 43522 33484
rect 40722 33444 40728 33456
rect 43516 33444 43522 33456
rect 43574 33444 43580 33496
rect 43976 33444 43982 33496
rect 44034 33484 44040 33496
rect 44071 33487 44129 33493
rect 44071 33484 44083 33487
rect 44034 33456 44083 33484
rect 44034 33444 44040 33456
rect 44071 33453 44083 33456
rect 44117 33453 44129 33487
rect 44071 33447 44129 33453
rect 45650 33456 47058 33484
rect 45650 33416 45678 33456
rect 46920 33416 46926 33428
rect 40038 33388 45678 33416
rect 46881 33388 46926 33416
rect 46920 33376 46926 33388
rect 46978 33376 46984 33428
rect 47030 33416 47058 33456
rect 47104 33444 47110 33496
rect 47162 33484 47168 33496
rect 48852 33484 48858 33496
rect 47162 33456 48858 33484
rect 47162 33444 47168 33456
rect 48852 33444 48858 33456
rect 48910 33444 48916 33496
rect 51155 33487 51213 33493
rect 51155 33453 51167 33487
rect 51201 33484 51213 33487
rect 52256 33484 52262 33496
rect 51201 33456 52262 33484
rect 51201 33453 51213 33456
rect 51155 33447 51213 33453
rect 52256 33444 52262 33456
rect 52314 33444 52320 33496
rect 52719 33487 52777 33493
rect 52719 33484 52731 33487
rect 52550 33456 52731 33484
rect 47472 33416 47478 33428
rect 47030 33388 47334 33416
rect 47433 33388 47478 33416
rect 32893 33320 35834 33348
rect 32893 33317 32905 33320
rect 32847 33311 32905 33317
rect 39560 33308 39566 33360
rect 39618 33348 39624 33360
rect 40207 33351 40265 33357
rect 40207 33348 40219 33351
rect 39618 33320 40219 33348
rect 39618 33308 39624 33320
rect 40207 33317 40219 33320
rect 40253 33317 40265 33351
rect 43976 33348 43982 33360
rect 43937 33320 43982 33348
rect 40207 33311 40265 33317
rect 43976 33308 43982 33320
rect 44034 33308 44040 33360
rect 44163 33351 44221 33357
rect 44163 33317 44175 33351
rect 44209 33348 44221 33351
rect 44712 33348 44718 33360
rect 44209 33320 44718 33348
rect 44209 33317 44221 33320
rect 44163 33311 44221 33317
rect 44712 33308 44718 33320
rect 44770 33308 44776 33360
rect 46644 33308 46650 33360
rect 46702 33348 46708 33360
rect 47012 33348 47018 33360
rect 46702 33320 47018 33348
rect 46702 33308 46708 33320
rect 47012 33308 47018 33320
rect 47070 33308 47076 33360
rect 47306 33348 47334 33388
rect 47472 33376 47478 33388
rect 47530 33376 47536 33428
rect 49680 33376 49686 33428
rect 49738 33416 49744 33428
rect 51247 33419 51305 33425
rect 51247 33416 51259 33419
rect 49738 33388 51259 33416
rect 49738 33376 49744 33388
rect 51247 33385 51259 33388
rect 51293 33385 51305 33419
rect 51247 33379 51305 33385
rect 52550 33416 52578 33456
rect 52719 33453 52731 33456
rect 52765 33453 52777 33487
rect 52900 33484 52906 33496
rect 52861 33456 52906 33484
rect 52719 33447 52777 33453
rect 52900 33444 52906 33456
rect 52958 33444 52964 33496
rect 53363 33487 53421 33493
rect 53363 33453 53375 33487
rect 53409 33453 53421 33487
rect 53363 33447 53421 33453
rect 53378 33416 53406 33447
rect 53452 33444 53458 33496
rect 53510 33484 53516 33496
rect 54283 33487 54341 33493
rect 54283 33484 54295 33487
rect 53510 33456 54295 33484
rect 53510 33444 53516 33456
rect 54283 33453 54295 33456
rect 54329 33484 54341 33487
rect 54467 33487 54525 33493
rect 54467 33484 54479 33487
rect 54329 33456 54479 33484
rect 54329 33453 54341 33456
rect 54283 33447 54341 33453
rect 54467 33453 54479 33456
rect 54513 33484 54525 33487
rect 57868 33484 57874 33496
rect 54513 33456 57874 33484
rect 54513 33453 54525 33456
rect 54467 33447 54525 33453
rect 57868 33444 57874 33456
rect 57926 33444 57932 33496
rect 57963 33487 58021 33493
rect 57963 33453 57975 33487
rect 58009 33453 58021 33487
rect 57963 33447 58021 33453
rect 58055 33487 58113 33493
rect 58055 33453 58067 33487
rect 58101 33453 58113 33487
rect 58420 33484 58426 33496
rect 58381 33456 58426 33484
rect 58055 33447 58113 33453
rect 52550 33388 53406 33416
rect 52550 33357 52578 33388
rect 57978 33360 58006 33447
rect 58070 33416 58098 33447
rect 58420 33444 58426 33456
rect 58478 33444 58484 33496
rect 58512 33444 58518 33496
rect 58570 33484 58576 33496
rect 58570 33456 58615 33484
rect 58570 33444 58576 33456
rect 59082 33416 59110 33524
rect 59251 33521 59263 33524
rect 59297 33552 59309 33555
rect 62836 33552 62842 33564
rect 59297 33524 62842 33552
rect 59297 33521 59309 33524
rect 59251 33515 59309 33521
rect 62836 33512 62842 33524
rect 62894 33512 62900 33564
rect 63575 33555 63633 33561
rect 63575 33521 63587 33555
rect 63621 33521 63633 33555
rect 65964 33552 65970 33564
rect 65925 33524 65970 33552
rect 63575 33515 63633 33521
rect 59340 33444 59346 33496
rect 59398 33484 59404 33496
rect 60326 33487 60384 33493
rect 60326 33484 60338 33487
rect 59398 33456 60338 33484
rect 59398 33444 59404 33456
rect 60326 33453 60338 33456
rect 60372 33453 60384 33487
rect 60904 33484 60910 33496
rect 60326 33447 60384 33453
rect 60462 33456 60910 33484
rect 58070 33388 59110 33416
rect 59156 33376 59162 33428
rect 59214 33416 59220 33428
rect 59987 33419 60045 33425
rect 59214 33388 59570 33416
rect 59214 33376 59220 33388
rect 52351 33351 52409 33357
rect 52351 33348 52363 33351
rect 47306 33320 52363 33348
rect 52351 33317 52363 33320
rect 52397 33348 52409 33351
rect 52535 33351 52593 33357
rect 52535 33348 52547 33351
rect 52397 33320 52547 33348
rect 52397 33317 52409 33320
rect 52351 33311 52409 33317
rect 52535 33317 52547 33320
rect 52581 33317 52593 33351
rect 57592 33348 57598 33360
rect 57553 33320 57598 33348
rect 52535 33311 52593 33317
rect 57592 33308 57598 33320
rect 57650 33308 57656 33360
rect 57960 33348 57966 33360
rect 57873 33320 57966 33348
rect 57960 33308 57966 33320
rect 58018 33348 58024 33360
rect 59432 33348 59438 33360
rect 58018 33320 59438 33348
rect 58018 33308 58024 33320
rect 59432 33308 59438 33320
rect 59490 33308 59496 33360
rect 59542 33348 59570 33388
rect 59987 33385 59999 33419
rect 60033 33416 60045 33419
rect 60462 33416 60490 33456
rect 60904 33444 60910 33456
rect 60962 33444 60968 33496
rect 63020 33444 63026 33496
rect 63078 33484 63084 33496
rect 63207 33487 63265 33493
rect 63207 33484 63219 33487
rect 63078 33456 63219 33484
rect 63078 33444 63084 33456
rect 63207 33453 63219 33456
rect 63253 33453 63265 33487
rect 63590 33484 63618 33515
rect 65964 33512 65970 33524
rect 66022 33512 66028 33564
rect 68724 33552 68730 33564
rect 68685 33524 68730 33552
rect 68724 33512 68730 33524
rect 68782 33512 68788 33564
rect 63940 33484 63946 33496
rect 63207 33447 63265 33453
rect 63314 33456 63618 33484
rect 63901 33456 63946 33484
rect 63115 33419 63173 33425
rect 63115 33416 63127 33419
rect 60033 33388 60490 33416
rect 60554 33388 63127 33416
rect 60033 33385 60045 33388
rect 59987 33379 60045 33385
rect 60554 33348 60582 33388
rect 63115 33385 63127 33388
rect 63161 33416 63173 33419
rect 63314 33416 63342 33456
rect 63940 33444 63946 33456
rect 63998 33444 64004 33496
rect 65746 33487 65804 33493
rect 65746 33453 65758 33487
rect 65792 33453 65804 33487
rect 67991 33487 68049 33493
rect 67991 33484 68003 33487
rect 65746 33447 65804 33453
rect 66258 33456 68003 33484
rect 63161 33388 63342 33416
rect 63161 33385 63173 33388
rect 63115 33379 63173 33385
rect 65504 33376 65510 33428
rect 65562 33416 65568 33428
rect 65599 33419 65657 33425
rect 65599 33416 65611 33419
rect 65562 33388 65611 33416
rect 65562 33376 65568 33388
rect 65599 33385 65611 33388
rect 65645 33385 65657 33419
rect 65761 33416 65789 33447
rect 66258 33416 66286 33456
rect 67991 33453 68003 33456
rect 68037 33453 68049 33487
rect 68632 33484 68638 33496
rect 68593 33456 68638 33484
rect 67991 33447 68049 33453
rect 68632 33444 68638 33456
rect 68690 33444 68696 33496
rect 69000 33484 69006 33496
rect 68961 33456 69006 33484
rect 69000 33444 69006 33456
rect 69058 33444 69064 33496
rect 69187 33487 69245 33493
rect 69187 33453 69199 33487
rect 69233 33484 69245 33487
rect 69233 33456 69414 33484
rect 69233 33453 69245 33456
rect 69187 33447 69245 33453
rect 65761 33388 66286 33416
rect 66335 33419 66393 33425
rect 65599 33379 65657 33385
rect 66335 33385 66347 33419
rect 66381 33416 66393 33419
rect 69092 33416 69098 33428
rect 66381 33388 69098 33416
rect 66381 33385 66393 33388
rect 66335 33379 66393 33385
rect 69092 33376 69098 33388
rect 69150 33376 69156 33428
rect 59542 33320 60582 33348
rect 61916 33308 61922 33360
rect 61974 33348 61980 33360
rect 65415 33351 65473 33357
rect 65415 33348 65427 33351
rect 61974 33320 65427 33348
rect 61974 33308 61980 33320
rect 65415 33317 65427 33320
rect 65461 33348 65473 33351
rect 65964 33348 65970 33360
rect 65461 33320 65970 33348
rect 65461 33317 65473 33320
rect 65415 33311 65473 33317
rect 65964 33308 65970 33320
rect 66022 33308 66028 33360
rect 67528 33308 67534 33360
rect 67586 33348 67592 33360
rect 67715 33351 67773 33357
rect 67715 33348 67727 33351
rect 67586 33320 67727 33348
rect 67586 33308 67592 33320
rect 67715 33317 67727 33320
rect 67761 33348 67773 33351
rect 68632 33348 68638 33360
rect 67761 33320 68638 33348
rect 67761 33317 67773 33320
rect 67715 33311 67773 33317
rect 68632 33308 68638 33320
rect 68690 33308 68696 33360
rect 69386 33357 69414 33456
rect 69662 33416 69690 33592
rect 81696 33580 81702 33592
rect 81754 33580 81760 33632
rect 86406 33620 86434 33660
rect 86406 33592 87354 33620
rect 73600 33552 73606 33564
rect 73561 33524 73606 33552
rect 73600 33512 73606 33524
rect 73658 33512 73664 33564
rect 74152 33552 74158 33564
rect 74113 33524 74158 33552
rect 74152 33512 74158 33524
rect 74210 33512 74216 33564
rect 78568 33512 78574 33564
rect 78626 33552 78632 33564
rect 78626 33524 79442 33552
rect 78626 33512 78632 33524
rect 73695 33487 73753 33493
rect 73695 33453 73707 33487
rect 73741 33484 73753 33487
rect 73876 33484 73882 33496
rect 73741 33456 73882 33484
rect 73741 33453 73753 33456
rect 73695 33447 73753 33453
rect 73876 33444 73882 33456
rect 73934 33444 73940 33496
rect 74428 33444 74434 33496
rect 74486 33484 74492 33496
rect 74983 33487 75041 33493
rect 74983 33484 74995 33487
rect 74486 33456 74995 33484
rect 74486 33444 74492 33456
rect 74983 33453 74995 33456
rect 75029 33484 75041 33487
rect 75348 33484 75354 33496
rect 75029 33456 75354 33484
rect 75029 33453 75041 33456
rect 74983 33447 75041 33453
rect 75348 33444 75354 33456
rect 75406 33444 75412 33496
rect 79215 33487 79273 33493
rect 79215 33453 79227 33487
rect 79261 33484 79273 33487
rect 79304 33484 79310 33496
rect 79261 33456 79310 33484
rect 79261 33453 79273 33456
rect 79215 33447 79273 33453
rect 79304 33444 79310 33456
rect 79362 33444 79368 33496
rect 79414 33493 79442 33524
rect 80408 33512 80414 33564
rect 80466 33552 80472 33564
rect 81423 33555 81481 33561
rect 81423 33552 81435 33555
rect 80466 33524 81435 33552
rect 80466 33512 80472 33524
rect 81423 33521 81435 33524
rect 81469 33521 81481 33555
rect 81423 33515 81481 33521
rect 79399 33487 79457 33493
rect 79399 33453 79411 33487
rect 79445 33453 79457 33487
rect 79856 33484 79862 33496
rect 79817 33456 79862 33484
rect 79399 33447 79457 33453
rect 79856 33444 79862 33456
rect 79914 33444 79920 33496
rect 79948 33444 79954 33496
rect 80006 33484 80012 33496
rect 80592 33484 80598 33496
rect 80006 33456 80598 33484
rect 80006 33444 80012 33456
rect 80592 33444 80598 33456
rect 80650 33484 80656 33496
rect 81607 33487 81665 33493
rect 81607 33484 81619 33487
rect 80650 33456 81619 33484
rect 80650 33444 80656 33456
rect 81607 33453 81619 33456
rect 81653 33453 81665 33487
rect 81607 33447 81665 33453
rect 82159 33487 82217 33493
rect 82159 33453 82171 33487
rect 82205 33453 82217 33487
rect 82340 33484 82346 33496
rect 82301 33456 82346 33484
rect 82159 33447 82217 33453
rect 80503 33419 80561 33425
rect 80503 33416 80515 33419
rect 69662 33388 80515 33416
rect 80503 33385 80515 33388
rect 80549 33385 80561 33419
rect 82174 33416 82202 33447
rect 82340 33444 82346 33456
rect 82398 33444 82404 33496
rect 86020 33484 86026 33496
rect 85981 33456 86026 33484
rect 86020 33444 86026 33456
rect 86078 33484 86084 33496
rect 86406 33493 86434 33592
rect 86207 33487 86265 33493
rect 86207 33484 86219 33487
rect 86078 33456 86219 33484
rect 86078 33444 86084 33456
rect 86207 33453 86219 33456
rect 86253 33453 86265 33487
rect 86207 33447 86265 33453
rect 86391 33487 86449 33493
rect 86391 33453 86403 33487
rect 86437 33453 86449 33487
rect 86391 33447 86449 33453
rect 86851 33487 86909 33493
rect 86851 33453 86863 33487
rect 86897 33453 86909 33487
rect 86851 33447 86909 33453
rect 86943 33487 87001 33493
rect 86943 33453 86955 33487
rect 86989 33484 87001 33487
rect 87326 33484 87354 33592
rect 90620 33580 90626 33632
rect 90678 33620 90684 33632
rect 91543 33623 91601 33629
rect 91543 33620 91555 33623
rect 90678 33592 91555 33620
rect 90678 33580 90684 33592
rect 91543 33589 91555 33592
rect 91589 33589 91601 33623
rect 91543 33583 91601 33589
rect 90344 33512 90350 33564
rect 90402 33552 90408 33564
rect 90531 33555 90589 33561
rect 90531 33552 90543 33555
rect 90402 33524 90543 33552
rect 90402 33512 90408 33524
rect 90531 33521 90543 33524
rect 90577 33552 90589 33555
rect 90577 33524 90758 33552
rect 90577 33521 90589 33524
rect 90531 33515 90589 33521
rect 86989 33456 87354 33484
rect 86989 33453 87001 33456
rect 86943 33447 87001 33453
rect 82248 33416 82254 33428
rect 82174 33388 82254 33416
rect 80503 33379 80561 33385
rect 82248 33376 82254 33388
rect 82306 33376 82312 33428
rect 82708 33416 82714 33428
rect 82669 33388 82714 33416
rect 82708 33376 82714 33388
rect 82766 33376 82772 33428
rect 86664 33376 86670 33428
rect 86722 33416 86728 33428
rect 86866 33416 86894 33447
rect 89792 33444 89798 33496
rect 89850 33484 89856 33496
rect 90623 33487 90681 33493
rect 90623 33484 90635 33487
rect 89850 33456 90635 33484
rect 89850 33444 89856 33456
rect 90623 33453 90635 33456
rect 90669 33453 90681 33487
rect 90730 33484 90758 33524
rect 91083 33487 91141 33493
rect 91083 33484 91095 33487
rect 90730 33456 91095 33484
rect 90623 33447 90681 33453
rect 91083 33453 91095 33456
rect 91129 33453 91141 33487
rect 91083 33447 91141 33453
rect 91175 33487 91233 33493
rect 91175 33453 91187 33487
rect 91221 33453 91233 33487
rect 91175 33447 91233 33453
rect 87679 33419 87737 33425
rect 87679 33416 87691 33419
rect 86722 33388 87691 33416
rect 86722 33376 86728 33388
rect 87679 33385 87691 33388
rect 87725 33385 87737 33419
rect 90638 33416 90666 33447
rect 91190 33416 91218 33447
rect 90638 33388 91218 33416
rect 87679 33379 87737 33385
rect 69371 33351 69429 33357
rect 69371 33317 69383 33351
rect 69417 33348 69429 33351
rect 69920 33348 69926 33360
rect 69417 33320 69926 33348
rect 69417 33317 69429 33320
rect 69371 33311 69429 33317
rect 69920 33308 69926 33320
rect 69978 33348 69984 33360
rect 72128 33348 72134 33360
rect 69978 33320 72134 33348
rect 69978 33308 69984 33320
rect 72128 33308 72134 33320
rect 72186 33308 72192 33360
rect 73876 33308 73882 33360
rect 73934 33348 73940 33360
rect 74339 33351 74397 33357
rect 74339 33348 74351 33351
rect 73934 33320 74351 33348
rect 73934 33308 73940 33320
rect 74339 33317 74351 33320
rect 74385 33348 74397 33351
rect 84180 33348 84186 33360
rect 74385 33320 84186 33348
rect 74385 33317 74397 33320
rect 74339 33311 74397 33317
rect 84180 33308 84186 33320
rect 84238 33308 84244 33360
rect 87403 33351 87461 33357
rect 87403 33317 87415 33351
rect 87449 33348 87461 33351
rect 87584 33348 87590 33360
rect 87449 33320 87590 33348
rect 87449 33317 87461 33320
rect 87403 33311 87461 33317
rect 87584 33308 87590 33320
rect 87642 33308 87648 33360
rect 538 33258 93642 33280
rect 538 33206 6344 33258
rect 6396 33206 6408 33258
rect 6460 33206 6472 33258
rect 6524 33206 6536 33258
rect 6588 33206 11672 33258
rect 11724 33206 11736 33258
rect 11788 33206 11800 33258
rect 11852 33206 11864 33258
rect 11916 33206 17000 33258
rect 17052 33206 17064 33258
rect 17116 33206 17128 33258
rect 17180 33206 17192 33258
rect 17244 33206 22328 33258
rect 22380 33206 22392 33258
rect 22444 33206 22456 33258
rect 22508 33206 22520 33258
rect 22572 33206 27656 33258
rect 27708 33206 27720 33258
rect 27772 33206 27784 33258
rect 27836 33206 27848 33258
rect 27900 33206 32984 33258
rect 33036 33206 33048 33258
rect 33100 33206 33112 33258
rect 33164 33206 33176 33258
rect 33228 33206 38312 33258
rect 38364 33206 38376 33258
rect 38428 33206 38440 33258
rect 38492 33206 38504 33258
rect 38556 33206 43640 33258
rect 43692 33206 43704 33258
rect 43756 33206 43768 33258
rect 43820 33206 43832 33258
rect 43884 33206 48968 33258
rect 49020 33206 49032 33258
rect 49084 33206 49096 33258
rect 49148 33206 49160 33258
rect 49212 33206 54296 33258
rect 54348 33206 54360 33258
rect 54412 33206 54424 33258
rect 54476 33206 54488 33258
rect 54540 33206 59624 33258
rect 59676 33206 59688 33258
rect 59740 33206 59752 33258
rect 59804 33206 59816 33258
rect 59868 33206 64952 33258
rect 65004 33206 65016 33258
rect 65068 33206 65080 33258
rect 65132 33206 65144 33258
rect 65196 33206 70280 33258
rect 70332 33206 70344 33258
rect 70396 33206 70408 33258
rect 70460 33206 70472 33258
rect 70524 33206 75608 33258
rect 75660 33206 75672 33258
rect 75724 33206 75736 33258
rect 75788 33206 75800 33258
rect 75852 33206 80936 33258
rect 80988 33206 81000 33258
rect 81052 33206 81064 33258
rect 81116 33206 81128 33258
rect 81180 33206 86264 33258
rect 86316 33206 86328 33258
rect 86380 33206 86392 33258
rect 86444 33206 86456 33258
rect 86508 33206 91592 33258
rect 91644 33206 91656 33258
rect 91708 33206 91720 33258
rect 91772 33206 91784 33258
rect 91836 33206 93642 33258
rect 538 33184 93642 33206
rect 6535 33147 6593 33153
rect 6535 33113 6547 33147
rect 6581 33144 6593 33147
rect 7084 33144 7090 33156
rect 6581 33116 7090 33144
rect 6581 33113 6593 33116
rect 6535 33107 6593 33113
rect 7084 33104 7090 33116
rect 7142 33104 7148 33156
rect 13435 33147 13493 33153
rect 13435 33113 13447 33147
rect 13481 33144 13493 33147
rect 15088 33144 15094 33156
rect 13481 33116 15094 33144
rect 13481 33113 13493 33116
rect 13435 33107 13493 33113
rect 4692 33008 4698 33020
rect 4653 32980 4698 33008
rect 4692 32968 4698 32980
rect 4750 32968 4756 33020
rect 4968 33008 4974 33020
rect 4929 32980 4974 33008
rect 4968 32968 4974 32980
rect 5026 32968 5032 33020
rect 10028 33008 10034 33020
rect 9989 32980 10034 33008
rect 10028 32968 10034 32980
rect 10086 33008 10092 33020
rect 11316 33008 11322 33020
rect 10086 32980 11322 33008
rect 10086 32968 10092 32980
rect 11316 32968 11322 32980
rect 11374 33008 11380 33020
rect 11779 33011 11837 33017
rect 11779 33008 11791 33011
rect 11374 32980 11791 33008
rect 11374 32968 11380 32980
rect 11779 32977 11791 32980
rect 11825 32977 11837 33011
rect 11779 32971 11837 32977
rect 12420 32968 12426 33020
rect 12478 33008 12484 33020
rect 12515 33011 12573 33017
rect 12515 33008 12527 33011
rect 12478 32980 12527 33008
rect 12478 32968 12484 32980
rect 12515 32977 12527 32980
rect 12561 32977 12573 33011
rect 12515 32971 12573 32977
rect 13156 32968 13162 33020
rect 13214 33008 13220 33020
rect 13542 33017 13570 33116
rect 15088 33104 15094 33116
rect 15146 33144 15152 33156
rect 15824 33144 15830 33156
rect 15146 33116 15830 33144
rect 15146 33104 15152 33116
rect 15824 33104 15830 33116
rect 15882 33104 15888 33156
rect 18676 33104 18682 33156
rect 18734 33144 18740 33156
rect 18863 33147 18921 33153
rect 18863 33144 18875 33147
rect 18734 33116 18875 33144
rect 18734 33104 18740 33116
rect 18863 33113 18875 33116
rect 18909 33113 18921 33147
rect 18863 33107 18921 33113
rect 21620 33104 21626 33156
rect 21678 33144 21684 33156
rect 21991 33147 22049 33153
rect 21991 33144 22003 33147
rect 21678 33116 22003 33144
rect 21678 33104 21684 33116
rect 21991 33113 22003 33116
rect 22037 33113 22049 33147
rect 21991 33107 22049 33113
rect 18771 33079 18829 33085
rect 18771 33076 18783 33079
rect 17958 33048 18783 33076
rect 17958 33017 17986 33048
rect 18771 33045 18783 33048
rect 18817 33076 18829 33079
rect 18952 33076 18958 33088
rect 18817 33048 18958 33076
rect 18817 33045 18829 33048
rect 18771 33039 18829 33045
rect 18952 33036 18958 33048
rect 19010 33076 19016 33088
rect 19320 33076 19326 33088
rect 19010 33048 19326 33076
rect 19010 33036 19016 33048
rect 19320 33036 19326 33048
rect 19378 33036 19384 33088
rect 13527 33011 13585 33017
rect 13527 33008 13539 33011
rect 13214 32980 13539 33008
rect 13214 32968 13220 32980
rect 13527 32977 13539 32980
rect 13573 32977 13585 33011
rect 13527 32971 13585 32977
rect 17391 33011 17449 33017
rect 17391 32977 17403 33011
rect 17437 32977 17449 33011
rect 17391 32971 17449 32977
rect 17943 33011 18001 33017
rect 17943 32977 17955 33011
rect 17989 32977 18001 33011
rect 17943 32971 18001 32977
rect 18127 33011 18185 33017
rect 18127 32977 18139 33011
rect 18173 33008 18185 33011
rect 18676 33008 18682 33020
rect 18173 32980 18682 33008
rect 18173 32977 18185 32980
rect 18127 32971 18185 32977
rect 10307 32943 10365 32949
rect 10307 32909 10319 32943
rect 10353 32940 10365 32943
rect 12607 32943 12665 32949
rect 12607 32940 12619 32943
rect 10353 32912 12619 32940
rect 10353 32909 10365 32912
rect 10307 32903 10365 32909
rect 12607 32909 12619 32912
rect 12653 32909 12665 32943
rect 17296 32940 17302 32952
rect 17257 32912 17302 32940
rect 12607 32903 12665 32909
rect 17296 32900 17302 32912
rect 17354 32900 17360 32952
rect 14168 32872 14174 32884
rect 10966 32844 14174 32872
rect 6256 32804 6262 32816
rect 6217 32776 6262 32804
rect 6256 32764 6262 32776
rect 6314 32764 6320 32816
rect 10396 32764 10402 32816
rect 10454 32804 10460 32816
rect 10966 32804 10994 32844
rect 14168 32832 14174 32844
rect 14226 32832 14232 32884
rect 17406 32872 17434 32971
rect 18676 32968 18682 32980
rect 18734 32968 18740 33020
rect 20887 33011 20945 33017
rect 20887 33008 20899 33011
rect 18878 32980 20899 33008
rect 18878 32884 18906 32980
rect 18860 32872 18866 32884
rect 17406 32844 18866 32872
rect 18860 32832 18866 32844
rect 18918 32832 18924 32884
rect 20718 32872 20746 32980
rect 20887 32977 20899 32980
rect 20933 32977 20945 33011
rect 22006 33008 22034 33107
rect 24288 33104 24294 33156
rect 24346 33144 24352 33156
rect 28796 33144 28802 33156
rect 24346 33116 28802 33144
rect 24346 33104 24352 33116
rect 28796 33104 28802 33116
rect 28854 33104 28860 33156
rect 28888 33104 28894 33156
rect 28946 33144 28952 33156
rect 28983 33147 29041 33153
rect 28983 33144 28995 33147
rect 28946 33116 28995 33144
rect 28946 33104 28952 33116
rect 28983 33113 28995 33116
rect 29029 33113 29041 33147
rect 33396 33144 33402 33156
rect 28983 33107 29041 33113
rect 31666 33116 33402 33144
rect 25944 33076 25950 33088
rect 25905 33048 25950 33076
rect 25944 33036 25950 33048
rect 26002 33036 26008 33088
rect 22175 33011 22233 33017
rect 22175 33008 22187 33011
rect 22006 32980 22187 33008
rect 20887 32971 20945 32977
rect 22175 32977 22187 32980
rect 22221 32977 22233 33011
rect 22175 32971 22233 32977
rect 25211 33011 25269 33017
rect 25211 32977 25223 33011
rect 25257 33008 25269 33011
rect 25257 32980 25530 33008
rect 25257 32977 25269 32980
rect 25211 32971 25269 32977
rect 20795 32943 20853 32949
rect 20795 32909 20807 32943
rect 20841 32940 20853 32943
rect 23368 32940 23374 32952
rect 20841 32912 23374 32940
rect 20841 32909 20853 32912
rect 20795 32903 20853 32909
rect 23368 32900 23374 32912
rect 23426 32900 23432 32952
rect 22267 32875 22325 32881
rect 22267 32872 22279 32875
rect 20718 32844 22279 32872
rect 22267 32841 22279 32844
rect 22313 32841 22325 32875
rect 22267 32835 22325 32841
rect 25027 32875 25085 32881
rect 25027 32841 25039 32875
rect 25073 32872 25085 32875
rect 25392 32872 25398 32884
rect 25073 32844 25398 32872
rect 25073 32841 25085 32844
rect 25027 32835 25085 32841
rect 25392 32832 25398 32844
rect 25450 32832 25456 32884
rect 10454 32776 10994 32804
rect 10454 32764 10460 32776
rect 11224 32764 11230 32816
rect 11282 32804 11288 32816
rect 11411 32807 11469 32813
rect 11411 32804 11423 32807
rect 11282 32776 11423 32804
rect 11282 32764 11288 32776
rect 11411 32773 11423 32776
rect 11457 32773 11469 32807
rect 13616 32804 13622 32816
rect 13577 32776 13622 32804
rect 11411 32767 11469 32773
rect 13616 32764 13622 32776
rect 13674 32764 13680 32816
rect 16100 32764 16106 32816
rect 16158 32804 16164 32816
rect 18403 32807 18461 32813
rect 18403 32804 18415 32807
rect 16158 32776 18415 32804
rect 16158 32764 16164 32776
rect 18403 32773 18415 32776
rect 18449 32773 18461 32807
rect 21068 32804 21074 32816
rect 21029 32776 21074 32804
rect 18403 32767 18461 32773
rect 21068 32764 21074 32776
rect 21126 32764 21132 32816
rect 25303 32807 25361 32813
rect 25303 32773 25315 32807
rect 25349 32804 25361 32807
rect 25502 32804 25530 32980
rect 25760 32968 25766 33020
rect 25818 33008 25824 33020
rect 26591 33011 26649 33017
rect 26591 33008 26603 33011
rect 25818 32980 26603 33008
rect 25818 32968 25824 32980
rect 26591 32977 26603 32980
rect 26637 32977 26649 33011
rect 26591 32971 26649 32977
rect 26128 32900 26134 32952
rect 26186 32940 26192 32952
rect 26407 32943 26465 32949
rect 26407 32940 26419 32943
rect 26186 32912 26419 32940
rect 26186 32900 26192 32912
rect 26407 32909 26419 32912
rect 26453 32909 26465 32943
rect 26407 32903 26465 32909
rect 26606 32872 26634 32971
rect 26772 32968 26778 33020
rect 26830 33008 26836 33020
rect 26959 33011 27017 33017
rect 26959 33008 26971 33011
rect 26830 32980 26971 33008
rect 26830 32968 26836 32980
rect 26959 32977 26971 32980
rect 27005 33008 27017 33011
rect 28891 33011 28949 33017
rect 27005 32980 27554 33008
rect 27005 32977 27017 32980
rect 26959 32971 27017 32977
rect 26864 32940 26870 32952
rect 26825 32912 26870 32940
rect 26864 32900 26870 32912
rect 26922 32900 26928 32952
rect 26606 32844 26818 32872
rect 26790 32816 26818 32844
rect 27526 32816 27554 32980
rect 28891 32977 28903 33011
rect 28937 33008 28949 33011
rect 29164 33008 29170 33020
rect 28937 32980 29170 33008
rect 28937 32977 28949 32980
rect 28891 32971 28949 32977
rect 29164 32968 29170 32980
rect 29222 32968 29228 33020
rect 31559 33011 31617 33017
rect 31559 32977 31571 33011
rect 31605 33008 31617 33011
rect 31666 33008 31694 33116
rect 33396 33104 33402 33116
rect 33454 33144 33460 33156
rect 33859 33147 33917 33153
rect 33859 33144 33871 33147
rect 33454 33116 33871 33144
rect 33454 33104 33460 33116
rect 33859 33113 33871 33116
rect 33905 33113 33917 33147
rect 35420 33144 35426 33156
rect 35381 33116 35426 33144
rect 33859 33107 33917 33113
rect 31832 33008 31838 33020
rect 31605 32980 31694 33008
rect 31793 32980 31838 33008
rect 31605 32977 31617 32980
rect 31559 32971 31617 32977
rect 31832 32968 31838 32980
rect 31890 32968 31896 33020
rect 33874 33008 33902 33107
rect 35420 33104 35426 33116
rect 35478 33104 35484 33156
rect 39284 33144 39290 33156
rect 39245 33116 39290 33144
rect 39284 33104 39290 33116
rect 39342 33104 39348 33156
rect 43703 33147 43761 33153
rect 43703 33113 43715 33147
rect 43749 33113 43761 33147
rect 43703 33107 43761 33113
rect 43718 33076 43746 33107
rect 43976 33104 43982 33156
rect 44034 33144 44040 33156
rect 44034 33116 49082 33144
rect 44034 33104 44040 33116
rect 44068 33076 44074 33088
rect 41418 33048 44074 33076
rect 34043 33011 34101 33017
rect 34043 33008 34055 33011
rect 33874 32980 34055 33008
rect 34043 32977 34055 32980
rect 34089 32977 34101 33011
rect 34043 32971 34101 32977
rect 34319 33011 34377 33017
rect 34319 32977 34331 33011
rect 34365 33008 34377 33011
rect 34408 33008 34414 33020
rect 34365 32980 34414 33008
rect 34365 32977 34377 32980
rect 34319 32971 34377 32977
rect 34408 32968 34414 32980
rect 34466 32968 34472 33020
rect 37812 32968 37818 33020
rect 37870 33008 37876 33020
rect 37907 33011 37965 33017
rect 37907 33008 37919 33011
rect 37870 32980 37919 33008
rect 37870 32968 37876 32980
rect 37907 32977 37919 32980
rect 37953 33008 37965 33011
rect 37953 32980 39882 33008
rect 37953 32977 37965 32980
rect 37907 32971 37965 32977
rect 38183 32943 38241 32949
rect 38183 32909 38195 32943
rect 38229 32940 38241 32943
rect 39744 32940 39750 32952
rect 38229 32912 39750 32940
rect 38229 32909 38241 32912
rect 38183 32903 38241 32909
rect 39744 32900 39750 32912
rect 39802 32900 39808 32952
rect 39854 32940 39882 32980
rect 40020 32968 40026 33020
rect 40078 33008 40084 33020
rect 41035 33011 41093 33017
rect 41035 33008 41047 33011
rect 40078 32980 41047 33008
rect 40078 32968 40084 32980
rect 41035 32977 41047 32980
rect 41081 32977 41093 33011
rect 41035 32971 41093 32977
rect 41124 32968 41130 33020
rect 41182 33008 41188 33020
rect 41418 33017 41446 33048
rect 44068 33036 44074 33048
rect 44126 33036 44132 33088
rect 46923 33079 46981 33085
rect 46923 33045 46935 33079
rect 46969 33076 46981 33079
rect 47472 33076 47478 33088
rect 46969 33048 47478 33076
rect 46969 33045 46981 33048
rect 46923 33039 46981 33045
rect 47472 33036 47478 33048
rect 47530 33076 47536 33088
rect 49054 33076 49082 33116
rect 49312 33104 49318 33156
rect 49370 33144 49376 33156
rect 57592 33144 57598 33156
rect 49370 33116 57598 33144
rect 49370 33104 49376 33116
rect 57592 33104 57598 33116
rect 57650 33144 57656 33156
rect 58420 33144 58426 33156
rect 57650 33116 58426 33144
rect 57650 33104 57656 33116
rect 58420 33104 58426 33116
rect 58478 33104 58484 33156
rect 58515 33147 58573 33153
rect 58515 33113 58527 33147
rect 58561 33144 58573 33147
rect 59340 33144 59346 33156
rect 58561 33116 59346 33144
rect 58561 33113 58573 33116
rect 58515 33107 58573 33113
rect 59340 33104 59346 33116
rect 59398 33104 59404 33156
rect 59772 33116 59938 33144
rect 59772 33076 59800 33116
rect 47530 33048 48990 33076
rect 49054 33048 59800 33076
rect 59910 33076 59938 33116
rect 60076 33104 60082 33156
rect 60134 33144 60140 33156
rect 60815 33147 60873 33153
rect 60815 33144 60827 33147
rect 60134 33116 60827 33144
rect 60134 33104 60140 33116
rect 60815 33113 60827 33116
rect 60861 33113 60873 33147
rect 60815 33107 60873 33113
rect 60904 33104 60910 33156
rect 60962 33144 60968 33156
rect 61183 33147 61241 33153
rect 61183 33144 61195 33147
rect 60962 33116 61195 33144
rect 60962 33104 60968 33116
rect 61183 33113 61195 33116
rect 61229 33144 61241 33147
rect 65412 33144 65418 33156
rect 61229 33116 65418 33144
rect 61229 33113 61241 33116
rect 61183 33107 61241 33113
rect 65412 33104 65418 33116
rect 65470 33104 65476 33156
rect 65504 33104 65510 33156
rect 65562 33144 65568 33156
rect 65875 33147 65933 33153
rect 65875 33144 65887 33147
rect 65562 33116 65887 33144
rect 65562 33104 65568 33116
rect 65875 33113 65887 33116
rect 65921 33113 65933 33147
rect 65875 33107 65933 33113
rect 65964 33104 65970 33156
rect 66022 33144 66028 33156
rect 66151 33147 66209 33153
rect 66151 33144 66163 33147
rect 66022 33116 66163 33144
rect 66022 33104 66028 33116
rect 66151 33113 66163 33116
rect 66197 33144 66209 33147
rect 82619 33147 82677 33153
rect 82619 33144 82631 33147
rect 66197 33116 82631 33144
rect 66197 33113 66209 33116
rect 66151 33107 66209 33113
rect 82619 33113 82631 33116
rect 82665 33113 82677 33147
rect 82892 33144 82898 33156
rect 82853 33116 82898 33144
rect 82619 33107 82677 33113
rect 82892 33104 82898 33116
rect 82950 33144 82956 33156
rect 82950 33116 84042 33144
rect 82950 33104 82956 33116
rect 61088 33076 61094 33088
rect 59910 33048 61094 33076
rect 47530 33036 47536 33048
rect 41403 33011 41461 33017
rect 41182 32980 41227 33008
rect 41182 32968 41188 32980
rect 41403 32977 41415 33011
rect 41449 32977 41461 33011
rect 41403 32971 41461 32977
rect 43525 33011 43583 33017
rect 43525 32977 43537 33011
rect 43571 32977 43583 33011
rect 43525 32971 43583 32977
rect 40664 32940 40670 32952
rect 39854 32912 40670 32940
rect 40664 32900 40670 32912
rect 40722 32900 40728 32952
rect 40756 32900 40762 32952
rect 40814 32940 40820 32952
rect 41418 32940 41446 32971
rect 40814 32912 41446 32940
rect 41495 32943 41553 32949
rect 40814 32900 40820 32912
rect 41495 32909 41507 32943
rect 41541 32940 41553 32943
rect 43534 32940 43562 32971
rect 44436 32968 44442 33020
rect 44494 33008 44500 33020
rect 44623 33011 44681 33017
rect 44623 33008 44635 33011
rect 44494 32980 44635 33008
rect 44494 32968 44500 32980
rect 44623 32977 44635 32980
rect 44669 32977 44681 33011
rect 44623 32971 44681 32977
rect 44712 32968 44718 33020
rect 44770 33017 44776 33020
rect 44770 33011 44828 33017
rect 44770 32977 44782 33011
rect 44816 32977 44828 33011
rect 44770 32971 44828 32977
rect 47015 33011 47073 33017
rect 47015 32977 47027 33011
rect 47061 33008 47073 33011
rect 47196 33008 47202 33020
rect 47061 32980 47202 33008
rect 47061 32977 47073 32980
rect 47015 32971 47073 32977
rect 44770 32968 44776 32971
rect 47196 32968 47202 32980
rect 47254 32968 47260 33020
rect 48962 33017 48990 33048
rect 61088 33036 61094 33048
rect 61146 33036 61152 33088
rect 61272 33036 61278 33088
rect 61330 33076 61336 33088
rect 77832 33076 77838 33088
rect 61330 33048 77838 33076
rect 61330 33036 61336 33048
rect 77832 33036 77838 33048
rect 77890 33036 77896 33088
rect 78568 33076 78574 33088
rect 78126 33048 78574 33076
rect 48947 33011 49005 33017
rect 48947 32977 48959 33011
rect 48993 32977 49005 33011
rect 49680 33008 49686 33020
rect 48947 32971 49005 32977
rect 49238 32980 49686 33008
rect 44730 32940 44758 32968
rect 44988 32940 44994 32952
rect 41541 32912 41998 32940
rect 43534 32912 44758 32940
rect 44949 32912 44994 32940
rect 41541 32909 41553 32912
rect 41495 32903 41553 32909
rect 37812 32872 37818 32884
rect 37773 32844 37818 32872
rect 37812 32832 37818 32844
rect 37870 32832 37876 32884
rect 40406 32844 40986 32872
rect 25760 32804 25766 32816
rect 25349 32776 25766 32804
rect 25349 32773 25361 32776
rect 25303 32767 25361 32773
rect 25760 32764 25766 32776
rect 25818 32764 25824 32816
rect 26772 32764 26778 32816
rect 26830 32804 26836 32816
rect 27235 32807 27293 32813
rect 27235 32804 27247 32807
rect 26830 32776 27247 32804
rect 26830 32764 26836 32776
rect 27235 32773 27247 32776
rect 27281 32773 27293 32807
rect 27508 32804 27514 32816
rect 27469 32776 27514 32804
rect 27235 32767 27293 32773
rect 27508 32764 27514 32776
rect 27566 32764 27572 32816
rect 33028 32764 33034 32816
rect 33086 32804 33092 32816
rect 33123 32807 33181 32813
rect 33123 32804 33135 32807
rect 33086 32776 33135 32804
rect 33086 32764 33092 32776
rect 33123 32773 33135 32776
rect 33169 32773 33181 32807
rect 33123 32767 33181 32773
rect 37720 32764 37726 32816
rect 37778 32804 37784 32816
rect 40406 32804 40434 32844
rect 37778 32776 40434 32804
rect 40483 32807 40541 32813
rect 37778 32764 37784 32776
rect 40483 32773 40495 32807
rect 40529 32804 40541 32807
rect 40848 32804 40854 32816
rect 40529 32776 40854 32804
rect 40529 32773 40541 32776
rect 40483 32767 40541 32773
rect 40848 32764 40854 32776
rect 40906 32764 40912 32816
rect 40958 32804 40986 32844
rect 41124 32832 41130 32884
rect 41182 32872 41188 32884
rect 41768 32872 41774 32884
rect 41182 32844 41774 32872
rect 41182 32832 41188 32844
rect 41768 32832 41774 32844
rect 41826 32832 41832 32884
rect 41970 32881 41998 32912
rect 44988 32900 44994 32912
rect 45046 32900 45052 32952
rect 47288 32900 47294 32952
rect 47346 32940 47352 32952
rect 49238 32940 49266 32980
rect 49680 32968 49686 32980
rect 49738 32968 49744 33020
rect 54743 33011 54801 33017
rect 54743 32977 54755 33011
rect 54789 33008 54801 33011
rect 57408 33008 57414 33020
rect 54789 32980 57414 33008
rect 54789 32977 54801 32980
rect 54743 32971 54801 32977
rect 47346 32912 49266 32940
rect 49315 32943 49373 32949
rect 47346 32900 47352 32912
rect 49315 32909 49327 32943
rect 49361 32940 49373 32943
rect 51428 32940 51434 32952
rect 49361 32912 51434 32940
rect 49361 32909 49373 32912
rect 49315 32903 49373 32909
rect 51428 32900 51434 32912
rect 51486 32900 51492 32952
rect 41955 32875 42013 32881
rect 41955 32841 41967 32875
rect 42001 32872 42013 32875
rect 42320 32872 42326 32884
rect 42001 32844 42326 32872
rect 42001 32841 42013 32844
rect 41955 32835 42013 32841
rect 42320 32832 42326 32844
rect 42378 32832 42384 32884
rect 44896 32872 44902 32884
rect 44857 32844 44902 32872
rect 44896 32832 44902 32844
rect 44954 32832 44960 32884
rect 45267 32875 45325 32881
rect 45267 32841 45279 32875
rect 45313 32872 45325 32875
rect 45313 32844 50554 32872
rect 45313 32841 45325 32844
rect 45267 32835 45325 32841
rect 44160 32804 44166 32816
rect 40958 32776 44166 32804
rect 44160 32764 44166 32776
rect 44218 32764 44224 32816
rect 44436 32804 44442 32816
rect 44397 32776 44442 32804
rect 44436 32764 44442 32776
rect 44494 32764 44500 32816
rect 44804 32764 44810 32816
rect 44862 32804 44868 32816
rect 46736 32804 46742 32816
rect 44862 32776 46742 32804
rect 44862 32764 44868 32776
rect 46736 32764 46742 32776
rect 46794 32764 46800 32816
rect 46828 32764 46834 32816
rect 46886 32804 46892 32816
rect 47199 32807 47257 32813
rect 47199 32804 47211 32807
rect 46886 32776 47211 32804
rect 46886 32764 46892 32776
rect 47199 32773 47211 32776
rect 47245 32773 47257 32807
rect 47564 32804 47570 32816
rect 47525 32776 47570 32804
rect 47199 32767 47257 32773
rect 47564 32764 47570 32776
rect 47622 32764 47628 32816
rect 47656 32764 47662 32816
rect 47714 32804 47720 32816
rect 48576 32804 48582 32816
rect 47714 32776 48582 32804
rect 47714 32764 47720 32776
rect 48576 32764 48582 32776
rect 48634 32764 48640 32816
rect 50526 32804 50554 32844
rect 50600 32832 50606 32884
rect 50658 32872 50664 32884
rect 50658 32844 53406 32872
rect 50658 32832 50664 32844
rect 52900 32804 52906 32816
rect 50526 32776 52906 32804
rect 52900 32764 52906 32776
rect 52958 32764 52964 32816
rect 53378 32804 53406 32844
rect 54188 32832 54194 32884
rect 54246 32872 54252 32884
rect 54758 32872 54786 32971
rect 57408 32968 57414 32980
rect 57466 32968 57472 33020
rect 57503 33011 57561 33017
rect 57503 32977 57515 33011
rect 57549 33008 57561 33011
rect 57960 33008 57966 33020
rect 57549 32980 57966 33008
rect 57549 32977 57561 32980
rect 57503 32971 57561 32977
rect 57960 32968 57966 32980
rect 58018 32968 58024 33020
rect 58052 32968 58058 33020
rect 58110 33008 58116 33020
rect 58236 33008 58242 33020
rect 58110 32980 58155 33008
rect 58197 32980 58242 33008
rect 58110 32968 58116 32980
rect 58236 32968 58242 32980
rect 58294 33008 58300 33020
rect 59067 33011 59125 33017
rect 58294 32980 58466 33008
rect 58294 32968 58300 32980
rect 56580 32900 56586 32952
rect 56638 32940 56644 32952
rect 57043 32943 57101 32949
rect 57043 32940 57055 32943
rect 56638 32912 57055 32940
rect 56638 32900 56644 32912
rect 57043 32909 57055 32912
rect 57089 32940 57101 32943
rect 57135 32943 57193 32949
rect 57135 32940 57147 32943
rect 57089 32912 57147 32940
rect 57089 32909 57101 32912
rect 57043 32903 57101 32909
rect 57135 32909 57147 32912
rect 57181 32909 57193 32943
rect 57316 32940 57322 32952
rect 57277 32912 57322 32940
rect 57135 32903 57193 32909
rect 57316 32900 57322 32912
rect 57374 32900 57380 32952
rect 58438 32940 58466 32980
rect 59067 32977 59079 33011
rect 59113 33008 59125 33011
rect 59432 33008 59438 33020
rect 59113 32980 59438 33008
rect 59113 32977 59125 32980
rect 59067 32971 59125 32977
rect 59432 32968 59438 32980
rect 59490 33008 59496 33020
rect 59803 33011 59861 33017
rect 59490 32980 59754 33008
rect 59490 32968 59496 32980
rect 59343 32943 59401 32949
rect 59343 32940 59355 32943
rect 58438 32912 59355 32940
rect 59343 32909 59355 32912
rect 59389 32940 59401 32943
rect 59619 32943 59677 32949
rect 59619 32940 59631 32943
rect 59389 32912 59631 32940
rect 59389 32909 59401 32912
rect 59343 32903 59401 32909
rect 59619 32909 59631 32912
rect 59665 32909 59677 32943
rect 59726 32940 59754 32980
rect 59803 32977 59815 33011
rect 59849 33008 59861 33011
rect 60168 33008 60174 33020
rect 59849 32980 60174 33008
rect 59849 32977 59861 32980
rect 59803 32971 59861 32977
rect 60168 32968 60174 32980
rect 60226 32968 60232 33020
rect 60352 33008 60358 33020
rect 60313 32980 60358 33008
rect 60352 32968 60358 32980
rect 60410 32968 60416 33020
rect 60539 33011 60597 33017
rect 60539 32977 60551 33011
rect 60585 33008 60597 33011
rect 60904 33008 60910 33020
rect 60585 32980 60910 33008
rect 60585 32977 60597 32980
rect 60539 32971 60597 32977
rect 60904 32968 60910 32980
rect 60962 32968 60968 33020
rect 62744 32968 62750 33020
rect 62802 33008 62808 33020
rect 62928 33008 62934 33020
rect 62802 32980 62934 33008
rect 62802 32968 62808 32980
rect 62928 32968 62934 32980
rect 62986 32968 62992 33020
rect 63115 33011 63173 33017
rect 63115 32977 63127 33011
rect 63161 32977 63173 33011
rect 63115 32971 63173 32977
rect 63130 32940 63158 32971
rect 63204 32968 63210 33020
rect 63262 33008 63268 33020
rect 63575 33011 63633 33017
rect 63575 33008 63587 33011
rect 63262 32980 63587 33008
rect 63262 32968 63268 32980
rect 63575 32977 63587 32980
rect 63621 32977 63633 33011
rect 63575 32971 63633 32977
rect 63667 33011 63725 33017
rect 63667 32977 63679 33011
rect 63713 33008 63725 33011
rect 65044 33008 65050 33020
rect 63713 32980 64078 33008
rect 63713 32977 63725 32980
rect 63667 32971 63725 32977
rect 59726 32912 59938 32940
rect 63130 32912 63250 32940
rect 59619 32903 59677 32909
rect 54246 32844 54786 32872
rect 54927 32875 54985 32881
rect 54246 32832 54252 32844
rect 54927 32841 54939 32875
rect 54973 32872 54985 32875
rect 59800 32872 59806 32884
rect 54973 32844 59806 32872
rect 54973 32841 54985 32844
rect 54927 32835 54985 32841
rect 54942 32804 54970 32835
rect 59800 32832 59806 32844
rect 59858 32832 59864 32884
rect 59910 32872 59938 32912
rect 63222 32872 63250 32912
rect 63848 32872 63854 32884
rect 59910 32844 61502 32872
rect 63222 32844 63854 32872
rect 53378 32776 54970 32804
rect 57043 32807 57101 32813
rect 57043 32773 57055 32807
rect 57089 32804 57101 32807
rect 58236 32804 58242 32816
rect 57089 32776 58242 32804
rect 57089 32773 57101 32776
rect 57043 32767 57101 32773
rect 58236 32764 58242 32776
rect 58294 32764 58300 32816
rect 58328 32764 58334 32816
rect 58386 32804 58392 32816
rect 58788 32804 58794 32816
rect 58386 32776 58794 32804
rect 58386 32764 58392 32776
rect 58788 32764 58794 32776
rect 58846 32764 58852 32816
rect 59340 32764 59346 32816
rect 59398 32804 59404 32816
rect 60352 32804 60358 32816
rect 59398 32776 60358 32804
rect 59398 32764 59404 32776
rect 60352 32764 60358 32776
rect 60410 32764 60416 32816
rect 61364 32804 61370 32816
rect 61325 32776 61370 32804
rect 61364 32764 61370 32776
rect 61422 32764 61428 32816
rect 61474 32804 61502 32844
rect 63848 32832 63854 32844
rect 63906 32832 63912 32884
rect 64050 32804 64078 32980
rect 64970 32980 65050 33008
rect 64219 32943 64277 32949
rect 64219 32909 64231 32943
rect 64265 32940 64277 32943
rect 64970 32940 64998 32980
rect 65044 32968 65050 32980
rect 65102 32968 65108 33020
rect 65231 33011 65289 33017
rect 65231 32977 65243 33011
rect 65277 33008 65289 33011
rect 65780 33008 65786 33020
rect 65277 32980 65786 33008
rect 65277 32977 65289 32980
rect 65231 32971 65289 32977
rect 65780 32968 65786 32980
rect 65838 32968 65844 33020
rect 66516 33008 66522 33020
rect 66477 32980 66522 33008
rect 66516 32968 66522 32980
rect 66574 32968 66580 33020
rect 67068 32968 67074 33020
rect 67126 33008 67132 33020
rect 67126 32980 67298 33008
rect 67126 32968 67132 32980
rect 64265 32912 64998 32940
rect 64265 32909 64277 32912
rect 64219 32903 64277 32909
rect 65596 32900 65602 32952
rect 65654 32940 65660 32952
rect 66534 32940 66562 32968
rect 66884 32940 66890 32952
rect 65654 32912 65699 32940
rect 66534 32912 66890 32940
rect 65654 32900 65660 32912
rect 66884 32900 66890 32912
rect 66942 32900 66948 32952
rect 64124 32832 64130 32884
rect 64182 32872 64188 32884
rect 64403 32875 64461 32881
rect 64403 32872 64415 32875
rect 64182 32844 64415 32872
rect 64182 32832 64188 32844
rect 64403 32841 64415 32844
rect 64449 32841 64461 32875
rect 64676 32872 64682 32884
rect 64637 32844 64682 32872
rect 64403 32835 64461 32841
rect 64676 32832 64682 32844
rect 64734 32832 64740 32884
rect 65044 32872 65050 32884
rect 65005 32844 65050 32872
rect 65044 32832 65050 32844
rect 65102 32872 65108 32884
rect 65507 32875 65565 32881
rect 65507 32872 65519 32875
rect 65102 32844 65519 32872
rect 65102 32832 65108 32844
rect 65507 32841 65519 32844
rect 65553 32841 65565 32875
rect 67270 32872 67298 32980
rect 67436 32968 67442 33020
rect 67494 33008 67500 33020
rect 67531 33011 67589 33017
rect 67531 33008 67543 33011
rect 67494 32980 67543 33008
rect 67494 32968 67500 32980
rect 67531 32977 67543 32980
rect 67577 32977 67589 33011
rect 67531 32971 67589 32977
rect 67623 33011 67681 33017
rect 67623 32977 67635 33011
rect 67669 33008 67681 33011
rect 68540 33008 68546 33020
rect 67669 32980 68546 33008
rect 67669 32977 67681 32980
rect 67623 32971 67681 32977
rect 68540 32968 68546 32980
rect 68598 32968 68604 33020
rect 69092 33008 69098 33020
rect 69053 32980 69098 33008
rect 69092 32968 69098 32980
rect 69150 32968 69156 33020
rect 74339 33011 74397 33017
rect 74339 32977 74351 33011
rect 74385 32977 74397 33011
rect 74339 32971 74397 32977
rect 74354 32940 74382 32971
rect 74428 32968 74434 33020
rect 74486 33008 74492 33020
rect 74486 32980 74531 33008
rect 74486 32968 74492 32980
rect 74704 32968 74710 33020
rect 74762 33008 74768 33020
rect 74799 33011 74857 33017
rect 74799 33008 74811 33011
rect 74762 32980 74811 33008
rect 74762 32968 74768 32980
rect 74799 32977 74811 32980
rect 74845 32977 74857 33011
rect 74799 32971 74857 32977
rect 74891 33011 74949 33017
rect 74891 32977 74903 33011
rect 74937 33008 74949 33011
rect 76820 33008 76826 33020
rect 74937 32980 76826 33008
rect 74937 32977 74949 32980
rect 74891 32971 74949 32977
rect 76820 32968 76826 32980
rect 76878 33008 76884 33020
rect 77467 33011 77525 33017
rect 77467 33008 77479 33011
rect 76878 32980 77479 33008
rect 76878 32968 76884 32980
rect 77467 32977 77479 32980
rect 77513 32977 77525 33011
rect 77924 33008 77930 33020
rect 77885 32980 77930 33008
rect 77467 32971 77525 32977
rect 77924 32968 77930 32980
rect 77982 32968 77988 33020
rect 78126 33017 78154 33048
rect 78568 33036 78574 33048
rect 78626 33036 78632 33088
rect 82818 33048 83858 33076
rect 82818 33020 82846 33048
rect 78107 33011 78165 33017
rect 78107 32977 78119 33011
rect 78153 32977 78165 33011
rect 78107 32971 78165 32977
rect 78200 32968 78206 33020
rect 78258 33008 78264 33020
rect 82711 33011 82769 33017
rect 82711 33008 82723 33011
rect 78258 32980 82723 33008
rect 78258 32968 78264 32980
rect 82711 32977 82723 32980
rect 82757 33008 82769 33011
rect 82800 33008 82806 33020
rect 82757 32980 82806 33008
rect 82757 32977 82769 32980
rect 82711 32971 82769 32977
rect 82800 32968 82806 32980
rect 82858 32968 82864 33020
rect 83260 33008 83266 33020
rect 83221 32980 83266 33008
rect 83260 32968 83266 32980
rect 83318 32968 83324 33020
rect 83355 33011 83413 33017
rect 83355 32977 83367 33011
rect 83401 33008 83413 33011
rect 83628 33008 83634 33020
rect 83401 32980 83634 33008
rect 83401 32977 83413 32980
rect 83355 32971 83413 32977
rect 83628 32968 83634 32980
rect 83686 32968 83692 33020
rect 83830 33017 83858 33048
rect 83815 33011 83873 33017
rect 83815 32977 83827 33011
rect 83861 33008 83873 33011
rect 83904 33008 83910 33020
rect 83861 32980 83910 33008
rect 83861 32977 83873 32980
rect 83815 32971 83873 32977
rect 83904 32968 83910 32980
rect 83962 32968 83968 33020
rect 84014 33017 84042 33116
rect 83999 33011 84057 33017
rect 83999 32977 84011 33011
rect 84045 32977 84057 33011
rect 86575 33011 86633 33017
rect 86575 33008 86587 33011
rect 83999 32971 84057 32977
rect 84198 32980 86587 33008
rect 75348 32940 75354 32952
rect 74354 32912 74474 32940
rect 75309 32912 75354 32940
rect 68359 32875 68417 32881
rect 68359 32872 68371 32875
rect 67270 32844 68371 32872
rect 65507 32835 65565 32841
rect 68359 32841 68371 32844
rect 68405 32841 68417 32875
rect 68359 32835 68417 32841
rect 64863 32807 64921 32813
rect 64863 32804 64875 32807
rect 61474 32776 64875 32804
rect 64863 32773 64875 32776
rect 64909 32804 64921 32807
rect 65228 32804 65234 32816
rect 64909 32776 65234 32804
rect 64909 32773 64921 32776
rect 64863 32767 64921 32773
rect 65228 32764 65234 32776
rect 65286 32764 65292 32816
rect 65396 32807 65454 32813
rect 65396 32773 65408 32807
rect 65442 32804 65454 32807
rect 65964 32804 65970 32816
rect 65442 32776 65970 32804
rect 65442 32773 65454 32776
rect 65396 32767 65454 32773
rect 65964 32764 65970 32776
rect 66022 32764 66028 32816
rect 66700 32804 66706 32816
rect 66661 32776 66706 32804
rect 66700 32764 66706 32776
rect 66758 32764 66764 32816
rect 68080 32804 68086 32816
rect 68041 32776 68086 32804
rect 68080 32764 68086 32776
rect 68138 32764 68144 32816
rect 68374 32804 68402 32835
rect 68540 32832 68546 32884
rect 68598 32872 68604 32884
rect 68635 32875 68693 32881
rect 68635 32872 68647 32875
rect 68598 32844 68647 32872
rect 68598 32832 68604 32844
rect 68635 32841 68647 32844
rect 68681 32872 68693 32875
rect 69276 32872 69282 32884
rect 68681 32844 69282 32872
rect 68681 32841 68693 32844
rect 68635 32835 68693 32841
rect 69276 32832 69282 32844
rect 69334 32832 69340 32884
rect 69368 32832 69374 32884
rect 69426 32872 69432 32884
rect 71208 32872 71214 32884
rect 69426 32844 71214 32872
rect 69426 32832 69432 32844
rect 71208 32832 71214 32844
rect 71266 32832 71272 32884
rect 74063 32875 74121 32881
rect 74063 32841 74075 32875
rect 74109 32872 74121 32875
rect 74336 32872 74342 32884
rect 74109 32844 74342 32872
rect 74109 32841 74121 32844
rect 74063 32835 74121 32841
rect 74336 32832 74342 32844
rect 74394 32832 74400 32884
rect 68724 32804 68730 32816
rect 68374 32776 68730 32804
rect 68724 32764 68730 32776
rect 68782 32764 68788 32816
rect 69187 32807 69245 32813
rect 69187 32773 69199 32807
rect 69233 32804 69245 32807
rect 69736 32804 69742 32816
rect 69233 32776 69742 32804
rect 69233 32773 69245 32776
rect 69187 32767 69245 32773
rect 69736 32764 69742 32776
rect 69794 32764 69800 32816
rect 74446 32804 74474 32912
rect 75348 32900 75354 32912
rect 75406 32900 75412 32952
rect 77007 32943 77065 32949
rect 77007 32909 77019 32943
rect 77053 32940 77065 32943
rect 77283 32943 77341 32949
rect 77283 32940 77295 32943
rect 77053 32912 77295 32940
rect 77053 32909 77065 32912
rect 77007 32903 77065 32909
rect 77283 32909 77295 32912
rect 77329 32909 77341 32943
rect 77283 32903 77341 32909
rect 74520 32832 74526 32884
rect 74578 32872 74584 32884
rect 81512 32872 81518 32884
rect 74578 32844 81518 32872
rect 74578 32832 74584 32844
rect 81512 32832 81518 32844
rect 81570 32832 81576 32884
rect 82619 32875 82677 32881
rect 82619 32841 82631 32875
rect 82665 32872 82677 32875
rect 83444 32872 83450 32884
rect 82665 32844 83450 32872
rect 82665 32841 82677 32844
rect 82619 32835 82677 32841
rect 83444 32832 83450 32844
rect 83502 32832 83508 32884
rect 83628 32832 83634 32884
rect 83686 32872 83692 32884
rect 84198 32872 84226 32980
rect 86575 32977 86587 32980
rect 86621 33008 86633 33011
rect 87492 33008 87498 33020
rect 86621 32980 87498 33008
rect 86621 32977 86633 32980
rect 86575 32971 86633 32977
rect 87492 32968 87498 32980
rect 87550 32968 87556 33020
rect 87952 33008 87958 33020
rect 87913 32980 87958 33008
rect 87952 32968 87958 32980
rect 88010 32968 88016 33020
rect 87400 32900 87406 32952
rect 87458 32940 87464 32952
rect 87679 32943 87737 32949
rect 87679 32940 87691 32943
rect 87458 32912 87691 32940
rect 87458 32900 87464 32912
rect 87679 32909 87691 32912
rect 87725 32909 87737 32943
rect 87679 32903 87737 32909
rect 83686 32844 84226 32872
rect 83686 32832 83692 32844
rect 86112 32832 86118 32884
rect 86170 32872 86176 32884
rect 86170 32844 87538 32872
rect 86170 32832 86176 32844
rect 75624 32804 75630 32816
rect 74446 32776 75630 32804
rect 75624 32764 75630 32776
rect 75682 32764 75688 32816
rect 75900 32764 75906 32816
rect 75958 32804 75964 32816
rect 76636 32804 76642 32816
rect 75958 32776 76642 32804
rect 75958 32764 75964 32776
rect 76636 32764 76642 32776
rect 76694 32804 76700 32816
rect 77007 32807 77065 32813
rect 77007 32804 77019 32807
rect 76694 32776 77019 32804
rect 76694 32764 76700 32776
rect 77007 32773 77019 32776
rect 77053 32804 77065 32807
rect 77099 32807 77157 32813
rect 77099 32804 77111 32807
rect 77053 32776 77111 32804
rect 77053 32773 77065 32776
rect 77007 32767 77065 32773
rect 77099 32773 77111 32776
rect 77145 32773 77157 32807
rect 77099 32767 77157 32773
rect 78479 32807 78537 32813
rect 78479 32773 78491 32807
rect 78525 32804 78537 32807
rect 81420 32804 81426 32816
rect 78525 32776 81426 32804
rect 78525 32773 78537 32776
rect 78479 32767 78537 32773
rect 81420 32764 81426 32776
rect 81478 32764 81484 32816
rect 83076 32764 83082 32816
rect 83134 32804 83140 32816
rect 84088 32804 84094 32816
rect 83134 32776 84094 32804
rect 83134 32764 83140 32776
rect 84088 32764 84094 32776
rect 84146 32764 84152 32816
rect 84272 32804 84278 32816
rect 84233 32776 84278 32804
rect 84272 32764 84278 32776
rect 84330 32764 84336 32816
rect 86664 32804 86670 32816
rect 86625 32776 86670 32804
rect 86664 32764 86670 32776
rect 86722 32764 86728 32816
rect 87400 32804 87406 32816
rect 87361 32776 87406 32804
rect 87400 32764 87406 32776
rect 87458 32764 87464 32816
rect 87510 32804 87538 32844
rect 89059 32807 89117 32813
rect 89059 32804 89071 32807
rect 87510 32776 89071 32804
rect 89059 32773 89071 32776
rect 89105 32773 89117 32807
rect 89059 32767 89117 32773
rect 538 32714 93642 32736
rect 538 32662 3680 32714
rect 3732 32662 3744 32714
rect 3796 32662 3808 32714
rect 3860 32662 3872 32714
rect 3924 32662 9008 32714
rect 9060 32662 9072 32714
rect 9124 32662 9136 32714
rect 9188 32662 9200 32714
rect 9252 32662 14336 32714
rect 14388 32662 14400 32714
rect 14452 32662 14464 32714
rect 14516 32662 14528 32714
rect 14580 32662 19664 32714
rect 19716 32662 19728 32714
rect 19780 32662 19792 32714
rect 19844 32662 19856 32714
rect 19908 32662 24992 32714
rect 25044 32662 25056 32714
rect 25108 32662 25120 32714
rect 25172 32662 25184 32714
rect 25236 32662 30320 32714
rect 30372 32662 30384 32714
rect 30436 32662 30448 32714
rect 30500 32662 30512 32714
rect 30564 32662 35648 32714
rect 35700 32662 35712 32714
rect 35764 32662 35776 32714
rect 35828 32662 35840 32714
rect 35892 32662 40976 32714
rect 41028 32662 41040 32714
rect 41092 32662 41104 32714
rect 41156 32662 41168 32714
rect 41220 32662 46304 32714
rect 46356 32662 46368 32714
rect 46420 32662 46432 32714
rect 46484 32662 46496 32714
rect 46548 32662 51632 32714
rect 51684 32662 51696 32714
rect 51748 32662 51760 32714
rect 51812 32662 51824 32714
rect 51876 32662 56960 32714
rect 57012 32662 57024 32714
rect 57076 32662 57088 32714
rect 57140 32662 57152 32714
rect 57204 32662 62288 32714
rect 62340 32662 62352 32714
rect 62404 32662 62416 32714
rect 62468 32662 62480 32714
rect 62532 32662 67616 32714
rect 67668 32662 67680 32714
rect 67732 32662 67744 32714
rect 67796 32662 67808 32714
rect 67860 32662 72944 32714
rect 72996 32662 73008 32714
rect 73060 32662 73072 32714
rect 73124 32662 73136 32714
rect 73188 32662 78272 32714
rect 78324 32662 78336 32714
rect 78388 32662 78400 32714
rect 78452 32662 78464 32714
rect 78516 32662 83600 32714
rect 83652 32662 83664 32714
rect 83716 32662 83728 32714
rect 83780 32662 83792 32714
rect 83844 32662 88928 32714
rect 88980 32662 88992 32714
rect 89044 32662 89056 32714
rect 89108 32662 89120 32714
rect 89172 32662 93642 32714
rect 538 32640 93642 32662
rect 4051 32603 4109 32609
rect 4051 32569 4063 32603
rect 4097 32600 4109 32603
rect 5152 32600 5158 32612
rect 4097 32572 5158 32600
rect 4097 32569 4109 32572
rect 4051 32563 4109 32569
rect 5152 32560 5158 32572
rect 5210 32560 5216 32612
rect 6256 32560 6262 32612
rect 6314 32600 6320 32612
rect 16100 32600 16106 32612
rect 6314 32572 13202 32600
rect 16061 32572 16106 32600
rect 6314 32560 6320 32572
rect 4327 32535 4385 32541
rect 4327 32532 4339 32535
rect 4250 32504 4339 32532
rect 2487 32467 2545 32473
rect 2487 32433 2499 32467
rect 2533 32464 2545 32467
rect 4250 32464 4278 32504
rect 4327 32501 4339 32504
rect 4373 32532 4385 32535
rect 4692 32532 4698 32544
rect 4373 32504 4698 32532
rect 4373 32501 4385 32504
rect 4327 32495 4385 32501
rect 4692 32492 4698 32504
rect 4750 32492 4756 32544
rect 5060 32532 5066 32544
rect 5021 32504 5066 32532
rect 5060 32492 5066 32504
rect 5118 32492 5124 32544
rect 7179 32535 7237 32541
rect 7179 32501 7191 32535
rect 7225 32532 7237 32535
rect 7912 32532 7918 32544
rect 7225 32504 7918 32532
rect 7225 32501 7237 32504
rect 7179 32495 7237 32501
rect 7912 32492 7918 32504
rect 7970 32492 7976 32544
rect 2533 32436 4278 32464
rect 2533 32433 2545 32436
rect 2487 32427 2545 32433
rect 1656 32288 1662 32340
rect 1714 32328 1720 32340
rect 2502 32328 2530 32427
rect 2760 32396 2766 32408
rect 2721 32368 2766 32396
rect 2760 32356 2766 32368
rect 2818 32356 2824 32408
rect 5078 32396 5106 32492
rect 5155 32399 5213 32405
rect 5155 32396 5167 32399
rect 5078 32368 5167 32396
rect 5155 32365 5167 32368
rect 5201 32365 5213 32399
rect 5155 32359 5213 32365
rect 5247 32399 5305 32405
rect 5247 32365 5259 32399
rect 5293 32396 5305 32399
rect 6624 32396 6630 32408
rect 5293 32368 6630 32396
rect 5293 32365 5305 32368
rect 5247 32359 5305 32365
rect 6624 32356 6630 32368
rect 6682 32356 6688 32408
rect 6992 32396 6998 32408
rect 6953 32368 6998 32396
rect 6992 32356 6998 32368
rect 7050 32356 7056 32408
rect 12791 32399 12849 32405
rect 12791 32365 12803 32399
rect 12837 32365 12849 32399
rect 12791 32359 12849 32365
rect 1714 32300 2530 32328
rect 12147 32331 12205 32337
rect 1714 32288 1720 32300
rect 12147 32297 12159 32331
rect 12193 32297 12205 32331
rect 12806 32328 12834 32359
rect 12880 32356 12886 32408
rect 12938 32396 12944 32408
rect 13174 32405 13202 32572
rect 16100 32560 16106 32572
rect 16158 32560 16164 32612
rect 16468 32600 16474 32612
rect 16429 32572 16474 32600
rect 16468 32560 16474 32572
rect 16526 32560 16532 32612
rect 18768 32560 18774 32612
rect 18826 32600 18832 32612
rect 18863 32603 18921 32609
rect 18863 32600 18875 32603
rect 18826 32572 18875 32600
rect 18826 32560 18832 32572
rect 18863 32569 18875 32572
rect 18909 32569 18921 32603
rect 18863 32563 18921 32569
rect 20424 32560 20430 32612
rect 20482 32600 20488 32612
rect 21163 32603 21221 32609
rect 21163 32600 21175 32603
rect 20482 32572 21175 32600
rect 20482 32560 20488 32572
rect 21163 32569 21175 32572
rect 21209 32569 21221 32603
rect 21163 32563 21221 32569
rect 26775 32603 26833 32609
rect 26775 32569 26787 32603
rect 26821 32600 26833 32603
rect 26864 32600 26870 32612
rect 26821 32572 26870 32600
rect 26821 32569 26833 32572
rect 26775 32563 26833 32569
rect 26864 32560 26870 32572
rect 26922 32560 26928 32612
rect 32568 32560 32574 32612
rect 32626 32600 32632 32612
rect 33123 32603 33181 32609
rect 33123 32600 33135 32603
rect 32626 32572 33135 32600
rect 32626 32560 32632 32572
rect 33123 32569 33135 32572
rect 33169 32569 33181 32603
rect 33123 32563 33181 32569
rect 34503 32603 34561 32609
rect 34503 32569 34515 32603
rect 34549 32600 34561 32603
rect 35144 32600 35150 32612
rect 34549 32572 35150 32600
rect 34549 32569 34561 32572
rect 34503 32563 34561 32569
rect 35144 32560 35150 32572
rect 35202 32600 35208 32612
rect 35239 32603 35297 32609
rect 35239 32600 35251 32603
rect 35202 32572 35251 32600
rect 35202 32560 35208 32572
rect 35239 32569 35251 32572
rect 35285 32569 35297 32603
rect 35239 32563 35297 32569
rect 39928 32560 39934 32612
rect 39986 32600 39992 32612
rect 40299 32603 40357 32609
rect 40299 32600 40311 32603
rect 39986 32572 40311 32600
rect 39986 32560 39992 32572
rect 40299 32569 40311 32572
rect 40345 32569 40357 32603
rect 40299 32563 40357 32569
rect 40572 32560 40578 32612
rect 40630 32600 40636 32612
rect 43703 32603 43761 32609
rect 43703 32600 43715 32603
rect 40630 32572 43715 32600
rect 40630 32560 40636 32572
rect 43703 32569 43715 32572
rect 43749 32600 43761 32603
rect 43749 32572 44022 32600
rect 43749 32569 43761 32572
rect 43703 32563 43761 32569
rect 15548 32492 15554 32544
rect 15606 32532 15612 32544
rect 17207 32535 17265 32541
rect 17207 32532 17219 32535
rect 15606 32504 17219 32532
rect 15606 32492 15612 32504
rect 17207 32501 17219 32504
rect 17253 32501 17265 32535
rect 17207 32495 17265 32501
rect 20979 32535 21037 32541
rect 20979 32501 20991 32535
rect 21025 32532 21037 32535
rect 22080 32532 22086 32544
rect 21025 32504 22086 32532
rect 21025 32501 21037 32504
rect 20979 32495 21037 32501
rect 14723 32467 14781 32473
rect 13358 32436 14306 32464
rect 13358 32408 13386 32436
rect 14278 32408 14306 32436
rect 14723 32433 14735 32467
rect 14769 32464 14781 32467
rect 16195 32467 16253 32473
rect 16195 32464 16207 32467
rect 14769 32436 16207 32464
rect 14769 32433 14781 32436
rect 14723 32427 14781 32433
rect 16195 32433 16207 32436
rect 16241 32433 16253 32467
rect 16195 32427 16253 32433
rect 13159 32399 13217 32405
rect 12938 32368 12983 32396
rect 12938 32356 12944 32368
rect 13159 32365 13171 32399
rect 13205 32365 13217 32399
rect 13340 32396 13346 32408
rect 13301 32368 13346 32396
rect 13159 32359 13217 32365
rect 13340 32356 13346 32368
rect 13398 32356 13404 32408
rect 14168 32396 14174 32408
rect 14129 32368 14174 32396
rect 14168 32356 14174 32368
rect 14226 32356 14232 32408
rect 14260 32356 14266 32408
rect 14318 32396 14324 32408
rect 15974 32399 16032 32405
rect 14318 32368 14411 32396
rect 14318 32356 14324 32368
rect 15974 32365 15986 32399
rect 16020 32396 16032 32399
rect 16284 32396 16290 32408
rect 16020 32368 16290 32396
rect 16020 32365 16032 32368
rect 15974 32359 16032 32365
rect 16284 32356 16290 32368
rect 16342 32356 16348 32408
rect 17222 32396 17250 32495
rect 22080 32492 22086 32504
rect 22138 32492 22144 32544
rect 28796 32492 28802 32544
rect 28854 32532 28860 32544
rect 34868 32532 34874 32544
rect 28854 32504 34874 32532
rect 28854 32492 28860 32504
rect 34868 32492 34874 32504
rect 34926 32492 34932 32544
rect 35052 32492 35058 32544
rect 35110 32532 35116 32544
rect 35607 32535 35665 32541
rect 35607 32532 35619 32535
rect 35110 32504 35619 32532
rect 35110 32492 35116 32504
rect 35607 32501 35619 32504
rect 35653 32532 35665 32535
rect 38088 32532 38094 32544
rect 35653 32504 38094 32532
rect 35653 32501 35665 32504
rect 35607 32495 35665 32501
rect 38088 32492 38094 32504
rect 38146 32492 38152 32544
rect 40664 32492 40670 32544
rect 40722 32532 40728 32544
rect 43994 32541 44022 32572
rect 44160 32560 44166 32612
rect 44218 32600 44224 32612
rect 60076 32600 60082 32612
rect 44218 32572 60082 32600
rect 44218 32560 44224 32572
rect 60076 32560 60082 32572
rect 60134 32560 60140 32612
rect 64311 32603 64369 32609
rect 64311 32569 64323 32603
rect 64357 32600 64369 32603
rect 65599 32603 65657 32609
rect 65599 32600 65611 32603
rect 64357 32572 65611 32600
rect 64357 32569 64369 32572
rect 64311 32563 64369 32569
rect 65599 32569 65611 32572
rect 65645 32569 65657 32603
rect 65780 32600 65786 32612
rect 65741 32572 65786 32600
rect 65599 32563 65657 32569
rect 65780 32560 65786 32572
rect 65838 32560 65844 32612
rect 74520 32600 74526 32612
rect 65890 32572 74526 32600
rect 41219 32535 41277 32541
rect 41219 32532 41231 32535
rect 40722 32504 41231 32532
rect 40722 32492 40728 32504
rect 41219 32501 41231 32504
rect 41265 32532 41277 32535
rect 43979 32535 44037 32541
rect 41265 32504 41446 32532
rect 41265 32501 41277 32504
rect 41219 32495 41277 32501
rect 21068 32464 21074 32476
rect 21029 32436 21074 32464
rect 21068 32424 21074 32436
rect 21126 32424 21132 32476
rect 25484 32464 25490 32476
rect 25445 32436 25490 32464
rect 25484 32424 25490 32436
rect 25542 32424 25548 32476
rect 39284 32464 39290 32476
rect 38658 32436 39290 32464
rect 17480 32396 17486 32408
rect 17222 32368 17486 32396
rect 17480 32356 17486 32368
rect 17538 32356 17544 32408
rect 17759 32399 17817 32405
rect 17759 32365 17771 32399
rect 17805 32396 17817 32399
rect 18216 32396 18222 32408
rect 17805 32368 18222 32396
rect 17805 32365 17817 32368
rect 17759 32359 17817 32365
rect 18216 32356 18222 32368
rect 18274 32356 18280 32408
rect 20850 32399 20908 32405
rect 20850 32365 20862 32399
rect 20896 32396 20908 32399
rect 21344 32396 21350 32408
rect 20896 32368 21350 32396
rect 20896 32365 20908 32368
rect 20850 32359 20908 32365
rect 21344 32356 21350 32368
rect 21402 32356 21408 32408
rect 25211 32399 25269 32405
rect 25211 32396 25223 32399
rect 25042 32368 25223 32396
rect 13616 32328 13622 32340
rect 12806 32300 13622 32328
rect 12147 32291 12205 32297
rect 12162 32260 12190 32291
rect 13616 32288 13622 32300
rect 13674 32288 13680 32340
rect 15827 32331 15885 32337
rect 15827 32297 15839 32331
rect 15873 32328 15885 32331
rect 16192 32328 16198 32340
rect 15873 32300 16198 32328
rect 15873 32297 15885 32300
rect 15827 32291 15885 32297
rect 16192 32288 16198 32300
rect 16250 32288 16256 32340
rect 20703 32331 20761 32337
rect 20703 32328 20715 32331
rect 16394 32300 17618 32328
rect 16394 32260 16422 32300
rect 12162 32232 16422 32260
rect 17590 32260 17618 32300
rect 18418 32300 20715 32328
rect 18418 32260 18446 32300
rect 20703 32297 20715 32300
rect 20749 32297 20761 32331
rect 23828 32328 23834 32340
rect 20703 32291 20761 32297
rect 20810 32300 23834 32328
rect 17590 32232 18446 32260
rect 19136 32220 19142 32272
rect 19194 32260 19200 32272
rect 20810 32260 20838 32300
rect 23828 32288 23834 32300
rect 23886 32288 23892 32340
rect 19194 32232 20838 32260
rect 19194 32220 19200 32232
rect 24840 32220 24846 32272
rect 24898 32260 24904 32272
rect 25042 32269 25070 32368
rect 25211 32365 25223 32368
rect 25257 32365 25269 32399
rect 33028 32396 33034 32408
rect 32989 32368 33034 32396
rect 25211 32359 25269 32365
rect 33028 32356 33034 32368
rect 33086 32356 33092 32408
rect 34319 32399 34377 32405
rect 34319 32365 34331 32399
rect 34365 32396 34377 32399
rect 34684 32396 34690 32408
rect 34365 32368 34690 32396
rect 34365 32365 34377 32368
rect 34319 32359 34377 32365
rect 34684 32356 34690 32368
rect 34742 32356 34748 32408
rect 35144 32356 35150 32408
rect 35202 32396 35208 32408
rect 38658 32405 38686 32436
rect 39284 32424 39290 32436
rect 39342 32424 39348 32476
rect 40020 32464 40026 32476
rect 39578 32436 40026 32464
rect 35423 32399 35481 32405
rect 35423 32396 35435 32399
rect 35202 32368 35435 32396
rect 35202 32356 35208 32368
rect 35423 32365 35435 32368
rect 35469 32365 35481 32399
rect 35423 32359 35481 32365
rect 38643 32399 38701 32405
rect 38643 32365 38655 32399
rect 38689 32365 38701 32399
rect 38643 32359 38701 32365
rect 39011 32399 39069 32405
rect 39011 32365 39023 32399
rect 39057 32396 39069 32399
rect 39468 32396 39474 32408
rect 39057 32368 39474 32396
rect 39057 32365 39069 32368
rect 39011 32359 39069 32365
rect 39468 32356 39474 32368
rect 39526 32356 39532 32408
rect 26956 32288 26962 32340
rect 27014 32328 27020 32340
rect 27508 32328 27514 32340
rect 27014 32300 27514 32328
rect 27014 32288 27020 32300
rect 27508 32288 27514 32300
rect 27566 32328 27572 32340
rect 38459 32331 38517 32337
rect 27566 32300 36018 32328
rect 27566 32288 27572 32300
rect 25027 32263 25085 32269
rect 25027 32260 25039 32263
rect 24898 32232 25039 32260
rect 24898 32220 24904 32232
rect 25027 32229 25039 32232
rect 25073 32229 25085 32263
rect 25027 32223 25085 32229
rect 26312 32220 26318 32272
rect 26370 32260 26376 32272
rect 34316 32260 34322 32272
rect 26370 32232 34322 32260
rect 26370 32220 26376 32232
rect 34316 32220 34322 32232
rect 34374 32220 34380 32272
rect 35990 32260 36018 32300
rect 38459 32297 38471 32331
rect 38505 32328 38517 32331
rect 39578 32328 39606 32436
rect 40020 32424 40026 32436
rect 40078 32424 40084 32476
rect 41418 32473 41446 32504
rect 43979 32501 43991 32535
rect 44025 32532 44037 32535
rect 44436 32532 44442 32544
rect 44025 32504 44442 32532
rect 44025 32501 44037 32504
rect 43979 32495 44037 32501
rect 44436 32492 44442 32504
rect 44494 32492 44500 32544
rect 44807 32535 44865 32541
rect 44807 32501 44819 32535
rect 44853 32532 44865 32535
rect 48392 32532 48398 32544
rect 44853 32504 48398 32532
rect 44853 32501 44865 32504
rect 44807 32495 44865 32501
rect 41403 32467 41461 32473
rect 41403 32433 41415 32467
rect 41449 32433 41461 32467
rect 42320 32464 42326 32476
rect 41403 32427 41461 32433
rect 41510 32436 42326 32464
rect 40207 32399 40265 32405
rect 40207 32365 40219 32399
rect 40253 32396 40265 32399
rect 40388 32396 40394 32408
rect 40253 32368 40394 32396
rect 40253 32365 40265 32368
rect 40207 32359 40265 32365
rect 40388 32356 40394 32368
rect 40446 32396 40452 32408
rect 40664 32396 40670 32408
rect 40446 32368 40670 32396
rect 40446 32356 40452 32368
rect 40664 32356 40670 32368
rect 40722 32356 40728 32408
rect 40759 32399 40817 32405
rect 40759 32365 40771 32399
rect 40805 32396 40817 32399
rect 41510 32396 41538 32436
rect 42320 32424 42326 32436
rect 42378 32464 42384 32476
rect 44822 32464 44850 32495
rect 48392 32492 48398 32504
rect 48450 32492 48456 32544
rect 48576 32532 48582 32544
rect 48544 32504 48582 32532
rect 48576 32492 48582 32504
rect 48634 32541 48640 32544
rect 48634 32535 48692 32541
rect 48634 32501 48646 32535
rect 48680 32532 48692 32535
rect 49407 32535 49465 32541
rect 49407 32532 49419 32535
rect 48680 32504 49419 32532
rect 48680 32501 48692 32504
rect 48634 32495 48692 32501
rect 49407 32501 49419 32504
rect 49453 32532 49465 32535
rect 50600 32532 50606 32544
rect 49453 32504 50606 32532
rect 49453 32501 49465 32504
rect 49407 32495 49465 32501
rect 48634 32492 48640 32495
rect 50600 32492 50606 32504
rect 50658 32492 50664 32544
rect 52256 32492 52262 32544
rect 52314 32532 52320 32544
rect 52627 32535 52685 32541
rect 52627 32532 52639 32535
rect 52314 32504 52639 32532
rect 52314 32492 52320 32504
rect 52627 32501 52639 32504
rect 52673 32532 52685 32535
rect 53176 32532 53182 32544
rect 52673 32504 53182 32532
rect 52673 32501 52685 32504
rect 52627 32495 52685 32501
rect 53176 32492 53182 32504
rect 53234 32492 53240 32544
rect 58420 32532 58426 32544
rect 58381 32504 58426 32532
rect 58420 32492 58426 32504
rect 58478 32532 58484 32544
rect 58478 32504 58650 32532
rect 58478 32492 58484 32504
rect 47567 32467 47625 32473
rect 47567 32464 47579 32467
rect 42378 32436 44850 32464
rect 46754 32436 47579 32464
rect 42378 32424 42384 32436
rect 41676 32396 41682 32408
rect 40805 32368 41538 32396
rect 41637 32368 41682 32396
rect 40805 32365 40817 32368
rect 40759 32359 40817 32365
rect 38505 32300 39606 32328
rect 40023 32331 40081 32337
rect 38505 32297 38517 32300
rect 38459 32291 38517 32297
rect 40023 32297 40035 32331
rect 40069 32328 40081 32331
rect 40774 32328 40802 32359
rect 41676 32356 41682 32368
rect 41734 32356 41740 32408
rect 43902 32405 43930 32436
rect 46754 32408 46782 32436
rect 47567 32433 47579 32436
rect 47613 32464 47625 32467
rect 48024 32464 48030 32476
rect 47613 32436 48030 32464
rect 47613 32433 47625 32436
rect 47567 32427 47625 32433
rect 48024 32424 48030 32436
rect 48082 32424 48088 32476
rect 48852 32464 48858 32476
rect 48813 32436 48858 32464
rect 48852 32424 48858 32436
rect 48910 32424 48916 32476
rect 49680 32464 49686 32476
rect 49146 32436 49686 32464
rect 43887 32399 43945 32405
rect 43887 32365 43899 32399
rect 43933 32365 43945 32399
rect 43887 32359 43945 32365
rect 44068 32356 44074 32408
rect 44126 32396 44132 32408
rect 44163 32399 44221 32405
rect 44163 32396 44175 32399
rect 44126 32368 44175 32396
rect 44126 32356 44132 32368
rect 44163 32365 44175 32368
rect 44209 32365 44221 32399
rect 44163 32359 44221 32365
rect 44623 32399 44681 32405
rect 44623 32365 44635 32399
rect 44669 32396 44681 32399
rect 46736 32396 46742 32408
rect 44669 32368 46742 32396
rect 44669 32365 44681 32368
rect 44623 32359 44681 32365
rect 46736 32356 46742 32368
rect 46794 32356 46800 32408
rect 47012 32356 47018 32408
rect 47070 32396 47076 32408
rect 47107 32399 47165 32405
rect 47107 32396 47119 32399
rect 47070 32368 47119 32396
rect 47070 32356 47076 32368
rect 47107 32365 47119 32368
rect 47153 32365 47165 32399
rect 47107 32359 47165 32365
rect 47196 32356 47202 32408
rect 47254 32396 47260 32408
rect 47472 32396 47478 32408
rect 47254 32368 47299 32396
rect 47433 32368 47478 32396
rect 47254 32356 47260 32368
rect 47472 32356 47478 32368
rect 47530 32356 47536 32408
rect 48717 32399 48775 32405
rect 47582 32368 48622 32396
rect 40069 32300 40802 32328
rect 43059 32331 43117 32337
rect 40069 32297 40081 32300
rect 40023 32291 40081 32297
rect 43059 32297 43071 32331
rect 43105 32328 43117 32331
rect 43976 32328 43982 32340
rect 43105 32300 43982 32328
rect 43105 32297 43117 32300
rect 43059 32291 43117 32297
rect 43976 32288 43982 32300
rect 44034 32288 44040 32340
rect 46460 32328 46466 32340
rect 46421 32300 46466 32328
rect 46460 32288 46466 32300
rect 46518 32288 46524 32340
rect 47582 32328 47610 32368
rect 48392 32328 48398 32340
rect 47490 32300 47610 32328
rect 47674 32300 48398 32328
rect 47490 32260 47518 32300
rect 35990 32232 47518 32260
rect 47564 32220 47570 32272
rect 47622 32260 47628 32272
rect 47674 32260 47702 32300
rect 48392 32288 48398 32300
rect 48450 32288 48456 32340
rect 48487 32331 48545 32337
rect 48487 32297 48499 32331
rect 48533 32297 48545 32331
rect 48487 32291 48545 32297
rect 47622 32232 47702 32260
rect 47622 32220 47628 32232
rect 47748 32220 47754 32272
rect 47806 32260 47812 32272
rect 47932 32260 47938 32272
rect 47806 32232 47851 32260
rect 47893 32232 47938 32260
rect 47806 32220 47812 32232
rect 47932 32220 47938 32232
rect 47990 32220 47996 32272
rect 48024 32220 48030 32272
rect 48082 32260 48088 32272
rect 48502 32260 48530 32291
rect 48082 32232 48530 32260
rect 48594 32260 48622 32368
rect 48717 32365 48729 32399
rect 48763 32396 48775 32399
rect 49146 32396 49174 32436
rect 49680 32424 49686 32436
rect 49738 32424 49744 32476
rect 51247 32467 51305 32473
rect 51247 32433 51259 32467
rect 51293 32464 51305 32467
rect 51293 32436 52026 32464
rect 51293 32433 51305 32436
rect 51247 32427 51305 32433
rect 51998 32408 52026 32436
rect 57316 32424 57322 32476
rect 57374 32464 57380 32476
rect 58328 32464 58334 32476
rect 57374 32436 58334 32464
rect 57374 32424 57380 32436
rect 58328 32424 58334 32436
rect 58386 32424 58392 32476
rect 58622 32473 58650 32504
rect 59524 32492 59530 32544
rect 59582 32532 59588 32544
rect 59711 32535 59769 32541
rect 59711 32532 59723 32535
rect 59582 32504 59723 32532
rect 59582 32492 59588 32504
rect 59711 32501 59723 32504
rect 59757 32501 59769 32535
rect 59711 32495 59769 32501
rect 62744 32492 62750 32544
rect 62802 32532 62808 32544
rect 62802 32504 64262 32532
rect 62802 32492 62808 32504
rect 58607 32467 58665 32473
rect 58607 32433 58619 32467
rect 58653 32433 58665 32467
rect 58607 32427 58665 32433
rect 60171 32467 60229 32473
rect 60171 32433 60183 32467
rect 60217 32464 60229 32467
rect 60217 32436 63434 32464
rect 60217 32433 60229 32436
rect 60171 32427 60229 32433
rect 48763 32368 49174 32396
rect 49223 32399 49281 32405
rect 48763 32365 48775 32368
rect 48717 32359 48775 32365
rect 49223 32365 49235 32399
rect 49269 32396 49281 32399
rect 51060 32396 51066 32408
rect 49269 32368 51066 32396
rect 49269 32365 49281 32368
rect 49223 32359 49281 32365
rect 51060 32356 51066 32368
rect 51118 32356 51124 32408
rect 51520 32396 51526 32408
rect 51481 32368 51526 32396
rect 51520 32356 51526 32368
rect 51578 32356 51584 32408
rect 51980 32356 51986 32408
rect 52038 32396 52044 32408
rect 52995 32399 53053 32405
rect 52995 32396 53007 32399
rect 52038 32368 53007 32396
rect 52038 32356 52044 32368
rect 52995 32365 53007 32368
rect 53041 32365 53053 32399
rect 52995 32359 53053 32365
rect 58052 32356 58058 32408
rect 58110 32396 58116 32408
rect 58512 32396 58518 32408
rect 58110 32368 58518 32396
rect 58110 32356 58116 32368
rect 58512 32356 58518 32368
rect 58570 32396 58576 32408
rect 58791 32399 58849 32405
rect 58791 32396 58803 32399
rect 58570 32368 58803 32396
rect 58570 32356 58576 32368
rect 58791 32365 58803 32368
rect 58837 32365 58849 32399
rect 59340 32396 59346 32408
rect 59301 32368 59346 32396
rect 58791 32359 58849 32365
rect 59340 32356 59346 32368
rect 59398 32356 59404 32408
rect 59527 32399 59585 32405
rect 59527 32365 59539 32399
rect 59573 32396 59585 32399
rect 60186 32396 60214 32427
rect 63406 32408 63434 32436
rect 60352 32396 60358 32408
rect 59573 32368 60214 32396
rect 60265 32368 60358 32396
rect 59573 32365 59585 32368
rect 59527 32359 59585 32365
rect 60352 32356 60358 32368
rect 60410 32396 60416 32408
rect 61364 32396 61370 32408
rect 60410 32368 61370 32396
rect 60410 32356 60416 32368
rect 61364 32356 61370 32368
rect 61422 32396 61428 32408
rect 63296 32396 63302 32408
rect 61422 32368 63302 32396
rect 61422 32356 61428 32368
rect 63296 32356 63302 32368
rect 63354 32356 63360 32408
rect 63388 32356 63394 32408
rect 63446 32396 63452 32408
rect 63848 32396 63854 32408
rect 63446 32368 63491 32396
rect 63761 32368 63854 32396
rect 63446 32356 63452 32368
rect 63848 32356 63854 32368
rect 63906 32356 63912 32408
rect 64035 32399 64093 32405
rect 64035 32365 64047 32399
rect 64081 32396 64093 32399
rect 64234 32396 64262 32504
rect 64492 32492 64498 32544
rect 64550 32532 64556 32544
rect 65139 32535 65197 32541
rect 65139 32532 65151 32535
rect 64550 32504 65151 32532
rect 64550 32492 64556 32504
rect 65139 32501 65151 32504
rect 65185 32532 65197 32535
rect 65461 32535 65519 32541
rect 65461 32532 65473 32535
rect 65185 32504 65473 32532
rect 65185 32501 65197 32504
rect 65139 32495 65197 32501
rect 65461 32501 65473 32504
rect 65507 32501 65519 32535
rect 65890 32532 65918 32572
rect 74520 32560 74526 32572
rect 74578 32560 74584 32612
rect 76268 32560 76274 32612
rect 76326 32600 76332 32612
rect 77651 32603 77709 32609
rect 77651 32600 77663 32603
rect 76326 32572 77663 32600
rect 76326 32560 76332 32572
rect 77651 32569 77663 32572
rect 77697 32600 77709 32603
rect 83076 32600 83082 32612
rect 77697 32572 83082 32600
rect 77697 32569 77709 32572
rect 77651 32563 77709 32569
rect 83076 32560 83082 32572
rect 83134 32560 83140 32612
rect 83244 32603 83302 32609
rect 83244 32569 83256 32603
rect 83290 32600 83302 32603
rect 84272 32600 84278 32612
rect 83290 32572 84278 32600
rect 83290 32569 83302 32572
rect 83244 32563 83302 32569
rect 84272 32560 84278 32572
rect 84330 32560 84336 32612
rect 65461 32495 65519 32501
rect 65611 32504 65918 32532
rect 64676 32424 64682 32476
rect 64734 32464 64740 32476
rect 65611 32464 65639 32504
rect 65964 32492 65970 32544
rect 66022 32532 66028 32544
rect 68540 32532 68546 32544
rect 66022 32504 68546 32532
rect 66022 32492 66028 32504
rect 68540 32492 68546 32504
rect 68598 32492 68604 32544
rect 71208 32532 71214 32544
rect 70766 32504 70978 32532
rect 71169 32504 71214 32532
rect 64734 32436 65639 32464
rect 65691 32467 65749 32473
rect 64734 32424 64740 32436
rect 65691 32433 65703 32467
rect 65737 32464 65749 32467
rect 70766 32464 70794 32504
rect 65737 32436 70794 32464
rect 70843 32467 70901 32473
rect 65737 32433 65749 32436
rect 65691 32427 65749 32433
rect 70843 32433 70855 32467
rect 70889 32433 70901 32467
rect 70950 32464 70978 32504
rect 71208 32492 71214 32504
rect 71266 32492 71272 32544
rect 77191 32535 77249 32541
rect 77191 32532 77203 32535
rect 74538 32504 77203 32532
rect 74538 32464 74566 32504
rect 77191 32501 77203 32504
rect 77237 32501 77249 32535
rect 77191 32495 77249 32501
rect 81420 32492 81426 32544
rect 81478 32532 81484 32544
rect 83355 32535 83413 32541
rect 83355 32532 83367 32535
rect 81478 32504 83367 32532
rect 81478 32492 81484 32504
rect 83355 32501 83367 32504
rect 83401 32501 83413 32535
rect 83536 32532 83542 32544
rect 83497 32504 83542 32532
rect 83355 32495 83413 32501
rect 83536 32492 83542 32504
rect 83594 32492 83600 32544
rect 86023 32535 86081 32541
rect 86023 32501 86035 32535
rect 86069 32532 86081 32535
rect 86572 32532 86578 32544
rect 86069 32504 86578 32532
rect 86069 32501 86081 32504
rect 86023 32495 86081 32501
rect 86572 32492 86578 32504
rect 86630 32492 86636 32544
rect 70950 32436 74566 32464
rect 70843 32427 70901 32433
rect 64081 32368 64262 32396
rect 64081 32365 64093 32368
rect 64035 32359 64093 32365
rect 65228 32356 65234 32408
rect 65286 32396 65292 32408
rect 65964 32396 65970 32408
rect 65286 32368 65970 32396
rect 65286 32356 65292 32368
rect 65964 32356 65970 32368
rect 66022 32356 66028 32408
rect 68816 32396 68822 32408
rect 66074 32368 68822 32396
rect 63866 32328 63894 32356
rect 64584 32328 64590 32340
rect 52182 32300 58558 32328
rect 63866 32300 64590 32328
rect 52182 32260 52210 32300
rect 48594 32232 52210 32260
rect 48082 32220 48088 32232
rect 52624 32220 52630 32272
rect 52682 32260 52688 32272
rect 58420 32260 58426 32272
rect 52682 32232 58426 32260
rect 52682 32220 52688 32232
rect 58420 32220 58426 32232
rect 58478 32220 58484 32272
rect 58530 32260 58558 32300
rect 64584 32288 64590 32300
rect 64642 32328 64648 32340
rect 64771 32331 64829 32337
rect 64771 32328 64783 32331
rect 64642 32300 64783 32328
rect 64642 32288 64648 32300
rect 64771 32297 64783 32300
rect 64817 32297 64829 32331
rect 64771 32291 64829 32297
rect 65136 32288 65142 32340
rect 65194 32328 65200 32340
rect 65323 32331 65381 32337
rect 65323 32328 65335 32331
rect 65194 32300 65335 32328
rect 65194 32288 65200 32300
rect 65323 32297 65335 32300
rect 65369 32297 65381 32331
rect 65323 32291 65381 32297
rect 65412 32288 65418 32340
rect 65470 32328 65476 32340
rect 66074 32328 66102 32368
rect 68816 32356 68822 32368
rect 68874 32356 68880 32408
rect 69368 32356 69374 32408
rect 69426 32396 69432 32408
rect 69463 32399 69521 32405
rect 69463 32396 69475 32399
rect 69426 32368 69475 32396
rect 69426 32356 69432 32368
rect 69463 32365 69475 32368
rect 69509 32365 69521 32399
rect 69736 32396 69742 32408
rect 69697 32368 69742 32396
rect 69463 32359 69521 32365
rect 69736 32356 69742 32368
rect 69794 32356 69800 32408
rect 69828 32356 69834 32408
rect 69886 32396 69892 32408
rect 70858 32396 70886 32427
rect 74612 32424 74618 32476
rect 74670 32464 74676 32476
rect 75443 32467 75501 32473
rect 75443 32464 75455 32467
rect 74670 32436 75455 32464
rect 74670 32424 74676 32436
rect 75443 32433 75455 32436
rect 75489 32433 75501 32467
rect 75900 32464 75906 32476
rect 75861 32436 75906 32464
rect 75443 32427 75501 32433
rect 75900 32424 75906 32436
rect 75958 32424 75964 32476
rect 76084 32464 76090 32476
rect 76045 32436 76090 32464
rect 76084 32424 76090 32436
rect 76142 32424 76148 32476
rect 79856 32424 79862 32476
rect 79914 32464 79920 32476
rect 80871 32467 80929 32473
rect 80871 32464 80883 32467
rect 79914 32436 80883 32464
rect 79914 32424 79920 32436
rect 80871 32433 80883 32436
rect 80917 32433 80929 32467
rect 80871 32427 80929 32433
rect 82159 32467 82217 32473
rect 82159 32433 82171 32467
rect 82205 32464 82217 32467
rect 82616 32464 82622 32476
rect 82205 32436 82622 32464
rect 82205 32433 82217 32436
rect 82159 32427 82217 32433
rect 82616 32424 82622 32436
rect 82674 32424 82680 32476
rect 83447 32467 83505 32473
rect 83447 32433 83459 32467
rect 83493 32464 83505 32467
rect 89056 32464 89062 32476
rect 83493 32436 89062 32464
rect 83493 32433 83505 32436
rect 83447 32427 83505 32433
rect 89056 32424 89062 32436
rect 89114 32424 89120 32476
rect 69886 32368 70886 32396
rect 69886 32356 69892 32368
rect 71208 32356 71214 32408
rect 71266 32396 71272 32408
rect 73603 32399 73661 32405
rect 73603 32396 73615 32399
rect 71266 32368 73615 32396
rect 71266 32356 71272 32368
rect 73603 32365 73615 32368
rect 73649 32396 73661 32399
rect 73692 32396 73698 32408
rect 73649 32368 73698 32396
rect 73649 32365 73661 32368
rect 73603 32359 73661 32365
rect 73692 32356 73698 32368
rect 73750 32356 73756 32408
rect 73879 32399 73937 32405
rect 73879 32365 73891 32399
rect 73925 32396 73937 32399
rect 73968 32396 73974 32408
rect 73925 32368 73974 32396
rect 73925 32365 73937 32368
rect 73879 32359 73937 32365
rect 73968 32356 73974 32368
rect 74026 32356 74032 32408
rect 74152 32356 74158 32408
rect 74210 32396 74216 32408
rect 75348 32396 75354 32408
rect 74210 32368 75354 32396
rect 74210 32356 74216 32368
rect 75348 32356 75354 32368
rect 75406 32356 75412 32408
rect 75624 32356 75630 32408
rect 75682 32396 75688 32408
rect 76268 32396 76274 32408
rect 75682 32368 76274 32396
rect 75682 32356 75688 32368
rect 76268 32356 76274 32368
rect 76326 32356 76332 32408
rect 76636 32356 76642 32408
rect 76694 32396 76700 32408
rect 76731 32399 76789 32405
rect 76731 32396 76743 32399
rect 76694 32368 76743 32396
rect 76694 32356 76700 32368
rect 76731 32365 76743 32368
rect 76777 32365 76789 32399
rect 76731 32359 76789 32365
rect 76820 32356 76826 32408
rect 76878 32396 76884 32408
rect 76878 32368 76923 32396
rect 76878 32356 76884 32368
rect 80408 32356 80414 32408
rect 80466 32396 80472 32408
rect 81055 32399 81113 32405
rect 81055 32396 81067 32399
rect 80466 32368 81067 32396
rect 80466 32356 80472 32368
rect 81055 32365 81067 32368
rect 81101 32365 81113 32399
rect 81055 32359 81113 32365
rect 81607 32399 81665 32405
rect 81607 32365 81619 32399
rect 81653 32396 81665 32399
rect 81791 32399 81849 32405
rect 81653 32368 81742 32396
rect 81653 32365 81665 32368
rect 81607 32359 81665 32365
rect 65470 32300 66102 32328
rect 65470 32288 65476 32300
rect 66884 32288 66890 32340
rect 66942 32328 66948 32340
rect 69184 32328 69190 32340
rect 66942 32300 69190 32328
rect 66942 32288 66948 32300
rect 69184 32288 69190 32300
rect 69242 32288 69248 32340
rect 81328 32328 81334 32340
rect 74630 32300 81334 32328
rect 62100 32260 62106 32272
rect 58530 32232 62106 32260
rect 62100 32220 62106 32232
rect 62158 32220 62164 32272
rect 64676 32220 64682 32272
rect 64734 32260 64740 32272
rect 64955 32263 65013 32269
rect 64955 32260 64967 32263
rect 64734 32232 64967 32260
rect 64734 32220 64740 32232
rect 64955 32229 64967 32232
rect 65001 32229 65013 32263
rect 64955 32223 65013 32229
rect 65504 32220 65510 32272
rect 65562 32260 65568 32272
rect 74630 32260 74658 32300
rect 81328 32288 81334 32300
rect 81386 32288 81392 32340
rect 81714 32328 81742 32368
rect 81791 32365 81803 32399
rect 81837 32396 81849 32399
rect 82524 32396 82530 32408
rect 81837 32368 82530 32396
rect 81837 32365 81849 32368
rect 81791 32359 81849 32365
rect 82524 32356 82530 32368
rect 82582 32356 82588 32408
rect 82708 32356 82714 32408
rect 82766 32396 82772 32408
rect 83079 32399 83137 32405
rect 83079 32396 83091 32399
rect 82766 32368 83091 32396
rect 82766 32356 82772 32368
rect 83079 32365 83091 32368
rect 83125 32365 83137 32399
rect 83079 32359 83137 32365
rect 83628 32356 83634 32408
rect 83686 32396 83692 32408
rect 86112 32396 86118 32408
rect 83686 32368 86118 32396
rect 83686 32356 83692 32368
rect 86112 32356 86118 32368
rect 86170 32356 86176 32408
rect 87311 32399 87369 32405
rect 87311 32365 87323 32399
rect 87357 32396 87369 32399
rect 87400 32396 87406 32408
rect 87357 32368 87406 32396
rect 87357 32365 87369 32368
rect 87311 32359 87369 32365
rect 82248 32328 82254 32340
rect 81714 32300 82254 32328
rect 82248 32288 82254 32300
rect 82306 32328 82312 32340
rect 82984 32328 82990 32340
rect 82306 32300 82990 32328
rect 82306 32288 82312 32300
rect 82984 32288 82990 32300
rect 83042 32288 83048 32340
rect 83444 32288 83450 32340
rect 83502 32328 83508 32340
rect 87326 32328 87354 32359
rect 87400 32356 87406 32368
rect 87458 32396 87464 32408
rect 87495 32399 87553 32405
rect 87495 32396 87507 32399
rect 87458 32368 87507 32396
rect 87458 32356 87464 32368
rect 87495 32365 87507 32368
rect 87541 32365 87553 32399
rect 87495 32359 87553 32365
rect 87584 32356 87590 32408
rect 87642 32396 87648 32408
rect 87771 32399 87829 32405
rect 87771 32396 87783 32399
rect 87642 32368 87783 32396
rect 87642 32356 87648 32368
rect 87771 32365 87783 32368
rect 87817 32365 87829 32399
rect 87771 32359 87829 32365
rect 83502 32300 87354 32328
rect 83502 32288 83508 32300
rect 74980 32260 74986 32272
rect 65562 32232 74658 32260
rect 74941 32232 74986 32260
rect 65562 32220 65568 32232
rect 74980 32220 74986 32232
rect 75038 32220 75044 32272
rect 76912 32220 76918 32272
rect 76970 32260 76976 32272
rect 86023 32263 86081 32269
rect 86023 32260 86035 32263
rect 76970 32232 86035 32260
rect 76970 32220 76976 32232
rect 86023 32229 86035 32232
rect 86069 32260 86081 32263
rect 86207 32263 86265 32269
rect 86207 32260 86219 32263
rect 86069 32232 86219 32260
rect 86069 32229 86081 32232
rect 86023 32223 86081 32229
rect 86207 32229 86219 32232
rect 86253 32229 86265 32263
rect 86207 32223 86265 32229
rect 87492 32220 87498 32272
rect 87550 32260 87556 32272
rect 88875 32263 88933 32269
rect 88875 32260 88887 32263
rect 87550 32232 88887 32260
rect 87550 32220 87556 32232
rect 88875 32229 88887 32232
rect 88921 32229 88933 32263
rect 88875 32223 88933 32229
rect 538 32170 93642 32192
rect 538 32118 6344 32170
rect 6396 32118 6408 32170
rect 6460 32118 6472 32170
rect 6524 32118 6536 32170
rect 6588 32118 11672 32170
rect 11724 32118 11736 32170
rect 11788 32118 11800 32170
rect 11852 32118 11864 32170
rect 11916 32118 17000 32170
rect 17052 32118 17064 32170
rect 17116 32118 17128 32170
rect 17180 32118 17192 32170
rect 17244 32118 22328 32170
rect 22380 32118 22392 32170
rect 22444 32118 22456 32170
rect 22508 32118 22520 32170
rect 22572 32118 27656 32170
rect 27708 32118 27720 32170
rect 27772 32118 27784 32170
rect 27836 32118 27848 32170
rect 27900 32118 32984 32170
rect 33036 32118 33048 32170
rect 33100 32118 33112 32170
rect 33164 32118 33176 32170
rect 33228 32118 38312 32170
rect 38364 32118 38376 32170
rect 38428 32118 38440 32170
rect 38492 32118 38504 32170
rect 38556 32118 43640 32170
rect 43692 32118 43704 32170
rect 43756 32118 43768 32170
rect 43820 32118 43832 32170
rect 43884 32118 48968 32170
rect 49020 32118 49032 32170
rect 49084 32118 49096 32170
rect 49148 32118 49160 32170
rect 49212 32118 54296 32170
rect 54348 32118 54360 32170
rect 54412 32118 54424 32170
rect 54476 32118 54488 32170
rect 54540 32118 59624 32170
rect 59676 32118 59688 32170
rect 59740 32118 59752 32170
rect 59804 32118 59816 32170
rect 59868 32118 64952 32170
rect 65004 32118 65016 32170
rect 65068 32118 65080 32170
rect 65132 32118 65144 32170
rect 65196 32118 70280 32170
rect 70332 32118 70344 32170
rect 70396 32118 70408 32170
rect 70460 32118 70472 32170
rect 70524 32118 75608 32170
rect 75660 32118 75672 32170
rect 75724 32118 75736 32170
rect 75788 32118 75800 32170
rect 75852 32118 80936 32170
rect 80988 32118 81000 32170
rect 81052 32118 81064 32170
rect 81116 32118 81128 32170
rect 81180 32118 86264 32170
rect 86316 32118 86328 32170
rect 86380 32118 86392 32170
rect 86444 32118 86456 32170
rect 86508 32118 91592 32170
rect 91644 32118 91656 32170
rect 91708 32118 91720 32170
rect 91772 32118 91784 32170
rect 91836 32118 93642 32170
rect 538 32096 93642 32118
rect 5247 32059 5305 32065
rect 5247 32025 5259 32059
rect 5293 32056 5305 32059
rect 5336 32056 5342 32068
rect 5293 32028 5342 32056
rect 5293 32025 5305 32028
rect 5247 32019 5305 32025
rect 5336 32016 5342 32028
rect 5394 32056 5400 32068
rect 5983 32059 6041 32065
rect 5983 32056 5995 32059
rect 5394 32028 5995 32056
rect 5394 32016 5400 32028
rect 5983 32025 5995 32028
rect 6029 32025 6041 32059
rect 5983 32019 6041 32025
rect 4968 31880 4974 31932
rect 5026 31920 5032 31932
rect 5354 31929 5382 32016
rect 5339 31923 5397 31929
rect 5339 31920 5351 31923
rect 5026 31892 5351 31920
rect 5026 31880 5032 31892
rect 5339 31889 5351 31892
rect 5385 31889 5397 31923
rect 5998 31920 6026 32019
rect 6072 32016 6078 32068
rect 6130 32056 6136 32068
rect 12880 32056 12886 32068
rect 6130 32028 12742 32056
rect 12841 32028 12886 32056
rect 6130 32016 6136 32028
rect 6164 31948 6170 32000
rect 6222 31988 6228 32000
rect 11963 31991 12021 31997
rect 6222 31960 6670 31988
rect 6222 31948 6228 31960
rect 6642 31929 6670 31960
rect 11963 31957 11975 31991
rect 12009 31988 12021 31991
rect 12512 31988 12518 32000
rect 12009 31960 12518 31988
rect 12009 31957 12021 31960
rect 11963 31951 12021 31957
rect 12512 31948 12518 31960
rect 12570 31948 12576 32000
rect 12714 31988 12742 32028
rect 12880 32016 12886 32028
rect 12938 32016 12944 32068
rect 26312 32056 26318 32068
rect 12990 32028 26318 32056
rect 12990 31988 13018 32028
rect 26312 32016 26318 32028
rect 26370 32016 26376 32068
rect 27511 32059 27569 32065
rect 27511 32025 27523 32059
rect 27557 32056 27569 32059
rect 28612 32056 28618 32068
rect 27557 32028 28618 32056
rect 27557 32025 27569 32028
rect 27511 32019 27569 32025
rect 28612 32016 28618 32028
rect 28670 32056 28676 32068
rect 28888 32056 28894 32068
rect 28670 32028 28894 32056
rect 28670 32016 28676 32028
rect 28888 32016 28894 32028
rect 28946 32016 28952 32068
rect 36064 32016 36070 32068
rect 36122 32056 36128 32068
rect 40756 32056 40762 32068
rect 36122 32028 40762 32056
rect 36122 32016 36128 32028
rect 40756 32016 40762 32028
rect 40814 32016 40820 32068
rect 41035 32059 41093 32065
rect 41035 32025 41047 32059
rect 41081 32056 41093 32059
rect 41676 32056 41682 32068
rect 41081 32028 41682 32056
rect 41081 32025 41093 32028
rect 41035 32019 41093 32025
rect 41676 32016 41682 32028
rect 41734 32016 41740 32068
rect 46920 32016 46926 32068
rect 46978 32056 46984 32068
rect 47015 32059 47073 32065
rect 47015 32056 47027 32059
rect 46978 32028 47027 32056
rect 46978 32016 46984 32028
rect 47015 32025 47027 32028
rect 47061 32025 47073 32059
rect 82895 32059 82953 32065
rect 82895 32056 82907 32059
rect 47015 32019 47073 32025
rect 47122 32028 82907 32056
rect 12714 31960 13018 31988
rect 16008 31948 16014 32000
rect 16066 31988 16072 32000
rect 16747 31991 16805 31997
rect 16747 31988 16759 31991
rect 16066 31960 16759 31988
rect 16066 31948 16072 31960
rect 16747 31957 16759 31960
rect 16793 31988 16805 31991
rect 18216 31988 18222 32000
rect 16793 31960 16974 31988
rect 16793 31957 16805 31960
rect 16747 31951 16805 31957
rect 6351 31923 6409 31929
rect 6351 31920 6363 31923
rect 5998 31892 6363 31920
rect 5339 31883 5397 31889
rect 6351 31889 6363 31892
rect 6397 31889 6409 31923
rect 6351 31883 6409 31889
rect 6627 31923 6685 31929
rect 6627 31889 6639 31923
rect 6673 31920 6685 31923
rect 7731 31923 7789 31929
rect 7731 31920 7743 31923
rect 6673 31892 7743 31920
rect 6673 31889 6685 31892
rect 6627 31883 6685 31889
rect 7731 31889 7743 31892
rect 7777 31920 7789 31923
rect 7915 31923 7973 31929
rect 7915 31920 7927 31923
rect 7777 31892 7927 31920
rect 7777 31889 7789 31892
rect 7731 31883 7789 31889
rect 7915 31889 7927 31892
rect 7961 31889 7973 31923
rect 7915 31883 7973 31889
rect 8464 31880 8470 31932
rect 8522 31920 8528 31932
rect 11040 31920 11046 31932
rect 8522 31892 11046 31920
rect 8522 31880 8528 31892
rect 11040 31880 11046 31892
rect 11098 31880 11104 31932
rect 11224 31920 11230 31932
rect 11185 31892 11230 31920
rect 11224 31880 11230 31892
rect 11282 31880 11288 31932
rect 11500 31880 11506 31932
rect 11558 31920 11564 31932
rect 11687 31923 11745 31929
rect 11687 31920 11699 31923
rect 11558 31892 11699 31920
rect 11558 31880 11564 31892
rect 11687 31889 11699 31892
rect 11733 31889 11745 31923
rect 11687 31883 11745 31889
rect 12699 31923 12757 31929
rect 12699 31889 12711 31923
rect 12745 31920 12757 31923
rect 12791 31923 12849 31929
rect 12791 31920 12803 31923
rect 12745 31892 12803 31920
rect 12745 31889 12757 31892
rect 12699 31883 12757 31889
rect 12791 31889 12803 31892
rect 12837 31920 12849 31923
rect 13064 31920 13070 31932
rect 12837 31892 13070 31920
rect 12837 31889 12849 31892
rect 12791 31883 12849 31889
rect 13064 31880 13070 31892
rect 13122 31880 13128 31932
rect 14260 31880 14266 31932
rect 14318 31920 14324 31932
rect 16946 31929 16974 31960
rect 17682 31960 17986 31988
rect 18177 31960 18222 31988
rect 17682 31929 17710 31960
rect 14723 31923 14781 31929
rect 14723 31920 14735 31923
rect 14318 31892 14735 31920
rect 14318 31880 14324 31892
rect 14723 31889 14735 31892
rect 14769 31889 14781 31923
rect 14723 31883 14781 31889
rect 16931 31923 16989 31929
rect 16931 31889 16943 31923
rect 16977 31889 16989 31923
rect 16931 31883 16989 31889
rect 17115 31923 17173 31929
rect 17115 31889 17127 31923
rect 17161 31920 17173 31923
rect 17667 31923 17725 31929
rect 17667 31920 17679 31923
rect 17161 31892 17679 31920
rect 17161 31889 17173 31892
rect 17115 31883 17173 31889
rect 17667 31889 17679 31892
rect 17713 31889 17725 31923
rect 17848 31920 17854 31932
rect 17809 31892 17854 31920
rect 17667 31883 17725 31889
rect 17848 31880 17854 31892
rect 17906 31880 17912 31932
rect 17958 31920 17986 31960
rect 18216 31948 18222 31960
rect 18274 31948 18280 32000
rect 18495 31991 18553 31997
rect 18495 31957 18507 31991
rect 18541 31988 18553 31991
rect 18676 31988 18682 32000
rect 18541 31960 18682 31988
rect 18541 31957 18553 31960
rect 18495 31951 18553 31957
rect 18676 31948 18682 31960
rect 18734 31948 18740 32000
rect 21730 31960 22126 31988
rect 18952 31920 18958 31932
rect 17958 31892 18958 31920
rect 18952 31880 18958 31892
rect 19010 31880 19016 31932
rect 19136 31920 19142 31932
rect 19097 31892 19142 31920
rect 19136 31880 19142 31892
rect 19194 31880 19200 31932
rect 21730 31920 21758 31960
rect 19246 31892 21758 31920
rect 5431 31855 5489 31861
rect 5431 31821 5443 31855
rect 5477 31852 5489 31855
rect 6992 31852 6998 31864
rect 5477 31824 6998 31852
rect 5477 31821 5489 31824
rect 5431 31815 5489 31821
rect 6992 31812 6998 31824
rect 7050 31812 7056 31864
rect 7087 31855 7145 31861
rect 7087 31821 7099 31855
rect 7133 31821 7145 31855
rect 11242 31852 11270 31880
rect 12055 31855 12113 31861
rect 12055 31852 12067 31855
rect 11242 31824 12067 31852
rect 7087 31815 7145 31821
rect 12055 31821 12067 31824
rect 12101 31821 12113 31855
rect 12055 31815 12113 31821
rect 3496 31744 3502 31796
rect 3554 31784 3560 31796
rect 6072 31784 6078 31796
rect 3554 31756 6078 31784
rect 3554 31744 3560 31756
rect 6072 31744 6078 31756
rect 6130 31744 6136 31796
rect 6443 31787 6501 31793
rect 6443 31753 6455 31787
rect 6489 31784 6501 31787
rect 6624 31784 6630 31796
rect 6489 31756 6630 31784
rect 6489 31753 6501 31756
rect 6443 31747 6501 31753
rect 6624 31744 6630 31756
rect 6682 31744 6688 31796
rect 7102 31784 7130 31815
rect 13524 31812 13530 31864
rect 13582 31852 13588 31864
rect 17296 31852 17302 31864
rect 13582 31824 17302 31852
rect 13582 31812 13588 31824
rect 17296 31812 17302 31824
rect 17354 31812 17360 31864
rect 18124 31812 18130 31864
rect 18182 31852 18188 31864
rect 19246 31852 19274 31892
rect 21804 31880 21810 31932
rect 21862 31920 21868 31932
rect 21991 31923 22049 31929
rect 21862 31892 21907 31920
rect 21862 31880 21868 31892
rect 21991 31889 22003 31923
rect 22037 31889 22049 31923
rect 21991 31883 22049 31889
rect 18182 31824 19274 31852
rect 18182 31812 18188 31824
rect 19412 31812 19418 31864
rect 19470 31852 19476 31864
rect 21528 31852 21534 31864
rect 19470 31824 21534 31852
rect 19470 31812 19476 31824
rect 21528 31812 21534 31824
rect 21586 31812 21592 31864
rect 21715 31855 21773 31861
rect 21715 31821 21727 31855
rect 21761 31852 21773 31855
rect 22006 31852 22034 31883
rect 21761 31824 22034 31852
rect 21761 31821 21773 31824
rect 21715 31815 21773 31821
rect 7102 31756 17802 31784
rect 6164 31716 6170 31728
rect 6125 31688 6170 31716
rect 6164 31676 6170 31688
rect 6222 31676 6228 31728
rect 8007 31719 8065 31725
rect 8007 31685 8019 31719
rect 8053 31716 8065 31719
rect 8188 31716 8194 31728
rect 8053 31688 8194 31716
rect 8053 31685 8065 31688
rect 8007 31679 8065 31685
rect 8188 31676 8194 31688
rect 8246 31676 8252 31728
rect 14907 31719 14965 31725
rect 14907 31685 14919 31719
rect 14953 31716 14965 31719
rect 16100 31716 16106 31728
rect 14953 31688 16106 31716
rect 14953 31685 14965 31688
rect 14907 31679 14965 31685
rect 16100 31676 16106 31688
rect 16158 31676 16164 31728
rect 17774 31716 17802 31756
rect 17848 31744 17854 31796
rect 17906 31784 17912 31796
rect 18676 31784 18682 31796
rect 17906 31756 18682 31784
rect 17906 31744 17912 31756
rect 18676 31744 18682 31756
rect 18734 31744 18740 31796
rect 20792 31784 20798 31796
rect 19154 31756 20798 31784
rect 19154 31716 19182 31756
rect 20792 31744 20798 31756
rect 20850 31784 20856 31796
rect 21730 31784 21758 31815
rect 20850 31756 21758 31784
rect 22098 31784 22126 31960
rect 24564 31948 24570 32000
rect 24622 31988 24628 32000
rect 35328 31988 35334 32000
rect 24622 31960 35334 31988
rect 24622 31948 24628 31960
rect 35328 31948 35334 31960
rect 35386 31948 35392 32000
rect 39468 31988 39474 32000
rect 39429 31960 39474 31988
rect 39468 31948 39474 31960
rect 39526 31948 39532 32000
rect 44804 31988 44810 32000
rect 40774 31960 44810 31988
rect 23736 31880 23742 31932
rect 23794 31920 23800 31932
rect 23831 31923 23889 31929
rect 23831 31920 23843 31923
rect 23794 31892 23843 31920
rect 23794 31880 23800 31892
rect 23831 31889 23843 31892
rect 23877 31889 23889 31923
rect 23831 31883 23889 31889
rect 26131 31923 26189 31929
rect 26131 31889 26143 31923
rect 26177 31920 26189 31923
rect 26864 31920 26870 31932
rect 26177 31892 26870 31920
rect 26177 31889 26189 31892
rect 26131 31883 26189 31889
rect 26864 31880 26870 31892
rect 26922 31880 26928 31932
rect 27879 31923 27937 31929
rect 27879 31889 27891 31923
rect 27925 31920 27937 31923
rect 28152 31920 28158 31932
rect 27925 31892 28158 31920
rect 27925 31889 27937 31892
rect 27879 31883 27937 31889
rect 28152 31880 28158 31892
rect 28210 31920 28216 31932
rect 28704 31929 28710 31932
rect 28385 31923 28443 31929
rect 28385 31920 28397 31923
rect 28210 31892 28397 31920
rect 28210 31880 28216 31892
rect 28385 31889 28397 31892
rect 28431 31889 28443 31923
rect 28385 31883 28443 31889
rect 28661 31923 28710 31929
rect 28661 31889 28673 31923
rect 28707 31889 28710 31923
rect 28661 31883 28710 31889
rect 28704 31880 28710 31883
rect 28762 31880 28768 31932
rect 28888 31920 28894 31932
rect 28849 31892 28894 31920
rect 28888 31880 28894 31892
rect 28946 31880 28952 31932
rect 29259 31923 29317 31929
rect 29259 31889 29271 31923
rect 29305 31920 29317 31923
rect 29535 31923 29593 31929
rect 29535 31920 29547 31923
rect 29305 31892 29547 31920
rect 29305 31889 29317 31892
rect 29259 31883 29317 31889
rect 29535 31889 29547 31892
rect 29581 31920 29593 31923
rect 30084 31920 30090 31932
rect 29581 31892 30090 31920
rect 29581 31889 29593 31892
rect 29535 31883 29593 31889
rect 30084 31880 30090 31892
rect 30142 31880 30148 31932
rect 39560 31920 39566 31932
rect 39521 31892 39566 31920
rect 39560 31880 39566 31892
rect 39618 31880 39624 31932
rect 40774 31920 40802 31960
rect 44804 31948 44810 31960
rect 44862 31948 44868 32000
rect 47122 31988 47150 32028
rect 82895 32025 82907 32028
rect 82941 32025 82953 32059
rect 82895 32019 82953 32025
rect 47472 31988 47478 32000
rect 44914 31960 47150 31988
rect 47433 31960 47478 31988
rect 40130 31892 40802 31920
rect 22359 31855 22417 31861
rect 22359 31821 22371 31855
rect 22405 31852 22417 31855
rect 24472 31852 24478 31864
rect 22405 31824 24478 31852
rect 22405 31821 22417 31824
rect 22359 31815 22417 31821
rect 24472 31812 24478 31824
rect 24530 31812 24536 31864
rect 25852 31812 25858 31864
rect 25910 31852 25916 31864
rect 27140 31852 27146 31864
rect 25910 31824 27146 31852
rect 25910 31812 25916 31824
rect 27140 31812 27146 31824
rect 27198 31812 27204 31864
rect 27971 31855 28029 31861
rect 27971 31821 27983 31855
rect 28017 31852 28029 31855
rect 28520 31852 28526 31864
rect 28017 31824 28526 31852
rect 28017 31821 28029 31824
rect 27971 31815 28029 31821
rect 28520 31812 28526 31824
rect 28578 31812 28584 31864
rect 29164 31812 29170 31864
rect 29222 31852 29228 31864
rect 40130 31861 40158 31892
rect 40848 31880 40854 31932
rect 40906 31920 40912 31932
rect 40943 31923 41001 31929
rect 40943 31920 40955 31923
rect 40906 31892 40955 31920
rect 40906 31880 40912 31892
rect 40943 31889 40955 31892
rect 40989 31889 41001 31923
rect 40943 31883 41001 31889
rect 43516 31880 43522 31932
rect 43574 31920 43580 31932
rect 44347 31923 44405 31929
rect 44347 31920 44359 31923
rect 43574 31892 44359 31920
rect 43574 31880 43580 31892
rect 44347 31889 44359 31892
rect 44393 31920 44405 31923
rect 44531 31923 44589 31929
rect 44531 31920 44543 31923
rect 44393 31892 44543 31920
rect 44393 31889 44405 31892
rect 44347 31883 44405 31889
rect 44531 31889 44543 31892
rect 44577 31889 44589 31923
rect 44712 31920 44718 31932
rect 44673 31892 44718 31920
rect 44531 31883 44589 31889
rect 44712 31880 44718 31892
rect 44770 31880 44776 31932
rect 29351 31855 29409 31861
rect 29351 31852 29363 31855
rect 29222 31824 29363 31852
rect 29222 31812 29228 31824
rect 29351 31821 29363 31824
rect 29397 31821 29409 31855
rect 29351 31815 29409 31821
rect 39287 31855 39345 31861
rect 39287 31821 39299 31855
rect 39333 31852 39345 31855
rect 40115 31855 40173 31861
rect 40115 31852 40127 31855
rect 39333 31824 40127 31852
rect 39333 31821 39345 31824
rect 39287 31815 39345 31821
rect 40115 31821 40127 31824
rect 40161 31821 40173 31855
rect 40115 31815 40173 31821
rect 40756 31812 40762 31864
rect 40814 31852 40820 31864
rect 44914 31852 44942 31960
rect 47472 31948 47478 31960
rect 47530 31948 47536 32000
rect 58604 31988 58610 32000
rect 50894 31960 58610 31988
rect 45172 31920 45178 31932
rect 45133 31892 45178 31920
rect 45172 31880 45178 31892
rect 45230 31880 45236 31932
rect 45267 31923 45325 31929
rect 45267 31889 45279 31923
rect 45313 31920 45325 31923
rect 46092 31920 46098 31932
rect 45313 31892 46098 31920
rect 45313 31889 45325 31892
rect 45267 31883 45325 31889
rect 46092 31880 46098 31892
rect 46150 31880 46156 31932
rect 46736 31920 46742 31932
rect 46697 31892 46742 31920
rect 46736 31880 46742 31892
rect 46794 31880 46800 31932
rect 46923 31923 46981 31929
rect 46923 31889 46935 31923
rect 46969 31920 46981 31923
rect 47490 31920 47518 31948
rect 48392 31920 48398 31932
rect 46969 31892 47518 31920
rect 48353 31892 48398 31920
rect 46969 31889 46981 31892
rect 46923 31883 46981 31889
rect 48392 31880 48398 31892
rect 48450 31880 48456 31932
rect 49867 31923 49925 31929
rect 49867 31889 49879 31923
rect 49913 31920 49925 31923
rect 50784 31920 50790 31932
rect 49913 31892 50790 31920
rect 49913 31889 49925 31892
rect 49867 31883 49925 31889
rect 50784 31880 50790 31892
rect 50842 31880 50848 31932
rect 40814 31824 44942 31852
rect 45819 31855 45877 31861
rect 40814 31812 40820 31824
rect 45819 31821 45831 31855
rect 45865 31852 45877 31855
rect 47656 31852 47662 31864
rect 45865 31824 47662 31852
rect 45865 31821 45877 31824
rect 45819 31815 45877 31821
rect 47656 31812 47662 31824
rect 47714 31812 47720 31864
rect 48487 31855 48545 31861
rect 48487 31821 48499 31855
rect 48533 31852 48545 31855
rect 50143 31855 50201 31861
rect 50143 31852 50155 31855
rect 48533 31824 50155 31852
rect 48533 31821 48545 31824
rect 48487 31815 48545 31821
rect 50143 31821 50155 31824
rect 50189 31821 50201 31855
rect 50143 31815 50201 31821
rect 32476 31784 32482 31796
rect 22098 31756 32482 31784
rect 20850 31744 20856 31756
rect 32476 31744 32482 31756
rect 32534 31744 32540 31796
rect 32568 31744 32574 31796
rect 32626 31784 32632 31796
rect 32626 31756 47518 31784
rect 32626 31744 32632 31756
rect 19320 31716 19326 31728
rect 17774 31688 19182 31716
rect 19281 31688 19326 31716
rect 19320 31676 19326 31688
rect 19378 31676 19384 31728
rect 21528 31676 21534 31728
rect 21586 31716 21592 31728
rect 21804 31716 21810 31728
rect 21586 31688 21810 31716
rect 21586 31676 21592 31688
rect 21804 31676 21810 31688
rect 21862 31676 21868 31728
rect 23736 31716 23742 31728
rect 23697 31688 23742 31716
rect 23736 31676 23742 31688
rect 23794 31676 23800 31728
rect 24012 31716 24018 31728
rect 23973 31688 24018 31716
rect 24012 31676 24018 31688
rect 24070 31676 24076 31728
rect 26128 31676 26134 31728
rect 26186 31716 26192 31728
rect 26223 31719 26281 31725
rect 26223 31716 26235 31719
rect 26186 31688 26235 31716
rect 26186 31676 26192 31688
rect 26223 31685 26235 31688
rect 26269 31685 26281 31719
rect 27692 31716 27698 31728
rect 27653 31688 27698 31716
rect 26223 31679 26281 31685
rect 27692 31676 27698 31688
rect 27750 31676 27756 31728
rect 28152 31676 28158 31728
rect 28210 31716 28216 31728
rect 37536 31716 37542 31728
rect 28210 31688 37542 31716
rect 28210 31676 28216 31688
rect 37536 31676 37542 31688
rect 37594 31676 37600 31728
rect 39744 31716 39750 31728
rect 39705 31688 39750 31716
rect 39744 31676 39750 31688
rect 39802 31676 39808 31728
rect 46092 31716 46098 31728
rect 46053 31688 46098 31716
rect 46092 31676 46098 31688
rect 46150 31676 46156 31728
rect 47490 31716 47518 31756
rect 50894 31716 50922 31960
rect 58604 31948 58610 31960
rect 58662 31948 58668 32000
rect 58696 31948 58702 32000
rect 58754 31988 58760 32000
rect 58754 31960 69598 31988
rect 58754 31948 58760 31960
rect 51523 31923 51581 31929
rect 51523 31889 51535 31923
rect 51569 31920 51581 31923
rect 52903 31923 52961 31929
rect 52903 31920 52915 31923
rect 51569 31892 52915 31920
rect 51569 31889 51581 31892
rect 51523 31883 51581 31889
rect 52903 31889 52915 31892
rect 52949 31889 52961 31923
rect 52903 31883 52961 31889
rect 53636 31880 53642 31932
rect 53694 31920 53700 31932
rect 54007 31923 54065 31929
rect 54007 31920 54019 31923
rect 53694 31892 54019 31920
rect 53694 31880 53700 31892
rect 54007 31889 54019 31892
rect 54053 31889 54065 31923
rect 54007 31883 54065 31889
rect 54096 31880 54102 31932
rect 54154 31920 54160 31932
rect 57592 31920 57598 31932
rect 54154 31892 57598 31920
rect 54154 31880 54160 31892
rect 57592 31880 57598 31892
rect 57650 31880 57656 31932
rect 57779 31923 57837 31929
rect 57779 31889 57791 31923
rect 57825 31889 57837 31923
rect 57779 31883 57837 31889
rect 58239 31923 58297 31929
rect 58239 31889 58251 31923
rect 58285 31920 58297 31923
rect 59619 31923 59677 31929
rect 58285 31892 58558 31920
rect 58285 31889 58297 31892
rect 58239 31883 58297 31889
rect 51060 31812 51066 31864
rect 51118 31852 51124 31864
rect 57684 31852 57690 31864
rect 51118 31824 57690 31852
rect 51118 31812 51124 31824
rect 57684 31812 57690 31824
rect 57742 31812 57748 31864
rect 57794 31852 57822 31883
rect 58530 31864 58558 31892
rect 59619 31889 59631 31923
rect 59665 31920 59677 31923
rect 60168 31920 60174 31932
rect 59665 31892 60174 31920
rect 59665 31889 59677 31892
rect 59619 31883 59677 31889
rect 60168 31880 60174 31892
rect 60226 31880 60232 31932
rect 63575 31923 63633 31929
rect 63575 31889 63587 31923
rect 63621 31920 63633 31923
rect 68356 31920 68362 31932
rect 63621 31892 68362 31920
rect 63621 31889 63633 31892
rect 63575 31883 63633 31889
rect 68356 31880 68362 31892
rect 68414 31880 68420 31932
rect 68635 31923 68693 31929
rect 68635 31920 68647 31923
rect 68466 31892 68647 31920
rect 57794 31824 58282 31852
rect 52995 31787 53053 31793
rect 52995 31753 53007 31787
rect 53041 31784 53053 31787
rect 53912 31784 53918 31796
rect 53041 31756 53918 31784
rect 53041 31753 53053 31756
rect 52995 31747 53053 31753
rect 53912 31744 53918 31756
rect 53970 31744 53976 31796
rect 57871 31787 57929 31793
rect 57871 31753 57883 31787
rect 57917 31784 57929 31787
rect 58144 31784 58150 31796
rect 57917 31756 58150 31784
rect 57917 31753 57929 31756
rect 57871 31747 57929 31753
rect 58144 31744 58150 31756
rect 58202 31744 58208 31796
rect 58254 31784 58282 31824
rect 58328 31812 58334 31864
rect 58386 31852 58392 31864
rect 58423 31855 58481 31861
rect 58423 31852 58435 31855
rect 58386 31824 58435 31852
rect 58386 31812 58392 31824
rect 58423 31821 58435 31824
rect 58469 31821 58481 31855
rect 58423 31815 58481 31821
rect 58512 31812 58518 31864
rect 58570 31852 58576 31864
rect 63940 31852 63946 31864
rect 58570 31824 59846 31852
rect 63901 31824 63946 31852
rect 58570 31812 58576 31824
rect 59818 31793 59846 31824
rect 63940 31812 63946 31824
rect 63998 31812 64004 31864
rect 64124 31852 64130 31864
rect 64085 31824 64130 31852
rect 64124 31812 64130 31824
rect 64182 31812 64188 31864
rect 64676 31812 64682 31864
rect 64734 31852 64740 31864
rect 68466 31852 68494 31892
rect 68635 31889 68647 31892
rect 68681 31920 68693 31923
rect 69000 31920 69006 31932
rect 68681 31892 69006 31920
rect 68681 31889 68693 31892
rect 68635 31883 68693 31889
rect 69000 31880 69006 31892
rect 69058 31880 69064 31932
rect 69184 31920 69190 31932
rect 69145 31892 69190 31920
rect 69184 31880 69190 31892
rect 69242 31880 69248 31932
rect 69368 31920 69374 31932
rect 69329 31892 69374 31920
rect 69368 31880 69374 31892
rect 69426 31880 69432 31932
rect 69570 31920 69598 31960
rect 69644 31948 69650 32000
rect 69702 31988 69708 32000
rect 69702 31960 70242 31988
rect 69702 31948 69708 31960
rect 69828 31920 69834 31932
rect 69570 31892 69834 31920
rect 69828 31880 69834 31892
rect 69886 31880 69892 31932
rect 70012 31920 70018 31932
rect 69973 31892 70018 31920
rect 70012 31880 70018 31892
rect 70070 31880 70076 31932
rect 64734 31824 68494 31852
rect 68543 31855 68601 31861
rect 64734 31812 64740 31824
rect 68543 31821 68555 31855
rect 68589 31852 68601 31855
rect 68816 31852 68822 31864
rect 68589 31824 68822 31852
rect 68589 31821 68601 31824
rect 68543 31815 68601 31821
rect 68816 31812 68822 31824
rect 68874 31812 68880 31864
rect 59803 31787 59861 31793
rect 58254 31756 58834 31784
rect 58806 31728 58834 31756
rect 59803 31753 59815 31787
rect 59849 31753 59861 31787
rect 63851 31787 63909 31793
rect 63851 31784 63863 31787
rect 59803 31747 59861 31753
rect 63406 31756 63863 31784
rect 63406 31728 63434 31756
rect 63851 31753 63863 31756
rect 63897 31753 63909 31787
rect 63851 31747 63909 31753
rect 64495 31787 64553 31793
rect 64495 31753 64507 31787
rect 64541 31784 64553 31787
rect 64541 31756 68402 31784
rect 64541 31753 64553 31756
rect 64495 31747 64553 31753
rect 47490 31688 50922 31716
rect 50968 31676 50974 31728
rect 51026 31716 51032 31728
rect 51707 31719 51765 31725
rect 51707 31716 51719 31719
rect 51026 31688 51719 31716
rect 51026 31676 51032 31688
rect 51707 31685 51719 31688
rect 51753 31716 51765 31719
rect 51980 31716 51986 31728
rect 51753 31688 51986 31716
rect 51753 31685 51765 31688
rect 51707 31679 51765 31685
rect 51980 31676 51986 31688
rect 52038 31676 52044 31728
rect 52716 31676 52722 31728
rect 52774 31716 52780 31728
rect 53820 31716 53826 31728
rect 52774 31688 53826 31716
rect 52774 31676 52780 31688
rect 53820 31676 53826 31688
rect 53878 31676 53884 31728
rect 54004 31676 54010 31728
rect 54062 31716 54068 31728
rect 54099 31719 54157 31725
rect 54099 31716 54111 31719
rect 54062 31688 54111 31716
rect 54062 31676 54068 31688
rect 54099 31685 54111 31688
rect 54145 31685 54157 31719
rect 54099 31679 54157 31685
rect 54188 31676 54194 31728
rect 54246 31716 54252 31728
rect 58604 31716 58610 31728
rect 54246 31688 58610 31716
rect 54246 31676 54252 31688
rect 58604 31676 58610 31688
rect 58662 31676 58668 31728
rect 58788 31716 58794 31728
rect 58749 31688 58794 31716
rect 58788 31676 58794 31688
rect 58846 31676 58852 31728
rect 58880 31676 58886 31728
rect 58938 31716 58944 31728
rect 63204 31716 63210 31728
rect 58938 31688 63210 31716
rect 58938 31676 58944 31688
rect 63204 31676 63210 31688
rect 63262 31676 63268 31728
rect 63388 31716 63394 31728
rect 63349 31688 63394 31716
rect 63388 31676 63394 31688
rect 63446 31676 63452 31728
rect 63740 31719 63798 31725
rect 63740 31685 63752 31719
rect 63786 31716 63798 31719
rect 64510 31716 64538 31747
rect 63786 31688 64538 31716
rect 63786 31685 63798 31688
rect 63740 31679 63798 31685
rect 66884 31676 66890 31728
rect 66942 31716 66948 31728
rect 68267 31719 68325 31725
rect 68267 31716 68279 31719
rect 66942 31688 68279 31716
rect 66942 31676 66948 31688
rect 68267 31685 68279 31688
rect 68313 31685 68325 31719
rect 68374 31716 68402 31756
rect 68632 31744 68638 31796
rect 68690 31784 68696 31796
rect 69555 31787 69613 31793
rect 69555 31784 69567 31787
rect 68690 31756 69567 31784
rect 68690 31744 68696 31756
rect 69555 31753 69567 31756
rect 69601 31753 69613 31787
rect 70030 31784 70058 31880
rect 70214 31793 70242 31960
rect 74704 31948 74710 32000
rect 74762 31988 74768 32000
rect 74762 31960 75118 31988
rect 74762 31948 74768 31960
rect 71760 31920 71766 31932
rect 71721 31892 71766 31920
rect 71760 31880 71766 31892
rect 71818 31920 71824 31932
rect 72039 31923 72097 31929
rect 72039 31920 72051 31923
rect 71818 31892 72051 31920
rect 71818 31880 71824 31892
rect 72039 31889 72051 31892
rect 72085 31889 72097 31923
rect 72039 31883 72097 31889
rect 72128 31880 72134 31932
rect 72186 31920 72192 31932
rect 74244 31920 74250 31932
rect 72186 31892 74014 31920
rect 74205 31892 74250 31920
rect 72186 31880 72192 31892
rect 73986 31852 74014 31892
rect 74244 31880 74250 31892
rect 74302 31920 74308 31932
rect 74523 31923 74581 31929
rect 74523 31920 74535 31923
rect 74302 31892 74535 31920
rect 74302 31880 74308 31892
rect 74523 31889 74535 31892
rect 74569 31920 74581 31923
rect 74980 31920 74986 31932
rect 74569 31892 74986 31920
rect 74569 31889 74581 31892
rect 74523 31883 74581 31889
rect 74980 31880 74986 31892
rect 75038 31880 75044 31932
rect 75090 31920 75118 31960
rect 76820 31948 76826 32000
rect 76878 31988 76884 32000
rect 77464 31988 77470 32000
rect 76878 31960 77470 31988
rect 76878 31948 76884 31960
rect 77464 31948 77470 31960
rect 77522 31988 77528 32000
rect 78568 31988 78574 32000
rect 77522 31960 77694 31988
rect 77522 31948 77528 31960
rect 77007 31923 77065 31929
rect 77007 31920 77019 31923
rect 75090 31892 77019 31920
rect 77007 31889 77019 31892
rect 77053 31889 77065 31923
rect 77372 31920 77378 31932
rect 77333 31892 77378 31920
rect 77007 31883 77065 31889
rect 75440 31852 75446 31864
rect 73986 31824 75446 31852
rect 75440 31812 75446 31824
rect 75498 31812 75504 31864
rect 77022 31852 77050 31883
rect 77372 31880 77378 31892
rect 77430 31880 77436 31932
rect 77666 31929 77694 31960
rect 78218 31960 78574 31988
rect 78218 31929 78246 31960
rect 78568 31948 78574 31960
rect 78626 31948 78632 32000
rect 82800 31988 82806 32000
rect 82761 31960 82806 31988
rect 82800 31948 82806 31960
rect 82858 31948 82864 32000
rect 82910 31988 82938 32019
rect 83260 32016 83266 32068
rect 83318 32056 83324 32068
rect 84824 32056 84830 32068
rect 83318 32028 84830 32056
rect 83318 32016 83324 32028
rect 84824 32016 84830 32028
rect 84882 32016 84888 32068
rect 87400 32016 87406 32068
rect 87458 32056 87464 32068
rect 88139 32059 88197 32065
rect 88139 32056 88151 32059
rect 87458 32028 88151 32056
rect 87458 32016 87464 32028
rect 88139 32025 88151 32028
rect 88185 32025 88197 32059
rect 88139 32019 88197 32025
rect 82910 31960 83766 31988
rect 77651 31923 77709 31929
rect 77651 31889 77663 31923
rect 77697 31889 77709 31923
rect 77651 31883 77709 31889
rect 78203 31923 78261 31929
rect 78203 31889 78215 31923
rect 78249 31889 78261 31923
rect 78203 31883 78261 31889
rect 78387 31923 78445 31929
rect 78387 31889 78399 31923
rect 78433 31920 78445 31923
rect 79304 31920 79310 31932
rect 78433 31892 79310 31920
rect 78433 31889 78445 31892
rect 78387 31883 78445 31889
rect 79304 31880 79310 31892
rect 79362 31880 79368 31932
rect 79672 31880 79678 31932
rect 79730 31920 79736 31932
rect 80408 31920 80414 31932
rect 79730 31892 80414 31920
rect 79730 31880 79736 31892
rect 80408 31880 80414 31892
rect 80466 31880 80472 31932
rect 83260 31920 83266 31932
rect 83221 31892 83266 31920
rect 83260 31880 83266 31892
rect 83318 31880 83324 31932
rect 83355 31923 83413 31929
rect 83355 31889 83367 31923
rect 83401 31920 83413 31923
rect 83628 31920 83634 31932
rect 83401 31892 83634 31920
rect 83401 31889 83413 31892
rect 83355 31883 83413 31889
rect 83628 31880 83634 31892
rect 83686 31880 83692 31932
rect 83738 31929 83766 31960
rect 83723 31923 83781 31929
rect 83723 31889 83735 31923
rect 83769 31889 83781 31923
rect 83723 31883 83781 31889
rect 83815 31923 83873 31929
rect 83815 31889 83827 31923
rect 83861 31920 83873 31923
rect 83904 31920 83910 31932
rect 83861 31892 83910 31920
rect 83861 31889 83873 31892
rect 83815 31883 83873 31889
rect 83904 31880 83910 31892
rect 83962 31880 83968 31932
rect 88154 31920 88182 32019
rect 89056 32016 89062 32068
rect 89114 32056 89120 32068
rect 92003 32059 92061 32065
rect 92003 32056 92015 32059
rect 89114 32028 92015 32056
rect 89114 32016 89120 32028
rect 92003 32025 92015 32028
rect 92049 32025 92061 32059
rect 92003 32019 92061 32025
rect 90822 31960 91494 31988
rect 88323 31923 88381 31929
rect 88323 31920 88335 31923
rect 88154 31892 88335 31920
rect 88323 31889 88335 31892
rect 88369 31889 88381 31923
rect 88323 31883 88381 31889
rect 90436 31880 90442 31932
rect 90494 31920 90500 31932
rect 90822 31929 90850 31960
rect 90807 31923 90865 31929
rect 90807 31920 90819 31923
rect 90494 31892 90819 31920
rect 90494 31880 90500 31892
rect 90807 31889 90819 31892
rect 90853 31889 90865 31923
rect 90807 31883 90865 31889
rect 90991 31923 91049 31929
rect 90991 31889 91003 31923
rect 91037 31920 91049 31923
rect 91356 31920 91362 31932
rect 91037 31892 91362 31920
rect 91037 31889 91049 31892
rect 90991 31883 91049 31889
rect 91356 31880 91362 31892
rect 91414 31880 91420 31932
rect 91466 31929 91494 31960
rect 91451 31923 91509 31929
rect 91451 31889 91463 31923
rect 91497 31889 91509 31923
rect 91451 31883 91509 31889
rect 91540 31880 91546 31932
rect 91598 31920 91604 31932
rect 91598 31892 91643 31920
rect 91598 31880 91604 31892
rect 77467 31855 77525 31861
rect 77467 31852 77479 31855
rect 77022 31824 77479 31852
rect 77467 31821 77479 31824
rect 77513 31821 77525 31855
rect 77467 31815 77525 31821
rect 78844 31812 78850 31864
rect 78902 31852 78908 31864
rect 83444 31852 83450 31864
rect 78902 31824 83450 31852
rect 78902 31812 78908 31824
rect 83444 31812 83450 31824
rect 83502 31812 83508 31864
rect 88599 31855 88657 31861
rect 88599 31821 88611 31855
rect 88645 31852 88657 31855
rect 89700 31852 89706 31864
rect 88645 31824 89706 31852
rect 88645 31821 88657 31824
rect 88599 31815 88657 31821
rect 89700 31812 89706 31824
rect 89758 31812 89764 31864
rect 69555 31747 69613 31753
rect 69662 31756 70058 31784
rect 70199 31787 70257 31793
rect 68816 31716 68822 31728
rect 68374 31688 68822 31716
rect 68267 31679 68325 31685
rect 68816 31676 68822 31688
rect 68874 31676 68880 31728
rect 68908 31676 68914 31728
rect 68966 31716 68972 31728
rect 69662 31716 69690 31756
rect 70199 31753 70211 31787
rect 70245 31784 70257 31787
rect 84364 31784 84370 31796
rect 70245 31756 84370 31784
rect 70245 31753 70257 31756
rect 70199 31747 70257 31753
rect 84364 31744 84370 31756
rect 84422 31744 84428 31796
rect 68966 31688 69690 31716
rect 68966 31676 68972 31688
rect 69828 31676 69834 31728
rect 69886 31716 69892 31728
rect 71855 31719 71913 31725
rect 71855 31716 71867 31719
rect 69886 31688 71867 31716
rect 69886 31676 69892 31688
rect 71855 31685 71867 31688
rect 71901 31716 71913 31719
rect 73876 31716 73882 31728
rect 71901 31688 73882 31716
rect 71901 31685 71913 31688
rect 71855 31679 71913 31685
rect 73876 31676 73882 31688
rect 73934 31676 73940 31728
rect 74339 31719 74397 31725
rect 74339 31685 74351 31719
rect 74385 31716 74397 31719
rect 75348 31716 75354 31728
rect 74385 31688 75354 31716
rect 74385 31685 74397 31688
rect 74339 31679 74397 31685
rect 75348 31676 75354 31688
rect 75406 31676 75412 31728
rect 77096 31676 77102 31728
rect 77154 31716 77160 31728
rect 77191 31719 77249 31725
rect 77191 31716 77203 31719
rect 77154 31688 77203 31716
rect 77154 31676 77160 31688
rect 77191 31685 77203 31688
rect 77237 31685 77249 31719
rect 78660 31716 78666 31728
rect 78621 31688 78666 31716
rect 77191 31679 77249 31685
rect 78660 31676 78666 31688
rect 78718 31676 78724 31728
rect 80592 31716 80598 31728
rect 80553 31688 80598 31716
rect 80592 31676 80598 31688
rect 80650 31676 80656 31728
rect 84272 31716 84278 31728
rect 84233 31688 84278 31716
rect 84272 31676 84278 31688
rect 84330 31676 84336 31728
rect 88320 31676 88326 31728
rect 88378 31716 88384 31728
rect 89703 31719 89761 31725
rect 89703 31716 89715 31719
rect 88378 31688 89715 31716
rect 88378 31676 88384 31688
rect 89703 31685 89715 31688
rect 89749 31685 89761 31719
rect 89703 31679 89761 31685
rect 538 31626 93642 31648
rect 538 31574 3680 31626
rect 3732 31574 3744 31626
rect 3796 31574 3808 31626
rect 3860 31574 3872 31626
rect 3924 31574 9008 31626
rect 9060 31574 9072 31626
rect 9124 31574 9136 31626
rect 9188 31574 9200 31626
rect 9252 31574 14336 31626
rect 14388 31574 14400 31626
rect 14452 31574 14464 31626
rect 14516 31574 14528 31626
rect 14580 31574 19664 31626
rect 19716 31574 19728 31626
rect 19780 31574 19792 31626
rect 19844 31574 19856 31626
rect 19908 31574 24992 31626
rect 25044 31574 25056 31626
rect 25108 31574 25120 31626
rect 25172 31574 25184 31626
rect 25236 31574 30320 31626
rect 30372 31574 30384 31626
rect 30436 31574 30448 31626
rect 30500 31574 30512 31626
rect 30564 31574 35648 31626
rect 35700 31574 35712 31626
rect 35764 31574 35776 31626
rect 35828 31574 35840 31626
rect 35892 31574 40976 31626
rect 41028 31574 41040 31626
rect 41092 31574 41104 31626
rect 41156 31574 41168 31626
rect 41220 31574 46304 31626
rect 46356 31574 46368 31626
rect 46420 31574 46432 31626
rect 46484 31574 46496 31626
rect 46548 31574 51632 31626
rect 51684 31574 51696 31626
rect 51748 31574 51760 31626
rect 51812 31574 51824 31626
rect 51876 31574 56960 31626
rect 57012 31574 57024 31626
rect 57076 31574 57088 31626
rect 57140 31574 57152 31626
rect 57204 31574 62288 31626
rect 62340 31574 62352 31626
rect 62404 31574 62416 31626
rect 62468 31574 62480 31626
rect 62532 31574 67616 31626
rect 67668 31574 67680 31626
rect 67732 31574 67744 31626
rect 67796 31574 67808 31626
rect 67860 31574 72944 31626
rect 72996 31574 73008 31626
rect 73060 31574 73072 31626
rect 73124 31574 73136 31626
rect 73188 31574 78272 31626
rect 78324 31574 78336 31626
rect 78388 31574 78400 31626
rect 78452 31574 78464 31626
rect 78516 31574 83600 31626
rect 83652 31574 83664 31626
rect 83716 31574 83728 31626
rect 83780 31574 83792 31626
rect 83844 31574 88928 31626
rect 88980 31574 88992 31626
rect 89044 31574 89056 31626
rect 89108 31574 89120 31626
rect 89172 31574 93642 31626
rect 538 31552 93642 31574
rect 828 31472 834 31524
rect 886 31512 892 31524
rect 886 31484 2714 31512
rect 886 31472 892 31484
rect 2686 31444 2714 31484
rect 2760 31472 2766 31524
rect 2818 31512 2824 31524
rect 3039 31515 3097 31521
rect 3039 31512 3051 31515
rect 2818 31484 3051 31512
rect 2818 31472 2824 31484
rect 3039 31481 3051 31484
rect 3085 31481 3097 31515
rect 3496 31512 3502 31524
rect 3457 31484 3502 31512
rect 3039 31475 3097 31481
rect 3496 31472 3502 31484
rect 3554 31472 3560 31524
rect 5152 31472 5158 31524
rect 5210 31512 5216 31524
rect 5983 31515 6041 31521
rect 5983 31512 5995 31515
rect 5210 31484 5995 31512
rect 5210 31472 5216 31484
rect 5983 31481 5995 31484
rect 6029 31512 6041 31515
rect 6440 31512 6446 31524
rect 6029 31484 6446 31512
rect 6029 31481 6041 31484
rect 5983 31475 6041 31481
rect 6440 31472 6446 31484
rect 6498 31472 6504 31524
rect 11040 31472 11046 31524
rect 11098 31512 11104 31524
rect 15275 31515 15333 31521
rect 15275 31512 15287 31515
rect 11098 31484 15287 31512
rect 11098 31472 11104 31484
rect 15275 31481 15287 31484
rect 15321 31481 15333 31515
rect 15275 31475 15333 31481
rect 15643 31515 15701 31521
rect 15643 31481 15655 31515
rect 15689 31512 15701 31515
rect 19136 31512 19142 31524
rect 15689 31484 19142 31512
rect 15689 31481 15701 31484
rect 15643 31475 15701 31481
rect 19136 31472 19142 31484
rect 19194 31472 19200 31524
rect 22080 31512 22086 31524
rect 22041 31484 22086 31512
rect 22080 31472 22086 31484
rect 22138 31472 22144 31524
rect 24564 31512 24570 31524
rect 24525 31484 24570 31512
rect 24564 31472 24570 31484
rect 24622 31472 24628 31524
rect 31835 31515 31893 31521
rect 31835 31512 31847 31515
rect 26238 31484 31847 31512
rect 4971 31447 5029 31453
rect 4971 31444 4983 31447
rect 2686 31416 4983 31444
rect 4971 31413 4983 31416
rect 5017 31444 5029 31447
rect 6164 31444 6170 31456
rect 5017 31416 6170 31444
rect 5017 31413 5029 31416
rect 4971 31407 5029 31413
rect 1656 31376 1662 31388
rect 1617 31348 1662 31376
rect 1656 31336 1662 31348
rect 1714 31336 1720 31388
rect 1935 31379 1993 31385
rect 1935 31345 1947 31379
rect 1981 31376 1993 31379
rect 3496 31376 3502 31388
rect 1981 31348 3502 31376
rect 1981 31345 1993 31348
rect 1935 31339 1993 31345
rect 3496 31336 3502 31348
rect 3554 31336 3560 31388
rect 1674 31308 1702 31336
rect 3591 31311 3649 31317
rect 3591 31308 3603 31311
rect 1674 31280 3603 31308
rect 3591 31277 3603 31280
rect 3637 31277 3649 31311
rect 4986 31308 5014 31407
rect 6164 31404 6170 31416
rect 6222 31404 6228 31456
rect 25852 31444 25858 31456
rect 6274 31416 25858 31444
rect 5063 31311 5121 31317
rect 5063 31308 5075 31311
rect 4986 31280 5075 31308
rect 3591 31271 3649 31277
rect 5063 31277 5075 31280
rect 5109 31277 5121 31311
rect 6274 31308 6302 31416
rect 25852 31404 25858 31416
rect 25910 31404 25916 31456
rect 6992 31376 6998 31388
rect 6366 31348 6998 31376
rect 6366 31317 6394 31348
rect 6992 31336 6998 31348
rect 7050 31336 7056 31388
rect 12328 31336 12334 31388
rect 12386 31376 12392 31388
rect 12975 31379 13033 31385
rect 12386 31348 12558 31376
rect 12386 31336 12392 31348
rect 5063 31271 5121 31277
rect 5170 31280 6302 31308
rect 6351 31311 6409 31317
rect 4876 31200 4882 31252
rect 4934 31240 4940 31252
rect 5170 31240 5198 31280
rect 6351 31277 6363 31311
rect 6397 31277 6409 31311
rect 6351 31271 6409 31277
rect 6440 31268 6446 31320
rect 6498 31308 6504 31320
rect 6627 31311 6685 31317
rect 6498 31280 6543 31308
rect 6498 31268 6504 31280
rect 6627 31277 6639 31311
rect 6673 31277 6685 31311
rect 6627 31271 6685 31277
rect 6642 31240 6670 31271
rect 6716 31268 6722 31320
rect 6774 31308 6780 31320
rect 7915 31311 7973 31317
rect 7915 31308 7927 31311
rect 6774 31280 7927 31308
rect 6774 31268 6780 31280
rect 7915 31277 7927 31280
rect 7961 31277 7973 31311
rect 7915 31271 7973 31277
rect 9292 31268 9298 31320
rect 9350 31308 9356 31320
rect 10491 31311 10549 31317
rect 10491 31308 10503 31311
rect 9350 31280 10503 31308
rect 9350 31268 9356 31280
rect 10491 31277 10503 31280
rect 10537 31277 10549 31311
rect 12420 31308 12426 31320
rect 12381 31280 12426 31308
rect 10491 31271 10549 31277
rect 12420 31268 12426 31280
rect 12478 31268 12484 31320
rect 12530 31317 12558 31348
rect 12975 31345 12987 31379
rect 13021 31376 13033 31379
rect 13340 31376 13346 31388
rect 13021 31348 13346 31376
rect 13021 31345 13033 31348
rect 12975 31339 13033 31345
rect 13340 31336 13346 31348
rect 13398 31336 13404 31388
rect 15275 31379 15333 31385
rect 15275 31345 15287 31379
rect 15321 31376 15333 31379
rect 15321 31348 15594 31376
rect 15321 31345 15333 31348
rect 15275 31339 15333 31345
rect 12515 31311 12573 31317
rect 12515 31277 12527 31311
rect 12561 31277 12573 31311
rect 15459 31311 15517 31317
rect 15459 31308 15471 31311
rect 12515 31271 12573 31277
rect 12898 31280 15471 31308
rect 6808 31240 6814 31252
rect 4934 31212 5198 31240
rect 5262 31212 6814 31240
rect 4934 31200 4940 31212
rect 5262 31181 5290 31212
rect 6808 31200 6814 31212
rect 6866 31200 6872 31252
rect 7087 31243 7145 31249
rect 7087 31209 7099 31243
rect 7133 31240 7145 31243
rect 12898 31240 12926 31280
rect 15459 31277 15471 31280
rect 15505 31277 15517 31311
rect 15566 31308 15594 31348
rect 16652 31336 16658 31388
rect 16710 31376 16716 31388
rect 17207 31379 17265 31385
rect 17207 31376 17219 31379
rect 16710 31348 17219 31376
rect 16710 31336 16716 31348
rect 17207 31345 17219 31348
rect 17253 31376 17265 31379
rect 17483 31379 17541 31385
rect 17483 31376 17495 31379
rect 17253 31348 17495 31376
rect 17253 31345 17265 31348
rect 17207 31339 17265 31345
rect 17483 31345 17495 31348
rect 17529 31345 17541 31379
rect 17483 31339 17541 31345
rect 18860 31336 18866 31388
rect 18918 31376 18924 31388
rect 23923 31379 23981 31385
rect 18918 31348 19734 31376
rect 18918 31336 18924 31348
rect 17667 31311 17725 31317
rect 15566 31280 16698 31308
rect 15459 31271 15517 31277
rect 7133 31212 12926 31240
rect 7133 31209 7145 31212
rect 7087 31203 7145 31209
rect 13064 31200 13070 31252
rect 13122 31240 13128 31252
rect 16670 31240 16698 31280
rect 17667 31277 17679 31311
rect 17713 31308 17725 31311
rect 17756 31308 17762 31320
rect 17713 31280 17762 31308
rect 17713 31277 17725 31280
rect 17667 31271 17725 31277
rect 17756 31268 17762 31280
rect 17814 31308 17820 31320
rect 18219 31311 18277 31317
rect 18219 31308 18231 31311
rect 17814 31280 18231 31308
rect 17814 31268 17820 31280
rect 18219 31277 18231 31280
rect 18265 31277 18277 31311
rect 18219 31271 18277 31277
rect 18403 31311 18461 31317
rect 18403 31277 18415 31311
rect 18449 31308 18461 31311
rect 18952 31308 18958 31320
rect 18449 31280 18958 31308
rect 18449 31277 18461 31280
rect 18403 31271 18461 31277
rect 18952 31268 18958 31280
rect 19010 31268 19016 31320
rect 19706 31317 19734 31348
rect 23923 31345 23935 31379
rect 23969 31376 23981 31379
rect 26128 31376 26134 31388
rect 23969 31348 26134 31376
rect 23969 31345 23981 31348
rect 23923 31339 23981 31345
rect 26128 31336 26134 31348
rect 26186 31336 26192 31388
rect 19691 31311 19749 31317
rect 19691 31277 19703 31311
rect 19737 31277 19749 31311
rect 19691 31271 19749 31277
rect 21991 31311 22049 31317
rect 21991 31277 22003 31311
rect 22037 31308 22049 31311
rect 23187 31311 23245 31317
rect 23187 31308 23199 31311
rect 22037 31280 23199 31308
rect 22037 31277 22049 31280
rect 21991 31271 22049 31277
rect 23187 31277 23199 31280
rect 23233 31277 23245 31311
rect 23187 31271 23245 31277
rect 23276 31268 23282 31320
rect 23334 31308 23340 31320
rect 23828 31308 23834 31320
rect 23334 31280 23834 31308
rect 23334 31268 23340 31280
rect 23828 31268 23834 31280
rect 23886 31268 23892 31320
rect 24104 31268 24110 31320
rect 24162 31308 24168 31320
rect 24199 31311 24257 31317
rect 24199 31308 24211 31311
rect 24162 31280 24211 31308
rect 24162 31268 24168 31280
rect 24199 31277 24211 31280
rect 24245 31277 24257 31311
rect 24199 31271 24257 31277
rect 24383 31311 24441 31317
rect 24383 31277 24395 31311
rect 24429 31308 24441 31311
rect 24564 31308 24570 31320
rect 24429 31280 24570 31308
rect 24429 31277 24441 31280
rect 24383 31271 24441 31277
rect 24564 31268 24570 31280
rect 24622 31268 24628 31320
rect 20700 31240 20706 31252
rect 13122 31212 16606 31240
rect 16670 31212 20706 31240
rect 13122 31200 13128 31212
rect 5247 31175 5305 31181
rect 5247 31141 5259 31175
rect 5293 31141 5305 31175
rect 8096 31172 8102 31184
rect 8057 31144 8102 31172
rect 5247 31135 5305 31141
rect 8096 31132 8102 31144
rect 8154 31132 8160 31184
rect 10675 31175 10733 31181
rect 10675 31141 10687 31175
rect 10721 31172 10733 31175
rect 12144 31172 12150 31184
rect 10721 31144 12150 31172
rect 10721 31141 10733 31144
rect 10675 31135 10733 31141
rect 12144 31132 12150 31144
rect 12202 31172 12208 31184
rect 13082 31172 13110 31200
rect 12202 31144 13110 31172
rect 16578 31172 16606 31212
rect 20700 31200 20706 31212
rect 20758 31240 20764 31252
rect 26238 31240 26266 31484
rect 31835 31481 31847 31484
rect 31881 31512 31893 31515
rect 32292 31512 32298 31524
rect 31881 31484 32298 31512
rect 31881 31481 31893 31484
rect 31835 31475 31893 31481
rect 32292 31472 32298 31484
rect 32350 31472 32356 31524
rect 32476 31472 32482 31524
rect 32534 31512 32540 31524
rect 39836 31512 39842 31524
rect 32534 31484 39842 31512
rect 32534 31472 32540 31484
rect 39836 31472 39842 31484
rect 39894 31472 39900 31524
rect 40020 31512 40026 31524
rect 39981 31484 40026 31512
rect 40020 31472 40026 31484
rect 40078 31472 40084 31524
rect 47012 31512 47018 31524
rect 46973 31484 47018 31512
rect 47012 31472 47018 31484
rect 47070 31472 47076 31524
rect 51520 31472 51526 31524
rect 51578 31512 51584 31524
rect 51615 31515 51673 31521
rect 51615 31512 51627 31515
rect 51578 31484 51627 31512
rect 51578 31472 51584 31484
rect 51615 31481 51627 31484
rect 51661 31481 51673 31515
rect 51615 31475 51673 31481
rect 52075 31515 52133 31521
rect 52075 31481 52087 31515
rect 52121 31512 52133 31515
rect 54096 31512 54102 31524
rect 52121 31484 54102 31512
rect 52121 31481 52133 31484
rect 52075 31475 52133 31481
rect 26867 31447 26925 31453
rect 26867 31413 26879 31447
rect 26913 31444 26925 31447
rect 26956 31444 26962 31456
rect 26913 31416 26962 31444
rect 26913 31413 26925 31416
rect 26867 31407 26925 31413
rect 26499 31311 26557 31317
rect 26499 31277 26511 31311
rect 26545 31308 26557 31311
rect 26882 31308 26910 31407
rect 26956 31404 26962 31416
rect 27014 31404 27020 31456
rect 27692 31404 27698 31456
rect 27750 31444 27756 31456
rect 28152 31444 28158 31456
rect 27750 31416 28158 31444
rect 27750 31404 27756 31416
rect 28152 31404 28158 31416
rect 28210 31444 28216 31456
rect 28428 31444 28434 31456
rect 28210 31416 28434 31444
rect 28210 31404 28216 31416
rect 28428 31404 28434 31416
rect 28486 31404 28492 31456
rect 30084 31444 30090 31456
rect 30045 31416 30090 31444
rect 30084 31404 30090 31416
rect 30142 31404 30148 31456
rect 44436 31404 44442 31456
rect 44494 31444 44500 31456
rect 44712 31444 44718 31456
rect 44494 31416 44718 31444
rect 44494 31404 44500 31416
rect 44712 31404 44718 31416
rect 44770 31444 44776 31456
rect 50876 31444 50882 31456
rect 44770 31416 50882 31444
rect 44770 31404 44776 31416
rect 50876 31404 50882 31416
rect 50934 31404 50940 31456
rect 51155 31447 51213 31453
rect 51155 31413 51167 31447
rect 51201 31444 51213 31447
rect 52090 31444 52118 31475
rect 54096 31472 54102 31484
rect 54154 31472 54160 31524
rect 63388 31512 63394 31524
rect 54206 31484 63394 31512
rect 51201 31416 52118 31444
rect 51201 31413 51213 31416
rect 51155 31407 51213 31413
rect 28520 31376 28526 31388
rect 26545 31280 26910 31308
rect 27066 31348 28526 31376
rect 26545 31277 26557 31280
rect 26499 31271 26557 31277
rect 20758 31212 26266 31240
rect 26591 31243 26649 31249
rect 20758 31200 20764 31212
rect 26591 31209 26603 31243
rect 26637 31240 26649 31243
rect 26772 31240 26778 31252
rect 26637 31212 26778 31240
rect 26637 31209 26649 31212
rect 26591 31203 26649 31209
rect 26772 31200 26778 31212
rect 26830 31240 26836 31252
rect 27066 31240 27094 31348
rect 28520 31336 28526 31348
rect 28578 31336 28584 31388
rect 28980 31376 28986 31388
rect 28941 31348 28986 31376
rect 28980 31336 28986 31348
rect 29038 31336 29044 31388
rect 46460 31376 46466 31388
rect 34242 31348 35926 31376
rect 28707 31311 28765 31317
rect 28707 31277 28719 31311
rect 28753 31277 28765 31311
rect 28707 31271 28765 31277
rect 26830 31212 27094 31240
rect 26830 31200 26836 31212
rect 18124 31172 18130 31184
rect 16578 31144 18130 31172
rect 12202 31132 12208 31144
rect 18124 31132 18130 31144
rect 18182 31132 18188 31184
rect 18676 31172 18682 31184
rect 18637 31144 18682 31172
rect 18676 31132 18682 31144
rect 18734 31132 18740 31184
rect 18952 31172 18958 31184
rect 18913 31144 18958 31172
rect 18952 31132 18958 31144
rect 19010 31132 19016 31184
rect 19872 31172 19878 31184
rect 19833 31144 19878 31172
rect 19872 31132 19878 31144
rect 19930 31132 19936 31184
rect 22908 31172 22914 31184
rect 22869 31144 22914 31172
rect 22908 31132 22914 31144
rect 22966 31172 22972 31184
rect 24104 31172 24110 31184
rect 22966 31144 24110 31172
rect 22966 31132 22972 31144
rect 24104 31132 24110 31144
rect 24162 31132 24168 31184
rect 28722 31172 28750 31271
rect 31464 31268 31470 31320
rect 31522 31308 31528 31320
rect 32200 31308 32206 31320
rect 31522 31280 32206 31308
rect 31522 31268 31528 31280
rect 32200 31268 32206 31280
rect 32258 31268 32264 31320
rect 32292 31268 32298 31320
rect 32350 31308 32356 31320
rect 32350 31280 32395 31308
rect 32350 31268 32356 31280
rect 32660 31268 32666 31320
rect 32718 31308 32724 31320
rect 32801 31311 32859 31317
rect 32801 31308 32813 31311
rect 32718 31280 32813 31308
rect 32718 31268 32724 31280
rect 32801 31277 32813 31280
rect 32847 31277 32859 31311
rect 32801 31271 32859 31277
rect 32939 31311 32997 31317
rect 32939 31277 32951 31311
rect 32985 31277 32997 31311
rect 32939 31271 32997 31277
rect 32954 31240 32982 31271
rect 33120 31240 33126 31252
rect 32954 31212 33126 31240
rect 33120 31200 33126 31212
rect 33178 31200 33184 31252
rect 33304 31240 33310 31252
rect 33265 31212 33310 31240
rect 33304 31200 33310 31212
rect 33362 31200 33368 31252
rect 34242 31240 34270 31348
rect 35898 31317 35926 31348
rect 46294 31348 46466 31376
rect 35699 31311 35757 31317
rect 35699 31308 35711 31311
rect 33414 31212 34270 31240
rect 35530 31280 35711 31308
rect 28796 31172 28802 31184
rect 28709 31144 28802 31172
rect 28796 31132 28802 31144
rect 28854 31172 28860 31184
rect 29256 31172 29262 31184
rect 28854 31144 29262 31172
rect 28854 31132 28860 31144
rect 29256 31132 29262 31144
rect 29314 31172 29320 31184
rect 30455 31175 30513 31181
rect 30455 31172 30467 31175
rect 29314 31144 30467 31172
rect 29314 31132 29320 31144
rect 30455 31141 30467 31144
rect 30501 31141 30513 31175
rect 30455 31135 30513 31141
rect 32200 31132 32206 31184
rect 32258 31172 32264 31184
rect 32660 31172 32666 31184
rect 32258 31144 32666 31172
rect 32258 31132 32264 31144
rect 32660 31132 32666 31144
rect 32718 31172 32724 31184
rect 33414 31172 33442 31212
rect 32718 31144 33442 31172
rect 32718 31132 32724 31144
rect 33488 31132 33494 31184
rect 33546 31172 33552 31184
rect 33583 31175 33641 31181
rect 33583 31172 33595 31175
rect 33546 31144 33595 31172
rect 33546 31132 33552 31144
rect 33583 31141 33595 31144
rect 33629 31172 33641 31175
rect 34408 31172 34414 31184
rect 33629 31144 34414 31172
rect 33629 31141 33641 31144
rect 33583 31135 33641 31141
rect 34408 31132 34414 31144
rect 34466 31132 34472 31184
rect 35420 31132 35426 31184
rect 35478 31172 35484 31184
rect 35530 31181 35558 31280
rect 35699 31277 35711 31280
rect 35745 31277 35757 31311
rect 35699 31271 35757 31277
rect 35883 31311 35941 31317
rect 35883 31277 35895 31311
rect 35929 31308 35941 31311
rect 36435 31311 36493 31317
rect 36435 31308 36447 31311
rect 35929 31280 36447 31308
rect 35929 31277 35941 31280
rect 35883 31271 35941 31277
rect 36435 31277 36447 31280
rect 36481 31277 36493 31311
rect 36435 31271 36493 31277
rect 36619 31311 36677 31317
rect 36619 31277 36631 31311
rect 36665 31308 36677 31311
rect 37352 31308 37358 31320
rect 36665 31280 37358 31308
rect 36665 31277 36677 31280
rect 36619 31271 36677 31277
rect 37352 31268 37358 31280
rect 37410 31268 37416 31320
rect 39928 31308 39934 31320
rect 39889 31280 39934 31308
rect 39928 31268 39934 31280
rect 39986 31268 39992 31320
rect 40848 31268 40854 31320
rect 40906 31308 40912 31320
rect 46294 31308 46322 31348
rect 46460 31336 46466 31348
rect 46518 31336 46524 31388
rect 48852 31336 48858 31388
rect 48910 31376 48916 31388
rect 54206 31376 54234 31484
rect 63388 31472 63394 31484
rect 63446 31472 63452 31524
rect 68632 31512 68638 31524
rect 68593 31484 68638 31512
rect 68632 31472 68638 31484
rect 68690 31472 68696 31524
rect 69003 31515 69061 31521
rect 69003 31512 69015 31515
rect 68742 31484 69015 31512
rect 54280 31404 54286 31456
rect 54338 31453 54344 31456
rect 54338 31447 54387 31453
rect 54338 31413 54341 31447
rect 54375 31413 54387 31447
rect 54338 31407 54387 31413
rect 54467 31447 54525 31453
rect 54467 31413 54479 31447
rect 54513 31413 54525 31447
rect 54467 31407 54525 31413
rect 54338 31404 54344 31407
rect 54482 31376 54510 31407
rect 54648 31404 54654 31456
rect 54706 31404 54712 31456
rect 62008 31404 62014 31456
rect 62066 31444 62072 31456
rect 62839 31447 62897 31453
rect 62839 31444 62851 31447
rect 62066 31416 62851 31444
rect 62066 31404 62072 31416
rect 62839 31413 62851 31416
rect 62885 31413 62897 31447
rect 67896 31444 67902 31456
rect 62839 31407 62897 31413
rect 63130 31416 67902 31444
rect 48910 31348 54234 31376
rect 54298 31348 54510 31376
rect 54556 31379 54614 31385
rect 48910 31336 48916 31348
rect 46920 31308 46926 31320
rect 40906 31280 46322 31308
rect 46881 31280 46926 31308
rect 40906 31268 40912 31280
rect 46920 31268 46926 31280
rect 46978 31268 46984 31320
rect 51428 31308 51434 31320
rect 51389 31280 51434 31308
rect 51428 31268 51434 31280
rect 51486 31268 51492 31320
rect 52995 31311 53053 31317
rect 52995 31277 53007 31311
rect 53041 31308 53053 31311
rect 53636 31308 53642 31320
rect 53041 31280 53642 31308
rect 53041 31277 53053 31280
rect 52995 31271 53053 31277
rect 53636 31268 53642 31280
rect 53694 31268 53700 31320
rect 54004 31268 54010 31320
rect 54062 31308 54068 31320
rect 54298 31308 54326 31348
rect 54556 31345 54568 31379
rect 54602 31376 54614 31379
rect 54666 31376 54694 31404
rect 54602 31348 54694 31376
rect 54602 31345 54614 31348
rect 54556 31339 54614 31345
rect 54740 31336 54746 31388
rect 54798 31376 54804 31388
rect 54798 31348 58558 31376
rect 54798 31336 54804 31348
rect 57500 31308 57506 31320
rect 54062 31280 54326 31308
rect 54574 31280 57506 31308
rect 54062 31268 54068 31280
rect 36984 31240 36990 31252
rect 36945 31212 36990 31240
rect 36984 31200 36990 31212
rect 37042 31200 37048 31252
rect 51060 31200 51066 31252
rect 51118 31240 51124 31252
rect 51339 31243 51397 31249
rect 51339 31240 51351 31243
rect 51118 31212 51351 31240
rect 51118 31200 51124 31212
rect 51339 31209 51351 31212
rect 51385 31209 51397 31243
rect 51339 31203 51397 31209
rect 54191 31243 54249 31249
rect 54191 31209 54203 31243
rect 54237 31240 54249 31243
rect 54574 31240 54602 31280
rect 57500 31268 57506 31280
rect 57558 31268 57564 31320
rect 57595 31311 57653 31317
rect 57595 31277 57607 31311
rect 57641 31277 57653 31311
rect 57868 31308 57874 31320
rect 57829 31280 57874 31308
rect 57595 31271 57653 31277
rect 54237 31212 54602 31240
rect 54237 31209 54249 31212
rect 54191 31203 54249 31209
rect 54648 31200 54654 31252
rect 54706 31240 54712 31252
rect 55019 31243 55077 31249
rect 55019 31240 55031 31243
rect 54706 31212 55031 31240
rect 54706 31200 54712 31212
rect 55019 31209 55031 31212
rect 55065 31209 55077 31243
rect 55019 31203 55077 31209
rect 35515 31175 35573 31181
rect 35515 31172 35527 31175
rect 35478 31144 35527 31172
rect 35478 31132 35484 31144
rect 35515 31141 35527 31144
rect 35561 31141 35573 31175
rect 35515 31135 35573 31141
rect 47380 31132 47386 31184
rect 47438 31172 47444 31184
rect 49772 31172 49778 31184
rect 47438 31144 49778 31172
rect 47438 31132 47444 31144
rect 49772 31132 49778 31144
rect 49830 31132 49836 31184
rect 50876 31132 50882 31184
rect 50934 31172 50940 31184
rect 53179 31175 53237 31181
rect 53179 31172 53191 31175
rect 50934 31144 53191 31172
rect 50934 31132 50940 31144
rect 53179 31141 53191 31144
rect 53225 31141 53237 31175
rect 53179 31135 53237 31141
rect 54096 31132 54102 31184
rect 54154 31172 54160 31184
rect 54666 31172 54694 31200
rect 54832 31172 54838 31184
rect 54154 31144 54694 31172
rect 54793 31144 54838 31172
rect 54154 31132 54160 31144
rect 54832 31132 54838 31144
rect 54890 31132 54896 31184
rect 57610 31172 57638 31271
rect 57868 31268 57874 31280
rect 57926 31268 57932 31320
rect 58530 31240 58558 31348
rect 58604 31336 58610 31388
rect 58662 31376 58668 31388
rect 63130 31376 63158 31416
rect 67896 31404 67902 31416
rect 67954 31404 67960 31456
rect 68356 31404 68362 31456
rect 68414 31444 68420 31456
rect 68742 31444 68770 31484
rect 69003 31481 69015 31484
rect 69049 31481 69061 31515
rect 69003 31475 69061 31481
rect 69184 31472 69190 31524
rect 69242 31512 69248 31524
rect 71668 31512 71674 31524
rect 69242 31484 71674 31512
rect 69242 31472 69248 31484
rect 71668 31472 71674 31484
rect 71726 31472 71732 31524
rect 73968 31472 73974 31524
rect 74026 31512 74032 31524
rect 74063 31515 74121 31521
rect 74063 31512 74075 31515
rect 74026 31484 74075 31512
rect 74026 31472 74032 31484
rect 74063 31481 74075 31484
rect 74109 31481 74121 31515
rect 74063 31475 74121 31481
rect 78660 31472 78666 31524
rect 78718 31512 78724 31524
rect 82895 31515 82953 31521
rect 82895 31512 82907 31515
rect 78718 31484 82907 31512
rect 78718 31472 78724 31484
rect 82895 31481 82907 31484
rect 82941 31481 82953 31515
rect 82895 31475 82953 31481
rect 82984 31472 82990 31524
rect 83042 31512 83048 31524
rect 88320 31512 88326 31524
rect 83042 31484 88326 31512
rect 83042 31472 83048 31484
rect 88320 31472 88326 31484
rect 88378 31472 88384 31524
rect 88412 31472 88418 31524
rect 88470 31512 88476 31524
rect 88470 31484 88515 31512
rect 88470 31472 88476 31484
rect 68414 31416 68770 31444
rect 68414 31404 68420 31416
rect 68816 31404 68822 31456
rect 68874 31444 68880 31456
rect 82784 31447 82842 31453
rect 68874 31416 82754 31444
rect 68874 31404 68880 31416
rect 58662 31348 63158 31376
rect 58662 31336 58668 31348
rect 63204 31336 63210 31388
rect 63262 31376 63268 31388
rect 68727 31379 68785 31385
rect 63262 31348 68678 31376
rect 63262 31336 63268 31348
rect 59251 31311 59309 31317
rect 59251 31277 59263 31311
rect 59297 31308 59309 31311
rect 60079 31311 60137 31317
rect 60079 31308 60091 31311
rect 59297 31280 60091 31308
rect 59297 31277 59309 31280
rect 59251 31271 59309 31277
rect 60079 31277 60091 31280
rect 60125 31277 60137 31311
rect 60079 31271 60137 31277
rect 60168 31268 60174 31320
rect 60226 31308 60232 31320
rect 62655 31311 62713 31317
rect 60226 31280 60271 31308
rect 60226 31268 60232 31280
rect 62655 31277 62667 31311
rect 62701 31308 62713 31311
rect 62744 31308 62750 31320
rect 62701 31280 62750 31308
rect 62701 31277 62713 31280
rect 62655 31271 62713 31277
rect 62744 31268 62750 31280
rect 62802 31268 62808 31320
rect 66243 31311 66301 31317
rect 66243 31308 66255 31311
rect 65890 31280 66255 31308
rect 61824 31240 61830 31252
rect 58530 31212 61830 31240
rect 61824 31200 61830 31212
rect 61882 31200 61888 31252
rect 65890 31184 65918 31280
rect 66243 31277 66255 31280
rect 66289 31277 66301 31311
rect 66243 31271 66301 31277
rect 68080 31268 68086 31320
rect 68138 31308 68144 31320
rect 68359 31311 68417 31317
rect 68359 31308 68371 31311
rect 68138 31280 68371 31308
rect 68138 31268 68144 31280
rect 68359 31277 68371 31280
rect 68405 31277 68417 31311
rect 68359 31271 68417 31277
rect 68506 31311 68564 31317
rect 68506 31277 68518 31311
rect 68552 31277 68564 31311
rect 68650 31308 68678 31348
rect 68727 31345 68739 31379
rect 68773 31376 68785 31379
rect 73784 31376 73790 31388
rect 68773 31348 73790 31376
rect 68773 31345 68785 31348
rect 68727 31339 68785 31345
rect 73784 31336 73790 31348
rect 73842 31336 73848 31388
rect 71760 31308 71766 31320
rect 68650 31280 71766 31308
rect 68506 31271 68564 31277
rect 68521 31240 68549 31271
rect 71760 31268 71766 31280
rect 71818 31268 71824 31320
rect 73603 31311 73661 31317
rect 73603 31308 73615 31311
rect 73342 31280 73615 31308
rect 68190 31212 68549 31240
rect 68190 31184 68218 31212
rect 60352 31172 60358 31184
rect 57610 31144 60358 31172
rect 60352 31132 60358 31144
rect 60410 31132 60416 31184
rect 65872 31172 65878 31184
rect 65833 31144 65878 31172
rect 65872 31132 65878 31144
rect 65930 31132 65936 31184
rect 66056 31172 66062 31184
rect 66017 31144 66062 31172
rect 66056 31132 66062 31144
rect 66114 31132 66120 31184
rect 68172 31172 68178 31184
rect 68133 31144 68178 31172
rect 68172 31132 68178 31144
rect 68230 31132 68236 31184
rect 73232 31132 73238 31184
rect 73290 31172 73296 31184
rect 73342 31181 73370 31280
rect 73603 31277 73615 31280
rect 73649 31277 73661 31311
rect 73603 31271 73661 31277
rect 73879 31311 73937 31317
rect 73879 31277 73891 31311
rect 73925 31308 73937 31311
rect 74152 31308 74158 31320
rect 73925 31280 74158 31308
rect 73925 31277 73937 31280
rect 73879 31271 73937 31277
rect 74152 31268 74158 31280
rect 74210 31268 74216 31320
rect 75348 31308 75354 31320
rect 75261 31280 75354 31308
rect 75348 31268 75354 31280
rect 75406 31308 75412 31320
rect 76544 31308 76550 31320
rect 75406 31280 76550 31308
rect 75406 31268 75412 31280
rect 76544 31268 76550 31280
rect 76602 31268 76608 31320
rect 80687 31311 80745 31317
rect 80687 31308 80699 31311
rect 80518 31280 80699 31308
rect 73787 31243 73845 31249
rect 73787 31209 73799 31243
rect 73833 31209 73845 31243
rect 73787 31203 73845 31209
rect 73327 31175 73385 31181
rect 73327 31172 73339 31175
rect 73290 31144 73339 31172
rect 73290 31132 73296 31144
rect 73327 31141 73339 31144
rect 73373 31141 73385 31175
rect 73802 31172 73830 31203
rect 74336 31200 74342 31252
rect 74394 31240 74400 31252
rect 75167 31243 75225 31249
rect 75167 31240 75179 31243
rect 74394 31212 75179 31240
rect 74394 31200 74400 31212
rect 75167 31209 75179 31212
rect 75213 31209 75225 31243
rect 75167 31203 75225 31209
rect 75719 31243 75777 31249
rect 75719 31209 75731 31243
rect 75765 31209 75777 31243
rect 75719 31203 75777 31209
rect 75734 31172 75762 31203
rect 80518 31184 80546 31280
rect 80687 31277 80699 31280
rect 80733 31277 80745 31311
rect 80687 31271 80745 31277
rect 81239 31311 81297 31317
rect 81239 31277 81251 31311
rect 81285 31277 81297 31311
rect 81512 31308 81518 31320
rect 81473 31280 81518 31308
rect 81239 31271 81297 31277
rect 80592 31200 80598 31252
rect 80650 31240 80656 31252
rect 81254 31240 81282 31271
rect 81512 31268 81518 31280
rect 81570 31268 81576 31320
rect 82616 31308 82622 31320
rect 82577 31280 82622 31308
rect 82616 31268 82622 31280
rect 82674 31268 82680 31320
rect 82726 31308 82754 31416
rect 82784 31413 82796 31447
rect 82830 31444 82842 31447
rect 84272 31444 84278 31456
rect 82830 31416 84278 31444
rect 82830 31413 82842 31416
rect 82784 31407 82842 31413
rect 84272 31404 84278 31416
rect 84330 31404 84336 31456
rect 84364 31404 84370 31456
rect 84422 31444 84428 31456
rect 89332 31444 89338 31456
rect 84422 31416 89338 31444
rect 84422 31404 84428 31416
rect 89332 31404 89338 31416
rect 89390 31404 89396 31456
rect 82987 31379 83045 31385
rect 82987 31345 82999 31379
rect 83033 31376 83045 31379
rect 90712 31376 90718 31388
rect 83033 31348 89010 31376
rect 90673 31348 90718 31376
rect 83033 31345 83045 31348
rect 82987 31339 83045 31345
rect 83355 31311 83413 31317
rect 83355 31308 83367 31311
rect 82726 31280 83367 31308
rect 83355 31277 83367 31280
rect 83401 31277 83413 31311
rect 88320 31308 88326 31320
rect 88281 31280 88326 31308
rect 83355 31271 83413 31277
rect 88320 31268 88326 31280
rect 88378 31268 88384 31320
rect 88982 31308 89010 31348
rect 90712 31336 90718 31348
rect 90770 31376 90776 31388
rect 90770 31348 91034 31376
rect 90770 31336 90776 31348
rect 90896 31308 90902 31320
rect 88982 31280 89194 31308
rect 90857 31280 90902 31308
rect 80650 31212 81282 31240
rect 89166 31240 89194 31280
rect 90896 31268 90902 31280
rect 90954 31268 90960 31320
rect 91006 31308 91034 31348
rect 91359 31311 91417 31317
rect 91359 31308 91371 31311
rect 91006 31280 91371 31308
rect 91359 31277 91371 31280
rect 91405 31277 91417 31311
rect 91359 31271 91417 31277
rect 91448 31268 91454 31320
rect 91506 31308 91512 31320
rect 91506 31280 91551 31308
rect 91506 31268 91512 31280
rect 92003 31243 92061 31249
rect 92003 31240 92015 31243
rect 89166 31212 92015 31240
rect 80650 31200 80656 31212
rect 92003 31209 92015 31212
rect 92049 31209 92061 31243
rect 92003 31203 92061 31209
rect 80316 31172 80322 31184
rect 73802 31144 80322 31172
rect 73327 31135 73385 31141
rect 80316 31132 80322 31144
rect 80374 31132 80380 31184
rect 80500 31172 80506 31184
rect 80461 31144 80506 31172
rect 80500 31132 80506 31144
rect 80558 31132 80564 31184
rect 80776 31172 80782 31184
rect 80737 31144 80782 31172
rect 80776 31132 80782 31144
rect 80834 31132 80840 31184
rect 538 31082 93642 31104
rect 538 31030 6344 31082
rect 6396 31030 6408 31082
rect 6460 31030 6472 31082
rect 6524 31030 6536 31082
rect 6588 31030 11672 31082
rect 11724 31030 11736 31082
rect 11788 31030 11800 31082
rect 11852 31030 11864 31082
rect 11916 31030 17000 31082
rect 17052 31030 17064 31082
rect 17116 31030 17128 31082
rect 17180 31030 17192 31082
rect 17244 31030 22328 31082
rect 22380 31030 22392 31082
rect 22444 31030 22456 31082
rect 22508 31030 22520 31082
rect 22572 31030 27656 31082
rect 27708 31030 27720 31082
rect 27772 31030 27784 31082
rect 27836 31030 27848 31082
rect 27900 31030 32984 31082
rect 33036 31030 33048 31082
rect 33100 31030 33112 31082
rect 33164 31030 33176 31082
rect 33228 31030 38312 31082
rect 38364 31030 38376 31082
rect 38428 31030 38440 31082
rect 38492 31030 38504 31082
rect 38556 31030 43640 31082
rect 43692 31030 43704 31082
rect 43756 31030 43768 31082
rect 43820 31030 43832 31082
rect 43884 31030 48968 31082
rect 49020 31030 49032 31082
rect 49084 31030 49096 31082
rect 49148 31030 49160 31082
rect 49212 31030 54296 31082
rect 54348 31030 54360 31082
rect 54412 31030 54424 31082
rect 54476 31030 54488 31082
rect 54540 31030 59624 31082
rect 59676 31030 59688 31082
rect 59740 31030 59752 31082
rect 59804 31030 59816 31082
rect 59868 31030 64952 31082
rect 65004 31030 65016 31082
rect 65068 31030 65080 31082
rect 65132 31030 65144 31082
rect 65196 31030 70280 31082
rect 70332 31030 70344 31082
rect 70396 31030 70408 31082
rect 70460 31030 70472 31082
rect 70524 31030 75608 31082
rect 75660 31030 75672 31082
rect 75724 31030 75736 31082
rect 75788 31030 75800 31082
rect 75852 31030 80936 31082
rect 80988 31030 81000 31082
rect 81052 31030 81064 31082
rect 81116 31030 81128 31082
rect 81180 31030 86264 31082
rect 86316 31030 86328 31082
rect 86380 31030 86392 31082
rect 86444 31030 86456 31082
rect 86508 31030 91592 31082
rect 91644 31030 91656 31082
rect 91708 31030 91720 31082
rect 91772 31030 91784 31082
rect 91836 31030 93642 31082
rect 538 31008 93642 31030
rect 4235 30971 4293 30977
rect 4235 30937 4247 30971
rect 4281 30968 4293 30971
rect 4968 30968 4974 30980
rect 4281 30940 4974 30968
rect 4281 30937 4293 30940
rect 4235 30931 4293 30937
rect 4342 30841 4370 30940
rect 4968 30928 4974 30940
rect 5026 30928 5032 30980
rect 5060 30928 5066 30980
rect 5118 30968 5124 30980
rect 5247 30971 5305 30977
rect 5247 30968 5259 30971
rect 5118 30940 5259 30968
rect 5118 30928 5124 30940
rect 5247 30937 5259 30940
rect 5293 30937 5305 30971
rect 14720 30968 14726 30980
rect 5247 30931 5305 30937
rect 10506 30940 14726 30968
rect 4327 30835 4385 30841
rect 4327 30801 4339 30835
rect 4373 30801 4385 30835
rect 5262 30832 5290 30931
rect 10506 30909 10534 30940
rect 14720 30928 14726 30940
rect 14778 30928 14784 30980
rect 15916 30968 15922 30980
rect 15877 30940 15922 30968
rect 15916 30928 15922 30940
rect 15974 30928 15980 30980
rect 17664 30928 17670 30980
rect 17722 30968 17728 30980
rect 29167 30971 29225 30977
rect 17722 30940 28290 30968
rect 17722 30928 17728 30940
rect 10031 30903 10089 30909
rect 10031 30869 10043 30903
rect 10077 30900 10089 30903
rect 10491 30903 10549 30909
rect 10491 30900 10503 30903
rect 10077 30872 10503 30900
rect 10077 30869 10089 30872
rect 10031 30863 10089 30869
rect 10491 30869 10503 30872
rect 10537 30869 10549 30903
rect 10491 30863 10549 30869
rect 10859 30903 10917 30909
rect 10859 30869 10871 30903
rect 10905 30900 10917 30903
rect 11500 30900 11506 30912
rect 10905 30872 11506 30900
rect 10905 30869 10917 30872
rect 10859 30863 10917 30869
rect 11500 30860 11506 30872
rect 11558 30860 11564 30912
rect 13343 30903 13401 30909
rect 13343 30900 13355 30903
rect 13174 30872 13355 30900
rect 5431 30835 5489 30841
rect 5431 30832 5443 30835
rect 5262 30804 5443 30832
rect 4327 30795 4385 30801
rect 5431 30801 5443 30804
rect 5477 30801 5489 30835
rect 5431 30795 5489 30801
rect 6535 30835 6593 30841
rect 6535 30801 6547 30835
rect 6581 30801 6593 30835
rect 6535 30795 6593 30801
rect 6256 30764 6262 30776
rect 4526 30736 6262 30764
rect 4526 30705 4554 30736
rect 6256 30724 6262 30736
rect 6314 30764 6320 30776
rect 6550 30764 6578 30795
rect 6624 30792 6630 30844
rect 6682 30832 6688 30844
rect 6811 30835 6869 30841
rect 6682 30804 6727 30832
rect 6682 30792 6688 30804
rect 6811 30801 6823 30835
rect 6857 30801 6869 30835
rect 6811 30795 6869 30801
rect 6826 30764 6854 30795
rect 6900 30792 6906 30844
rect 6958 30832 6964 30844
rect 10304 30832 10310 30844
rect 6958 30804 10310 30832
rect 6958 30792 6964 30804
rect 10304 30792 10310 30804
rect 10362 30792 10368 30844
rect 10396 30792 10402 30844
rect 10454 30832 10460 30844
rect 10454 30804 10499 30832
rect 10454 30792 10460 30804
rect 11408 30792 11414 30844
rect 11466 30832 11472 30844
rect 12147 30835 12205 30841
rect 12147 30832 12159 30835
rect 11466 30804 12159 30832
rect 11466 30792 11472 30804
rect 12147 30801 12159 30804
rect 12193 30801 12205 30835
rect 12328 30832 12334 30844
rect 12289 30804 12334 30832
rect 12147 30795 12205 30801
rect 12328 30792 12334 30804
rect 12386 30792 12392 30844
rect 12420 30792 12426 30844
rect 12478 30832 12484 30844
rect 12607 30835 12665 30841
rect 12607 30832 12619 30835
rect 12478 30804 12619 30832
rect 12478 30792 12484 30804
rect 12607 30801 12619 30804
rect 12653 30832 12665 30835
rect 12788 30832 12794 30844
rect 12653 30804 12794 30832
rect 12653 30801 12665 30804
rect 12607 30795 12665 30801
rect 12788 30792 12794 30804
rect 12846 30792 12852 30844
rect 13174 30841 13202 30872
rect 13343 30869 13355 30872
rect 13389 30900 13401 30903
rect 19872 30900 19878 30912
rect 13389 30872 19878 30900
rect 13389 30869 13401 30872
rect 13343 30863 13401 30869
rect 19872 30860 19878 30872
rect 19930 30860 19936 30912
rect 21899 30903 21957 30909
rect 21899 30900 21911 30903
rect 21454 30872 21911 30900
rect 13159 30835 13217 30841
rect 13159 30801 13171 30835
rect 13205 30801 13217 30835
rect 13159 30795 13217 30801
rect 14812 30792 14818 30844
rect 14870 30832 14876 30844
rect 15916 30832 15922 30844
rect 14870 30804 15922 30832
rect 14870 30792 14876 30804
rect 15916 30792 15922 30804
rect 15974 30832 15980 30844
rect 16011 30835 16069 30841
rect 16011 30832 16023 30835
rect 15974 30804 16023 30832
rect 15974 30792 15980 30804
rect 16011 30801 16023 30804
rect 16057 30801 16069 30835
rect 16011 30795 16069 30801
rect 16195 30835 16253 30841
rect 16195 30801 16207 30835
rect 16241 30832 16253 30835
rect 16744 30832 16750 30844
rect 16241 30804 16750 30832
rect 16241 30801 16253 30804
rect 16195 30795 16253 30801
rect 16744 30792 16750 30804
rect 16802 30792 16808 30844
rect 16931 30835 16989 30841
rect 16931 30801 16943 30835
rect 16977 30832 16989 30835
rect 17572 30832 17578 30844
rect 16977 30804 17578 30832
rect 16977 30801 16989 30804
rect 16931 30795 16989 30801
rect 17572 30792 17578 30804
rect 17630 30792 17636 30844
rect 18495 30835 18553 30841
rect 18495 30801 18507 30835
rect 18541 30832 18553 30835
rect 18860 30832 18866 30844
rect 18541 30804 18866 30832
rect 18541 30801 18553 30804
rect 18495 30795 18553 30801
rect 18860 30792 18866 30804
rect 18918 30792 18924 30844
rect 6314 30736 6578 30764
rect 6734 30736 6854 30764
rect 7271 30767 7329 30773
rect 6314 30724 6320 30736
rect 4511 30699 4569 30705
rect 4511 30665 4523 30699
rect 4557 30665 4569 30699
rect 4511 30659 4569 30665
rect 5060 30656 5066 30708
rect 5118 30696 5124 30708
rect 6734 30696 6762 30736
rect 7271 30733 7283 30767
rect 7317 30764 7329 30767
rect 9476 30764 9482 30776
rect 7317 30736 9482 30764
rect 7317 30733 7329 30736
rect 7271 30727 7329 30733
rect 9476 30724 9482 30736
rect 9534 30724 9540 30776
rect 10120 30764 10126 30776
rect 10081 30736 10126 30764
rect 10120 30724 10126 30736
rect 10178 30724 10184 30776
rect 11500 30724 11506 30776
rect 11558 30764 11564 30776
rect 11687 30767 11745 30773
rect 11687 30764 11699 30767
rect 11558 30736 11699 30764
rect 11558 30724 11564 30736
rect 11687 30733 11699 30736
rect 11733 30733 11745 30767
rect 11687 30727 11745 30733
rect 12975 30767 13033 30773
rect 12975 30733 12987 30767
rect 13021 30764 13033 30767
rect 13435 30767 13493 30773
rect 13435 30764 13447 30767
rect 13021 30736 13447 30764
rect 13021 30733 13033 30736
rect 12975 30727 13033 30733
rect 13435 30733 13447 30736
rect 13481 30733 13493 30767
rect 13435 30727 13493 30733
rect 8188 30696 8194 30708
rect 5118 30668 8194 30696
rect 5118 30656 5124 30668
rect 8188 30656 8194 30668
rect 8246 30656 8252 30708
rect 5615 30631 5673 30637
rect 5615 30597 5627 30631
rect 5661 30628 5673 30631
rect 6900 30628 6906 30640
rect 5661 30600 6906 30628
rect 5661 30597 5673 30600
rect 5615 30591 5673 30597
rect 6900 30588 6906 30600
rect 6958 30588 6964 30640
rect 7084 30588 7090 30640
rect 7142 30628 7148 30640
rect 13156 30628 13162 30640
rect 7142 30600 13162 30628
rect 7142 30588 7148 30600
rect 13156 30588 13162 30600
rect 13214 30588 13220 30640
rect 13450 30628 13478 30727
rect 18032 30724 18038 30776
rect 18090 30764 18096 30776
rect 21454 30764 21482 30872
rect 21899 30869 21911 30872
rect 21945 30900 21957 30903
rect 28262 30900 28290 30940
rect 29167 30937 29179 30971
rect 29213 30968 29225 30971
rect 29256 30968 29262 30980
rect 29213 30940 29262 30968
rect 29213 30937 29225 30940
rect 29167 30931 29225 30937
rect 29256 30928 29262 30940
rect 29314 30928 29320 30980
rect 29348 30928 29354 30980
rect 29406 30968 29412 30980
rect 29406 30940 38134 30968
rect 29406 30928 29412 30940
rect 30912 30900 30918 30912
rect 21945 30872 22126 30900
rect 28262 30872 30918 30900
rect 21945 30869 21957 30872
rect 21899 30863 21957 30869
rect 22098 30841 22126 30872
rect 30912 30860 30918 30872
rect 30970 30860 30976 30912
rect 38106 30900 38134 30940
rect 38640 30928 38646 30980
rect 38698 30968 38704 30980
rect 68172 30968 68178 30980
rect 38698 30940 68178 30968
rect 38698 30928 38704 30940
rect 68172 30928 68178 30940
rect 68230 30928 68236 30980
rect 68926 30940 79626 30968
rect 52164 30900 52170 30912
rect 38106 30872 52170 30900
rect 52164 30860 52170 30872
rect 52222 30860 52228 30912
rect 53820 30900 53826 30912
rect 52366 30872 53826 30900
rect 22083 30835 22141 30841
rect 22083 30801 22095 30835
rect 22129 30832 22141 30835
rect 23920 30832 23926 30844
rect 22129 30804 23926 30832
rect 22129 30801 22141 30804
rect 22083 30795 22141 30801
rect 23920 30792 23926 30804
rect 23978 30832 23984 30844
rect 24840 30832 24846 30844
rect 23978 30804 24846 30832
rect 23978 30792 23984 30804
rect 24840 30792 24846 30804
rect 24898 30792 24904 30844
rect 27327 30835 27385 30841
rect 27327 30801 27339 30835
rect 27373 30832 27385 30835
rect 28796 30832 28802 30844
rect 27373 30804 28802 30832
rect 27373 30801 27385 30804
rect 27327 30795 27385 30801
rect 28796 30792 28802 30804
rect 28854 30792 28860 30844
rect 32939 30835 32997 30841
rect 32586 30804 32798 30832
rect 18090 30736 21482 30764
rect 22359 30767 22417 30773
rect 18090 30724 18096 30736
rect 22359 30733 22371 30767
rect 22405 30764 22417 30767
rect 23092 30764 23098 30776
rect 22405 30736 23098 30764
rect 22405 30733 22417 30736
rect 22359 30727 22417 30733
rect 23092 30724 23098 30736
rect 23150 30724 23156 30776
rect 27508 30724 27514 30776
rect 27566 30764 27572 30776
rect 27603 30767 27661 30773
rect 27603 30764 27615 30767
rect 27566 30736 27615 30764
rect 27566 30724 27572 30736
rect 27603 30733 27615 30736
rect 27649 30733 27661 30767
rect 27603 30727 27661 30733
rect 27692 30724 27698 30776
rect 27750 30764 27756 30776
rect 32586 30764 32614 30804
rect 27750 30736 32614 30764
rect 32663 30767 32721 30773
rect 27750 30724 27756 30736
rect 32663 30733 32675 30767
rect 32709 30733 32721 30767
rect 32770 30764 32798 30804
rect 32939 30801 32951 30835
rect 32985 30832 32997 30835
rect 33304 30832 33310 30844
rect 32985 30804 33310 30832
rect 32985 30801 32997 30804
rect 32939 30795 32997 30801
rect 33304 30792 33310 30804
rect 33362 30792 33368 30844
rect 35147 30835 35205 30841
rect 35147 30832 35159 30835
rect 34978 30804 35159 30832
rect 34500 30764 34506 30776
rect 32770 30736 34506 30764
rect 32663 30727 32721 30733
rect 16376 30656 16382 30708
rect 16434 30696 16440 30708
rect 17115 30699 17173 30705
rect 17115 30696 17127 30699
rect 16434 30668 17127 30696
rect 16434 30656 16440 30668
rect 17115 30665 17127 30668
rect 17161 30665 17173 30699
rect 19504 30696 19510 30708
rect 17115 30659 17173 30665
rect 17406 30668 19510 30696
rect 17406 30628 17434 30668
rect 19504 30656 19510 30668
rect 19562 30656 19568 30708
rect 23736 30656 23742 30708
rect 23794 30696 23800 30708
rect 27324 30696 27330 30708
rect 23794 30668 27330 30696
rect 23794 30656 23800 30668
rect 27324 30656 27330 30668
rect 27382 30656 27388 30708
rect 17572 30628 17578 30640
rect 13450 30600 17434 30628
rect 17533 30600 17578 30628
rect 17572 30588 17578 30600
rect 17630 30588 17636 30640
rect 18679 30631 18737 30637
rect 18679 30597 18691 30631
rect 18725 30628 18737 30631
rect 18860 30628 18866 30640
rect 18725 30600 18866 30628
rect 18725 30597 18737 30600
rect 18679 30591 18737 30597
rect 18860 30588 18866 30600
rect 18918 30588 18924 30640
rect 23644 30628 23650 30640
rect 23605 30600 23650 30628
rect 23644 30588 23650 30600
rect 23702 30588 23708 30640
rect 28704 30628 28710 30640
rect 28665 30600 28710 30628
rect 28704 30588 28710 30600
rect 28762 30588 28768 30640
rect 32678 30628 32706 30727
rect 34500 30724 34506 30736
rect 34558 30724 34564 30776
rect 33874 30668 34178 30696
rect 33874 30628 33902 30668
rect 34040 30628 34046 30640
rect 32678 30600 33902 30628
rect 34001 30600 34046 30628
rect 34040 30588 34046 30600
rect 34098 30588 34104 30640
rect 34150 30628 34178 30668
rect 34224 30656 34230 30708
rect 34282 30696 34288 30708
rect 34684 30696 34690 30708
rect 34282 30668 34690 30696
rect 34282 30656 34288 30668
rect 34684 30656 34690 30668
rect 34742 30696 34748 30708
rect 34978 30705 35006 30804
rect 35147 30801 35159 30804
rect 35193 30801 35205 30835
rect 35147 30795 35205 30801
rect 36984 30792 36990 30844
rect 37042 30832 37048 30844
rect 37447 30835 37505 30841
rect 37447 30832 37459 30835
rect 37042 30804 37459 30832
rect 37042 30792 37048 30804
rect 37447 30801 37459 30804
rect 37493 30801 37505 30835
rect 37447 30795 37505 30801
rect 43608 30792 43614 30844
rect 43666 30832 43672 30844
rect 44436 30832 44442 30844
rect 43666 30804 44442 30832
rect 43666 30792 43672 30804
rect 44436 30792 44442 30804
rect 44494 30792 44500 30844
rect 44620 30792 44626 30844
rect 44678 30832 44684 30844
rect 52366 30841 52394 30872
rect 53820 30860 53826 30872
rect 53878 30900 53884 30912
rect 57595 30903 57653 30909
rect 53878 30872 54326 30900
rect 53878 30860 53884 30872
rect 44899 30835 44957 30841
rect 44899 30832 44911 30835
rect 44678 30804 44911 30832
rect 44678 30792 44684 30804
rect 44899 30801 44911 30804
rect 44945 30801 44957 30835
rect 44899 30795 44957 30801
rect 44991 30835 45049 30841
rect 44991 30801 45003 30835
rect 45037 30832 45049 30835
rect 48395 30835 48453 30841
rect 45037 30804 45862 30832
rect 45037 30801 45049 30804
rect 44991 30795 45049 30801
rect 37171 30767 37229 30773
rect 37171 30764 37183 30767
rect 36910 30736 37183 30764
rect 34963 30699 35021 30705
rect 34963 30696 34975 30699
rect 34742 30668 34975 30696
rect 34742 30656 34748 30668
rect 34963 30665 34975 30668
rect 35009 30665 35021 30699
rect 34963 30659 35021 30665
rect 35052 30656 35058 30708
rect 35110 30696 35116 30708
rect 35331 30699 35389 30705
rect 35331 30696 35343 30699
rect 35110 30668 35343 30696
rect 35110 30656 35116 30668
rect 35331 30665 35343 30668
rect 35377 30665 35389 30699
rect 35331 30659 35389 30665
rect 36910 30637 36938 30736
rect 37171 30733 37183 30736
rect 37217 30764 37229 30767
rect 37812 30764 37818 30776
rect 37217 30736 37818 30764
rect 37217 30733 37229 30736
rect 37171 30727 37229 30733
rect 37812 30724 37818 30736
rect 37870 30724 37876 30776
rect 42872 30724 42878 30776
rect 42930 30764 42936 30776
rect 43424 30764 43430 30776
rect 42930 30736 43430 30764
rect 42930 30724 42936 30736
rect 43424 30724 43430 30736
rect 43482 30764 43488 30776
rect 44071 30767 44129 30773
rect 44071 30764 44083 30767
rect 43482 30736 44083 30764
rect 43482 30724 43488 30736
rect 44071 30733 44083 30736
rect 44117 30764 44129 30767
rect 44255 30767 44313 30773
rect 44255 30764 44267 30767
rect 44117 30736 44267 30764
rect 44117 30733 44129 30736
rect 44071 30727 44129 30733
rect 44255 30733 44267 30736
rect 44301 30733 44313 30767
rect 44255 30727 44313 30733
rect 45834 30705 45862 30804
rect 48395 30801 48407 30835
rect 48441 30832 48453 30835
rect 52259 30835 52317 30841
rect 52259 30832 52271 30835
rect 48441 30804 52271 30832
rect 48441 30801 48453 30804
rect 48395 30795 48453 30801
rect 52259 30801 52271 30804
rect 52305 30801 52317 30835
rect 52259 30795 52317 30801
rect 52351 30835 52409 30841
rect 52351 30801 52363 30835
rect 52397 30801 52409 30835
rect 52351 30795 52409 30801
rect 52627 30835 52685 30841
rect 52627 30801 52639 30835
rect 52673 30832 52685 30835
rect 53179 30835 53237 30841
rect 53179 30832 53191 30835
rect 52673 30804 53191 30832
rect 52673 30801 52685 30804
rect 52627 30795 52685 30801
rect 53179 30801 53191 30804
rect 53225 30832 53237 30835
rect 54096 30832 54102 30844
rect 53225 30804 54102 30832
rect 53225 30801 53237 30804
rect 53179 30795 53237 30801
rect 47656 30724 47662 30776
rect 47714 30764 47720 30776
rect 48763 30767 48821 30773
rect 48763 30764 48775 30767
rect 47714 30736 48775 30764
rect 47714 30724 47720 30736
rect 48763 30733 48775 30736
rect 48809 30733 48821 30767
rect 48763 30727 48821 30733
rect 48852 30724 48858 30776
rect 48910 30764 48916 30776
rect 48910 30736 48955 30764
rect 48910 30724 48916 30736
rect 50692 30724 50698 30776
rect 50750 30764 50756 30776
rect 52642 30764 52670 30795
rect 54096 30792 54102 30804
rect 54154 30792 54160 30844
rect 54298 30841 54326 30872
rect 57595 30869 57607 30903
rect 57641 30900 57653 30903
rect 57868 30900 57874 30912
rect 57641 30872 57874 30900
rect 57641 30869 57653 30872
rect 57595 30863 57653 30869
rect 57868 30860 57874 30872
rect 57926 30860 57932 30912
rect 62100 30860 62106 30912
rect 62158 30900 62164 30912
rect 63115 30903 63173 30909
rect 63115 30900 63127 30903
rect 62158 30872 63127 30900
rect 62158 30860 62164 30872
rect 54283 30835 54341 30841
rect 54283 30801 54295 30835
rect 54329 30801 54341 30835
rect 54283 30795 54341 30801
rect 54559 30835 54617 30841
rect 54559 30801 54571 30835
rect 54605 30832 54617 30835
rect 54832 30832 54838 30844
rect 54605 30804 54838 30832
rect 54605 30801 54617 30804
rect 54559 30795 54617 30801
rect 54832 30792 54838 30804
rect 54890 30792 54896 30844
rect 55019 30835 55077 30841
rect 55019 30801 55031 30835
rect 55065 30832 55077 30835
rect 58144 30832 58150 30844
rect 55065 30804 58006 30832
rect 58105 30804 58150 30832
rect 55065 30801 55077 30804
rect 55019 30795 55077 30801
rect 52808 30764 52814 30776
rect 50750 30736 52670 30764
rect 52769 30736 52814 30764
rect 50750 30724 50756 30736
rect 52808 30724 52814 30736
rect 52866 30724 52872 30776
rect 52900 30724 52906 30776
rect 52958 30764 52964 30776
rect 54375 30767 54433 30773
rect 54375 30764 54387 30767
rect 52958 30736 54387 30764
rect 52958 30724 52964 30736
rect 54375 30733 54387 30736
rect 54421 30733 54433 30767
rect 57978 30764 58006 30804
rect 58144 30792 58150 30804
rect 58202 30792 58208 30844
rect 58328 30792 58334 30844
rect 58386 30832 58392 30844
rect 58423 30835 58481 30841
rect 58423 30832 58435 30835
rect 58386 30804 58435 30832
rect 58386 30792 58392 30804
rect 58423 30801 58435 30804
rect 58469 30801 58481 30835
rect 58423 30795 58481 30801
rect 58512 30792 58518 30844
rect 58570 30832 58576 30844
rect 58607 30835 58665 30841
rect 58607 30832 58619 30835
rect 58570 30804 58619 30832
rect 58570 30792 58576 30804
rect 58607 30801 58619 30804
rect 58653 30801 58665 30835
rect 58607 30795 58665 30801
rect 62008 30792 62014 30844
rect 62066 30832 62072 30844
rect 62486 30841 62514 30872
rect 63115 30869 63127 30872
rect 63161 30900 63173 30903
rect 63388 30900 63394 30912
rect 63161 30872 63394 30900
rect 63161 30869 63173 30872
rect 63115 30863 63173 30869
rect 63388 30860 63394 30872
rect 63446 30860 63452 30912
rect 62287 30835 62345 30841
rect 62287 30832 62299 30835
rect 62066 30804 62299 30832
rect 62066 30792 62072 30804
rect 62287 30801 62299 30804
rect 62333 30801 62345 30835
rect 62287 30795 62345 30801
rect 62471 30835 62529 30841
rect 62471 30801 62483 30835
rect 62517 30801 62529 30835
rect 62471 30795 62529 30801
rect 62302 30764 62330 30795
rect 62652 30792 62658 30844
rect 62710 30832 62716 30844
rect 62839 30835 62897 30841
rect 62839 30832 62851 30835
rect 62710 30804 62851 30832
rect 62710 30792 62716 30804
rect 62839 30801 62851 30804
rect 62885 30801 62897 30835
rect 62839 30795 62897 30801
rect 63020 30792 63026 30844
rect 63078 30832 63084 30844
rect 68926 30832 68954 30940
rect 75256 30900 75262 30912
rect 72882 30872 74474 30900
rect 63078 30804 68954 30832
rect 69003 30835 69061 30841
rect 63078 30792 63084 30804
rect 69003 30801 69015 30835
rect 69049 30832 69061 30835
rect 69920 30832 69926 30844
rect 69049 30804 69926 30832
rect 69049 30801 69061 30804
rect 69003 30795 69061 30801
rect 69920 30792 69926 30804
rect 69978 30792 69984 30844
rect 71119 30835 71177 30841
rect 71119 30801 71131 30835
rect 71165 30832 71177 30835
rect 71208 30832 71214 30844
rect 71165 30804 71214 30832
rect 71165 30801 71177 30804
rect 71119 30795 71177 30801
rect 71208 30792 71214 30804
rect 71266 30832 71272 30844
rect 72882 30841 72910 30872
rect 72867 30835 72925 30841
rect 72867 30832 72879 30835
rect 71266 30804 72879 30832
rect 71266 30792 71272 30804
rect 72867 30801 72879 30804
rect 72913 30801 72925 30835
rect 72867 30795 72925 30801
rect 73971 30835 74029 30841
rect 73971 30801 73983 30835
rect 74017 30801 74029 30835
rect 74152 30832 74158 30844
rect 74113 30804 74158 30832
rect 73971 30795 74029 30801
rect 62931 30767 62989 30773
rect 62931 30764 62943 30767
rect 57978 30736 59754 30764
rect 62302 30736 62943 30764
rect 54375 30727 54433 30733
rect 45819 30699 45877 30705
rect 45819 30665 45831 30699
rect 45865 30696 45877 30699
rect 46092 30696 46098 30708
rect 45865 30668 46098 30696
rect 45865 30665 45877 30668
rect 45819 30659 45877 30665
rect 46092 30656 46098 30668
rect 46150 30696 46156 30708
rect 52443 30699 52501 30705
rect 46150 30668 48898 30696
rect 46150 30656 46156 30668
rect 34411 30631 34469 30637
rect 34411 30628 34423 30631
rect 34150 30600 34423 30628
rect 34411 30597 34423 30600
rect 34457 30628 34469 30631
rect 36895 30631 36953 30637
rect 36895 30628 36907 30631
rect 34457 30600 36907 30628
rect 34457 30597 34469 30600
rect 34411 30591 34469 30597
rect 36895 30597 36907 30600
rect 36941 30597 36953 30631
rect 36895 30591 36953 30597
rect 36984 30588 36990 30640
rect 37042 30628 37048 30640
rect 38551 30631 38609 30637
rect 38551 30628 38563 30631
rect 37042 30600 38563 30628
rect 37042 30588 37048 30600
rect 38551 30597 38563 30600
rect 38597 30597 38609 30631
rect 45448 30628 45454 30640
rect 45409 30600 45454 30628
rect 38551 30591 38609 30597
rect 45448 30588 45454 30600
rect 45506 30588 45512 30640
rect 48300 30588 48306 30640
rect 48358 30628 48364 30640
rect 48533 30631 48591 30637
rect 48533 30628 48545 30631
rect 48358 30600 48545 30628
rect 48358 30588 48364 30600
rect 48533 30597 48545 30600
rect 48579 30597 48591 30631
rect 48533 30591 48591 30597
rect 48668 30588 48674 30640
rect 48726 30628 48732 30640
rect 48870 30628 48898 30668
rect 52443 30665 52455 30699
rect 52489 30696 52501 30699
rect 54004 30696 54010 30708
rect 52489 30668 54010 30696
rect 52489 30665 52501 30668
rect 52443 30659 52501 30665
rect 54004 30656 54010 30668
rect 54062 30656 54068 30708
rect 49404 30628 49410 30640
rect 48726 30600 48771 30628
rect 48870 30600 49410 30628
rect 48726 30588 48732 30600
rect 49404 30588 49410 30600
rect 49462 30588 49468 30640
rect 52259 30631 52317 30637
rect 52259 30597 52271 30631
rect 52305 30628 52317 30631
rect 59616 30628 59622 30640
rect 52305 30600 59622 30628
rect 52305 30597 52317 30600
rect 52259 30591 52317 30597
rect 59616 30588 59622 30600
rect 59674 30588 59680 30640
rect 59726 30628 59754 30736
rect 62931 30733 62943 30736
rect 62977 30733 62989 30767
rect 66516 30764 66522 30776
rect 66477 30736 66522 30764
rect 62931 30727 62989 30733
rect 66516 30724 66522 30736
rect 66574 30724 66580 30776
rect 66792 30764 66798 30776
rect 66753 30736 66798 30764
rect 66792 30724 66798 30736
rect 66850 30724 66856 30776
rect 66976 30724 66982 30776
rect 67034 30764 67040 30776
rect 67899 30767 67957 30773
rect 67899 30764 67911 30767
rect 67034 30736 67911 30764
rect 67034 30724 67040 30736
rect 67899 30733 67911 30736
rect 67945 30733 67957 30767
rect 71392 30764 71398 30776
rect 71353 30736 71398 30764
rect 67899 30727 67957 30733
rect 71392 30724 71398 30736
rect 71450 30724 71456 30776
rect 71760 30724 71766 30776
rect 71818 30764 71824 30776
rect 72312 30764 72318 30776
rect 71818 30736 72318 30764
rect 71818 30724 71824 30736
rect 72312 30724 72318 30736
rect 72370 30764 72376 30776
rect 72499 30767 72557 30773
rect 72499 30764 72511 30767
rect 72370 30736 72511 30764
rect 72370 30724 72376 30736
rect 72499 30733 72511 30736
rect 72545 30733 72557 30767
rect 73986 30764 74014 30795
rect 74152 30792 74158 30804
rect 74210 30792 74216 30844
rect 74446 30764 74474 30872
rect 74538 30872 75262 30900
rect 74538 30841 74566 30872
rect 75256 30860 75262 30872
rect 75314 30860 75320 30912
rect 79598 30900 79626 30940
rect 79672 30928 79678 30980
rect 79730 30968 79736 30980
rect 82159 30971 82217 30977
rect 82159 30968 82171 30971
rect 79730 30940 82171 30968
rect 79730 30928 79736 30940
rect 82159 30937 82171 30940
rect 82205 30937 82217 30971
rect 84824 30968 84830 30980
rect 84785 30940 84830 30968
rect 82159 30931 82217 30937
rect 84824 30928 84830 30940
rect 84882 30928 84888 30980
rect 87676 30968 87682 30980
rect 85762 30940 87682 30968
rect 79598 30872 84778 30900
rect 74523 30835 74581 30841
rect 74523 30801 74535 30835
rect 74569 30801 74581 30835
rect 74523 30795 74581 30801
rect 75072 30792 75078 30844
rect 75130 30832 75136 30844
rect 75351 30835 75409 30841
rect 75351 30832 75363 30835
rect 75130 30804 75363 30832
rect 75130 30792 75136 30804
rect 75351 30801 75363 30804
rect 75397 30801 75409 30835
rect 75351 30795 75409 30801
rect 75443 30835 75501 30841
rect 75443 30801 75455 30835
rect 75489 30832 75501 30835
rect 75532 30832 75538 30844
rect 75489 30804 75538 30832
rect 75489 30801 75501 30804
rect 75443 30795 75501 30801
rect 75532 30792 75538 30804
rect 75590 30792 75596 30844
rect 77464 30792 77470 30844
rect 77522 30832 77528 30844
rect 80687 30835 80745 30841
rect 77522 30804 78522 30832
rect 77522 30792 77528 30804
rect 77096 30764 77102 30776
rect 73986 30736 74382 30764
rect 74446 30736 77102 30764
rect 72499 30727 72557 30733
rect 74354 30708 74382 30736
rect 77096 30724 77102 30736
rect 77154 30724 77160 30776
rect 77375 30767 77433 30773
rect 77375 30733 77387 30767
rect 77421 30764 77433 30767
rect 78108 30764 78114 30776
rect 77421 30736 78114 30764
rect 77421 30733 77433 30736
rect 77375 30727 77433 30733
rect 78108 30724 78114 30736
rect 78166 30724 78172 30776
rect 78494 30773 78522 30804
rect 80687 30801 80699 30835
rect 80733 30832 80745 30835
rect 80776 30832 80782 30844
rect 80733 30804 80782 30832
rect 80733 30801 80745 30804
rect 80687 30795 80745 30801
rect 80776 30792 80782 30804
rect 80834 30792 80840 30844
rect 80960 30832 80966 30844
rect 80921 30804 80966 30832
rect 80960 30792 80966 30804
rect 81018 30832 81024 30844
rect 81512 30832 81518 30844
rect 81018 30804 81518 30832
rect 81018 30792 81024 30804
rect 81512 30792 81518 30804
rect 81570 30792 81576 30844
rect 82064 30832 82070 30844
rect 82025 30804 82070 30832
rect 82064 30792 82070 30804
rect 82122 30792 82128 30844
rect 84750 30841 84778 30872
rect 84735 30835 84793 30841
rect 84735 30801 84747 30835
rect 84781 30801 84793 30835
rect 84842 30832 84870 30928
rect 85762 30909 85790 30940
rect 87676 30928 87682 30940
rect 87734 30968 87740 30980
rect 88507 30971 88565 30977
rect 88507 30968 88519 30971
rect 87734 30940 88519 30968
rect 87734 30928 87740 30940
rect 88507 30937 88519 30940
rect 88553 30937 88565 30971
rect 89700 30968 89706 30980
rect 89661 30940 89706 30968
rect 88507 30931 88565 30937
rect 89700 30928 89706 30940
rect 89758 30928 89764 30980
rect 85747 30903 85805 30909
rect 85747 30869 85759 30903
rect 85793 30869 85805 30903
rect 85747 30863 85805 30869
rect 88231 30903 88289 30909
rect 88231 30869 88243 30903
rect 88277 30900 88289 30903
rect 89240 30900 89246 30912
rect 88277 30872 89246 30900
rect 88277 30869 88289 30872
rect 88231 30863 88289 30869
rect 89240 30860 89246 30872
rect 89298 30860 89304 30912
rect 85931 30835 85989 30841
rect 85931 30832 85943 30835
rect 84842 30804 85943 30832
rect 84735 30795 84793 30801
rect 85931 30801 85943 30804
rect 85977 30801 85989 30835
rect 88412 30832 88418 30844
rect 88373 30804 88418 30832
rect 85931 30795 85989 30801
rect 78479 30767 78537 30773
rect 78479 30733 78491 30767
rect 78525 30733 78537 30767
rect 78479 30727 78537 30733
rect 80135 30767 80193 30773
rect 80135 30733 80147 30767
rect 80181 30764 80193 30767
rect 81052 30764 81058 30776
rect 80181 30736 81058 30764
rect 80181 30733 80193 30736
rect 80135 30727 80193 30733
rect 81052 30724 81058 30736
rect 81110 30724 81116 30776
rect 81147 30767 81205 30773
rect 81147 30733 81159 30767
rect 81193 30733 81205 30767
rect 84750 30764 84778 30795
rect 88412 30792 88418 30804
rect 88470 30832 88476 30844
rect 88780 30832 88786 30844
rect 88470 30804 88786 30832
rect 88470 30792 88476 30804
rect 88780 30792 88786 30804
rect 88838 30832 88844 30844
rect 88875 30835 88933 30841
rect 88875 30832 88887 30835
rect 88838 30804 88887 30832
rect 88838 30792 88844 30804
rect 88875 30801 88887 30804
rect 88921 30801 88933 30835
rect 89608 30832 89614 30844
rect 89569 30804 89614 30832
rect 88875 30795 88933 30801
rect 89608 30792 89614 30804
rect 89666 30792 89672 30844
rect 90896 30792 90902 30844
rect 90954 30832 90960 30844
rect 91356 30832 91362 30844
rect 90954 30804 91362 30832
rect 90954 30792 90960 30804
rect 91356 30792 91362 30804
rect 91414 30792 91420 30844
rect 85011 30767 85069 30773
rect 85011 30764 85023 30767
rect 84750 30736 85023 30764
rect 81147 30727 81205 30733
rect 85011 30733 85023 30736
rect 85057 30764 85069 30767
rect 86756 30764 86762 30776
rect 85057 30736 86762 30764
rect 85057 30733 85069 30736
rect 85011 30727 85069 30733
rect 61272 30656 61278 30708
rect 61330 30696 61336 30708
rect 66056 30696 66062 30708
rect 61330 30668 66062 30696
rect 61330 30656 61336 30668
rect 66056 30656 66062 30668
rect 66114 30656 66120 30708
rect 74336 30656 74342 30708
rect 74394 30656 74400 30708
rect 74428 30656 74434 30708
rect 74486 30696 74492 30708
rect 74486 30668 75302 30696
rect 74486 30656 74492 30668
rect 67252 30628 67258 30640
rect 59726 30600 67258 30628
rect 67252 30588 67258 30600
rect 67310 30588 67316 30640
rect 69184 30628 69190 30640
rect 69145 30600 69190 30628
rect 69184 30588 69190 30600
rect 69242 30588 69248 30640
rect 75274 30628 75302 30668
rect 75440 30656 75446 30708
rect 75498 30696 75504 30708
rect 77004 30696 77010 30708
rect 75498 30668 77010 30696
rect 75498 30656 75504 30668
rect 77004 30656 77010 30668
rect 77062 30656 77068 30708
rect 80592 30656 80598 30708
rect 80650 30696 80656 30708
rect 81162 30696 81190 30727
rect 86756 30724 86762 30736
rect 86814 30724 86820 30776
rect 80650 30668 81190 30696
rect 80650 30656 80656 30668
rect 77740 30628 77746 30640
rect 75274 30600 77746 30628
rect 77740 30588 77746 30600
rect 77798 30588 77804 30640
rect 78016 30588 78022 30640
rect 78074 30628 78080 30640
rect 78844 30628 78850 30640
rect 78074 30600 78850 30628
rect 78074 30588 78080 30600
rect 78844 30588 78850 30600
rect 78902 30588 78908 30640
rect 86023 30631 86081 30637
rect 86023 30597 86035 30631
rect 86069 30628 86081 30631
rect 86112 30628 86118 30640
rect 86069 30600 86118 30628
rect 86069 30597 86081 30600
rect 86023 30591 86081 30597
rect 86112 30588 86118 30600
rect 86170 30588 86176 30640
rect 91448 30588 91454 30640
rect 91506 30628 91512 30640
rect 91543 30631 91601 30637
rect 91543 30628 91555 30631
rect 91506 30600 91555 30628
rect 91506 30588 91512 30600
rect 91543 30597 91555 30600
rect 91589 30597 91601 30631
rect 91543 30591 91601 30597
rect 538 30538 93642 30560
rect 538 30486 3680 30538
rect 3732 30486 3744 30538
rect 3796 30486 3808 30538
rect 3860 30486 3872 30538
rect 3924 30486 9008 30538
rect 9060 30486 9072 30538
rect 9124 30486 9136 30538
rect 9188 30486 9200 30538
rect 9252 30486 14336 30538
rect 14388 30486 14400 30538
rect 14452 30486 14464 30538
rect 14516 30486 14528 30538
rect 14580 30486 19664 30538
rect 19716 30486 19728 30538
rect 19780 30486 19792 30538
rect 19844 30486 19856 30538
rect 19908 30486 24992 30538
rect 25044 30486 25056 30538
rect 25108 30486 25120 30538
rect 25172 30486 25184 30538
rect 25236 30486 30320 30538
rect 30372 30486 30384 30538
rect 30436 30486 30448 30538
rect 30500 30486 30512 30538
rect 30564 30486 35648 30538
rect 35700 30486 35712 30538
rect 35764 30486 35776 30538
rect 35828 30486 35840 30538
rect 35892 30486 40976 30538
rect 41028 30486 41040 30538
rect 41092 30486 41104 30538
rect 41156 30486 41168 30538
rect 41220 30486 46304 30538
rect 46356 30486 46368 30538
rect 46420 30486 46432 30538
rect 46484 30486 46496 30538
rect 46548 30486 51632 30538
rect 51684 30486 51696 30538
rect 51748 30486 51760 30538
rect 51812 30486 51824 30538
rect 51876 30486 56960 30538
rect 57012 30486 57024 30538
rect 57076 30486 57088 30538
rect 57140 30486 57152 30538
rect 57204 30486 62288 30538
rect 62340 30486 62352 30538
rect 62404 30486 62416 30538
rect 62468 30486 62480 30538
rect 62532 30486 67616 30538
rect 67668 30486 67680 30538
rect 67732 30486 67744 30538
rect 67796 30486 67808 30538
rect 67860 30486 72944 30538
rect 72996 30486 73008 30538
rect 73060 30486 73072 30538
rect 73124 30486 73136 30538
rect 73188 30486 78272 30538
rect 78324 30486 78336 30538
rect 78388 30486 78400 30538
rect 78452 30486 78464 30538
rect 78516 30486 83600 30538
rect 83652 30486 83664 30538
rect 83716 30486 83728 30538
rect 83780 30486 83792 30538
rect 83844 30486 88928 30538
rect 88980 30486 88992 30538
rect 89044 30486 89056 30538
rect 89108 30486 89120 30538
rect 89172 30486 93642 30538
rect 538 30464 93642 30486
rect 3220 30424 3226 30436
rect 3181 30396 3226 30424
rect 3220 30384 3226 30396
rect 3278 30384 3284 30436
rect 5704 30384 5710 30436
rect 5762 30424 5768 30436
rect 18860 30424 18866 30436
rect 5762 30396 13202 30424
rect 5762 30384 5768 30396
rect 8007 30359 8065 30365
rect 8007 30325 8019 30359
rect 8053 30356 8065 30359
rect 8096 30356 8102 30368
rect 8053 30328 8102 30356
rect 8053 30325 8065 30328
rect 8007 30319 8065 30325
rect 8096 30316 8102 30328
rect 8154 30316 8160 30368
rect 8280 30316 8286 30368
rect 8338 30356 8344 30368
rect 9663 30359 9721 30365
rect 8338 30328 9430 30356
rect 8338 30316 8344 30328
rect 2392 30248 2398 30300
rect 2450 30288 2456 30300
rect 6443 30291 6501 30297
rect 2450 30260 3542 30288
rect 2450 30248 2456 30260
rect 1659 30223 1717 30229
rect 1659 30189 1671 30223
rect 1705 30189 1717 30223
rect 1659 30183 1717 30189
rect 1935 30223 1993 30229
rect 1935 30189 1947 30223
rect 1981 30220 1993 30223
rect 3036 30220 3042 30232
rect 1981 30192 3042 30220
rect 1981 30189 1993 30192
rect 1935 30183 1993 30189
rect 1674 30084 1702 30183
rect 3036 30180 3042 30192
rect 3094 30180 3100 30232
rect 3407 30155 3465 30161
rect 3407 30152 3419 30155
rect 2870 30124 3419 30152
rect 2870 30084 2898 30124
rect 3407 30121 3419 30124
rect 3453 30121 3465 30155
rect 3514 30152 3542 30260
rect 6443 30257 6455 30291
rect 6489 30288 6501 30291
rect 6900 30288 6906 30300
rect 6489 30260 6906 30288
rect 6489 30257 6501 30260
rect 6443 30251 6501 30257
rect 6900 30248 6906 30260
rect 6958 30248 6964 30300
rect 7084 30288 7090 30300
rect 7045 30260 7090 30288
rect 7084 30248 7090 30260
rect 7142 30248 7148 30300
rect 8651 30291 8709 30297
rect 8651 30257 8663 30291
rect 8697 30288 8709 30291
rect 9292 30288 9298 30300
rect 8697 30260 9298 30288
rect 8697 30257 8709 30260
rect 8651 30251 8709 30257
rect 9292 30248 9298 30260
rect 9350 30248 9356 30300
rect 9402 30288 9430 30328
rect 9663 30325 9675 30359
rect 9709 30356 9721 30359
rect 12604 30356 12610 30368
rect 9709 30328 12610 30356
rect 9709 30325 9721 30328
rect 9663 30319 9721 30325
rect 12604 30316 12610 30328
rect 12662 30316 12668 30368
rect 12328 30288 12334 30300
rect 9402 30260 12334 30288
rect 12328 30248 12334 30260
rect 12386 30288 12392 30300
rect 12386 30260 12650 30288
rect 12386 30248 12392 30260
rect 5060 30220 5066 30232
rect 5021 30192 5066 30220
rect 5060 30180 5066 30192
rect 5118 30180 5124 30232
rect 6256 30180 6262 30232
rect 6314 30220 6320 30232
rect 6351 30223 6409 30229
rect 6351 30220 6363 30223
rect 6314 30192 6363 30220
rect 6314 30180 6320 30192
rect 6351 30189 6363 30192
rect 6397 30189 6409 30223
rect 6351 30183 6409 30189
rect 6627 30223 6685 30229
rect 6627 30189 6639 30223
rect 6673 30220 6685 30223
rect 6808 30220 6814 30232
rect 6673 30192 6814 30220
rect 6673 30189 6685 30192
rect 6627 30183 6685 30189
rect 6808 30180 6814 30192
rect 6866 30220 6872 30232
rect 7728 30220 7734 30232
rect 6866 30192 7734 30220
rect 6866 30180 6872 30192
rect 7728 30180 7734 30192
rect 7786 30180 7792 30232
rect 7912 30220 7918 30232
rect 7873 30192 7918 30220
rect 7912 30180 7918 30192
rect 7970 30180 7976 30232
rect 8188 30220 8194 30232
rect 8149 30192 8194 30220
rect 8188 30180 8194 30192
rect 8246 30180 8252 30232
rect 9476 30220 9482 30232
rect 9437 30192 9482 30220
rect 9476 30180 9482 30192
rect 9534 30180 9540 30232
rect 12512 30220 12518 30232
rect 12473 30192 12518 30220
rect 12512 30180 12518 30192
rect 12570 30180 12576 30232
rect 12622 30229 12650 30260
rect 12607 30223 12665 30229
rect 12607 30189 12619 30223
rect 12653 30189 12665 30223
rect 12788 30220 12794 30232
rect 12749 30192 12794 30220
rect 12607 30183 12665 30189
rect 12788 30180 12794 30192
rect 12846 30180 12852 30232
rect 7930 30152 7958 30180
rect 11408 30152 11414 30164
rect 3514 30124 6854 30152
rect 7930 30124 11414 30152
rect 3407 30115 3465 30121
rect 2944 30084 2950 30096
rect 1674 30056 2950 30084
rect 2944 30044 2950 30056
rect 3002 30044 3008 30096
rect 5247 30087 5305 30093
rect 5247 30053 5259 30087
rect 5293 30084 5305 30087
rect 6716 30084 6722 30096
rect 5293 30056 6722 30084
rect 5293 30053 5305 30056
rect 5247 30047 5305 30053
rect 6716 30044 6722 30056
rect 6774 30044 6780 30096
rect 6826 30084 6854 30124
rect 11408 30112 11414 30124
rect 11466 30112 11472 30164
rect 11960 30152 11966 30164
rect 11921 30124 11966 30152
rect 11960 30112 11966 30124
rect 12018 30112 12024 30164
rect 13174 30152 13202 30396
rect 17590 30396 18866 30424
rect 13343 30291 13401 30297
rect 13343 30257 13355 30291
rect 13389 30288 13401 30291
rect 13619 30291 13677 30297
rect 13619 30288 13631 30291
rect 13389 30260 13631 30288
rect 13389 30257 13401 30260
rect 13343 30251 13401 30257
rect 13619 30257 13631 30260
rect 13665 30288 13677 30291
rect 17590 30288 17618 30396
rect 18860 30384 18866 30396
rect 18918 30424 18924 30436
rect 22359 30427 22417 30433
rect 22359 30424 22371 30427
rect 18918 30396 22371 30424
rect 18918 30384 18924 30396
rect 22359 30393 22371 30396
rect 22405 30424 22417 30427
rect 23828 30424 23834 30436
rect 22405 30396 23834 30424
rect 22405 30393 22417 30396
rect 22359 30387 22417 30393
rect 23828 30384 23834 30396
rect 23886 30384 23892 30436
rect 27140 30384 27146 30436
rect 27198 30424 27204 30436
rect 27419 30427 27477 30433
rect 27419 30424 27431 30427
rect 27198 30396 27431 30424
rect 27198 30384 27204 30396
rect 27419 30393 27431 30396
rect 27465 30393 27477 30427
rect 27419 30387 27477 30393
rect 27968 30384 27974 30436
rect 28026 30424 28032 30436
rect 36800 30424 36806 30436
rect 28026 30396 36806 30424
rect 28026 30384 28032 30396
rect 36800 30384 36806 30396
rect 36858 30384 36864 30436
rect 38091 30427 38149 30433
rect 38091 30393 38103 30427
rect 38137 30424 38149 30427
rect 38640 30424 38646 30436
rect 38137 30396 38646 30424
rect 38137 30393 38149 30396
rect 38091 30387 38149 30393
rect 38640 30384 38646 30396
rect 38698 30384 38704 30436
rect 42780 30384 42786 30436
rect 42838 30424 42844 30436
rect 48303 30427 48361 30433
rect 42838 30396 44206 30424
rect 42838 30384 42844 30396
rect 23644 30316 23650 30368
rect 23702 30356 23708 30368
rect 24012 30356 24018 30368
rect 23702 30328 24018 30356
rect 23702 30316 23708 30328
rect 24012 30316 24018 30328
rect 24070 30356 24076 30368
rect 24751 30359 24809 30365
rect 24751 30356 24763 30359
rect 24070 30328 24763 30356
rect 24070 30316 24076 30328
rect 13665 30260 17618 30288
rect 18219 30291 18277 30297
rect 13665 30257 13677 30260
rect 13619 30251 13677 30257
rect 18219 30257 18231 30291
rect 18265 30288 18277 30291
rect 18676 30288 18682 30300
rect 18265 30260 18682 30288
rect 18265 30257 18277 30260
rect 18219 30251 18277 30257
rect 18676 30248 18682 30260
rect 18734 30248 18740 30300
rect 19596 30288 19602 30300
rect 19557 30260 19602 30288
rect 19596 30248 19602 30260
rect 19654 30248 19660 30300
rect 23092 30288 23098 30300
rect 23053 30260 23098 30288
rect 23092 30248 23098 30260
rect 23150 30248 23156 30300
rect 24398 30297 24426 30328
rect 24751 30325 24763 30328
rect 24797 30356 24809 30359
rect 27692 30356 27698 30368
rect 24797 30328 27698 30356
rect 24797 30325 24809 30328
rect 24751 30319 24809 30325
rect 27692 30316 27698 30328
rect 27750 30316 27756 30368
rect 28336 30316 28342 30368
rect 28394 30356 28400 30368
rect 29348 30356 29354 30368
rect 28394 30328 29354 30356
rect 28394 30316 28400 30328
rect 29348 30316 29354 30328
rect 29406 30316 29412 30368
rect 30084 30316 30090 30368
rect 30142 30356 30148 30368
rect 30142 30328 40894 30356
rect 30142 30316 30148 30328
rect 24383 30291 24441 30297
rect 24383 30257 24395 30291
rect 24429 30257 24441 30291
rect 24383 30251 24441 30257
rect 27143 30291 27201 30297
rect 27143 30257 27155 30291
rect 27189 30288 27201 30291
rect 34040 30288 34046 30300
rect 27189 30260 34046 30288
rect 27189 30257 27201 30260
rect 27143 30251 27201 30257
rect 34040 30248 34046 30260
rect 34098 30288 34104 30300
rect 40866 30288 40894 30328
rect 40940 30316 40946 30368
rect 40998 30356 41004 30368
rect 43700 30356 43706 30368
rect 40998 30328 43706 30356
rect 40998 30316 41004 30328
rect 43700 30316 43706 30328
rect 43758 30316 43764 30368
rect 43976 30316 43982 30368
rect 44034 30356 44040 30368
rect 44034 30328 44079 30356
rect 44034 30316 44040 30328
rect 41127 30291 41185 30297
rect 41127 30288 41139 30291
rect 34098 30260 34362 30288
rect 34098 30248 34104 30260
rect 13251 30223 13309 30229
rect 13251 30189 13263 30223
rect 13297 30220 13309 30223
rect 17480 30220 17486 30232
rect 13297 30192 17486 30220
rect 13297 30189 13309 30192
rect 13251 30183 13309 30189
rect 17480 30180 17486 30192
rect 17538 30180 17544 30232
rect 17943 30223 18001 30229
rect 17943 30220 17955 30223
rect 17774 30192 17955 30220
rect 17774 30164 17802 30192
rect 17943 30189 17955 30192
rect 17989 30220 18001 30223
rect 18032 30220 18038 30232
rect 17989 30192 18038 30220
rect 17989 30189 18001 30192
rect 17943 30183 18001 30189
rect 18032 30180 18038 30192
rect 18090 30180 18096 30232
rect 23555 30223 23613 30229
rect 23555 30220 23567 30223
rect 22558 30192 23567 30220
rect 14720 30152 14726 30164
rect 13174 30124 14726 30152
rect 14720 30112 14726 30124
rect 14778 30112 14784 30164
rect 17756 30152 17762 30164
rect 17717 30124 17762 30152
rect 17756 30112 17762 30124
rect 17814 30112 17820 30164
rect 13156 30084 13162 30096
rect 6826 30056 13162 30084
rect 13156 30044 13162 30056
rect 13214 30044 13220 30096
rect 15916 30044 15922 30096
rect 15974 30084 15980 30096
rect 17388 30084 17394 30096
rect 15974 30056 17394 30084
rect 15974 30044 15980 30056
rect 17388 30044 17394 30056
rect 17446 30084 17452 30096
rect 22558 30093 22586 30192
rect 23555 30189 23567 30192
rect 23601 30220 23613 30223
rect 23644 30220 23650 30232
rect 23601 30192 23650 30220
rect 23601 30189 23613 30192
rect 23555 30183 23613 30189
rect 23644 30180 23650 30192
rect 23702 30180 23708 30232
rect 23739 30223 23797 30229
rect 23739 30189 23751 30223
rect 23785 30189 23797 30223
rect 23739 30183 23797 30189
rect 22816 30152 22822 30164
rect 22729 30124 22822 30152
rect 22816 30112 22822 30124
rect 22874 30152 22880 30164
rect 23754 30152 23782 30183
rect 23828 30180 23834 30232
rect 23886 30220 23892 30232
rect 23923 30223 23981 30229
rect 23923 30220 23935 30223
rect 23886 30192 23935 30220
rect 23886 30180 23892 30192
rect 23923 30189 23935 30192
rect 23969 30220 23981 30223
rect 24288 30220 24294 30232
rect 23969 30192 24294 30220
rect 23969 30189 23981 30192
rect 23923 30183 23981 30189
rect 24288 30180 24294 30192
rect 24346 30180 24352 30232
rect 24472 30220 24478 30232
rect 24433 30192 24478 30220
rect 24472 30180 24478 30192
rect 24530 30180 24536 30232
rect 27048 30220 27054 30232
rect 24582 30192 27054 30220
rect 24582 30152 24610 30192
rect 27048 30180 27054 30192
rect 27106 30180 27112 30232
rect 27235 30223 27293 30229
rect 27235 30220 27247 30223
rect 27158 30192 27247 30220
rect 27158 30152 27186 30192
rect 27235 30189 27247 30192
rect 27281 30189 27293 30223
rect 27235 30183 27293 30189
rect 27324 30180 27330 30232
rect 27382 30220 27388 30232
rect 34224 30220 34230 30232
rect 27382 30192 34230 30220
rect 27382 30180 27388 30192
rect 34224 30180 34230 30192
rect 34282 30180 34288 30232
rect 34334 30229 34362 30260
rect 36726 30260 37214 30288
rect 40866 30260 41139 30288
rect 34319 30223 34377 30229
rect 34319 30189 34331 30223
rect 34365 30189 34377 30223
rect 34319 30183 34377 30189
rect 22874 30124 24610 30152
rect 26974 30124 27186 30152
rect 22874 30112 22880 30124
rect 22543 30087 22601 30093
rect 22543 30084 22555 30087
rect 17446 30056 22555 30084
rect 17446 30044 17452 30056
rect 22543 30053 22555 30056
rect 22589 30053 22601 30087
rect 22543 30047 22601 30053
rect 23000 30044 23006 30096
rect 23058 30084 23064 30096
rect 26974 30093 27002 30124
rect 27416 30112 27422 30164
rect 27474 30152 27480 30164
rect 36726 30161 36754 30260
rect 36892 30220 36898 30232
rect 36853 30192 36898 30220
rect 36892 30180 36898 30192
rect 36950 30180 36956 30232
rect 37079 30223 37137 30229
rect 37079 30189 37091 30223
rect 37125 30189 37137 30223
rect 37186 30220 37214 30260
rect 41127 30257 41139 30260
rect 41173 30288 41185 30291
rect 41311 30291 41369 30297
rect 41311 30288 41323 30291
rect 41173 30260 41323 30288
rect 41173 30257 41185 30260
rect 41127 30251 41185 30257
rect 41311 30257 41323 30260
rect 41357 30288 41369 30291
rect 41495 30291 41553 30297
rect 41495 30288 41507 30291
rect 41357 30260 41507 30288
rect 41357 30257 41369 30260
rect 41311 30251 41369 30257
rect 41495 30257 41507 30260
rect 41541 30288 41553 30291
rect 42783 30291 42841 30297
rect 41541 30260 41814 30288
rect 41541 30257 41553 30260
rect 41495 30251 41553 30257
rect 37539 30223 37597 30229
rect 37539 30220 37551 30223
rect 37186 30192 37551 30220
rect 37079 30183 37137 30189
rect 37539 30189 37551 30192
rect 37585 30189 37597 30223
rect 37539 30183 37597 30189
rect 37631 30223 37689 30229
rect 37631 30189 37643 30223
rect 37677 30220 37689 30223
rect 41679 30223 41737 30229
rect 37677 30192 38686 30220
rect 37677 30189 37689 30192
rect 37631 30183 37689 30189
rect 36711 30155 36769 30161
rect 36711 30152 36723 30155
rect 27474 30124 36723 30152
rect 27474 30112 27480 30124
rect 36711 30121 36723 30124
rect 36757 30121 36769 30155
rect 36711 30115 36769 30121
rect 26959 30087 27017 30093
rect 26959 30084 26971 30087
rect 23058 30056 26971 30084
rect 23058 30044 23064 30056
rect 26959 30053 26971 30056
rect 27005 30084 27017 30087
rect 28888 30084 28894 30096
rect 27005 30056 28894 30084
rect 27005 30053 27017 30056
rect 26959 30047 27017 30053
rect 28888 30044 28894 30056
rect 28946 30044 28952 30096
rect 34408 30084 34414 30096
rect 34369 30056 34414 30084
rect 34408 30044 34414 30056
rect 34466 30044 34472 30096
rect 37094 30084 37122 30183
rect 38658 30096 38686 30192
rect 41679 30189 41691 30223
rect 41725 30189 41737 30223
rect 41786 30220 41814 30260
rect 42783 30257 42795 30291
rect 42829 30288 42841 30291
rect 44071 30291 44129 30297
rect 44071 30288 44083 30291
rect 42829 30260 44083 30288
rect 42829 30257 42841 30260
rect 42783 30251 42841 30257
rect 44071 30257 44083 30260
rect 44117 30257 44129 30291
rect 44178 30288 44206 30396
rect 48303 30393 48315 30427
rect 48349 30424 48361 30427
rect 48668 30424 48674 30436
rect 48349 30396 48674 30424
rect 48349 30393 48361 30396
rect 48303 30387 48361 30393
rect 48668 30384 48674 30396
rect 48726 30384 48732 30436
rect 62100 30424 62106 30436
rect 52274 30396 62106 30424
rect 44347 30359 44405 30365
rect 44347 30325 44359 30359
rect 44393 30356 44405 30359
rect 52274 30356 52302 30396
rect 62100 30384 62106 30396
rect 62158 30384 62164 30436
rect 62195 30427 62253 30433
rect 62195 30393 62207 30427
rect 62241 30424 62253 30427
rect 66979 30427 67037 30433
rect 66979 30424 66991 30427
rect 62241 30396 66991 30424
rect 62241 30393 62253 30396
rect 62195 30387 62253 30393
rect 66979 30393 66991 30396
rect 67025 30424 67037 30427
rect 67344 30424 67350 30436
rect 67025 30396 67350 30424
rect 67025 30393 67037 30396
rect 66979 30387 67037 30393
rect 67344 30384 67350 30396
rect 67402 30384 67408 30436
rect 70748 30424 70754 30436
rect 67454 30396 70754 30424
rect 53636 30356 53642 30368
rect 44393 30328 52302 30356
rect 53597 30328 53642 30356
rect 44393 30325 44405 30328
rect 44347 30319 44405 30325
rect 53636 30316 53642 30328
rect 53694 30316 53700 30368
rect 60168 30356 60174 30368
rect 58530 30328 60030 30356
rect 60081 30328 60174 30356
rect 47015 30291 47073 30297
rect 47015 30288 47027 30291
rect 44178 30260 47027 30288
rect 44071 30251 44129 30257
rect 47015 30257 47027 30260
rect 47061 30288 47073 30291
rect 47061 30260 47426 30288
rect 47061 30257 47073 30260
rect 47015 30251 47073 30257
rect 42139 30223 42197 30229
rect 42139 30220 42151 30223
rect 41786 30192 42151 30220
rect 41679 30183 41737 30189
rect 42139 30189 42151 30192
rect 42185 30189 42197 30223
rect 42139 30183 42197 30189
rect 42231 30223 42289 30229
rect 42231 30189 42243 30223
rect 42277 30220 42289 30223
rect 43700 30220 43706 30232
rect 42277 30192 43286 30220
rect 43661 30192 43706 30220
rect 42277 30189 42289 30192
rect 42231 30183 42289 30189
rect 41694 30152 41722 30183
rect 41694 30124 43102 30152
rect 43074 30096 43102 30124
rect 38180 30084 38186 30096
rect 37094 30056 38186 30084
rect 38180 30044 38186 30056
rect 38238 30084 38244 30096
rect 38367 30087 38425 30093
rect 38367 30084 38379 30087
rect 38238 30056 38379 30084
rect 38238 30044 38244 30056
rect 38367 30053 38379 30056
rect 38413 30053 38425 30087
rect 38640 30084 38646 30096
rect 38553 30056 38646 30084
rect 38367 30047 38425 30053
rect 38640 30044 38646 30056
rect 38698 30084 38704 30096
rect 39744 30084 39750 30096
rect 38698 30056 39750 30084
rect 38698 30044 38704 30056
rect 39744 30044 39750 30056
rect 39802 30044 39808 30096
rect 43056 30084 43062 30096
rect 43017 30056 43062 30084
rect 43056 30044 43062 30056
rect 43114 30044 43120 30096
rect 43258 30093 43286 30192
rect 43700 30180 43706 30192
rect 43758 30180 43764 30232
rect 43850 30223 43908 30229
rect 43850 30189 43862 30223
rect 43896 30220 43908 30223
rect 47107 30223 47165 30229
rect 47107 30220 47119 30223
rect 43896 30192 44114 30220
rect 43896 30189 43908 30192
rect 43850 30183 43908 30189
rect 44086 30164 44114 30192
rect 46754 30192 47119 30220
rect 44068 30112 44074 30164
rect 44126 30112 44132 30164
rect 43243 30087 43301 30093
rect 43243 30053 43255 30087
rect 43289 30084 43301 30087
rect 44160 30084 44166 30096
rect 43289 30056 44166 30084
rect 43289 30053 43301 30056
rect 43243 30047 43301 30053
rect 44160 30044 44166 30056
rect 44218 30044 44224 30096
rect 45356 30044 45362 30096
rect 45414 30084 45420 30096
rect 46754 30093 46782 30192
rect 47107 30189 47119 30192
rect 47153 30189 47165 30223
rect 47107 30183 47165 30189
rect 47291 30223 47349 30229
rect 47291 30189 47303 30223
rect 47337 30189 47349 30223
rect 47398 30220 47426 30260
rect 53912 30248 53918 30300
rect 53970 30288 53976 30300
rect 58530 30297 58558 30328
rect 58239 30291 58297 30297
rect 58239 30288 58251 30291
rect 53970 30260 58251 30288
rect 53970 30248 53976 30260
rect 58239 30257 58251 30260
rect 58285 30257 58297 30291
rect 58239 30251 58297 30257
rect 58515 30291 58573 30297
rect 58515 30257 58527 30291
rect 58561 30257 58573 30291
rect 59616 30288 59622 30300
rect 59577 30260 59622 30288
rect 58515 30251 58573 30257
rect 47751 30223 47809 30229
rect 47751 30220 47763 30223
rect 47398 30192 47763 30220
rect 47291 30183 47349 30189
rect 47751 30189 47763 30192
rect 47797 30189 47809 30223
rect 47751 30183 47809 30189
rect 47306 30152 47334 30183
rect 47840 30180 47846 30232
rect 47898 30220 47904 30232
rect 47898 30192 47943 30220
rect 47898 30180 47904 30192
rect 51060 30180 51066 30232
rect 51118 30220 51124 30232
rect 51980 30220 51986 30232
rect 51118 30192 51986 30220
rect 51118 30180 51124 30192
rect 51980 30180 51986 30192
rect 52038 30220 52044 30232
rect 52259 30223 52317 30229
rect 52259 30220 52271 30223
rect 52038 30192 52271 30220
rect 52038 30180 52044 30192
rect 52259 30189 52271 30192
rect 52305 30189 52317 30223
rect 52259 30183 52317 30189
rect 52535 30223 52593 30229
rect 52535 30189 52547 30223
rect 52581 30220 52593 30223
rect 52624 30220 52630 30232
rect 52581 30192 52630 30220
rect 52581 30189 52593 30192
rect 52535 30183 52593 30189
rect 48852 30152 48858 30164
rect 47306 30124 48858 30152
rect 48852 30112 48858 30124
rect 48910 30112 48916 30164
rect 46739 30087 46797 30093
rect 46739 30084 46751 30087
rect 45414 30056 46751 30084
rect 45414 30044 45420 30056
rect 46739 30053 46751 30056
rect 46785 30053 46797 30087
rect 52274 30084 52302 30183
rect 52624 30180 52630 30192
rect 52682 30180 52688 30232
rect 54004 30180 54010 30232
rect 54062 30220 54068 30232
rect 54927 30223 54985 30229
rect 54927 30220 54939 30223
rect 54062 30192 54939 30220
rect 54062 30180 54068 30192
rect 54927 30189 54939 30192
rect 54973 30189 54985 30223
rect 54927 30183 54985 30189
rect 54188 30112 54194 30164
rect 54246 30152 54252 30164
rect 54743 30155 54801 30161
rect 54743 30152 54755 30155
rect 54246 30124 54755 30152
rect 54246 30112 54252 30124
rect 54743 30121 54755 30124
rect 54789 30121 54801 30155
rect 58254 30152 58282 30251
rect 59616 30248 59622 30260
rect 59674 30248 59680 30300
rect 60002 30232 60030 30328
rect 60168 30316 60174 30328
rect 60226 30356 60232 30368
rect 63020 30356 63026 30368
rect 60226 30328 63026 30356
rect 60226 30316 60232 30328
rect 63020 30316 63026 30328
rect 63078 30316 63084 30368
rect 66056 30316 66062 30368
rect 66114 30356 66120 30368
rect 67454 30356 67482 30396
rect 70748 30384 70754 30396
rect 70806 30384 70812 30436
rect 70935 30427 70993 30433
rect 70935 30393 70947 30427
rect 70981 30424 70993 30427
rect 71024 30424 71030 30436
rect 70981 30396 71030 30424
rect 70981 30393 70993 30396
rect 70935 30387 70993 30393
rect 71024 30384 71030 30396
rect 71082 30424 71088 30436
rect 74428 30424 74434 30436
rect 71082 30396 74434 30424
rect 71082 30384 71088 30396
rect 74428 30384 74434 30396
rect 74486 30384 74492 30436
rect 74520 30384 74526 30436
rect 74578 30424 74584 30436
rect 76912 30424 76918 30436
rect 74578 30396 76918 30424
rect 74578 30384 74584 30396
rect 76912 30384 76918 30396
rect 76970 30384 76976 30436
rect 77096 30384 77102 30436
rect 77154 30424 77160 30436
rect 78016 30424 78022 30436
rect 77154 30396 78022 30424
rect 77154 30384 77160 30396
rect 78016 30384 78022 30396
rect 78074 30384 78080 30436
rect 82064 30384 82070 30436
rect 82122 30424 82128 30436
rect 82159 30427 82217 30433
rect 82159 30424 82171 30427
rect 82122 30396 82171 30424
rect 82122 30384 82128 30396
rect 82159 30393 82171 30396
rect 82205 30393 82217 30427
rect 86756 30424 86762 30436
rect 86717 30396 86762 30424
rect 82159 30387 82217 30393
rect 86756 30384 86762 30396
rect 86814 30384 86820 30436
rect 87955 30427 88013 30433
rect 87955 30393 87967 30427
rect 88001 30424 88013 30427
rect 89608 30424 89614 30436
rect 88001 30396 89614 30424
rect 88001 30393 88013 30396
rect 87955 30387 88013 30393
rect 89608 30384 89614 30396
rect 89666 30384 89672 30436
rect 91356 30384 91362 30436
rect 91414 30424 91420 30436
rect 92095 30427 92153 30433
rect 92095 30424 92107 30427
rect 91414 30396 92107 30424
rect 91414 30384 91420 30396
rect 92095 30393 92107 30396
rect 92141 30393 92153 30427
rect 92095 30387 92153 30393
rect 66114 30328 67482 30356
rect 66114 30316 66120 30328
rect 62284 30248 62290 30300
rect 62342 30288 62348 30300
rect 64403 30291 64461 30297
rect 64403 30288 64415 30291
rect 62342 30260 64415 30288
rect 62342 30248 62348 30260
rect 64403 30257 64415 30260
rect 64449 30288 64461 30291
rect 66516 30288 66522 30300
rect 64449 30260 66522 30288
rect 64449 30257 64461 30260
rect 64403 30251 64461 30257
rect 66516 30248 66522 30260
rect 66574 30248 66580 30300
rect 66608 30248 66614 30300
rect 66666 30288 66672 30300
rect 69828 30288 69834 30300
rect 66666 30260 69834 30288
rect 66666 30248 66672 30260
rect 69828 30248 69834 30260
rect 69886 30248 69892 30300
rect 70840 30288 70846 30300
rect 69938 30260 70846 30288
rect 69938 30232 69966 30260
rect 70840 30248 70846 30260
rect 70898 30288 70904 30300
rect 71119 30291 71177 30297
rect 71119 30288 71131 30291
rect 70898 30260 71131 30288
rect 70898 30248 70904 30260
rect 71119 30257 71131 30260
rect 71165 30257 71177 30291
rect 75532 30288 75538 30300
rect 71119 30251 71177 30257
rect 72146 30260 75538 30288
rect 58604 30220 58610 30232
rect 58565 30192 58610 30220
rect 58604 30180 58610 30192
rect 58662 30180 58668 30232
rect 59067 30223 59125 30229
rect 59067 30220 59079 30223
rect 58714 30192 59079 30220
rect 58714 30152 58742 30192
rect 59067 30189 59079 30192
rect 59113 30189 59125 30223
rect 59067 30183 59125 30189
rect 59156 30180 59162 30232
rect 59214 30220 59220 30232
rect 59984 30220 59990 30232
rect 59214 30192 59259 30220
rect 59945 30192 59990 30220
rect 59214 30180 59220 30192
rect 59984 30180 59990 30192
rect 60042 30180 60048 30232
rect 62379 30223 62437 30229
rect 62379 30189 62391 30223
rect 62425 30189 62437 30223
rect 62652 30220 62658 30232
rect 62613 30192 62658 30220
rect 62379 30183 62437 30189
rect 54743 30115 54801 30121
rect 54850 30124 55154 30152
rect 58254 30124 58742 30152
rect 54004 30084 54010 30096
rect 52274 30056 54010 30084
rect 46739 30047 46797 30053
rect 54004 30044 54010 30056
rect 54062 30044 54068 30096
rect 54096 30044 54102 30096
rect 54154 30084 54160 30096
rect 54850 30084 54878 30124
rect 55016 30084 55022 30096
rect 54154 30056 54878 30084
rect 54977 30056 55022 30084
rect 54154 30044 54160 30056
rect 55016 30044 55022 30056
rect 55074 30044 55080 30096
rect 55126 30084 55154 30124
rect 59524 30112 59530 30164
rect 59582 30152 59588 30164
rect 62394 30152 62422 30183
rect 62652 30180 62658 30192
rect 62710 30180 62716 30232
rect 64679 30223 64737 30229
rect 64679 30189 64691 30223
rect 64725 30220 64737 30223
rect 65780 30220 65786 30232
rect 64725 30192 65786 30220
rect 64725 30189 64737 30192
rect 64679 30183 64737 30189
rect 65780 30180 65786 30192
rect 65838 30180 65844 30232
rect 66884 30220 66890 30232
rect 66845 30192 66890 30220
rect 66884 30180 66890 30192
rect 66942 30180 66948 30232
rect 68819 30223 68877 30229
rect 68819 30189 68831 30223
rect 68865 30189 68877 30223
rect 69920 30220 69926 30232
rect 69881 30192 69926 30220
rect 68819 30183 68877 30189
rect 62560 30152 62566 30164
rect 59582 30124 62422 30152
rect 62521 30124 62566 30152
rect 59582 30112 59588 30124
rect 62195 30087 62253 30093
rect 62195 30084 62207 30087
rect 55126 30056 62207 30084
rect 62195 30053 62207 30056
rect 62241 30053 62253 30087
rect 62394 30084 62422 30124
rect 62560 30112 62566 30124
rect 62618 30112 62624 30164
rect 63112 30152 63118 30164
rect 63073 30124 63118 30152
rect 63112 30112 63118 30124
rect 63170 30112 63176 30164
rect 63940 30152 63946 30164
rect 63222 30124 63946 30152
rect 63222 30084 63250 30124
rect 63940 30112 63946 30124
rect 63998 30112 64004 30164
rect 65412 30112 65418 30164
rect 65470 30152 65476 30164
rect 67160 30152 67166 30164
rect 65470 30124 67166 30152
rect 65470 30112 65476 30124
rect 67160 30112 67166 30124
rect 67218 30112 67224 30164
rect 67252 30112 67258 30164
rect 67310 30152 67316 30164
rect 68632 30152 68638 30164
rect 67310 30124 68638 30152
rect 67310 30112 67316 30124
rect 68632 30112 68638 30124
rect 68690 30112 68696 30164
rect 68727 30155 68785 30161
rect 68727 30121 68739 30155
rect 68773 30152 68785 30155
rect 68834 30152 68862 30183
rect 69920 30180 69926 30192
rect 69978 30180 69984 30232
rect 71024 30220 71030 30232
rect 70985 30192 71030 30220
rect 71024 30180 71030 30192
rect 71082 30180 71088 30232
rect 72146 30229 72174 30260
rect 75532 30248 75538 30260
rect 75590 30288 75596 30300
rect 76912 30288 76918 30300
rect 75590 30260 76130 30288
rect 75590 30248 75596 30260
rect 72131 30223 72189 30229
rect 72131 30189 72143 30223
rect 72177 30189 72189 30223
rect 72312 30220 72318 30232
rect 72273 30192 72318 30220
rect 72131 30183 72189 30189
rect 72312 30180 72318 30192
rect 72370 30180 72376 30232
rect 72683 30223 72741 30229
rect 72683 30189 72695 30223
rect 72729 30220 72741 30223
rect 72772 30220 72778 30232
rect 72729 30192 72778 30220
rect 72729 30189 72741 30192
rect 72683 30183 72741 30189
rect 72772 30180 72778 30192
rect 72830 30180 72836 30232
rect 73876 30220 73882 30232
rect 73837 30192 73882 30220
rect 73876 30180 73882 30192
rect 73934 30220 73940 30232
rect 74247 30223 74305 30229
rect 74247 30220 74259 30223
rect 73934 30192 74259 30220
rect 73934 30180 73940 30192
rect 74247 30189 74259 30192
rect 74293 30220 74305 30223
rect 75992 30220 75998 30232
rect 74293 30192 75998 30220
rect 74293 30189 74305 30192
rect 74247 30183 74305 30189
rect 75992 30180 75998 30192
rect 76050 30180 76056 30232
rect 76102 30229 76130 30260
rect 76470 30260 76918 30288
rect 76087 30223 76145 30229
rect 76087 30189 76099 30223
rect 76133 30189 76145 30223
rect 76087 30183 76145 30189
rect 76176 30180 76182 30232
rect 76234 30220 76240 30232
rect 76470 30229 76498 30260
rect 76912 30248 76918 30260
rect 76970 30288 76976 30300
rect 77559 30291 77617 30297
rect 77559 30288 77571 30291
rect 76970 30260 77571 30288
rect 76970 30248 76976 30260
rect 77559 30257 77571 30260
rect 77605 30257 77617 30291
rect 77559 30251 77617 30257
rect 77740 30248 77746 30300
rect 77798 30288 77804 30300
rect 93288 30288 93294 30300
rect 77798 30260 93294 30288
rect 77798 30248 77804 30260
rect 93288 30248 93294 30260
rect 93346 30248 93352 30300
rect 76455 30223 76513 30229
rect 76234 30192 76279 30220
rect 76234 30180 76240 30192
rect 76455 30189 76467 30223
rect 76501 30189 76513 30223
rect 76636 30220 76642 30232
rect 76597 30192 76642 30220
rect 76455 30183 76513 30189
rect 76636 30180 76642 30192
rect 76694 30180 76700 30232
rect 77464 30220 77470 30232
rect 77425 30192 77470 30220
rect 77464 30180 77470 30192
rect 77522 30180 77528 30232
rect 80779 30223 80837 30229
rect 80779 30189 80791 30223
rect 80825 30189 80837 30223
rect 81052 30220 81058 30232
rect 81013 30192 81058 30220
rect 80779 30183 80837 30189
rect 71042 30152 71070 30180
rect 68773 30124 71070 30152
rect 72330 30152 72358 30180
rect 72867 30155 72925 30161
rect 72867 30152 72879 30155
rect 72330 30124 72879 30152
rect 68773 30121 68785 30124
rect 68727 30115 68785 30121
rect 72867 30121 72879 30124
rect 72913 30121 72925 30155
rect 72867 30115 72925 30121
rect 74063 30155 74121 30161
rect 74063 30121 74075 30155
rect 74109 30152 74121 30155
rect 75072 30152 75078 30164
rect 74109 30124 75078 30152
rect 74109 30121 74121 30124
rect 74063 30115 74121 30121
rect 75072 30112 75078 30124
rect 75130 30112 75136 30164
rect 75443 30155 75501 30161
rect 75443 30121 75455 30155
rect 75489 30152 75501 30155
rect 78016 30152 78022 30164
rect 75489 30124 78022 30152
rect 75489 30121 75501 30124
rect 75443 30115 75501 30121
rect 78016 30112 78022 30124
rect 78074 30112 78080 30164
rect 79764 30152 79770 30164
rect 78126 30124 79770 30152
rect 62394 30056 63250 30084
rect 62195 30047 62253 30053
rect 63388 30044 63394 30096
rect 63446 30084 63452 30096
rect 65783 30087 65841 30093
rect 65783 30084 65795 30087
rect 63446 30056 65795 30084
rect 63446 30044 63452 30056
rect 65783 30053 65795 30056
rect 65829 30053 65841 30087
rect 65783 30047 65841 30053
rect 67712 30044 67718 30096
rect 67770 30084 67776 30096
rect 69003 30087 69061 30093
rect 69003 30084 69015 30087
rect 67770 30056 69015 30084
rect 67770 30044 67776 30056
rect 69003 30053 69015 30056
rect 69049 30053 69061 30087
rect 69003 30047 69061 30053
rect 70012 30044 70018 30096
rect 70070 30084 70076 30096
rect 70107 30087 70165 30093
rect 70107 30084 70119 30087
rect 70070 30056 70119 30084
rect 70070 30044 70076 30056
rect 70107 30053 70119 30056
rect 70153 30053 70165 30087
rect 70107 30047 70165 30053
rect 70748 30044 70754 30096
rect 70806 30084 70812 30096
rect 74152 30084 74158 30096
rect 70806 30056 74158 30084
rect 70806 30044 70812 30056
rect 74152 30044 74158 30056
rect 74210 30044 74216 30096
rect 74336 30084 74342 30096
rect 74297 30056 74342 30084
rect 74336 30044 74342 30056
rect 74394 30044 74400 30096
rect 74704 30044 74710 30096
rect 74762 30084 74768 30096
rect 75348 30084 75354 30096
rect 74762 30056 75354 30084
rect 74762 30044 74768 30056
rect 75348 30044 75354 30056
rect 75406 30044 75412 30096
rect 75900 30044 75906 30096
rect 75958 30084 75964 30096
rect 78126 30084 78154 30124
rect 79764 30112 79770 30124
rect 79822 30112 79828 30164
rect 75958 30056 78154 30084
rect 75958 30044 75964 30056
rect 79488 30044 79494 30096
rect 79546 30084 79552 30096
rect 80687 30087 80745 30093
rect 80687 30084 80699 30087
rect 79546 30056 80699 30084
rect 79546 30044 79552 30056
rect 80687 30053 80699 30056
rect 80733 30084 80745 30087
rect 80794 30084 80822 30183
rect 81052 30180 81058 30192
rect 81110 30180 81116 30232
rect 85379 30223 85437 30229
rect 85379 30220 85391 30223
rect 85210 30192 85391 30220
rect 85210 30096 85238 30192
rect 85379 30189 85391 30192
rect 85425 30189 85437 30223
rect 85379 30183 85437 30189
rect 85655 30223 85713 30229
rect 85655 30189 85667 30223
rect 85701 30220 85713 30223
rect 86020 30220 86026 30232
rect 85701 30192 86026 30220
rect 85701 30189 85713 30192
rect 85655 30183 85713 30189
rect 86020 30180 86026 30192
rect 86078 30180 86084 30232
rect 88504 30220 88510 30232
rect 88465 30192 88510 30220
rect 88504 30180 88510 30192
rect 88562 30180 88568 30232
rect 88599 30223 88657 30229
rect 88599 30189 88611 30223
rect 88645 30189 88657 30223
rect 88599 30183 88657 30189
rect 85192 30084 85198 30096
rect 80733 30056 85198 30084
rect 80733 30053 80745 30056
rect 80687 30047 80745 30053
rect 85192 30044 85198 30056
rect 85250 30044 85256 30096
rect 87584 30044 87590 30096
rect 87642 30084 87648 30096
rect 87679 30087 87737 30093
rect 87679 30084 87691 30087
rect 87642 30056 87691 30084
rect 87642 30044 87648 30056
rect 87679 30053 87691 30056
rect 87725 30084 87737 30087
rect 88614 30084 88642 30183
rect 88780 30180 88786 30232
rect 88838 30220 88844 30232
rect 88875 30223 88933 30229
rect 88875 30220 88887 30223
rect 88838 30192 88887 30220
rect 88838 30180 88844 30192
rect 88875 30189 88887 30192
rect 88921 30189 88933 30223
rect 88875 30183 88933 30189
rect 89059 30223 89117 30229
rect 89059 30189 89071 30223
rect 89105 30220 89117 30223
rect 89240 30220 89246 30232
rect 89105 30192 89246 30220
rect 89105 30189 89117 30192
rect 89059 30183 89117 30189
rect 88890 30152 88918 30183
rect 89240 30180 89246 30192
rect 89298 30180 89304 30232
rect 90436 30180 90442 30232
rect 90494 30220 90500 30232
rect 90623 30223 90681 30229
rect 90623 30220 90635 30223
rect 90494 30192 90635 30220
rect 90494 30180 90500 30192
rect 90623 30189 90635 30192
rect 90669 30220 90681 30223
rect 90715 30223 90773 30229
rect 90715 30220 90727 30223
rect 90669 30192 90727 30220
rect 90669 30189 90681 30192
rect 90623 30183 90681 30189
rect 90715 30189 90727 30192
rect 90761 30189 90773 30223
rect 90988 30220 90994 30232
rect 90949 30192 90994 30220
rect 90715 30183 90773 30189
rect 90988 30180 90994 30192
rect 91046 30180 91052 30232
rect 89151 30155 89209 30161
rect 89151 30152 89163 30155
rect 88890 30124 89163 30152
rect 89151 30121 89163 30124
rect 89197 30121 89209 30155
rect 89151 30115 89209 30121
rect 87725 30056 88642 30084
rect 87725 30053 87737 30056
rect 87679 30047 87737 30053
rect 538 29994 93642 30016
rect 538 29942 6344 29994
rect 6396 29942 6408 29994
rect 6460 29942 6472 29994
rect 6524 29942 6536 29994
rect 6588 29942 11672 29994
rect 11724 29942 11736 29994
rect 11788 29942 11800 29994
rect 11852 29942 11864 29994
rect 11916 29942 17000 29994
rect 17052 29942 17064 29994
rect 17116 29942 17128 29994
rect 17180 29942 17192 29994
rect 17244 29942 22328 29994
rect 22380 29942 22392 29994
rect 22444 29942 22456 29994
rect 22508 29942 22520 29994
rect 22572 29942 27656 29994
rect 27708 29942 27720 29994
rect 27772 29942 27784 29994
rect 27836 29942 27848 29994
rect 27900 29942 32984 29994
rect 33036 29942 33048 29994
rect 33100 29942 33112 29994
rect 33164 29942 33176 29994
rect 33228 29942 38312 29994
rect 38364 29942 38376 29994
rect 38428 29942 38440 29994
rect 38492 29942 38504 29994
rect 38556 29942 43640 29994
rect 43692 29942 43704 29994
rect 43756 29942 43768 29994
rect 43820 29942 43832 29994
rect 43884 29942 48968 29994
rect 49020 29942 49032 29994
rect 49084 29942 49096 29994
rect 49148 29942 49160 29994
rect 49212 29942 54296 29994
rect 54348 29942 54360 29994
rect 54412 29942 54424 29994
rect 54476 29942 54488 29994
rect 54540 29942 59624 29994
rect 59676 29942 59688 29994
rect 59740 29942 59752 29994
rect 59804 29942 59816 29994
rect 59868 29942 64952 29994
rect 65004 29942 65016 29994
rect 65068 29942 65080 29994
rect 65132 29942 65144 29994
rect 65196 29942 70280 29994
rect 70332 29942 70344 29994
rect 70396 29942 70408 29994
rect 70460 29942 70472 29994
rect 70524 29942 75608 29994
rect 75660 29942 75672 29994
rect 75724 29942 75736 29994
rect 75788 29942 75800 29994
rect 75852 29942 80936 29994
rect 80988 29942 81000 29994
rect 81052 29942 81064 29994
rect 81116 29942 81128 29994
rect 81180 29942 86264 29994
rect 86316 29942 86328 29994
rect 86380 29942 86392 29994
rect 86444 29942 86456 29994
rect 86508 29942 91592 29994
rect 91644 29942 91656 29994
rect 91708 29942 91720 29994
rect 91772 29942 91784 29994
rect 91836 29942 93642 29994
rect 538 29920 93642 29942
rect 11408 29840 11414 29892
rect 11466 29880 11472 29892
rect 11595 29883 11653 29889
rect 11595 29880 11607 29883
rect 11466 29852 11607 29880
rect 11466 29840 11472 29852
rect 11595 29849 11607 29852
rect 11641 29849 11653 29883
rect 12239 29883 12297 29889
rect 12239 29880 12251 29883
rect 11595 29843 11653 29849
rect 11702 29852 12251 29880
rect 5704 29812 5710 29824
rect 5665 29784 5710 29812
rect 5704 29772 5710 29784
rect 5762 29772 5768 29824
rect 8096 29772 8102 29824
rect 8154 29812 8160 29824
rect 9295 29815 9353 29821
rect 9295 29812 9307 29815
rect 8154 29784 9307 29812
rect 8154 29772 8160 29784
rect 9295 29781 9307 29784
rect 9341 29781 9353 29815
rect 9476 29812 9482 29824
rect 9437 29784 9482 29812
rect 9295 29775 9353 29781
rect 9476 29772 9482 29784
rect 9534 29772 9540 29824
rect 10304 29772 10310 29824
rect 10362 29812 10368 29824
rect 11503 29815 11561 29821
rect 11503 29812 11515 29815
rect 10362 29784 11515 29812
rect 10362 29772 10368 29784
rect 11503 29781 11515 29784
rect 11549 29781 11561 29815
rect 11503 29775 11561 29781
rect 6164 29744 6170 29756
rect 6125 29716 6170 29744
rect 6164 29704 6170 29716
rect 6222 29704 6228 29756
rect 6348 29744 6354 29756
rect 6309 29716 6354 29744
rect 6348 29704 6354 29716
rect 6406 29704 6412 29756
rect 6440 29704 6446 29756
rect 6498 29744 6504 29756
rect 6627 29747 6685 29753
rect 6627 29744 6639 29747
rect 6498 29716 6639 29744
rect 6498 29704 6504 29716
rect 6627 29713 6639 29716
rect 6673 29744 6685 29747
rect 6716 29744 6722 29756
rect 6673 29716 6722 29744
rect 6673 29713 6685 29716
rect 6627 29707 6685 29713
rect 6716 29704 6722 29716
rect 6774 29744 6780 29756
rect 7179 29747 7237 29753
rect 6774 29716 7130 29744
rect 6774 29704 6780 29716
rect 6182 29676 6210 29704
rect 6811 29679 6869 29685
rect 6811 29676 6823 29679
rect 6182 29648 6823 29676
rect 6811 29645 6823 29648
rect 6857 29645 6869 29679
rect 7102 29676 7130 29716
rect 7179 29713 7191 29747
rect 7225 29744 7237 29747
rect 8004 29744 8010 29756
rect 7225 29716 8010 29744
rect 7225 29713 7237 29716
rect 7179 29707 7237 29713
rect 8004 29704 8010 29716
rect 8062 29704 8068 29756
rect 8188 29704 8194 29756
rect 8246 29744 8252 29756
rect 9384 29744 9390 29756
rect 8246 29716 9154 29744
rect 9345 29716 9390 29744
rect 8246 29704 8252 29716
rect 9126 29685 9154 29716
rect 9384 29704 9390 29716
rect 9442 29704 9448 29756
rect 11319 29747 11377 29753
rect 11319 29744 11331 29747
rect 9586 29716 11331 29744
rect 9111 29679 9169 29685
rect 7102 29648 9062 29676
rect 6811 29639 6869 29645
rect 9034 29608 9062 29648
rect 9111 29645 9123 29679
rect 9157 29676 9169 29679
rect 9586 29676 9614 29716
rect 11319 29713 11331 29716
rect 11365 29713 11377 29747
rect 11610 29744 11638 29843
rect 11702 29821 11730 29852
rect 12239 29849 12251 29852
rect 12285 29880 12297 29883
rect 13067 29883 13125 29889
rect 13067 29880 13079 29883
rect 12285 29852 13079 29880
rect 12285 29849 12297 29852
rect 12239 29843 12297 29849
rect 13067 29849 13079 29852
rect 13113 29880 13125 29883
rect 17480 29880 17486 29892
rect 13113 29852 17066 29880
rect 17441 29852 17486 29880
rect 13113 29849 13125 29852
rect 13067 29843 13125 29849
rect 11687 29815 11745 29821
rect 11687 29781 11699 29815
rect 11733 29781 11745 29815
rect 11687 29775 11745 29781
rect 12055 29815 12113 29821
rect 12055 29781 12067 29815
rect 12101 29812 12113 29815
rect 17038 29812 17066 29852
rect 17480 29840 17486 29852
rect 17538 29840 17544 29892
rect 18771 29883 18829 29889
rect 18771 29849 18783 29883
rect 18817 29880 18829 29883
rect 18952 29880 18958 29892
rect 18817 29852 18958 29880
rect 18817 29849 18829 29852
rect 18771 29843 18829 29849
rect 18952 29840 18958 29852
rect 19010 29880 19016 29892
rect 22724 29880 22730 29892
rect 19010 29852 22730 29880
rect 19010 29840 19016 29852
rect 22724 29840 22730 29852
rect 22782 29840 22788 29892
rect 27066 29852 28382 29880
rect 22816 29812 22822 29824
rect 12101 29784 16238 29812
rect 17038 29784 22822 29812
rect 12101 29781 12113 29784
rect 12055 29775 12113 29781
rect 12788 29744 12794 29756
rect 11610 29716 12794 29744
rect 11319 29707 11377 29713
rect 12788 29704 12794 29716
rect 12846 29704 12852 29756
rect 12883 29747 12941 29753
rect 12883 29713 12895 29747
rect 12929 29713 12941 29747
rect 12883 29707 12941 29713
rect 9844 29676 9850 29688
rect 9157 29648 9614 29676
rect 9805 29648 9850 29676
rect 9157 29645 9169 29648
rect 9111 29639 9169 29645
rect 9844 29636 9850 29648
rect 9902 29636 9908 29688
rect 9292 29608 9298 29620
rect 9034 29580 9298 29608
rect 9292 29568 9298 29580
rect 9350 29608 9356 29620
rect 10120 29608 10126 29620
rect 9350 29580 10126 29608
rect 9350 29568 9356 29580
rect 10120 29568 10126 29580
rect 10178 29568 10184 29620
rect 12898 29552 12926 29707
rect 13156 29704 13162 29756
rect 13214 29744 13220 29756
rect 15916 29744 15922 29756
rect 13214 29716 15922 29744
rect 13214 29704 13220 29716
rect 15916 29704 15922 29716
rect 15974 29704 15980 29756
rect 16103 29679 16161 29685
rect 16103 29676 16115 29679
rect 15934 29648 16115 29676
rect 4324 29500 4330 29552
rect 4382 29540 4388 29552
rect 8464 29540 8470 29552
rect 4382 29512 8470 29540
rect 4382 29500 4388 29512
rect 8464 29500 8470 29512
rect 8522 29500 8528 29552
rect 9476 29500 9482 29552
rect 9534 29540 9540 29552
rect 12880 29540 12886 29552
rect 9534 29512 12886 29540
rect 9534 29500 9540 29512
rect 12880 29500 12886 29512
rect 12938 29500 12944 29552
rect 15824 29500 15830 29552
rect 15882 29540 15888 29552
rect 15934 29549 15962 29648
rect 16103 29645 16115 29648
rect 16149 29645 16161 29679
rect 16210 29676 16238 29784
rect 22816 29772 22822 29784
rect 22874 29772 22880 29824
rect 23294 29784 23966 29812
rect 16376 29744 16382 29756
rect 16337 29716 16382 29744
rect 16376 29704 16382 29716
rect 16434 29704 16440 29756
rect 18679 29747 18737 29753
rect 18679 29713 18691 29747
rect 18725 29744 18737 29747
rect 19047 29747 19105 29753
rect 19047 29744 19059 29747
rect 18725 29716 19059 29744
rect 18725 29713 18737 29716
rect 18679 29707 18737 29713
rect 19047 29713 19059 29716
rect 19093 29744 19105 29747
rect 19596 29744 19602 29756
rect 19093 29716 19602 29744
rect 19093 29713 19105 29716
rect 19047 29707 19105 29713
rect 19596 29704 19602 29716
rect 19654 29704 19660 29756
rect 23294 29753 23322 29784
rect 23279 29747 23337 29753
rect 23279 29713 23291 29747
rect 23325 29713 23337 29747
rect 23279 29707 23337 29713
rect 23463 29747 23521 29753
rect 23463 29713 23475 29747
rect 23509 29713 23521 29747
rect 23736 29744 23742 29756
rect 23697 29716 23742 29744
rect 23463 29707 23521 29713
rect 17664 29676 17670 29688
rect 16210 29648 17670 29676
rect 16103 29639 16161 29645
rect 17664 29636 17670 29648
rect 17722 29636 17728 29688
rect 21804 29636 21810 29688
rect 21862 29676 21868 29688
rect 22911 29679 22969 29685
rect 22911 29676 22923 29679
rect 21862 29648 22923 29676
rect 21862 29636 21868 29648
rect 22911 29645 22923 29648
rect 22957 29676 22969 29679
rect 23478 29676 23506 29707
rect 23736 29704 23742 29716
rect 23794 29704 23800 29756
rect 23938 29685 23966 29784
rect 24288 29772 24294 29824
rect 24346 29812 24352 29824
rect 27066 29821 27094 29852
rect 27051 29815 27109 29821
rect 27051 29812 27063 29815
rect 24346 29784 27063 29812
rect 24346 29772 24352 29784
rect 27051 29781 27063 29784
rect 27097 29781 27109 29815
rect 27508 29812 27514 29824
rect 27469 29784 27514 29812
rect 27051 29775 27109 29781
rect 27508 29772 27514 29784
rect 27566 29772 27572 29824
rect 27600 29772 27606 29824
rect 27658 29812 27664 29824
rect 28354 29812 28382 29852
rect 28888 29840 28894 29892
rect 28946 29880 28952 29892
rect 33951 29883 34009 29889
rect 28946 29852 30590 29880
rect 28946 29840 28952 29852
rect 28612 29812 28618 29824
rect 27658 29784 28198 29812
rect 27658 29772 27664 29784
rect 28170 29756 28198 29784
rect 28354 29784 28618 29812
rect 24472 29704 24478 29756
rect 24530 29744 24536 29756
rect 24530 29716 27922 29744
rect 24530 29704 24536 29716
rect 22957 29648 23506 29676
rect 23923 29679 23981 29685
rect 22957 29645 22969 29648
rect 22911 29639 22969 29645
rect 23923 29645 23935 29679
rect 23969 29676 23981 29679
rect 24104 29676 24110 29688
rect 23969 29648 24110 29676
rect 23969 29645 23981 29648
rect 23923 29639 23981 29645
rect 24104 29636 24110 29648
rect 24162 29636 24168 29688
rect 27048 29636 27054 29688
rect 27106 29676 27112 29688
rect 27235 29679 27293 29685
rect 27235 29676 27247 29679
rect 27106 29648 27247 29676
rect 27106 29636 27112 29648
rect 27235 29645 27247 29648
rect 27281 29676 27293 29679
rect 27600 29676 27606 29688
rect 27281 29648 27606 29676
rect 27281 29645 27293 29648
rect 27235 29639 27293 29645
rect 27600 29636 27606 29648
rect 27658 29636 27664 29688
rect 27894 29676 27922 29716
rect 27968 29704 27974 29756
rect 28026 29744 28032 29756
rect 28152 29744 28158 29756
rect 28026 29716 28071 29744
rect 28113 29716 28158 29744
rect 28026 29704 28032 29716
rect 28152 29704 28158 29716
rect 28210 29704 28216 29756
rect 28354 29753 28382 29784
rect 28612 29772 28618 29784
rect 28670 29812 28676 29824
rect 29627 29815 29685 29821
rect 29627 29812 29639 29815
rect 28670 29784 29639 29812
rect 28670 29772 28676 29784
rect 29627 29781 29639 29784
rect 29673 29781 29685 29815
rect 30084 29812 30090 29824
rect 29627 29775 29685 29781
rect 29826 29784 30090 29812
rect 28339 29747 28397 29753
rect 28339 29713 28351 29747
rect 28385 29713 28397 29747
rect 28704 29744 28710 29756
rect 28665 29716 28710 29744
rect 28339 29707 28397 29713
rect 28704 29704 28710 29716
rect 28762 29744 28768 29756
rect 29072 29744 29078 29756
rect 28762 29716 29078 29744
rect 28762 29704 28768 29716
rect 29072 29704 29078 29716
rect 29130 29704 29136 29756
rect 28891 29679 28949 29685
rect 28891 29676 28903 29679
rect 27894 29648 28903 29676
rect 28891 29645 28903 29648
rect 28937 29676 28949 29679
rect 29164 29676 29170 29688
rect 28937 29648 29170 29676
rect 28937 29645 28949 29648
rect 28891 29639 28949 29645
rect 29164 29636 29170 29648
rect 29222 29636 29228 29688
rect 29642 29676 29670 29775
rect 29826 29753 29854 29784
rect 30084 29772 30090 29784
rect 30142 29812 30148 29824
rect 30455 29815 30513 29821
rect 30455 29812 30467 29815
rect 30142 29784 30467 29812
rect 30142 29772 30148 29784
rect 30455 29781 30467 29784
rect 30501 29781 30513 29815
rect 30455 29775 30513 29781
rect 29811 29747 29869 29753
rect 29811 29713 29823 29747
rect 29857 29713 29869 29747
rect 29811 29707 29869 29713
rect 29903 29747 29961 29753
rect 29903 29713 29915 29747
rect 29949 29713 29961 29747
rect 30562 29744 30590 29852
rect 33951 29849 33963 29883
rect 33997 29880 34009 29883
rect 34224 29880 34230 29892
rect 33997 29852 34230 29880
rect 33997 29849 34009 29852
rect 33951 29843 34009 29849
rect 34224 29840 34230 29852
rect 34282 29840 34288 29892
rect 34960 29880 34966 29892
rect 34334 29852 34966 29880
rect 30820 29772 30826 29824
rect 30878 29812 30884 29824
rect 32111 29815 32169 29821
rect 32111 29812 32123 29815
rect 30878 29784 32123 29812
rect 30878 29772 30884 29784
rect 32111 29781 32123 29784
rect 32157 29781 32169 29815
rect 34135 29815 34193 29821
rect 34135 29812 34147 29815
rect 32111 29775 32169 29781
rect 33782 29784 34147 29812
rect 33782 29753 33810 29784
rect 34135 29781 34147 29784
rect 34181 29812 34193 29815
rect 34334 29812 34362 29852
rect 34960 29840 34966 29852
rect 35018 29840 35024 29892
rect 37352 29880 37358 29892
rect 37313 29852 37358 29880
rect 37352 29840 37358 29852
rect 37410 29840 37416 29892
rect 39747 29883 39805 29889
rect 39747 29849 39759 29883
rect 39793 29880 39805 29883
rect 40940 29880 40946 29892
rect 39793 29852 40946 29880
rect 39793 29849 39805 29852
rect 39747 29843 39805 29849
rect 40940 29840 40946 29852
rect 40998 29840 41004 29892
rect 43056 29840 43062 29892
rect 43114 29880 43120 29892
rect 43976 29880 43982 29892
rect 43114 29852 43746 29880
rect 43937 29852 43982 29880
rect 43114 29840 43120 29852
rect 34181 29784 34362 29812
rect 34181 29781 34193 29784
rect 34135 29775 34193 29781
rect 34408 29772 34414 29824
rect 34466 29812 34472 29824
rect 34466 29784 38962 29812
rect 34466 29772 34472 29784
rect 31651 29747 31709 29753
rect 31651 29744 31663 29747
rect 30562 29716 31663 29744
rect 29903 29707 29961 29713
rect 31651 29713 31663 29716
rect 31697 29744 31709 29747
rect 32203 29747 32261 29753
rect 32203 29744 32215 29747
rect 31697 29716 32215 29744
rect 31697 29713 31709 29716
rect 31651 29707 31709 29713
rect 32203 29713 32215 29716
rect 32249 29713 32261 29747
rect 32203 29707 32261 29713
rect 33767 29747 33825 29753
rect 33767 29713 33779 29747
rect 33813 29713 33825 29747
rect 36892 29744 36898 29756
rect 33767 29707 33825 29713
rect 34058 29716 36898 29744
rect 29918 29676 29946 29707
rect 29642 29648 29946 29676
rect 30084 29636 30090 29688
rect 30142 29676 30148 29688
rect 30363 29679 30421 29685
rect 30363 29676 30375 29679
rect 30142 29648 30375 29676
rect 30142 29636 30148 29648
rect 30363 29645 30375 29648
rect 30409 29645 30421 29679
rect 30363 29639 30421 29645
rect 31559 29679 31617 29685
rect 31559 29645 31571 29679
rect 31605 29676 31617 29679
rect 34058 29676 34086 29716
rect 36892 29704 36898 29716
rect 36950 29744 36956 29756
rect 37263 29747 37321 29753
rect 37263 29744 37275 29747
rect 36950 29716 37275 29744
rect 36950 29704 36956 29716
rect 37263 29713 37275 29716
rect 37309 29713 37321 29747
rect 37263 29707 37321 29713
rect 37352 29704 37358 29756
rect 37410 29744 37416 29756
rect 38551 29747 38609 29753
rect 38551 29744 38563 29747
rect 37410 29716 38563 29744
rect 37410 29704 37416 29716
rect 38551 29713 38563 29716
rect 38597 29713 38609 29747
rect 38551 29707 38609 29713
rect 38735 29747 38793 29753
rect 38735 29713 38747 29747
rect 38781 29744 38793 29747
rect 38824 29744 38830 29756
rect 38781 29716 38830 29744
rect 38781 29713 38793 29716
rect 38735 29707 38793 29713
rect 38824 29704 38830 29716
rect 38882 29704 38888 29756
rect 31605 29648 34086 29676
rect 31605 29645 31617 29648
rect 31559 29639 31617 29645
rect 34500 29636 34506 29688
rect 34558 29676 34564 29688
rect 34558 29648 38502 29676
rect 34558 29636 34564 29648
rect 17296 29568 17302 29620
rect 17354 29608 17360 29620
rect 22816 29608 22822 29620
rect 17354 29580 22822 29608
rect 17354 29568 17360 29580
rect 22816 29568 22822 29580
rect 22874 29568 22880 29620
rect 23184 29568 23190 29620
rect 23242 29608 23248 29620
rect 24656 29608 24662 29620
rect 23242 29580 24662 29608
rect 23242 29568 23248 29580
rect 24656 29568 24662 29580
rect 24714 29568 24720 29620
rect 25852 29568 25858 29620
rect 25910 29608 25916 29620
rect 27327 29611 27385 29617
rect 27327 29608 27339 29611
rect 25910 29580 27339 29608
rect 25910 29568 25916 29580
rect 27327 29577 27339 29580
rect 27373 29608 27385 29611
rect 27968 29608 27974 29620
rect 27373 29580 27974 29608
rect 27373 29577 27385 29580
rect 27327 29571 27385 29577
rect 27968 29568 27974 29580
rect 28026 29568 28032 29620
rect 28152 29568 28158 29620
rect 28210 29608 28216 29620
rect 36340 29608 36346 29620
rect 28210 29580 36346 29608
rect 28210 29568 28216 29580
rect 36340 29568 36346 29580
rect 36398 29568 36404 29620
rect 15919 29543 15977 29549
rect 15919 29540 15931 29543
rect 15882 29512 15931 29540
rect 15882 29500 15888 29512
rect 15919 29509 15931 29512
rect 15965 29509 15977 29543
rect 15919 29503 15977 29509
rect 18308 29500 18314 29552
rect 18366 29540 18372 29552
rect 28980 29540 28986 29552
rect 18366 29512 28986 29540
rect 18366 29500 18372 29512
rect 28980 29500 28986 29512
rect 29038 29500 29044 29552
rect 29072 29500 29078 29552
rect 29130 29540 29136 29552
rect 29167 29543 29225 29549
rect 29167 29540 29179 29543
rect 29130 29512 29179 29540
rect 29130 29500 29136 29512
rect 29167 29509 29179 29512
rect 29213 29540 29225 29543
rect 37812 29540 37818 29552
rect 29213 29512 37818 29540
rect 29213 29509 29225 29512
rect 29167 29503 29225 29509
rect 37812 29500 37818 29512
rect 37870 29500 37876 29552
rect 38474 29549 38502 29648
rect 38934 29608 38962 29784
rect 39192 29744 39198 29756
rect 39153 29716 39198 29744
rect 39192 29704 39198 29716
rect 39250 29704 39256 29756
rect 39287 29747 39345 29753
rect 39287 29713 39299 29747
rect 39333 29744 39345 29747
rect 39468 29744 39474 29756
rect 39333 29716 39474 29744
rect 39333 29713 39345 29716
rect 39287 29707 39345 29713
rect 39468 29704 39474 29716
rect 39526 29704 39532 29756
rect 42415 29747 42473 29753
rect 42415 29713 42427 29747
rect 42461 29744 42473 29747
rect 42780 29744 42786 29756
rect 42461 29716 42786 29744
rect 42461 29713 42473 29716
rect 42415 29707 42473 29713
rect 42430 29676 42458 29707
rect 42780 29704 42786 29716
rect 42838 29704 42844 29756
rect 42967 29747 43025 29753
rect 42967 29713 42979 29747
rect 43013 29744 43025 29747
rect 43056 29744 43062 29756
rect 43013 29716 43062 29744
rect 43013 29713 43025 29716
rect 42967 29707 43025 29713
rect 43056 29704 43062 29716
rect 43114 29704 43120 29756
rect 43424 29744 43430 29756
rect 43166 29716 43430 29744
rect 39670 29648 42458 29676
rect 42599 29679 42657 29685
rect 39670 29608 39698 29648
rect 42599 29645 42611 29679
rect 42645 29676 42657 29679
rect 43166 29676 43194 29716
rect 43424 29704 43430 29716
rect 43482 29704 43488 29756
rect 43516 29704 43522 29756
rect 43574 29744 43580 29756
rect 43718 29744 43746 29852
rect 43976 29840 43982 29852
rect 44034 29840 44040 29892
rect 44160 29840 44166 29892
rect 44218 29880 44224 29892
rect 48763 29883 48821 29889
rect 48763 29880 48775 29883
rect 44218 29852 48775 29880
rect 44218 29840 44224 29852
rect 48763 29849 48775 29852
rect 48809 29849 48821 29883
rect 48763 29843 48821 29849
rect 48778 29812 48806 29843
rect 49404 29840 49410 29892
rect 49462 29880 49468 29892
rect 54096 29880 54102 29892
rect 49462 29852 54102 29880
rect 49462 29840 49468 29852
rect 54096 29840 54102 29852
rect 54154 29840 54160 29892
rect 54188 29840 54194 29892
rect 54246 29880 54252 29892
rect 54283 29883 54341 29889
rect 54283 29880 54295 29883
rect 54246 29852 54295 29880
rect 54246 29840 54252 29852
rect 54283 29849 54295 29852
rect 54329 29849 54341 29883
rect 54283 29843 54341 29849
rect 54648 29840 54654 29892
rect 54706 29880 54712 29892
rect 55847 29883 55905 29889
rect 55847 29880 55859 29883
rect 54706 29852 55859 29880
rect 54706 29840 54712 29852
rect 55847 29849 55859 29852
rect 55893 29849 55905 29883
rect 55847 29843 55905 29849
rect 57503 29883 57561 29889
rect 57503 29849 57515 29883
rect 57549 29849 57561 29883
rect 57503 29843 57561 29849
rect 50784 29812 50790 29824
rect 48778 29784 50790 29812
rect 50784 29772 50790 29784
rect 50842 29772 50848 29824
rect 50971 29815 51029 29821
rect 50971 29781 50983 29815
rect 51017 29812 51029 29815
rect 52440 29812 52446 29824
rect 51017 29784 52446 29812
rect 51017 29781 51029 29784
rect 50971 29775 51029 29781
rect 52440 29772 52446 29784
rect 52498 29772 52504 29824
rect 55016 29812 55022 29824
rect 52642 29784 55022 29812
rect 48579 29747 48637 29753
rect 48579 29744 48591 29747
rect 43574 29716 43619 29744
rect 43718 29716 48591 29744
rect 43574 29704 43580 29716
rect 48579 29713 48591 29716
rect 48625 29744 48637 29747
rect 48947 29747 49005 29753
rect 48947 29744 48959 29747
rect 48625 29716 48959 29744
rect 48625 29713 48637 29716
rect 48579 29707 48637 29713
rect 48947 29713 48959 29716
rect 48993 29744 49005 29747
rect 50692 29744 50698 29756
rect 48993 29716 50698 29744
rect 48993 29713 49005 29716
rect 48947 29707 49005 29713
rect 50692 29704 50698 29716
rect 50750 29704 50756 29756
rect 50876 29704 50882 29756
rect 50934 29744 50940 29756
rect 52642 29753 52670 29784
rect 55016 29772 55022 29784
rect 55074 29772 55080 29824
rect 57518 29812 57546 29843
rect 58604 29840 58610 29892
rect 58662 29880 58668 29892
rect 60168 29880 60174 29892
rect 58662 29852 60174 29880
rect 58662 29840 58668 29852
rect 60168 29840 60174 29852
rect 60226 29840 60232 29892
rect 60352 29880 60358 29892
rect 60313 29852 60358 29880
rect 60352 29840 60358 29852
rect 60410 29880 60416 29892
rect 61180 29880 61186 29892
rect 60410 29852 61186 29880
rect 60410 29840 60416 29852
rect 61180 29840 61186 29852
rect 61238 29840 61244 29892
rect 66792 29880 66798 29892
rect 66753 29852 66798 29880
rect 66792 29840 66798 29852
rect 66850 29840 66856 29892
rect 67899 29883 67957 29889
rect 67899 29849 67911 29883
rect 67945 29880 67957 29883
rect 74707 29883 74765 29889
rect 67945 29852 74658 29880
rect 67945 29849 67957 29852
rect 67899 29843 67957 29849
rect 65780 29812 65786 29824
rect 55586 29784 60582 29812
rect 65741 29784 65786 29812
rect 51155 29747 51213 29753
rect 51155 29744 51167 29747
rect 50934 29716 51167 29744
rect 50934 29704 50940 29716
rect 51155 29713 51167 29716
rect 51201 29713 51213 29747
rect 51155 29707 51213 29713
rect 51523 29747 51581 29753
rect 51523 29713 51535 29747
rect 51569 29744 51581 29747
rect 52535 29747 52593 29753
rect 52535 29744 52547 29747
rect 51569 29716 52547 29744
rect 51569 29713 51581 29716
rect 51523 29707 51581 29713
rect 52535 29713 52547 29716
rect 52581 29713 52593 29747
rect 52535 29707 52593 29713
rect 52627 29747 52685 29753
rect 52627 29713 52639 29747
rect 52673 29713 52685 29747
rect 52627 29707 52685 29713
rect 52808 29704 52814 29756
rect 52866 29744 52872 29756
rect 53820 29744 53826 29756
rect 52866 29716 53826 29744
rect 52866 29704 52872 29716
rect 53820 29704 53826 29716
rect 53878 29744 53884 29756
rect 54007 29747 54065 29753
rect 54007 29744 54019 29747
rect 53878 29716 54019 29744
rect 53878 29704 53884 29716
rect 54007 29713 54019 29716
rect 54053 29713 54065 29747
rect 54007 29707 54065 29713
rect 42645 29648 43194 29676
rect 42645 29645 42657 29648
rect 42599 29639 42657 29645
rect 38934 29580 39698 29608
rect 39744 29568 39750 29620
rect 39802 29608 39808 29620
rect 52256 29608 52262 29620
rect 39802 29580 52262 29608
rect 39802 29568 39808 29580
rect 52256 29568 52262 29580
rect 52314 29568 52320 29620
rect 53179 29611 53237 29617
rect 53179 29608 53191 29611
rect 52458 29580 53191 29608
rect 52458 29552 52486 29580
rect 53179 29577 53191 29580
rect 53225 29608 53237 29611
rect 53912 29608 53918 29620
rect 53225 29580 53918 29608
rect 53225 29577 53237 29580
rect 53179 29571 53237 29577
rect 53912 29568 53918 29580
rect 53970 29568 53976 29620
rect 54022 29608 54050 29707
rect 54096 29704 54102 29756
rect 54154 29744 54160 29756
rect 55586 29753 55614 29784
rect 54191 29747 54249 29753
rect 54191 29744 54203 29747
rect 54154 29716 54203 29744
rect 54154 29704 54160 29716
rect 54191 29713 54203 29716
rect 54237 29744 54249 29747
rect 54651 29747 54709 29753
rect 54651 29744 54663 29747
rect 54237 29716 54663 29744
rect 54237 29713 54249 29716
rect 54191 29707 54249 29713
rect 54651 29713 54663 29716
rect 54697 29713 54709 29747
rect 54651 29707 54709 29713
rect 55571 29747 55629 29753
rect 55571 29713 55583 29747
rect 55617 29713 55629 29747
rect 55571 29707 55629 29713
rect 55755 29747 55813 29753
rect 55755 29713 55767 29747
rect 55801 29744 55813 29747
rect 56396 29744 56402 29756
rect 55801 29716 56402 29744
rect 55801 29713 55813 29716
rect 55755 29707 55813 29713
rect 56396 29704 56402 29716
rect 56454 29704 56460 29756
rect 60554 29753 60582 29784
rect 65780 29772 65786 29784
rect 65838 29772 65844 29824
rect 66151 29815 66209 29821
rect 66151 29781 66163 29815
rect 66197 29812 66209 29815
rect 67914 29812 67942 29843
rect 66197 29784 67942 29812
rect 66197 29781 66209 29784
rect 66151 29775 66209 29781
rect 57687 29747 57745 29753
rect 57687 29713 57699 29747
rect 57733 29713 57745 29747
rect 57687 29707 57745 29713
rect 60539 29747 60597 29753
rect 60539 29713 60551 29747
rect 60585 29713 60597 29747
rect 60539 29707 60597 29713
rect 61367 29747 61425 29753
rect 61367 29713 61379 29747
rect 61413 29744 61425 29747
rect 62655 29747 62713 29753
rect 61413 29716 62606 29744
rect 61413 29713 61425 29716
rect 61367 29707 61425 29713
rect 57702 29676 57730 29707
rect 57871 29679 57929 29685
rect 57871 29676 57883 29679
rect 57702 29648 57883 29676
rect 57871 29645 57883 29648
rect 57917 29676 57929 29679
rect 61272 29676 61278 29688
rect 57917 29648 61278 29676
rect 57917 29645 57929 29648
rect 57871 29639 57929 29645
rect 61272 29636 61278 29648
rect 61330 29636 61336 29688
rect 62379 29679 62437 29685
rect 62379 29645 62391 29679
rect 62425 29645 62437 29679
rect 62578 29676 62606 29716
rect 62655 29713 62667 29747
rect 62701 29744 62713 29747
rect 63112 29744 63118 29756
rect 62701 29716 63118 29744
rect 62701 29713 62713 29716
rect 62655 29707 62713 29713
rect 63112 29704 63118 29716
rect 63170 29704 63176 29756
rect 65320 29744 65326 29756
rect 65233 29716 65326 29744
rect 65320 29704 65326 29716
rect 65378 29744 65384 29756
rect 65875 29747 65933 29753
rect 65875 29744 65887 29747
rect 65378 29716 65887 29744
rect 65378 29704 65384 29716
rect 65875 29713 65887 29716
rect 65921 29713 65933 29747
rect 65875 29707 65933 29713
rect 62744 29676 62750 29688
rect 62578 29648 62750 29676
rect 62379 29639 62437 29645
rect 54372 29608 54378 29620
rect 54022 29580 54378 29608
rect 54372 29568 54378 29580
rect 54430 29568 54436 29620
rect 54464 29568 54470 29620
rect 54522 29608 54528 29620
rect 60444 29608 60450 29620
rect 54522 29580 60450 29608
rect 54522 29568 54528 29580
rect 60444 29568 60450 29580
rect 60502 29568 60508 29620
rect 61180 29568 61186 29620
rect 61238 29608 61244 29620
rect 62284 29608 62290 29620
rect 61238 29580 62290 29608
rect 61238 29568 61244 29580
rect 62284 29568 62290 29580
rect 62342 29608 62348 29620
rect 62394 29608 62422 29639
rect 62744 29636 62750 29648
rect 62802 29676 62808 29688
rect 63759 29679 63817 29685
rect 63759 29676 63771 29679
rect 62802 29648 63771 29676
rect 62802 29636 62808 29648
rect 63759 29645 63771 29648
rect 63805 29645 63817 29679
rect 63759 29639 63817 29645
rect 65231 29679 65289 29685
rect 65231 29645 65243 29679
rect 65277 29676 65289 29679
rect 66166 29676 66194 29775
rect 68632 29772 68638 29824
rect 68690 29812 68696 29824
rect 68727 29815 68785 29821
rect 68727 29812 68739 29815
rect 68690 29784 68739 29812
rect 68690 29772 68696 29784
rect 68727 29781 68739 29784
rect 68773 29781 68785 29815
rect 68727 29775 68785 29781
rect 68926 29784 69322 29812
rect 66703 29747 66761 29753
rect 66703 29713 66715 29747
rect 66749 29744 66761 29747
rect 67436 29744 67442 29756
rect 66749 29716 67442 29744
rect 66749 29713 66761 29716
rect 66703 29707 66761 29713
rect 67436 29704 67442 29716
rect 67494 29704 67500 29756
rect 67712 29744 67718 29756
rect 67673 29716 67718 29744
rect 67712 29704 67718 29716
rect 67770 29704 67776 29756
rect 68926 29753 68954 29784
rect 68911 29747 68969 29753
rect 68911 29744 68923 29747
rect 67822 29716 68923 29744
rect 65277 29648 66194 29676
rect 65277 29645 65289 29648
rect 65231 29639 65289 29645
rect 67730 29608 67758 29704
rect 62342 29580 62422 29608
rect 67270 29580 67758 29608
rect 67822 29608 67850 29716
rect 68911 29713 68923 29716
rect 68957 29744 68969 29747
rect 69000 29744 69006 29756
rect 68957 29716 69006 29744
rect 68957 29713 68969 29716
rect 68911 29707 68969 29713
rect 69000 29704 69006 29716
rect 69058 29704 69064 29756
rect 69092 29704 69098 29756
rect 69150 29744 69156 29756
rect 69294 29753 69322 29784
rect 71392 29772 71398 29824
rect 71450 29812 71456 29824
rect 73235 29815 73293 29821
rect 73235 29812 73247 29815
rect 71450 29784 73247 29812
rect 71450 29772 71456 29784
rect 73235 29781 73247 29784
rect 73281 29781 73293 29815
rect 73235 29775 73293 29781
rect 74152 29772 74158 29824
rect 74210 29812 74216 29824
rect 74523 29815 74581 29821
rect 74523 29812 74535 29815
rect 74210 29784 74535 29812
rect 74210 29772 74216 29784
rect 74523 29781 74535 29784
rect 74569 29781 74581 29815
rect 74630 29812 74658 29852
rect 74707 29849 74719 29883
rect 74753 29880 74765 29883
rect 77372 29880 77378 29892
rect 74753 29852 77378 29880
rect 74753 29849 74765 29852
rect 74707 29843 74765 29849
rect 77372 29840 77378 29852
rect 77430 29880 77436 29892
rect 77740 29880 77746 29892
rect 77430 29852 77746 29880
rect 77430 29840 77436 29852
rect 77740 29840 77746 29852
rect 77798 29840 77804 29892
rect 78108 29880 78114 29892
rect 78069 29852 78114 29880
rect 78108 29840 78114 29852
rect 78166 29840 78172 29892
rect 79120 29840 79126 29892
rect 79178 29880 79184 29892
rect 79859 29883 79917 29889
rect 79859 29880 79871 29883
rect 79178 29852 79871 29880
rect 79178 29840 79184 29852
rect 79859 29849 79871 29852
rect 79905 29849 79917 29883
rect 79859 29843 79917 29849
rect 75900 29812 75906 29824
rect 74630 29784 75906 29812
rect 74523 29775 74581 29781
rect 69279 29747 69337 29753
rect 69150 29716 69243 29744
rect 69150 29704 69156 29716
rect 68632 29636 68638 29688
rect 68690 29676 68696 29688
rect 69202 29676 69230 29716
rect 69279 29713 69291 29747
rect 69325 29713 69337 29747
rect 70840 29744 70846 29756
rect 70801 29716 70846 29744
rect 69279 29707 69337 29713
rect 70840 29704 70846 29716
rect 70898 29704 70904 29756
rect 72683 29747 72741 29753
rect 72683 29713 72695 29747
rect 72729 29713 72741 29747
rect 72683 29707 72741 29713
rect 69644 29676 69650 29688
rect 68690 29648 69230 29676
rect 69605 29648 69650 29676
rect 68690 29636 68696 29648
rect 69644 29636 69650 29648
rect 69702 29636 69708 29688
rect 70012 29636 70018 29688
rect 70070 29676 70076 29688
rect 72698 29676 72726 29707
rect 72772 29704 72778 29756
rect 72830 29744 72836 29756
rect 74336 29744 74342 29756
rect 72830 29716 72875 29744
rect 72974 29716 74342 29744
rect 72830 29704 72836 29716
rect 72974 29676 73002 29716
rect 74336 29704 74342 29716
rect 74394 29704 74400 29756
rect 74538 29744 74566 29775
rect 75900 29772 75906 29784
rect 75958 29772 75964 29824
rect 75992 29772 75998 29824
rect 76050 29812 76056 29824
rect 76179 29815 76237 29821
rect 76179 29812 76191 29815
rect 76050 29784 76191 29812
rect 76050 29772 76056 29784
rect 76179 29781 76191 29784
rect 76225 29812 76237 29815
rect 76268 29812 76274 29824
rect 76225 29784 76274 29812
rect 76225 29781 76237 29784
rect 76179 29775 76237 29781
rect 76268 29772 76274 29784
rect 76326 29772 76332 29824
rect 76455 29815 76513 29821
rect 76455 29781 76467 29815
rect 76501 29812 76513 29815
rect 79672 29812 79678 29824
rect 76501 29784 79678 29812
rect 76501 29781 76513 29784
rect 76455 29775 76513 29781
rect 79672 29772 79678 29784
rect 79730 29772 79736 29824
rect 74867 29747 74925 29753
rect 74867 29744 74879 29747
rect 74538 29716 74879 29744
rect 74867 29713 74879 29716
rect 74913 29713 74925 29747
rect 74867 29707 74925 29713
rect 74980 29704 74986 29756
rect 75038 29744 75044 29756
rect 75038 29716 75083 29744
rect 75038 29704 75044 29716
rect 75164 29704 75170 29756
rect 75222 29744 75228 29756
rect 78016 29744 78022 29756
rect 75222 29716 75267 29744
rect 77977 29716 78022 29744
rect 75222 29704 75228 29716
rect 78016 29704 78022 29716
rect 78074 29704 78080 29756
rect 78936 29704 78942 29756
rect 78994 29744 79000 29756
rect 79031 29747 79089 29753
rect 79031 29744 79043 29747
rect 78994 29716 79043 29744
rect 78994 29704 79000 29716
rect 79031 29713 79043 29716
rect 79077 29744 79089 29747
rect 79307 29747 79365 29753
rect 79307 29744 79319 29747
rect 79077 29716 79319 29744
rect 79077 29713 79089 29716
rect 79031 29707 79089 29713
rect 79307 29713 79319 29716
rect 79353 29713 79365 29747
rect 79874 29744 79902 29843
rect 84088 29840 84094 29892
rect 84146 29880 84152 29892
rect 84275 29883 84333 29889
rect 84275 29880 84287 29883
rect 84146 29852 84287 29880
rect 84146 29840 84152 29852
rect 84275 29849 84287 29852
rect 84321 29880 84333 29883
rect 84548 29880 84554 29892
rect 84321 29852 84554 29880
rect 84321 29849 84333 29852
rect 84275 29843 84333 29849
rect 84548 29840 84554 29852
rect 84606 29840 84612 29892
rect 87768 29880 87774 29892
rect 87681 29852 87774 29880
rect 87768 29840 87774 29852
rect 87826 29880 87832 29892
rect 88504 29880 88510 29892
rect 87826 29852 88510 29880
rect 87826 29840 87832 29852
rect 88504 29840 88510 29852
rect 88562 29840 88568 29892
rect 80043 29815 80101 29821
rect 80043 29781 80055 29815
rect 80089 29812 80101 29815
rect 80316 29812 80322 29824
rect 80089 29784 80322 29812
rect 80089 29781 80101 29784
rect 80043 29775 80101 29781
rect 80316 29772 80322 29784
rect 80374 29772 80380 29824
rect 86023 29815 86081 29821
rect 86023 29781 86035 29815
rect 86069 29812 86081 29815
rect 86664 29812 86670 29824
rect 86069 29784 86670 29812
rect 86069 29781 86081 29784
rect 86023 29775 86081 29781
rect 86664 29772 86670 29784
rect 86722 29772 86728 29824
rect 80227 29747 80285 29753
rect 80227 29744 80239 29747
rect 79874 29716 80239 29744
rect 79307 29707 79365 29713
rect 80227 29713 80239 29716
rect 80273 29713 80285 29747
rect 84180 29744 84186 29756
rect 84141 29716 84186 29744
rect 80227 29707 80285 29713
rect 84180 29704 84186 29716
rect 84238 29744 84244 29756
rect 84459 29747 84517 29753
rect 84459 29744 84471 29747
rect 84238 29716 84471 29744
rect 84238 29704 84244 29716
rect 84459 29713 84471 29716
rect 84505 29713 84517 29747
rect 84459 29707 84517 29713
rect 86112 29704 86118 29756
rect 86170 29744 86176 29756
rect 87676 29744 87682 29756
rect 86170 29716 86215 29744
rect 87637 29716 87682 29744
rect 86170 29704 86176 29716
rect 87676 29704 87682 29716
rect 87734 29704 87740 29756
rect 90528 29744 90534 29756
rect 90489 29716 90534 29744
rect 90528 29704 90534 29716
rect 90586 29704 90592 29756
rect 90620 29704 90626 29756
rect 90678 29744 90684 29756
rect 90715 29747 90773 29753
rect 90715 29744 90727 29747
rect 90678 29716 90727 29744
rect 90678 29704 90684 29716
rect 90715 29713 90727 29716
rect 90761 29713 90773 29747
rect 90715 29707 90773 29713
rect 74704 29676 74710 29688
rect 70070 29648 72634 29676
rect 72698 29648 73002 29676
rect 73066 29648 74710 29676
rect 70070 29636 70076 29648
rect 68080 29608 68086 29620
rect 67822 29580 68086 29608
rect 62342 29568 62348 29580
rect 38459 29543 38517 29549
rect 38459 29509 38471 29543
rect 38505 29540 38517 29543
rect 39192 29540 39198 29552
rect 38505 29512 39198 29540
rect 38505 29509 38517 29512
rect 38459 29503 38517 29509
rect 39192 29500 39198 29512
rect 39250 29540 39256 29552
rect 46828 29540 46834 29552
rect 39250 29512 46834 29540
rect 39250 29500 39256 29512
rect 46828 29500 46834 29512
rect 46886 29500 46892 29552
rect 47840 29500 47846 29552
rect 47898 29540 47904 29552
rect 48392 29540 48398 29552
rect 47898 29512 48398 29540
rect 47898 29500 47904 29512
rect 48392 29500 48398 29512
rect 48450 29500 48456 29552
rect 52351 29543 52409 29549
rect 52351 29509 52363 29543
rect 52397 29540 52409 29543
rect 52440 29540 52446 29552
rect 52397 29512 52446 29540
rect 52397 29509 52409 29512
rect 52351 29503 52409 29509
rect 52440 29500 52446 29512
rect 52498 29500 52504 29552
rect 52624 29500 52630 29552
rect 52682 29540 52688 29552
rect 52811 29543 52869 29549
rect 52811 29540 52823 29543
rect 52682 29512 52823 29540
rect 52682 29500 52688 29512
rect 52811 29509 52823 29512
rect 52857 29509 52869 29543
rect 52811 29503 52869 29509
rect 54004 29500 54010 29552
rect 54062 29540 54068 29552
rect 55387 29543 55445 29549
rect 55387 29540 55399 29543
rect 54062 29512 55399 29540
rect 54062 29500 54068 29512
rect 55387 29509 55399 29512
rect 55433 29509 55445 29543
rect 55387 29503 55445 29509
rect 61459 29543 61517 29549
rect 61459 29509 61471 29543
rect 61505 29540 61517 29543
rect 62836 29540 62842 29552
rect 61505 29512 62842 29540
rect 61505 29509 61517 29512
rect 61459 29503 61517 29509
rect 62836 29500 62842 29512
rect 62894 29500 62900 29552
rect 63940 29500 63946 29552
rect 63998 29540 64004 29552
rect 67160 29540 67166 29552
rect 63998 29512 67166 29540
rect 63998 29500 64004 29512
rect 67160 29500 67166 29512
rect 67218 29540 67224 29552
rect 67270 29540 67298 29580
rect 67218 29512 67298 29540
rect 67218 29500 67224 29512
rect 67344 29500 67350 29552
rect 67402 29540 67408 29552
rect 67822 29540 67850 29580
rect 68080 29568 68086 29580
rect 68138 29568 68144 29620
rect 68172 29568 68178 29620
rect 68230 29608 68236 29620
rect 72315 29611 72373 29617
rect 72315 29608 72327 29611
rect 68230 29580 72327 29608
rect 68230 29568 68236 29580
rect 72315 29577 72327 29580
rect 72361 29608 72373 29611
rect 72499 29611 72557 29617
rect 72499 29608 72511 29611
rect 72361 29580 72511 29608
rect 72361 29577 72373 29580
rect 72315 29571 72373 29577
rect 72499 29577 72511 29580
rect 72545 29577 72557 29611
rect 72606 29608 72634 29648
rect 73066 29608 73094 29648
rect 74704 29636 74710 29648
rect 74762 29636 74768 29688
rect 75072 29636 75078 29688
rect 75130 29676 75136 29688
rect 75443 29679 75501 29685
rect 75443 29676 75455 29679
rect 75130 29648 75455 29676
rect 75130 29636 75136 29648
rect 75443 29645 75455 29648
rect 75489 29645 75501 29679
rect 75443 29639 75501 29645
rect 75532 29636 75538 29688
rect 75590 29676 75596 29688
rect 75992 29676 75998 29688
rect 75590 29648 75998 29676
rect 75590 29636 75596 29648
rect 75992 29636 75998 29648
rect 76050 29636 76056 29688
rect 76823 29679 76881 29685
rect 76823 29676 76835 29679
rect 76102 29648 76835 29676
rect 72606 29580 73094 29608
rect 72499 29571 72557 29577
rect 67402 29512 67850 29540
rect 67402 29500 67408 29512
rect 69552 29500 69558 29552
rect 69610 29540 69616 29552
rect 69736 29540 69742 29552
rect 69610 29512 69742 29540
rect 69610 29500 69616 29512
rect 69736 29500 69742 29512
rect 69794 29500 69800 29552
rect 71024 29540 71030 29552
rect 70985 29512 71030 29540
rect 71024 29500 71030 29512
rect 71082 29500 71088 29552
rect 72514 29540 72542 29571
rect 75164 29568 75170 29620
rect 75222 29608 75228 29620
rect 76102 29608 76130 29648
rect 76823 29645 76835 29648
rect 76869 29676 76881 29679
rect 76912 29676 76918 29688
rect 76869 29648 76918 29676
rect 76869 29645 76881 29648
rect 76823 29639 76881 29645
rect 76912 29636 76918 29648
rect 76970 29636 76976 29688
rect 77004 29636 77010 29688
rect 77062 29676 77068 29688
rect 79120 29676 79126 29688
rect 77062 29648 79126 29676
rect 77062 29636 77068 29648
rect 79120 29636 79126 29648
rect 79178 29636 79184 29688
rect 80592 29676 80598 29688
rect 80553 29648 80598 29676
rect 80592 29636 80598 29648
rect 80650 29636 80656 29688
rect 85747 29679 85805 29685
rect 85747 29676 85759 29679
rect 85670 29648 85759 29676
rect 75222 29580 76130 29608
rect 75222 29568 75228 29580
rect 76544 29568 76550 29620
rect 76602 29617 76608 29620
rect 76602 29611 76651 29617
rect 76602 29577 76605 29611
rect 76639 29577 76651 29611
rect 76602 29571 76651 29577
rect 76602 29568 76608 29571
rect 83168 29568 83174 29620
rect 83226 29608 83232 29620
rect 85670 29608 85698 29648
rect 85747 29645 85759 29648
rect 85793 29676 85805 29679
rect 85836 29676 85842 29688
rect 85793 29648 85842 29676
rect 85793 29645 85805 29648
rect 85747 29639 85805 29645
rect 85836 29636 85842 29648
rect 85894 29636 85900 29688
rect 86020 29636 86026 29688
rect 86078 29676 86084 29688
rect 86575 29679 86633 29685
rect 86575 29676 86587 29679
rect 86078 29648 86587 29676
rect 86078 29636 86084 29648
rect 86575 29645 86587 29648
rect 86621 29645 86633 29679
rect 86575 29639 86633 29645
rect 83226 29580 85698 29608
rect 83226 29568 83232 29580
rect 73232 29540 73238 29552
rect 72514 29512 73238 29540
rect 73232 29500 73238 29512
rect 73290 29500 73296 29552
rect 76268 29500 76274 29552
rect 76326 29540 76332 29552
rect 76731 29543 76789 29549
rect 76731 29540 76743 29543
rect 76326 29512 76743 29540
rect 76326 29500 76332 29512
rect 76731 29509 76743 29512
rect 76777 29509 76789 29543
rect 76912 29540 76918 29552
rect 76873 29512 76918 29540
rect 76731 29503 76789 29509
rect 76912 29500 76918 29512
rect 76970 29500 76976 29552
rect 90804 29540 90810 29552
rect 90765 29512 90810 29540
rect 90804 29500 90810 29512
rect 90862 29500 90868 29552
rect 538 29450 93642 29472
rect 538 29398 3680 29450
rect 3732 29398 3744 29450
rect 3796 29398 3808 29450
rect 3860 29398 3872 29450
rect 3924 29398 9008 29450
rect 9060 29398 9072 29450
rect 9124 29398 9136 29450
rect 9188 29398 9200 29450
rect 9252 29398 14336 29450
rect 14388 29398 14400 29450
rect 14452 29398 14464 29450
rect 14516 29398 14528 29450
rect 14580 29398 19664 29450
rect 19716 29398 19728 29450
rect 19780 29398 19792 29450
rect 19844 29398 19856 29450
rect 19908 29398 24992 29450
rect 25044 29398 25056 29450
rect 25108 29398 25120 29450
rect 25172 29398 25184 29450
rect 25236 29398 30320 29450
rect 30372 29398 30384 29450
rect 30436 29398 30448 29450
rect 30500 29398 30512 29450
rect 30564 29398 35648 29450
rect 35700 29398 35712 29450
rect 35764 29398 35776 29450
rect 35828 29398 35840 29450
rect 35892 29398 40976 29450
rect 41028 29398 41040 29450
rect 41092 29398 41104 29450
rect 41156 29398 41168 29450
rect 41220 29398 46304 29450
rect 46356 29398 46368 29450
rect 46420 29398 46432 29450
rect 46484 29398 46496 29450
rect 46548 29398 51632 29450
rect 51684 29398 51696 29450
rect 51748 29398 51760 29450
rect 51812 29398 51824 29450
rect 51876 29398 56960 29450
rect 57012 29398 57024 29450
rect 57076 29398 57088 29450
rect 57140 29398 57152 29450
rect 57204 29398 62288 29450
rect 62340 29398 62352 29450
rect 62404 29398 62416 29450
rect 62468 29398 62480 29450
rect 62532 29398 67616 29450
rect 67668 29398 67680 29450
rect 67732 29398 67744 29450
rect 67796 29398 67808 29450
rect 67860 29398 72944 29450
rect 72996 29398 73008 29450
rect 73060 29398 73072 29450
rect 73124 29398 73136 29450
rect 73188 29398 78272 29450
rect 78324 29398 78336 29450
rect 78388 29398 78400 29450
rect 78452 29398 78464 29450
rect 78516 29398 83600 29450
rect 83652 29398 83664 29450
rect 83716 29398 83728 29450
rect 83780 29398 83792 29450
rect 83844 29398 88928 29450
rect 88980 29398 88992 29450
rect 89044 29398 89056 29450
rect 89108 29398 89120 29450
rect 89172 29398 93642 29450
rect 538 29376 93642 29398
rect 3036 29336 3042 29348
rect 2997 29308 3042 29336
rect 3036 29296 3042 29308
rect 3094 29296 3100 29348
rect 8004 29296 8010 29348
rect 8062 29336 8068 29348
rect 8280 29336 8286 29348
rect 8062 29308 8286 29336
rect 8062 29296 8068 29308
rect 8280 29296 8286 29308
rect 8338 29296 8344 29348
rect 9384 29296 9390 29348
rect 9442 29336 9448 29348
rect 10396 29336 10402 29348
rect 9442 29308 10402 29336
rect 9442 29296 9448 29308
rect 10396 29296 10402 29308
rect 10454 29296 10460 29348
rect 12880 29296 12886 29348
rect 12938 29336 12944 29348
rect 12975 29339 13033 29345
rect 12975 29336 12987 29339
rect 12938 29308 12987 29336
rect 12938 29296 12944 29308
rect 12975 29305 12987 29308
rect 13021 29305 13033 29339
rect 12975 29299 13033 29305
rect 13251 29339 13309 29345
rect 13251 29305 13263 29339
rect 13297 29336 13309 29339
rect 13524 29336 13530 29348
rect 13297 29308 13530 29336
rect 13297 29305 13309 29308
rect 13251 29299 13309 29305
rect 4692 29228 4698 29280
rect 4750 29268 4756 29280
rect 4750 29240 7222 29268
rect 4750 29228 4756 29240
rect 6440 29200 6446 29212
rect 6401 29172 6446 29200
rect 6440 29160 6446 29172
rect 6498 29160 6504 29212
rect 7194 29209 7222 29240
rect 7179 29203 7237 29209
rect 7179 29169 7191 29203
rect 7225 29169 7237 29203
rect 7179 29163 7237 29169
rect 7728 29160 7734 29212
rect 7786 29200 7792 29212
rect 8007 29203 8065 29209
rect 8007 29200 8019 29203
rect 7786 29172 8019 29200
rect 7786 29160 7792 29172
rect 8007 29169 8019 29172
rect 8053 29200 8065 29203
rect 8188 29200 8194 29212
rect 8053 29172 8194 29200
rect 8053 29169 8065 29172
rect 8007 29163 8065 29169
rect 8188 29160 8194 29172
rect 8246 29160 8252 29212
rect 10120 29160 10126 29212
rect 10178 29200 10184 29212
rect 10215 29203 10273 29209
rect 10215 29200 10227 29203
rect 10178 29172 10227 29200
rect 10178 29160 10184 29172
rect 10215 29169 10227 29172
rect 10261 29169 10273 29203
rect 10414 29200 10442 29296
rect 10414 29172 10534 29200
rect 10215 29163 10273 29169
rect 1659 29135 1717 29141
rect 1659 29101 1671 29135
rect 1705 29101 1717 29135
rect 1659 29095 1717 29101
rect 1935 29135 1993 29141
rect 1935 29101 1947 29135
rect 1981 29132 1993 29135
rect 3036 29132 3042 29144
rect 1981 29104 3042 29132
rect 1981 29101 1993 29104
rect 1935 29095 1993 29101
rect 1674 28996 1702 29095
rect 3036 29092 3042 29104
rect 3094 29092 3100 29144
rect 6348 29092 6354 29144
rect 6406 29132 6412 29144
rect 6627 29135 6685 29141
rect 6627 29132 6639 29135
rect 6406 29104 6639 29132
rect 6406 29092 6412 29104
rect 6627 29101 6639 29104
rect 6673 29132 6685 29135
rect 6900 29132 6906 29144
rect 6673 29104 6906 29132
rect 6673 29101 6685 29104
rect 6627 29095 6685 29101
rect 6900 29092 6906 29104
rect 6958 29092 6964 29144
rect 8096 29132 8102 29144
rect 8057 29104 8102 29132
rect 8096 29092 8102 29104
rect 8154 29132 8160 29144
rect 10506 29141 10534 29172
rect 10399 29135 10457 29141
rect 10399 29132 10411 29135
rect 8154 29104 10411 29132
rect 8154 29092 8160 29104
rect 10399 29101 10411 29104
rect 10445 29101 10457 29135
rect 10399 29095 10457 29101
rect 10491 29135 10549 29141
rect 10491 29101 10503 29135
rect 10537 29101 10549 29135
rect 12883 29135 12941 29141
rect 10491 29095 10549 29101
rect 10598 29104 11178 29132
rect 6811 29067 6869 29073
rect 6811 29033 6823 29067
rect 6857 29064 6869 29067
rect 9476 29064 9482 29076
rect 6857 29036 9482 29064
rect 6857 29033 6869 29036
rect 6811 29027 6869 29033
rect 9476 29024 9482 29036
rect 9534 29024 9540 29076
rect 10598 29073 10626 29104
rect 10583 29067 10641 29073
rect 10583 29033 10595 29067
rect 10629 29033 10641 29067
rect 10948 29064 10954 29076
rect 10909 29036 10954 29064
rect 10583 29027 10641 29033
rect 10948 29024 10954 29036
rect 11006 29024 11012 29076
rect 11150 29073 11178 29104
rect 12883 29101 12895 29135
rect 12929 29132 12941 29135
rect 13266 29132 13294 29299
rect 13524 29296 13530 29308
rect 13582 29296 13588 29348
rect 19139 29339 19197 29345
rect 19139 29336 19151 29339
rect 18786 29308 19151 29336
rect 18786 29280 18814 29308
rect 19139 29305 19151 29308
rect 19185 29336 19197 29339
rect 19320 29336 19326 29348
rect 19185 29308 19326 29336
rect 19185 29305 19197 29308
rect 19139 29299 19197 29305
rect 19320 29296 19326 29308
rect 19378 29296 19384 29348
rect 19964 29296 19970 29348
rect 20022 29336 20028 29348
rect 22819 29339 22877 29345
rect 22819 29336 22831 29339
rect 20022 29308 22831 29336
rect 20022 29296 20028 29308
rect 22819 29305 22831 29308
rect 22865 29336 22877 29339
rect 23000 29336 23006 29348
rect 22865 29308 23006 29336
rect 22865 29305 22877 29308
rect 22819 29299 22877 29305
rect 23000 29296 23006 29308
rect 23058 29336 23064 29348
rect 23095 29339 23153 29345
rect 23095 29336 23107 29339
rect 23058 29308 23107 29336
rect 23058 29296 23064 29308
rect 23095 29305 23107 29308
rect 23141 29305 23153 29339
rect 23460 29336 23466 29348
rect 23421 29308 23466 29336
rect 23095 29299 23153 29305
rect 23460 29296 23466 29308
rect 23518 29296 23524 29348
rect 23736 29296 23742 29348
rect 23794 29336 23800 29348
rect 24383 29339 24441 29345
rect 24383 29336 24395 29339
rect 23794 29308 24395 29336
rect 23794 29296 23800 29308
rect 24383 29305 24395 29308
rect 24429 29305 24441 29339
rect 24383 29299 24441 29305
rect 24840 29296 24846 29348
rect 24898 29336 24904 29348
rect 36340 29336 36346 29348
rect 24898 29308 36202 29336
rect 36301 29308 36346 29336
rect 24898 29296 24904 29308
rect 18768 29268 18774 29280
rect 12929 29104 13294 29132
rect 13450 29240 18774 29268
rect 12929 29101 12941 29104
rect 12883 29095 12941 29101
rect 11135 29067 11193 29073
rect 11135 29033 11147 29067
rect 11181 29064 11193 29067
rect 13450 29064 13478 29240
rect 18768 29228 18774 29240
rect 18826 29228 18832 29280
rect 18952 29268 18958 29280
rect 18865 29240 18958 29268
rect 18952 29228 18958 29240
rect 19010 29268 19016 29280
rect 28152 29268 28158 29280
rect 19010 29240 28158 29268
rect 19010 29228 19016 29240
rect 28152 29228 28158 29240
rect 28210 29228 28216 29280
rect 28888 29268 28894 29280
rect 28849 29240 28894 29268
rect 28888 29228 28894 29240
rect 28946 29228 28952 29280
rect 28980 29228 28986 29280
rect 29038 29268 29044 29280
rect 31835 29271 31893 29277
rect 31835 29268 31847 29271
rect 29038 29240 31847 29268
rect 29038 29228 29044 29240
rect 31835 29237 31847 29240
rect 31881 29237 31893 29271
rect 31835 29231 31893 29237
rect 32292 29228 32298 29280
rect 32350 29268 32356 29280
rect 34132 29268 34138 29280
rect 32350 29240 34138 29268
rect 32350 29228 32356 29240
rect 34132 29228 34138 29240
rect 34190 29228 34196 29280
rect 36174 29268 36202 29308
rect 36340 29296 36346 29308
rect 36398 29296 36404 29348
rect 37720 29336 37726 29348
rect 37681 29308 37726 29336
rect 37720 29296 37726 29308
rect 37778 29296 37784 29348
rect 37812 29296 37818 29348
rect 37870 29336 37876 29348
rect 41219 29339 41277 29345
rect 41219 29336 41231 29339
rect 37870 29308 41231 29336
rect 37870 29296 37876 29308
rect 41219 29305 41231 29308
rect 41265 29336 41277 29339
rect 42228 29336 42234 29348
rect 41265 29308 42234 29336
rect 41265 29305 41277 29308
rect 41219 29299 41277 29305
rect 42228 29296 42234 29308
rect 42286 29296 42292 29348
rect 42783 29339 42841 29345
rect 42783 29305 42795 29339
rect 42829 29336 42841 29339
rect 44068 29336 44074 29348
rect 42829 29308 44074 29336
rect 42829 29305 42841 29308
rect 42783 29299 42841 29305
rect 44068 29296 44074 29308
rect 44126 29296 44132 29348
rect 47288 29296 47294 29348
rect 47346 29336 47352 29348
rect 48116 29336 48122 29348
rect 47346 29308 48122 29336
rect 47346 29296 47352 29308
rect 48116 29296 48122 29308
rect 48174 29296 48180 29348
rect 48300 29336 48306 29348
rect 48261 29308 48306 29336
rect 48300 29296 48306 29308
rect 48358 29296 48364 29348
rect 48392 29296 48398 29348
rect 48450 29336 48456 29348
rect 48576 29336 48582 29348
rect 48450 29308 48582 29336
rect 48450 29296 48456 29308
rect 48576 29296 48582 29308
rect 48634 29336 48640 29348
rect 50876 29336 50882 29348
rect 48634 29308 50882 29336
rect 48634 29296 48640 29308
rect 50876 29296 50882 29308
rect 50934 29296 50940 29348
rect 50968 29296 50974 29348
rect 51026 29336 51032 29348
rect 52811 29339 52869 29345
rect 52811 29336 52823 29339
rect 51026 29308 52823 29336
rect 51026 29296 51032 29308
rect 52811 29305 52823 29308
rect 52857 29336 52869 29339
rect 54096 29336 54102 29348
rect 52857 29308 54102 29336
rect 52857 29305 52869 29308
rect 52811 29299 52869 29305
rect 54096 29296 54102 29308
rect 54154 29296 54160 29348
rect 54280 29296 54286 29348
rect 54338 29336 54344 29348
rect 60352 29336 60358 29348
rect 54338 29308 60358 29336
rect 54338 29296 54344 29308
rect 60352 29296 60358 29308
rect 60410 29296 60416 29348
rect 60720 29296 60726 29348
rect 60778 29336 60784 29348
rect 62701 29339 62759 29345
rect 62701 29336 62713 29339
rect 60778 29308 62713 29336
rect 60778 29296 60784 29308
rect 62701 29305 62713 29308
rect 62747 29336 62759 29339
rect 62928 29336 62934 29348
rect 62747 29308 62934 29336
rect 62747 29305 62759 29308
rect 62701 29299 62759 29305
rect 62928 29296 62934 29308
rect 62986 29296 62992 29348
rect 67252 29296 67258 29348
rect 67310 29336 67316 29348
rect 67531 29339 67589 29345
rect 67531 29336 67543 29339
rect 67310 29308 67543 29336
rect 67310 29296 67316 29308
rect 67531 29305 67543 29308
rect 67577 29305 67589 29339
rect 67531 29299 67589 29305
rect 67807 29339 67865 29345
rect 67807 29305 67819 29339
rect 67853 29336 67865 29339
rect 68080 29336 68086 29348
rect 67853 29308 68086 29336
rect 67853 29305 67865 29308
rect 67807 29299 67865 29305
rect 68080 29296 68086 29308
rect 68138 29296 68144 29348
rect 86388 29336 86394 29348
rect 68190 29308 86394 29336
rect 36248 29268 36254 29280
rect 36174 29240 36254 29268
rect 36248 29228 36254 29240
rect 36306 29228 36312 29280
rect 16100 29160 16106 29212
rect 16158 29200 16164 29212
rect 22724 29200 22730 29212
rect 16158 29172 22730 29200
rect 16158 29160 16164 29172
rect 22724 29160 22730 29172
rect 22782 29160 22788 29212
rect 23095 29203 23153 29209
rect 23095 29169 23107 29203
rect 23141 29200 23153 29203
rect 23141 29172 23322 29200
rect 23141 29169 23153 29172
rect 23095 29163 23153 29169
rect 17480 29132 17486 29144
rect 17441 29104 17486 29132
rect 17480 29092 17486 29104
rect 17538 29092 17544 29144
rect 18768 29092 18774 29144
rect 18826 29132 18832 29144
rect 18863 29135 18921 29141
rect 18863 29132 18875 29135
rect 18826 29104 18875 29132
rect 18826 29092 18832 29104
rect 18863 29101 18875 29104
rect 18909 29101 18921 29135
rect 23000 29132 23006 29144
rect 18863 29095 18921 29101
rect 18970 29104 23006 29132
rect 18970 29064 18998 29104
rect 23000 29092 23006 29104
rect 23058 29092 23064 29144
rect 23184 29132 23190 29144
rect 23145 29104 23190 29132
rect 23184 29092 23190 29104
rect 23242 29092 23248 29144
rect 23294 29141 23322 29172
rect 23368 29160 23374 29212
rect 23426 29200 23432 29212
rect 23923 29203 23981 29209
rect 23923 29200 23935 29203
rect 23426 29172 23935 29200
rect 23426 29160 23432 29172
rect 23923 29169 23935 29172
rect 23969 29200 23981 29203
rect 24012 29200 24018 29212
rect 23969 29172 24018 29200
rect 23969 29169 23981 29172
rect 23923 29163 23981 29169
rect 24012 29160 24018 29172
rect 24070 29160 24076 29212
rect 24196 29160 24202 29212
rect 24254 29200 24260 29212
rect 28704 29200 28710 29212
rect 24254 29172 28710 29200
rect 24254 29160 24260 29172
rect 28704 29160 28710 29172
rect 28762 29160 28768 29212
rect 28906 29200 28934 29228
rect 28906 29172 29210 29200
rect 23279 29135 23337 29141
rect 23279 29101 23291 29135
rect 23325 29101 23337 29135
rect 23279 29095 23337 29101
rect 23736 29092 23742 29144
rect 23794 29132 23800 29144
rect 24567 29135 24625 29141
rect 24567 29132 24579 29135
rect 23794 29104 24579 29132
rect 23794 29092 23800 29104
rect 24567 29101 24579 29104
rect 24613 29101 24625 29135
rect 24567 29095 24625 29101
rect 24656 29092 24662 29144
rect 24714 29132 24720 29144
rect 28520 29132 28526 29144
rect 24714 29104 28526 29132
rect 24714 29092 24720 29104
rect 28520 29092 28526 29104
rect 28578 29092 28584 29144
rect 28799 29135 28857 29141
rect 28799 29101 28811 29135
rect 28845 29132 28857 29135
rect 29072 29132 29078 29144
rect 28845 29104 29078 29132
rect 28845 29101 28857 29104
rect 28799 29095 28857 29101
rect 29072 29092 29078 29104
rect 29130 29092 29136 29144
rect 29182 29141 29210 29172
rect 29532 29160 29538 29212
rect 29590 29200 29596 29212
rect 30087 29203 30145 29209
rect 30087 29200 30099 29203
rect 29590 29172 30099 29200
rect 29590 29160 29596 29172
rect 30087 29169 30099 29172
rect 30133 29200 30145 29203
rect 30176 29200 30182 29212
rect 30133 29172 30182 29200
rect 30133 29169 30145 29172
rect 30087 29163 30145 29169
rect 30176 29160 30182 29172
rect 30234 29200 30240 29212
rect 32016 29200 32022 29212
rect 30234 29172 31050 29200
rect 30234 29160 30240 29172
rect 29167 29135 29225 29141
rect 29167 29101 29179 29135
rect 29213 29101 29225 29135
rect 29167 29095 29225 29101
rect 29627 29135 29685 29141
rect 29627 29101 29639 29135
rect 29673 29132 29685 29135
rect 29992 29132 29998 29144
rect 29673 29104 29998 29132
rect 29673 29101 29685 29104
rect 29627 29095 29685 29101
rect 29992 29092 29998 29104
rect 30050 29092 30056 29144
rect 30452 29132 30458 29144
rect 30413 29104 30458 29132
rect 30452 29092 30458 29104
rect 30510 29092 30516 29144
rect 30820 29132 30826 29144
rect 30781 29104 30826 29132
rect 30820 29092 30826 29104
rect 30878 29092 30884 29144
rect 31022 29141 31050 29172
rect 31206 29172 32022 29200
rect 31206 29141 31234 29172
rect 32016 29160 32022 29172
rect 32074 29160 32080 29212
rect 36358 29200 36386 29296
rect 37260 29228 37266 29280
rect 37318 29268 37324 29280
rect 38275 29271 38333 29277
rect 38275 29268 38287 29271
rect 37318 29240 38287 29268
rect 37318 29228 37324 29240
rect 38275 29237 38287 29240
rect 38321 29268 38333 29271
rect 38640 29268 38646 29280
rect 38321 29240 38646 29268
rect 38321 29237 38333 29240
rect 38275 29231 38333 29237
rect 38640 29228 38646 29240
rect 38698 29228 38704 29280
rect 41602 29240 43378 29268
rect 36358 29172 36846 29200
rect 31007 29135 31065 29141
rect 31007 29101 31019 29135
rect 31053 29101 31065 29135
rect 31007 29095 31065 29101
rect 31191 29135 31249 29141
rect 31191 29101 31203 29135
rect 31237 29101 31249 29135
rect 31191 29095 31249 29101
rect 31280 29092 31286 29144
rect 31338 29132 31344 29144
rect 31375 29135 31433 29141
rect 31375 29132 31387 29135
rect 31338 29104 31387 29132
rect 31338 29092 31344 29104
rect 31375 29101 31387 29104
rect 31421 29101 31433 29135
rect 31375 29095 31433 29101
rect 33948 29092 33954 29144
rect 34006 29132 34012 29144
rect 35880 29132 35886 29144
rect 34006 29104 35886 29132
rect 34006 29092 34012 29104
rect 35880 29092 35886 29104
rect 35938 29092 35944 29144
rect 36156 29092 36162 29144
rect 36214 29132 36220 29144
rect 36527 29135 36585 29141
rect 36527 29132 36539 29135
rect 36214 29104 36539 29132
rect 36214 29092 36220 29104
rect 36527 29101 36539 29104
rect 36573 29101 36585 29135
rect 36708 29132 36714 29144
rect 36669 29104 36714 29132
rect 36527 29095 36585 29101
rect 36708 29092 36714 29104
rect 36766 29092 36772 29144
rect 36818 29132 36846 29172
rect 37812 29160 37818 29212
rect 37870 29200 37876 29212
rect 41602 29209 41630 29240
rect 41403 29203 41461 29209
rect 41403 29200 41415 29203
rect 37870 29172 41415 29200
rect 37870 29160 37876 29172
rect 41403 29169 41415 29172
rect 41449 29200 41461 29203
rect 41587 29203 41645 29209
rect 41587 29200 41599 29203
rect 41449 29172 41599 29200
rect 41449 29169 41461 29172
rect 41403 29163 41461 29169
rect 41587 29169 41599 29172
rect 41633 29169 41645 29203
rect 41587 29163 41645 29169
rect 37171 29135 37229 29141
rect 37171 29132 37183 29135
rect 36818 29104 37183 29132
rect 37171 29101 37183 29104
rect 37217 29101 37229 29135
rect 37171 29095 37229 29101
rect 37260 29092 37266 29144
rect 37318 29132 37324 29144
rect 38735 29135 38793 29141
rect 37318 29104 37363 29132
rect 37318 29092 37324 29104
rect 38735 29101 38747 29135
rect 38781 29132 38793 29135
rect 38824 29132 38830 29144
rect 38781 29104 38830 29132
rect 38781 29101 38793 29104
rect 38735 29095 38793 29101
rect 38824 29092 38830 29104
rect 38882 29092 38888 29144
rect 41768 29132 41774 29144
rect 41729 29104 41774 29132
rect 41768 29092 41774 29104
rect 41826 29092 41832 29144
rect 42228 29132 42234 29144
rect 42189 29104 42234 29132
rect 42228 29092 42234 29104
rect 42286 29092 42292 29144
rect 42320 29092 42326 29144
rect 42378 29132 42384 29144
rect 42378 29104 42423 29132
rect 42378 29092 42384 29104
rect 42964 29092 42970 29144
rect 43022 29132 43028 29144
rect 43243 29135 43301 29141
rect 43243 29132 43255 29135
rect 43022 29104 43255 29132
rect 43022 29092 43028 29104
rect 43243 29101 43255 29104
rect 43289 29101 43301 29135
rect 43350 29132 43378 29240
rect 44988 29228 44994 29280
rect 45046 29268 45052 29280
rect 45681 29271 45739 29277
rect 45681 29268 45693 29271
rect 45046 29240 45693 29268
rect 45046 29228 45052 29240
rect 45681 29237 45693 29240
rect 45727 29237 45739 29271
rect 45816 29268 45822 29280
rect 45777 29240 45822 29268
rect 45681 29231 45739 29237
rect 45816 29228 45822 29240
rect 45874 29228 45880 29280
rect 46000 29228 46006 29280
rect 46058 29268 46064 29280
rect 46058 29240 54510 29268
rect 46058 29228 46064 29240
rect 45448 29160 45454 29212
rect 45506 29200 45512 29212
rect 45911 29203 45969 29209
rect 45911 29200 45923 29203
rect 45506 29172 45923 29200
rect 45506 29160 45512 29172
rect 45911 29169 45923 29172
rect 45957 29169 45969 29203
rect 46828 29200 46834 29212
rect 46741 29172 46834 29200
rect 45911 29163 45969 29169
rect 46828 29160 46834 29172
rect 46886 29200 46892 29212
rect 47107 29203 47165 29209
rect 47107 29200 47119 29203
rect 46886 29172 47119 29200
rect 46886 29160 46892 29172
rect 47107 29169 47119 29172
rect 47153 29169 47165 29203
rect 47107 29163 47165 29169
rect 47214 29172 47518 29200
rect 46923 29135 46981 29141
rect 46923 29132 46935 29135
rect 43350 29104 46935 29132
rect 43243 29095 43301 29101
rect 46923 29101 46935 29104
rect 46969 29132 46981 29135
rect 47214 29132 47242 29172
rect 46969 29104 47242 29132
rect 46969 29101 46981 29104
rect 46923 29095 46981 29101
rect 47288 29092 47294 29144
rect 47346 29132 47352 29144
rect 47490 29132 47518 29172
rect 48300 29160 48306 29212
rect 48358 29200 48364 29212
rect 48484 29200 48490 29212
rect 48358 29172 48490 29200
rect 48358 29160 48364 29172
rect 48484 29160 48490 29172
rect 48542 29200 48548 29212
rect 52348 29200 52354 29212
rect 48542 29172 52354 29200
rect 48542 29160 48548 29172
rect 47751 29135 47809 29141
rect 47751 29132 47763 29135
rect 47346 29104 47391 29132
rect 47490 29104 47763 29132
rect 47346 29092 47352 29104
rect 47751 29101 47763 29104
rect 47797 29101 47809 29135
rect 47751 29095 47809 29101
rect 47843 29135 47901 29141
rect 47843 29101 47855 29135
rect 47889 29132 47901 29135
rect 48668 29132 48674 29144
rect 47889 29104 48674 29132
rect 47889 29101 47901 29104
rect 47843 29095 47901 29101
rect 48668 29092 48674 29104
rect 48726 29092 48732 29144
rect 49330 29141 49358 29172
rect 52348 29160 52354 29172
rect 52406 29160 52412 29212
rect 53547 29203 53605 29209
rect 53547 29200 53559 29203
rect 52458 29172 53559 29200
rect 49315 29135 49373 29141
rect 49315 29101 49327 29135
rect 49361 29101 49373 29135
rect 51152 29132 51158 29144
rect 51113 29104 51158 29132
rect 49315 29095 49373 29101
rect 51152 29092 51158 29104
rect 51210 29092 51216 29144
rect 51796 29092 51802 29144
rect 51854 29132 51860 29144
rect 52458 29132 52486 29172
rect 53547 29169 53559 29172
rect 53593 29200 53605 29203
rect 54280 29200 54286 29212
rect 53593 29172 54286 29200
rect 53593 29169 53605 29172
rect 53547 29163 53605 29169
rect 54280 29160 54286 29172
rect 54338 29160 54344 29212
rect 54482 29200 54510 29240
rect 54924 29228 54930 29280
rect 54982 29268 54988 29280
rect 59343 29271 59401 29277
rect 59343 29268 59355 29271
rect 54982 29240 59355 29268
rect 54982 29228 54988 29240
rect 59343 29237 59355 29240
rect 59389 29237 59401 29271
rect 59343 29231 59401 29237
rect 59987 29271 60045 29277
rect 59987 29237 59999 29271
rect 60033 29268 60045 29271
rect 60168 29268 60174 29280
rect 60033 29240 60174 29268
rect 60033 29237 60045 29240
rect 59987 29231 60045 29237
rect 60168 29228 60174 29240
rect 60226 29228 60232 29280
rect 68190 29268 68218 29308
rect 86388 29296 86394 29308
rect 86446 29296 86452 29348
rect 86664 29336 86670 29348
rect 86625 29308 86670 29336
rect 86664 29296 86670 29308
rect 86722 29296 86728 29348
rect 86756 29296 86762 29348
rect 86814 29336 86820 29348
rect 87035 29339 87093 29345
rect 87035 29336 87047 29339
rect 86814 29308 87047 29336
rect 86814 29296 86820 29308
rect 87035 29305 87047 29308
rect 87081 29305 87093 29339
rect 90988 29336 90994 29348
rect 90949 29308 90994 29336
rect 87035 29299 87093 29305
rect 90988 29296 90994 29308
rect 91046 29296 91052 29348
rect 61750 29240 68218 29268
rect 68650 29240 69230 29268
rect 58604 29200 58610 29212
rect 54482 29172 58190 29200
rect 51854 29104 52486 29132
rect 51854 29092 51860 29104
rect 52532 29092 52538 29144
rect 52590 29132 52596 29144
rect 53636 29132 53642 29144
rect 52590 29104 53642 29132
rect 52590 29092 52596 29104
rect 53636 29092 53642 29104
rect 53694 29092 53700 29144
rect 54007 29135 54065 29141
rect 54007 29101 54019 29135
rect 54053 29132 54065 29135
rect 54096 29132 54102 29144
rect 54053 29104 54102 29132
rect 54053 29101 54065 29104
rect 54007 29095 54065 29101
rect 54096 29092 54102 29104
rect 54154 29092 54160 29144
rect 54191 29135 54249 29141
rect 54191 29101 54203 29135
rect 54237 29132 54249 29135
rect 54372 29132 54378 29144
rect 54237 29104 54378 29132
rect 54237 29101 54249 29104
rect 54191 29095 54249 29101
rect 54372 29092 54378 29104
rect 54430 29092 54436 29144
rect 55019 29135 55077 29141
rect 55019 29101 55031 29135
rect 55065 29101 55077 29135
rect 55019 29095 55077 29101
rect 55111 29135 55169 29141
rect 55111 29101 55123 29135
rect 55157 29132 55169 29135
rect 55292 29132 55298 29144
rect 55157 29104 55298 29132
rect 55157 29101 55169 29104
rect 55111 29095 55169 29101
rect 33212 29064 33218 29076
rect 11181 29036 13478 29064
rect 13542 29036 18998 29064
rect 19062 29036 33218 29064
rect 11181 29033 11193 29036
rect 11135 29027 11193 29033
rect 2300 28996 2306 29008
rect 1674 28968 2306 28996
rect 2300 28956 2306 28968
rect 2358 28996 2364 29008
rect 2944 28996 2950 29008
rect 2358 28968 2950 28996
rect 2358 28956 2364 28968
rect 2944 28956 2950 28968
rect 3002 28996 3008 29008
rect 3407 28999 3465 29005
rect 3407 28996 3419 28999
rect 3002 28968 3419 28996
rect 3002 28956 3008 28968
rect 3407 28965 3419 28968
rect 3453 28965 3465 28999
rect 6716 28996 6722 29008
rect 6677 28968 6722 28996
rect 3407 28959 3465 28965
rect 6716 28956 6722 28968
rect 6774 28956 6780 29008
rect 11316 28956 11322 29008
rect 11374 28996 11380 29008
rect 13542 28996 13570 29036
rect 17572 28996 17578 29008
rect 11374 28968 13570 28996
rect 17485 28968 17578 28996
rect 11374 28956 11380 28968
rect 17572 28956 17578 28968
rect 17630 28996 17636 29008
rect 19062 28996 19090 29036
rect 33212 29024 33218 29036
rect 33270 29024 33276 29076
rect 37720 29024 37726 29076
rect 37778 29064 37784 29076
rect 38272 29064 38278 29076
rect 37778 29036 38278 29064
rect 37778 29024 37784 29036
rect 38272 29024 38278 29036
rect 38330 29024 38336 29076
rect 42246 29064 42274 29092
rect 45356 29064 45362 29076
rect 42246 29036 45362 29064
rect 45356 29024 45362 29036
rect 45414 29024 45420 29076
rect 45540 29064 45546 29076
rect 45501 29036 45546 29064
rect 45540 29024 45546 29036
rect 45598 29024 45604 29076
rect 46279 29067 46337 29073
rect 46279 29033 46291 29067
rect 46325 29064 46337 29067
rect 52624 29064 52630 29076
rect 46325 29036 52630 29064
rect 46325 29033 46337 29036
rect 46279 29027 46337 29033
rect 52624 29024 52630 29036
rect 52682 29024 52688 29076
rect 52995 29067 53053 29073
rect 52995 29033 53007 29067
rect 53041 29064 53053 29067
rect 55034 29064 55062 29095
rect 55292 29092 55298 29104
rect 55350 29092 55356 29144
rect 57500 29064 57506 29076
rect 53041 29036 55062 29064
rect 55126 29036 57506 29064
rect 53041 29033 53053 29036
rect 52995 29027 53053 29033
rect 17630 28968 19090 28996
rect 17630 28956 17636 28968
rect 19320 28956 19326 29008
rect 19378 28996 19384 29008
rect 24656 28996 24662 29008
rect 19378 28968 24662 28996
rect 19378 28956 19384 28968
rect 24656 28956 24662 28968
rect 24714 28956 24720 29008
rect 24748 28956 24754 29008
rect 24806 28996 24812 29008
rect 30268 28996 30274 29008
rect 24806 28968 24851 28996
rect 30229 28968 30274 28996
rect 24806 28956 24812 28968
rect 30268 28956 30274 28968
rect 30326 28956 30332 29008
rect 30360 28956 30366 29008
rect 30418 28996 30424 29008
rect 34040 28996 34046 29008
rect 30418 28968 34046 28996
rect 30418 28956 30424 28968
rect 34040 28956 34046 28968
rect 34098 28996 34104 29008
rect 35420 28996 35426 29008
rect 34098 28968 35426 28996
rect 34098 28956 34104 28968
rect 35420 28956 35426 28968
rect 35478 28956 35484 29008
rect 36708 28956 36714 29008
rect 36766 28996 36772 29008
rect 38091 28999 38149 29005
rect 38091 28996 38103 28999
rect 36766 28968 38103 28996
rect 36766 28956 36772 28968
rect 38091 28965 38103 28968
rect 38137 28996 38149 28999
rect 38180 28996 38186 29008
rect 38137 28968 38186 28996
rect 38137 28965 38149 28968
rect 38091 28959 38149 28965
rect 38180 28956 38186 28968
rect 38238 28996 38244 29008
rect 38827 28999 38885 29005
rect 38827 28996 38839 28999
rect 38238 28968 38839 28996
rect 38238 28956 38244 28968
rect 38827 28965 38839 28968
rect 38873 28996 38885 28999
rect 39008 28996 39014 29008
rect 38873 28968 39014 28996
rect 38873 28965 38885 28968
rect 38827 28959 38885 28965
rect 39008 28956 39014 28968
rect 39066 28956 39072 29008
rect 42320 28956 42326 29008
rect 42378 28996 42384 29008
rect 43151 28999 43209 29005
rect 43151 28996 43163 28999
rect 42378 28968 43163 28996
rect 42378 28956 42384 28968
rect 43151 28965 43163 28968
rect 43197 28996 43209 28999
rect 43424 28996 43430 29008
rect 43197 28968 43430 28996
rect 43197 28965 43209 28968
rect 43151 28959 43209 28965
rect 43424 28956 43430 28968
rect 43482 28956 43488 29008
rect 48668 28996 48674 29008
rect 48629 28968 48674 28996
rect 48668 28956 48674 28968
rect 48726 28956 48732 29008
rect 49499 28999 49557 29005
rect 49499 28965 49511 28999
rect 49545 28996 49557 28999
rect 49680 28996 49686 29008
rect 49545 28968 49686 28996
rect 49545 28965 49557 28968
rect 49499 28959 49557 28965
rect 49680 28956 49686 28968
rect 49738 28956 49744 29008
rect 49956 28956 49962 29008
rect 50014 28996 50020 29008
rect 51247 28999 51305 29005
rect 51247 28996 51259 28999
rect 50014 28968 51259 28996
rect 50014 28956 50020 28968
rect 51247 28965 51259 28968
rect 51293 28965 51305 28999
rect 51247 28959 51305 28965
rect 53820 28956 53826 29008
rect 53878 28996 53884 29008
rect 55126 28996 55154 29036
rect 57500 29024 57506 29036
rect 57558 29024 57564 29076
rect 58162 29005 58190 29172
rect 58438 29172 58610 29200
rect 58438 29141 58466 29172
rect 58604 29160 58610 29172
rect 58662 29160 58668 29212
rect 59432 29160 59438 29212
rect 59490 29200 59496 29212
rect 59803 29203 59861 29209
rect 59803 29200 59815 29203
rect 59490 29172 59815 29200
rect 59490 29160 59496 29172
rect 59803 29169 59815 29172
rect 59849 29200 59861 29203
rect 61750 29200 61778 29240
rect 59849 29172 61778 29200
rect 59849 29169 59861 29172
rect 59803 29163 59861 29169
rect 61824 29160 61830 29212
rect 61882 29200 61888 29212
rect 62471 29203 62529 29209
rect 62471 29200 62483 29203
rect 61882 29172 62483 29200
rect 61882 29160 61888 29172
rect 62471 29169 62483 29172
rect 62517 29200 62529 29203
rect 62931 29203 62989 29209
rect 62931 29200 62943 29203
rect 62517 29172 62943 29200
rect 62517 29169 62529 29172
rect 62471 29163 62529 29169
rect 62931 29169 62943 29172
rect 62977 29200 62989 29203
rect 64035 29203 64093 29209
rect 64035 29200 64047 29203
rect 62977 29172 64047 29200
rect 62977 29169 62989 29172
rect 62931 29163 62989 29169
rect 64035 29169 64047 29172
rect 64081 29200 64093 29203
rect 64081 29172 64354 29200
rect 64081 29169 64093 29172
rect 64035 29163 64093 29169
rect 58423 29135 58481 29141
rect 58423 29101 58435 29135
rect 58469 29101 58481 29135
rect 58423 29095 58481 29101
rect 58515 29135 58573 29141
rect 58515 29101 58527 29135
rect 58561 29101 58573 29135
rect 58880 29132 58886 29144
rect 58841 29104 58886 29132
rect 58515 29095 58573 29101
rect 58530 29064 58558 29095
rect 58880 29092 58886 29104
rect 58938 29092 58944 29144
rect 58975 29135 59033 29141
rect 58975 29101 58987 29135
rect 59021 29132 59033 29135
rect 59156 29132 59162 29144
rect 59021 29104 59162 29132
rect 59021 29101 59033 29104
rect 58975 29095 59033 29101
rect 59156 29092 59162 29104
rect 59214 29132 59220 29144
rect 60444 29132 60450 29144
rect 59214 29104 60306 29132
rect 60357 29104 60450 29132
rect 59214 29092 59220 29104
rect 59432 29064 59438 29076
rect 58530 29036 59438 29064
rect 59432 29024 59438 29036
rect 59490 29024 59496 29076
rect 60278 29064 60306 29104
rect 60444 29092 60450 29104
rect 60502 29132 60508 29144
rect 62836 29141 62842 29144
rect 62793 29135 62842 29141
rect 62793 29132 62805 29135
rect 60502 29104 60858 29132
rect 62749 29104 62805 29132
rect 60502 29092 60508 29104
rect 60539 29067 60597 29073
rect 60539 29064 60551 29067
rect 60278 29036 60551 29064
rect 60539 29033 60551 29036
rect 60585 29064 60597 29067
rect 60720 29064 60726 29076
rect 60585 29036 60726 29064
rect 60585 29033 60597 29036
rect 60539 29027 60597 29033
rect 60720 29024 60726 29036
rect 60778 29024 60784 29076
rect 53878 28968 55154 28996
rect 58147 28999 58205 29005
rect 53878 28956 53884 28968
rect 58147 28965 58159 28999
rect 58193 28996 58205 28999
rect 58880 28996 58886 29008
rect 58193 28968 58886 28996
rect 58193 28965 58205 28968
rect 58147 28959 58205 28965
rect 58880 28956 58886 28968
rect 58938 28956 58944 29008
rect 60830 29005 60858 29104
rect 62793 29101 62805 29104
rect 62839 29101 62842 29135
rect 62793 29095 62842 29101
rect 62836 29092 62842 29095
rect 62894 29132 62900 29144
rect 64326 29141 64354 29172
rect 67436 29160 67442 29212
rect 67494 29200 67500 29212
rect 67991 29203 68049 29209
rect 67991 29200 68003 29203
rect 67494 29172 68003 29200
rect 67494 29160 67500 29172
rect 67991 29169 68003 29172
rect 68037 29169 68049 29203
rect 67991 29163 68049 29169
rect 68650 29144 68678 29240
rect 69092 29200 69098 29212
rect 69053 29172 69098 29200
rect 69092 29160 69098 29172
rect 69150 29160 69156 29212
rect 69202 29200 69230 29240
rect 69460 29228 69466 29280
rect 69518 29268 69524 29280
rect 76087 29271 76145 29277
rect 69518 29240 71530 29268
rect 69518 29228 69524 29240
rect 70107 29203 70165 29209
rect 70107 29200 70119 29203
rect 69202 29172 70119 29200
rect 70107 29169 70119 29172
rect 70153 29169 70165 29203
rect 70107 29163 70165 29169
rect 64127 29135 64185 29141
rect 64127 29132 64139 29135
rect 62894 29104 64139 29132
rect 62894 29092 62900 29104
rect 64127 29101 64139 29104
rect 64173 29101 64185 29135
rect 64127 29095 64185 29101
rect 64311 29135 64369 29141
rect 64311 29101 64323 29135
rect 64357 29132 64369 29135
rect 65320 29132 65326 29144
rect 64357 29104 65326 29132
rect 64357 29101 64369 29104
rect 64311 29095 64369 29101
rect 65320 29092 65326 29104
rect 65378 29092 65384 29144
rect 67896 29092 67902 29144
rect 67954 29132 67960 29144
rect 68172 29132 68178 29144
rect 67954 29104 68178 29132
rect 67954 29092 67960 29104
rect 68172 29092 68178 29104
rect 68230 29092 68236 29144
rect 68632 29132 68638 29144
rect 68593 29104 68638 29132
rect 68632 29092 68638 29104
rect 68690 29092 68696 29144
rect 68727 29135 68785 29141
rect 68727 29101 68739 29135
rect 68773 29101 68785 29135
rect 69000 29132 69006 29144
rect 68961 29104 69006 29132
rect 68727 29095 68785 29101
rect 62100 29024 62106 29076
rect 62158 29064 62164 29076
rect 62563 29067 62621 29073
rect 62563 29064 62575 29067
rect 62158 29036 62575 29064
rect 62158 29024 62164 29036
rect 62563 29033 62575 29036
rect 62609 29033 62621 29067
rect 62563 29027 62621 29033
rect 64492 29024 64498 29076
rect 64550 29064 64556 29076
rect 68742 29064 68770 29095
rect 69000 29092 69006 29104
rect 69058 29092 69064 29144
rect 64550 29036 68770 29064
rect 69110 29064 69138 29160
rect 69552 29092 69558 29144
rect 69610 29132 69616 29144
rect 70015 29135 70073 29141
rect 70015 29132 70027 29135
rect 69610 29104 70027 29132
rect 69610 29092 69616 29104
rect 70015 29101 70027 29104
rect 70061 29101 70073 29135
rect 70015 29095 70073 29101
rect 71027 29135 71085 29141
rect 71027 29101 71039 29135
rect 71073 29101 71085 29135
rect 71027 29095 71085 29101
rect 69110 29036 69414 29064
rect 64550 29024 64556 29036
rect 60815 28999 60873 29005
rect 60815 28965 60827 28999
rect 60861 28996 60873 28999
rect 62652 28996 62658 29008
rect 60861 28968 62658 28996
rect 60861 28965 60873 28968
rect 60815 28959 60873 28965
rect 62652 28956 62658 28968
rect 62710 28956 62716 29008
rect 63204 28996 63210 29008
rect 63165 28968 63210 28996
rect 63204 28956 63210 28968
rect 63262 28956 63268 29008
rect 64400 28996 64406 29008
rect 64361 28968 64406 28996
rect 64400 28956 64406 28968
rect 64458 28956 64464 29008
rect 68742 28996 68770 29036
rect 69184 28996 69190 29008
rect 68742 28968 69190 28996
rect 69184 28956 69190 28968
rect 69242 28996 69248 29008
rect 69279 28999 69337 29005
rect 69279 28996 69291 28999
rect 69242 28968 69291 28996
rect 69242 28956 69248 28968
rect 69279 28965 69291 28968
rect 69325 28965 69337 28999
rect 69386 28996 69414 29036
rect 69460 29024 69466 29076
rect 69518 29064 69524 29076
rect 70843 29067 70901 29073
rect 70843 29064 70855 29067
rect 69518 29036 70855 29064
rect 69518 29024 69524 29036
rect 70843 29033 70855 29036
rect 70889 29064 70901 29067
rect 71042 29064 71070 29095
rect 71116 29092 71122 29144
rect 71174 29132 71180 29144
rect 71502 29132 71530 29240
rect 71594 29240 76038 29268
rect 71594 29209 71622 29240
rect 71579 29203 71637 29209
rect 71579 29169 71591 29203
rect 71625 29169 71637 29203
rect 71579 29163 71637 29169
rect 74980 29160 74986 29212
rect 75038 29200 75044 29212
rect 75075 29203 75133 29209
rect 75075 29200 75087 29203
rect 75038 29172 75087 29200
rect 75038 29160 75044 29172
rect 75075 29169 75087 29172
rect 75121 29169 75133 29203
rect 76010 29200 76038 29240
rect 76087 29237 76099 29271
rect 76133 29268 76145 29271
rect 76912 29268 76918 29280
rect 76133 29240 76918 29268
rect 76133 29237 76145 29240
rect 76087 29231 76145 29237
rect 76912 29228 76918 29240
rect 76970 29228 76976 29280
rect 84916 29268 84922 29280
rect 77114 29240 84318 29268
rect 84877 29240 84922 29268
rect 77114 29200 77142 29240
rect 76010 29172 77142 29200
rect 75075 29163 75133 29169
rect 78936 29160 78942 29212
rect 78994 29200 79000 29212
rect 80871 29203 80929 29209
rect 80871 29200 80883 29203
rect 78994 29172 80883 29200
rect 78994 29160 79000 29172
rect 80871 29169 80883 29172
rect 80917 29200 80929 29203
rect 84290 29200 84318 29240
rect 84916 29228 84922 29240
rect 84974 29228 84980 29280
rect 85836 29228 85842 29280
rect 85894 29268 85900 29280
rect 90163 29271 90221 29277
rect 90163 29268 90175 29271
rect 85894 29240 90175 29268
rect 85894 29228 85900 29240
rect 90163 29237 90175 29240
rect 90209 29268 90221 29271
rect 90531 29271 90589 29277
rect 90531 29268 90543 29271
rect 90209 29240 90543 29268
rect 90209 29237 90221 29240
rect 90163 29231 90221 29237
rect 90531 29237 90543 29240
rect 90577 29237 90589 29271
rect 90531 29231 90589 29237
rect 91080 29200 91086 29212
rect 80917 29172 81282 29200
rect 84290 29172 91086 29200
rect 80917 29169 80929 29172
rect 80871 29163 80929 29169
rect 81254 29144 81282 29172
rect 91080 29160 91086 29172
rect 91138 29160 91144 29212
rect 73603 29135 73661 29141
rect 73603 29132 73615 29135
rect 71174 29104 71219 29132
rect 71502 29104 73615 29132
rect 71174 29092 71180 29104
rect 73603 29101 73615 29104
rect 73649 29132 73661 29135
rect 73879 29135 73937 29141
rect 73879 29132 73891 29135
rect 73649 29104 73891 29132
rect 73649 29101 73661 29104
rect 73603 29095 73661 29101
rect 73879 29101 73891 29104
rect 73925 29132 73937 29135
rect 74244 29132 74250 29144
rect 73925 29104 74250 29132
rect 73925 29101 73937 29104
rect 73879 29095 73937 29101
rect 74244 29092 74250 29104
rect 74302 29092 74308 29144
rect 74799 29135 74857 29141
rect 74799 29132 74811 29135
rect 74446 29104 74811 29132
rect 74446 29073 74474 29104
rect 74799 29101 74811 29104
rect 74845 29132 74857 29135
rect 75811 29135 75869 29141
rect 75811 29132 75823 29135
rect 74845 29104 75823 29132
rect 74845 29101 74857 29104
rect 74799 29095 74857 29101
rect 75811 29101 75823 29104
rect 75857 29132 75869 29135
rect 75995 29135 76053 29141
rect 75995 29132 76007 29135
rect 75857 29104 76007 29132
rect 75857 29101 75869 29104
rect 75811 29095 75869 29101
rect 75995 29101 76007 29104
rect 76041 29101 76053 29135
rect 75995 29095 76053 29101
rect 76271 29135 76329 29141
rect 76271 29101 76283 29135
rect 76317 29101 76329 29135
rect 77740 29132 77746 29144
rect 77701 29104 77746 29132
rect 76271 29095 76329 29101
rect 74431 29067 74489 29073
rect 74431 29064 74443 29067
rect 70889 29036 71070 29064
rect 71410 29036 74443 29064
rect 70889 29033 70901 29036
rect 70843 29027 70901 29033
rect 71410 28996 71438 29036
rect 74431 29033 74443 29036
rect 74477 29033 74489 29067
rect 74612 29064 74618 29076
rect 74573 29036 74618 29064
rect 74431 29027 74489 29033
rect 74612 29024 74618 29036
rect 74670 29064 74676 29076
rect 76286 29064 76314 29095
rect 77740 29092 77746 29104
rect 77798 29092 77804 29144
rect 79856 29132 79862 29144
rect 79817 29104 79862 29132
rect 79856 29092 79862 29104
rect 79914 29092 79920 29144
rect 81236 29132 81242 29144
rect 81149 29104 81242 29132
rect 81236 29092 81242 29104
rect 81294 29092 81300 29144
rect 84824 29092 84830 29144
rect 84882 29132 84888 29144
rect 85011 29135 85069 29141
rect 85011 29132 85023 29135
rect 84882 29104 85023 29132
rect 84882 29092 84888 29104
rect 85011 29101 85023 29104
rect 85057 29101 85069 29135
rect 85011 29095 85069 29101
rect 85379 29135 85437 29141
rect 85379 29101 85391 29135
rect 85425 29101 85437 29135
rect 85379 29095 85437 29101
rect 86575 29135 86633 29141
rect 86575 29101 86587 29135
rect 86621 29132 86633 29135
rect 86756 29132 86762 29144
rect 86621 29104 86762 29132
rect 86621 29101 86633 29104
rect 86575 29095 86633 29101
rect 74670 29036 76314 29064
rect 76731 29067 76789 29073
rect 74670 29024 74676 29036
rect 76731 29033 76743 29067
rect 76777 29064 76789 29067
rect 79675 29067 79733 29073
rect 79675 29064 79687 29067
rect 76777 29036 79687 29064
rect 76777 29033 76789 29036
rect 76731 29027 76789 29033
rect 79675 29033 79687 29036
rect 79721 29064 79733 29067
rect 80132 29064 80138 29076
rect 79721 29036 80138 29064
rect 79721 29033 79733 29036
rect 79675 29027 79733 29033
rect 80132 29024 80138 29036
rect 80190 29024 80196 29076
rect 80227 29067 80285 29073
rect 80227 29033 80239 29067
rect 80273 29064 80285 29067
rect 80316 29064 80322 29076
rect 80273 29036 80322 29064
rect 80273 29033 80285 29036
rect 80227 29027 80285 29033
rect 80316 29024 80322 29036
rect 80374 29024 80380 29076
rect 81055 29067 81113 29073
rect 81055 29033 81067 29067
rect 81101 29064 81113 29067
rect 81420 29064 81426 29076
rect 81101 29036 81426 29064
rect 81101 29033 81113 29036
rect 81055 29027 81113 29033
rect 81420 29024 81426 29036
rect 81478 29024 81484 29076
rect 84088 29024 84094 29076
rect 84146 29064 84152 29076
rect 84548 29064 84554 29076
rect 84146 29036 84554 29064
rect 84146 29024 84152 29036
rect 84548 29024 84554 29036
rect 84606 29064 84612 29076
rect 85394 29064 85422 29095
rect 86756 29092 86762 29104
rect 86814 29092 86820 29144
rect 90804 29132 90810 29144
rect 90765 29104 90810 29132
rect 90804 29092 90810 29104
rect 90862 29092 90868 29144
rect 91448 29092 91454 29144
rect 91506 29132 91512 29144
rect 91908 29132 91914 29144
rect 91506 29104 91914 29132
rect 91506 29092 91512 29104
rect 91908 29092 91914 29104
rect 91966 29132 91972 29144
rect 92095 29135 92153 29141
rect 92095 29132 92107 29135
rect 91966 29104 92107 29132
rect 91966 29092 91972 29104
rect 92095 29101 92107 29104
rect 92141 29101 92153 29135
rect 92095 29095 92153 29101
rect 84606 29036 85422 29064
rect 86391 29067 86449 29073
rect 84606 29024 84612 29036
rect 86391 29033 86403 29067
rect 86437 29064 86449 29067
rect 87768 29064 87774 29076
rect 86437 29036 87774 29064
rect 86437 29033 86449 29036
rect 86391 29027 86449 29033
rect 87768 29024 87774 29036
rect 87826 29024 87832 29076
rect 90712 29064 90718 29076
rect 90673 29036 90718 29064
rect 90712 29024 90718 29036
rect 90770 29024 90776 29076
rect 69386 28968 71438 28996
rect 69279 28959 69337 28965
rect 73692 28956 73698 29008
rect 73750 28996 73756 29008
rect 77556 28996 77562 29008
rect 73750 28968 73795 28996
rect 77469 28968 77562 28996
rect 73750 28956 73756 28968
rect 77556 28956 77562 28968
rect 77614 28996 77620 29008
rect 79488 28996 79494 29008
rect 77614 28968 79494 28996
rect 77614 28956 77620 28968
rect 79488 28956 79494 28968
rect 79546 28956 79552 29008
rect 81328 28996 81334 29008
rect 81289 28968 81334 28996
rect 81328 28956 81334 28968
rect 81386 28956 81392 29008
rect 90620 28956 90626 29008
rect 90678 28996 90684 29008
rect 92187 28999 92245 29005
rect 92187 28996 92199 28999
rect 90678 28968 92199 28996
rect 90678 28956 90684 28968
rect 92187 28965 92199 28968
rect 92233 28965 92245 28999
rect 92187 28959 92245 28965
rect 538 28906 93642 28928
rect 538 28854 6344 28906
rect 6396 28854 6408 28906
rect 6460 28854 6472 28906
rect 6524 28854 6536 28906
rect 6588 28854 11672 28906
rect 11724 28854 11736 28906
rect 11788 28854 11800 28906
rect 11852 28854 11864 28906
rect 11916 28854 17000 28906
rect 17052 28854 17064 28906
rect 17116 28854 17128 28906
rect 17180 28854 17192 28906
rect 17244 28854 22328 28906
rect 22380 28854 22392 28906
rect 22444 28854 22456 28906
rect 22508 28854 22520 28906
rect 22572 28854 27656 28906
rect 27708 28854 27720 28906
rect 27772 28854 27784 28906
rect 27836 28854 27848 28906
rect 27900 28854 32984 28906
rect 33036 28854 33048 28906
rect 33100 28854 33112 28906
rect 33164 28854 33176 28906
rect 33228 28854 38312 28906
rect 38364 28854 38376 28906
rect 38428 28854 38440 28906
rect 38492 28854 38504 28906
rect 38556 28854 43640 28906
rect 43692 28854 43704 28906
rect 43756 28854 43768 28906
rect 43820 28854 43832 28906
rect 43884 28854 48968 28906
rect 49020 28854 49032 28906
rect 49084 28854 49096 28906
rect 49148 28854 49160 28906
rect 49212 28854 54296 28906
rect 54348 28854 54360 28906
rect 54412 28854 54424 28906
rect 54476 28854 54488 28906
rect 54540 28854 59624 28906
rect 59676 28854 59688 28906
rect 59740 28854 59752 28906
rect 59804 28854 59816 28906
rect 59868 28854 64952 28906
rect 65004 28854 65016 28906
rect 65068 28854 65080 28906
rect 65132 28854 65144 28906
rect 65196 28854 70280 28906
rect 70332 28854 70344 28906
rect 70396 28854 70408 28906
rect 70460 28854 70472 28906
rect 70524 28854 75608 28906
rect 75660 28854 75672 28906
rect 75724 28854 75736 28906
rect 75788 28854 75800 28906
rect 75852 28854 80936 28906
rect 80988 28854 81000 28906
rect 81052 28854 81064 28906
rect 81116 28854 81128 28906
rect 81180 28854 86264 28906
rect 86316 28854 86328 28906
rect 86380 28854 86392 28906
rect 86444 28854 86456 28906
rect 86508 28854 91592 28906
rect 91644 28854 91656 28906
rect 91708 28854 91720 28906
rect 91772 28854 91784 28906
rect 91836 28854 93642 28906
rect 538 28832 93642 28854
rect 6716 28792 6722 28804
rect 6677 28764 6722 28792
rect 6716 28752 6722 28764
rect 6774 28752 6780 28804
rect 9292 28792 9298 28804
rect 9126 28764 9298 28792
rect 6164 28616 6170 28668
rect 6222 28656 6228 28668
rect 6535 28659 6593 28665
rect 6535 28656 6547 28659
rect 6222 28628 6547 28656
rect 6222 28616 6228 28628
rect 6535 28625 6547 28628
rect 6581 28625 6593 28659
rect 6535 28619 6593 28625
rect 6734 28588 6762 28752
rect 9126 28733 9154 28764
rect 9292 28752 9298 28764
rect 9350 28752 9356 28804
rect 13159 28795 13217 28801
rect 13159 28761 13171 28795
rect 13205 28792 13217 28795
rect 13524 28792 13530 28804
rect 13205 28764 13530 28792
rect 13205 28761 13217 28764
rect 13159 28755 13217 28761
rect 9111 28727 9169 28733
rect 9111 28693 9123 28727
rect 9157 28693 9169 28727
rect 9476 28724 9482 28736
rect 9437 28696 9482 28724
rect 9111 28687 9169 28693
rect 9476 28684 9482 28696
rect 9534 28684 9540 28736
rect 10948 28684 10954 28736
rect 11006 28724 11012 28736
rect 12972 28724 12978 28736
rect 11006 28696 11730 28724
rect 12933 28696 12978 28724
rect 11006 28684 11012 28696
rect 8096 28616 8102 28668
rect 8154 28656 8160 28668
rect 9295 28659 9353 28665
rect 9295 28656 9307 28659
rect 8154 28628 9307 28656
rect 8154 28616 8160 28628
rect 9295 28625 9307 28628
rect 9341 28625 9353 28659
rect 9295 28619 9353 28625
rect 9384 28616 9390 28668
rect 9442 28656 9448 28668
rect 11500 28656 11506 28668
rect 9442 28628 9535 28656
rect 11461 28628 11506 28656
rect 9442 28616 9448 28628
rect 11500 28616 11506 28628
rect 11558 28616 11564 28668
rect 11702 28665 11730 28696
rect 12972 28684 12978 28696
rect 13030 28684 13036 28736
rect 11687 28659 11745 28665
rect 11687 28625 11699 28659
rect 11733 28625 11745 28659
rect 12052 28656 12058 28668
rect 12013 28628 12058 28656
rect 11687 28619 11745 28625
rect 12052 28616 12058 28628
rect 12110 28616 12116 28668
rect 12239 28659 12297 28665
rect 12239 28625 12251 28659
rect 12285 28625 12297 28659
rect 12239 28619 12297 28625
rect 12515 28659 12573 28665
rect 12515 28625 12527 28659
rect 12561 28656 12573 28659
rect 13174 28656 13202 28755
rect 13524 28752 13530 28764
rect 13582 28792 13588 28804
rect 14907 28795 14965 28801
rect 14907 28792 14919 28795
rect 13582 28764 14919 28792
rect 13582 28752 13588 28764
rect 14907 28761 14919 28764
rect 14953 28792 14965 28795
rect 17296 28792 17302 28804
rect 14953 28764 17302 28792
rect 14953 28761 14965 28764
rect 14907 28755 14965 28761
rect 17296 28752 17302 28764
rect 17354 28752 17360 28804
rect 17848 28752 17854 28804
rect 17906 28792 17912 28804
rect 24475 28795 24533 28801
rect 24475 28792 24487 28795
rect 17906 28764 24487 28792
rect 17906 28752 17912 28764
rect 24475 28761 24487 28764
rect 24521 28761 24533 28795
rect 24475 28755 24533 28761
rect 24656 28752 24662 28804
rect 24714 28792 24720 28804
rect 24714 28764 28474 28792
rect 24714 28752 24720 28764
rect 16652 28684 16658 28736
rect 16710 28724 16716 28736
rect 17207 28727 17265 28733
rect 17207 28724 17219 28727
rect 16710 28696 17219 28724
rect 16710 28684 16716 28696
rect 17207 28693 17219 28696
rect 17253 28693 17265 28727
rect 17207 28687 17265 28693
rect 14720 28656 14726 28668
rect 12561 28628 13202 28656
rect 14681 28628 14726 28656
rect 12561 28625 12573 28628
rect 12515 28619 12573 28625
rect 9402 28588 9430 28616
rect 6734 28560 9430 28588
rect 9847 28591 9905 28597
rect 9847 28557 9859 28591
rect 9893 28588 9905 28591
rect 10948 28588 10954 28600
rect 9893 28560 10954 28588
rect 9893 28557 9905 28560
rect 9847 28551 9905 28557
rect 10948 28548 10954 28560
rect 11006 28548 11012 28600
rect 5980 28480 5986 28532
rect 6038 28520 6044 28532
rect 11316 28520 11322 28532
rect 6038 28492 11322 28520
rect 6038 28480 6044 28492
rect 11316 28480 11322 28492
rect 11374 28480 11380 28532
rect 11411 28523 11469 28529
rect 11411 28489 11423 28523
rect 11457 28520 11469 28523
rect 11500 28520 11506 28532
rect 11457 28492 11506 28520
rect 11457 28489 11469 28492
rect 11411 28483 11469 28489
rect 11500 28480 11506 28492
rect 11558 28520 11564 28532
rect 12254 28520 12282 28619
rect 14720 28616 14726 28628
rect 14778 28656 14784 28668
rect 15091 28659 15149 28665
rect 15091 28656 15103 28659
rect 14778 28628 15103 28656
rect 14778 28616 14784 28628
rect 15091 28625 15103 28628
rect 15137 28656 15149 28659
rect 15827 28659 15885 28665
rect 15827 28656 15839 28659
rect 15137 28628 15839 28656
rect 15137 28625 15149 28628
rect 15091 28619 15149 28625
rect 15827 28625 15839 28628
rect 15873 28656 15885 28659
rect 15916 28656 15922 28668
rect 15873 28628 15922 28656
rect 15873 28625 15885 28628
rect 15827 28619 15885 28625
rect 15916 28616 15922 28628
rect 15974 28656 15980 28668
rect 16103 28659 16161 28665
rect 16103 28656 16115 28659
rect 15974 28628 16115 28656
rect 15974 28616 15980 28628
rect 16103 28625 16115 28628
rect 16149 28625 16161 28659
rect 16103 28619 16161 28625
rect 15735 28591 15793 28597
rect 15735 28557 15747 28591
rect 15781 28588 15793 28591
rect 16011 28591 16069 28597
rect 16011 28588 16023 28591
rect 15781 28560 16023 28588
rect 15781 28557 15793 28560
rect 15735 28551 15793 28557
rect 16011 28557 16023 28560
rect 16057 28588 16069 28591
rect 16744 28588 16750 28600
rect 16057 28560 16750 28588
rect 16057 28557 16069 28560
rect 16011 28551 16069 28557
rect 16744 28548 16750 28560
rect 16802 28548 16808 28600
rect 17222 28588 17250 28687
rect 18584 28684 18590 28736
rect 18642 28724 18648 28736
rect 25484 28724 25490 28736
rect 18642 28696 25490 28724
rect 18642 28684 18648 28696
rect 25484 28684 25490 28696
rect 25542 28684 25548 28736
rect 25760 28724 25766 28736
rect 25594 28696 25766 28724
rect 17296 28616 17302 28668
rect 17354 28656 17360 28668
rect 17575 28659 17633 28665
rect 17575 28656 17587 28659
rect 17354 28628 17587 28656
rect 17354 28616 17360 28628
rect 17575 28625 17587 28628
rect 17621 28656 17633 28659
rect 18127 28659 18185 28665
rect 18127 28656 18139 28659
rect 17621 28628 18139 28656
rect 17621 28625 17633 28628
rect 17575 28619 17633 28625
rect 17391 28591 17449 28597
rect 17391 28588 17403 28591
rect 17222 28560 17403 28588
rect 17391 28557 17403 28560
rect 17437 28588 17449 28591
rect 17664 28588 17670 28600
rect 17437 28560 17670 28588
rect 17437 28557 17449 28560
rect 17391 28551 17449 28557
rect 17664 28548 17670 28560
rect 17722 28548 17728 28600
rect 11558 28492 12282 28520
rect 11558 28480 11564 28492
rect 15088 28412 15094 28464
rect 15146 28452 15152 28464
rect 16100 28452 16106 28464
rect 15146 28424 16106 28452
rect 15146 28412 15152 28424
rect 16100 28412 16106 28424
rect 16158 28412 16164 28464
rect 16284 28452 16290 28464
rect 16245 28424 16290 28452
rect 16284 28412 16290 28424
rect 16342 28412 16348 28464
rect 17774 28452 17802 28628
rect 18127 28625 18139 28628
rect 18173 28625 18185 28659
rect 18127 28619 18185 28625
rect 18311 28659 18369 28665
rect 18311 28625 18323 28659
rect 18357 28656 18369 28659
rect 18952 28656 18958 28668
rect 18357 28628 18958 28656
rect 18357 28625 18369 28628
rect 18311 28619 18369 28625
rect 18952 28616 18958 28628
rect 19010 28616 19016 28668
rect 22724 28656 22730 28668
rect 22685 28628 22730 28656
rect 22724 28616 22730 28628
rect 22782 28656 22788 28668
rect 23460 28656 23466 28668
rect 22782 28628 23322 28656
rect 23421 28628 23466 28656
rect 22782 28616 22788 28628
rect 23092 28588 23098 28600
rect 23053 28560 23098 28588
rect 23092 28548 23098 28560
rect 23150 28548 23156 28600
rect 23294 28588 23322 28628
rect 23460 28616 23466 28628
rect 23518 28616 23524 28668
rect 23647 28659 23705 28665
rect 23647 28625 23659 28659
rect 23693 28625 23705 28659
rect 23828 28656 23834 28668
rect 23789 28628 23834 28656
rect 23647 28619 23705 28625
rect 23662 28588 23690 28619
rect 23828 28616 23834 28628
rect 23886 28616 23892 28668
rect 24107 28659 24165 28665
rect 24107 28656 24119 28659
rect 24030 28628 24119 28656
rect 23736 28588 23742 28600
rect 23294 28560 23742 28588
rect 23736 28548 23742 28560
rect 23794 28548 23800 28600
rect 18216 28480 18222 28532
rect 18274 28520 18280 28532
rect 18495 28523 18553 28529
rect 18495 28520 18507 28523
rect 18274 28492 18507 28520
rect 18274 28480 18280 28492
rect 18495 28489 18507 28492
rect 18541 28489 18553 28523
rect 18495 28483 18553 28489
rect 20976 28480 20982 28532
rect 21034 28520 21040 28532
rect 23003 28523 23061 28529
rect 23003 28520 23015 28523
rect 21034 28492 23015 28520
rect 21034 28480 21040 28492
rect 23003 28489 23015 28492
rect 23049 28520 23061 28523
rect 24030 28520 24058 28628
rect 24107 28625 24119 28628
rect 24153 28625 24165 28659
rect 24107 28619 24165 28625
rect 24751 28659 24809 28665
rect 24751 28625 24763 28659
rect 24797 28656 24809 28659
rect 24840 28656 24846 28668
rect 24797 28628 24846 28656
rect 24797 28625 24809 28628
rect 24751 28619 24809 28625
rect 24840 28616 24846 28628
rect 24898 28616 24904 28668
rect 25594 28665 25622 28696
rect 25760 28684 25766 28696
rect 25818 28684 25824 28736
rect 26496 28684 26502 28736
rect 26554 28724 26560 28736
rect 27416 28724 27422 28736
rect 26554 28696 27422 28724
rect 26554 28684 26560 28696
rect 25579 28659 25637 28665
rect 25579 28625 25591 28659
rect 25625 28625 25637 28659
rect 25579 28619 25637 28625
rect 26959 28659 27017 28665
rect 26959 28625 26971 28659
rect 27005 28656 27017 28659
rect 27140 28656 27146 28668
rect 27005 28628 27146 28656
rect 27005 28625 27017 28628
rect 26959 28619 27017 28625
rect 27140 28616 27146 28628
rect 27198 28616 27204 28668
rect 27250 28665 27278 28696
rect 27416 28684 27422 28696
rect 27474 28684 27480 28736
rect 28336 28724 28342 28736
rect 27526 28696 28342 28724
rect 27526 28665 27554 28696
rect 28336 28684 28342 28696
rect 28394 28684 28400 28736
rect 28446 28724 28474 28764
rect 28520 28752 28526 28804
rect 28578 28792 28584 28804
rect 30360 28792 30366 28804
rect 28578 28764 30366 28792
rect 28578 28752 28584 28764
rect 30360 28752 30366 28764
rect 30418 28752 30424 28804
rect 30452 28752 30458 28804
rect 30510 28792 30516 28804
rect 31651 28795 31709 28801
rect 31651 28792 31663 28795
rect 30510 28764 31663 28792
rect 30510 28752 30516 28764
rect 31651 28761 31663 28764
rect 31697 28761 31709 28795
rect 31651 28755 31709 28761
rect 34040 28752 34046 28804
rect 34098 28792 34104 28804
rect 34135 28795 34193 28801
rect 34135 28792 34147 28795
rect 34098 28764 34147 28792
rect 34098 28752 34104 28764
rect 34135 28761 34147 28764
rect 34181 28792 34193 28795
rect 34500 28792 34506 28804
rect 34181 28764 34506 28792
rect 34181 28761 34193 28764
rect 34135 28755 34193 28761
rect 34500 28752 34506 28764
rect 34558 28752 34564 28804
rect 37720 28792 37726 28804
rect 34610 28764 37726 28792
rect 34610 28724 34638 28764
rect 37720 28752 37726 28764
rect 37778 28752 37784 28804
rect 42872 28792 42878 28804
rect 42833 28764 42878 28792
rect 42872 28752 42878 28764
rect 42930 28792 42936 28804
rect 42930 28764 43930 28792
rect 42930 28752 42936 28764
rect 36156 28724 36162 28736
rect 28446 28696 34638 28724
rect 36117 28696 36162 28724
rect 36156 28684 36162 28696
rect 36214 28684 36220 28736
rect 36248 28684 36254 28736
rect 36306 28724 36312 28736
rect 39560 28724 39566 28736
rect 36306 28696 39566 28724
rect 36306 28684 36312 28696
rect 39560 28684 39566 28696
rect 39618 28684 39624 28736
rect 43056 28684 43062 28736
rect 43114 28724 43120 28736
rect 43792 28724 43798 28736
rect 43114 28696 43798 28724
rect 43114 28684 43120 28696
rect 27235 28659 27293 28665
rect 27235 28625 27247 28659
rect 27281 28625 27293 28659
rect 27235 28619 27293 28625
rect 27511 28659 27569 28665
rect 27511 28625 27523 28659
rect 27557 28625 27569 28659
rect 27511 28619 27569 28625
rect 27603 28659 27661 28665
rect 27603 28625 27615 28659
rect 27649 28656 27661 28659
rect 27649 28628 27830 28656
rect 27649 28625 27661 28628
rect 27603 28619 27661 28625
rect 26683 28591 26741 28597
rect 24214 28560 26634 28588
rect 24214 28520 24242 28560
rect 26315 28523 26373 28529
rect 26315 28520 26327 28523
rect 23049 28492 24242 28520
rect 24490 28492 26327 28520
rect 23049 28489 23061 28492
rect 23003 28483 23061 28489
rect 19047 28455 19105 28461
rect 19047 28452 19059 28455
rect 17774 28424 19059 28452
rect 19047 28421 19059 28424
rect 19093 28452 19105 28455
rect 19231 28455 19289 28461
rect 19231 28452 19243 28455
rect 19093 28424 19243 28452
rect 19093 28421 19105 28424
rect 19047 28415 19105 28421
rect 19231 28421 19243 28424
rect 19277 28452 19289 28455
rect 22632 28452 22638 28464
rect 19277 28424 22638 28452
rect 19277 28421 19289 28424
rect 19231 28415 19289 28421
rect 22632 28412 22638 28424
rect 22690 28412 22696 28464
rect 23736 28412 23742 28464
rect 23794 28452 23800 28464
rect 24490 28452 24518 28492
rect 26315 28489 26327 28492
rect 26361 28520 26373 28523
rect 26496 28520 26502 28532
rect 26361 28492 26502 28520
rect 26361 28489 26373 28492
rect 26315 28483 26373 28489
rect 26496 28480 26502 28492
rect 26554 28480 26560 28532
rect 26606 28529 26634 28560
rect 26683 28557 26695 28591
rect 26729 28588 26741 28591
rect 27692 28588 27698 28600
rect 26729 28560 27698 28588
rect 26729 28557 26741 28560
rect 26683 28551 26741 28557
rect 27692 28548 27698 28560
rect 27750 28548 27756 28600
rect 26591 28523 26649 28529
rect 26591 28489 26603 28523
rect 26637 28520 26649 28523
rect 27802 28520 27830 28628
rect 28704 28616 28710 28668
rect 28762 28656 28768 28668
rect 29167 28659 29225 28665
rect 29167 28656 29179 28659
rect 28762 28628 29179 28656
rect 28762 28616 28768 28628
rect 29167 28625 29179 28628
rect 29213 28625 29225 28659
rect 29808 28656 29814 28668
rect 29769 28628 29814 28656
rect 29167 28619 29225 28625
rect 29808 28616 29814 28628
rect 29866 28616 29872 28668
rect 29903 28659 29961 28665
rect 29903 28625 29915 28659
rect 29949 28656 29961 28659
rect 30084 28656 30090 28668
rect 29949 28628 30090 28656
rect 29949 28625 29961 28628
rect 29903 28619 29961 28625
rect 30084 28616 30090 28628
rect 30142 28616 30148 28668
rect 30179 28659 30237 28665
rect 30179 28625 30191 28659
rect 30225 28656 30237 28659
rect 31556 28656 31562 28668
rect 30225 28628 30590 28656
rect 31517 28628 31562 28656
rect 30225 28625 30237 28628
rect 30179 28619 30237 28625
rect 27876 28548 27882 28600
rect 27934 28588 27940 28600
rect 29532 28588 29538 28600
rect 27934 28560 29538 28588
rect 27934 28548 27940 28560
rect 29532 28548 29538 28560
rect 29590 28548 29596 28600
rect 29716 28548 29722 28600
rect 29774 28588 29780 28600
rect 30268 28588 30274 28600
rect 29774 28560 30274 28588
rect 29774 28548 29780 28560
rect 30268 28548 30274 28560
rect 30326 28548 30332 28600
rect 30562 28597 30590 28628
rect 31556 28616 31562 28628
rect 31614 28616 31620 28668
rect 32016 28616 32022 28668
rect 32074 28656 32080 28668
rect 38735 28659 38793 28665
rect 32074 28628 38686 28656
rect 32074 28616 32080 28628
rect 30547 28591 30605 28597
rect 30547 28557 30559 28591
rect 30593 28588 30605 28591
rect 33948 28588 33954 28600
rect 30593 28560 33954 28588
rect 30593 28557 30605 28560
rect 30547 28551 30605 28557
rect 33948 28548 33954 28560
rect 34006 28548 34012 28600
rect 34408 28588 34414 28600
rect 34369 28560 34414 28588
rect 34408 28548 34414 28560
rect 34466 28588 34472 28600
rect 34503 28591 34561 28597
rect 34503 28588 34515 28591
rect 34466 28560 34515 28588
rect 34466 28548 34472 28560
rect 34503 28557 34515 28560
rect 34549 28557 34561 28591
rect 34503 28551 34561 28557
rect 34779 28591 34837 28597
rect 34779 28557 34791 28591
rect 34825 28588 34837 28591
rect 35420 28588 35426 28600
rect 34825 28560 35426 28588
rect 34825 28557 34837 28560
rect 34779 28551 34837 28557
rect 35420 28548 35426 28560
rect 35478 28548 35484 28600
rect 35512 28548 35518 28600
rect 35570 28588 35576 28600
rect 37444 28588 37450 28600
rect 35570 28560 37450 28588
rect 35570 28548 35576 28560
rect 37444 28548 37450 28560
rect 37502 28548 37508 28600
rect 38548 28588 38554 28600
rect 38509 28560 38554 28588
rect 38548 28548 38554 28560
rect 38606 28548 38612 28600
rect 38658 28588 38686 28628
rect 38735 28625 38747 28659
rect 38781 28656 38793 28659
rect 38824 28656 38830 28668
rect 38781 28628 38830 28656
rect 38781 28625 38793 28628
rect 38735 28619 38793 28625
rect 38824 28616 38830 28628
rect 38882 28616 38888 28668
rect 39192 28656 39198 28668
rect 39153 28628 39198 28656
rect 39192 28616 39198 28628
rect 39250 28616 39256 28668
rect 39287 28659 39345 28665
rect 39287 28625 39299 28659
rect 39333 28656 39345 28659
rect 39468 28656 39474 28668
rect 39333 28628 39474 28656
rect 39333 28625 39345 28628
rect 39287 28619 39345 28625
rect 39468 28616 39474 28628
rect 39526 28656 39532 28668
rect 40664 28656 40670 28668
rect 39526 28628 40670 28656
rect 39526 28616 39532 28628
rect 40664 28616 40670 28628
rect 40722 28656 40728 28668
rect 43166 28665 43194 28696
rect 43792 28684 43798 28696
rect 43850 28684 43856 28736
rect 43151 28659 43209 28665
rect 40722 28628 43102 28656
rect 40722 28616 40728 28628
rect 42967 28591 43025 28597
rect 42967 28588 42979 28591
rect 38658 28560 38962 28588
rect 26637 28492 27830 28520
rect 26637 28489 26649 28492
rect 26591 28483 26649 28489
rect 27968 28480 27974 28532
rect 28026 28520 28032 28532
rect 31096 28520 31102 28532
rect 28026 28492 31102 28520
rect 28026 28480 28032 28492
rect 31096 28480 31102 28492
rect 31154 28480 31160 28532
rect 35880 28480 35886 28532
rect 35938 28520 35944 28532
rect 36892 28520 36898 28532
rect 35938 28492 36898 28520
rect 35938 28480 35944 28492
rect 36892 28480 36898 28492
rect 36950 28480 36956 28532
rect 38934 28520 38962 28560
rect 42890 28560 42979 28588
rect 39836 28520 39842 28532
rect 38934 28492 39842 28520
rect 39836 28480 39842 28492
rect 39894 28480 39900 28532
rect 42890 28464 42918 28560
rect 42967 28557 42979 28560
rect 43013 28557 43025 28591
rect 42967 28551 43025 28557
rect 43074 28520 43102 28628
rect 43151 28625 43163 28659
rect 43197 28625 43209 28659
rect 43151 28619 43209 28625
rect 43516 28616 43522 28668
rect 43574 28656 43580 28668
rect 43902 28665 43930 28764
rect 45540 28752 45546 28804
rect 45598 28792 45604 28804
rect 54924 28792 54930 28804
rect 45598 28764 54930 28792
rect 45598 28752 45604 28764
rect 54924 28752 54930 28764
rect 54982 28752 54988 28804
rect 56396 28792 56402 28804
rect 55126 28764 55982 28792
rect 56357 28764 56402 28792
rect 50143 28727 50201 28733
rect 50143 28724 50155 28727
rect 49514 28696 50155 28724
rect 43703 28659 43761 28665
rect 43703 28656 43715 28659
rect 43574 28628 43715 28656
rect 43574 28616 43580 28628
rect 43703 28625 43715 28628
rect 43749 28625 43761 28659
rect 43703 28619 43761 28625
rect 43887 28659 43945 28665
rect 43887 28625 43899 28659
rect 43933 28625 43945 28659
rect 49312 28656 49318 28668
rect 49273 28628 49318 28656
rect 43887 28619 43945 28625
rect 49312 28616 49318 28628
rect 49370 28616 49376 28668
rect 47932 28548 47938 28600
rect 47990 28588 47996 28600
rect 49223 28591 49281 28597
rect 49223 28588 49235 28591
rect 47990 28560 49235 28588
rect 47990 28548 47996 28560
rect 49223 28557 49235 28560
rect 49269 28588 49281 28591
rect 49514 28588 49542 28696
rect 50143 28693 50155 28696
rect 50189 28693 50201 28727
rect 50143 28687 50201 28693
rect 49680 28656 49686 28668
rect 49593 28628 49686 28656
rect 49680 28616 49686 28628
rect 49738 28656 49744 28668
rect 50048 28656 50054 28668
rect 49738 28628 50054 28656
rect 49738 28616 49744 28628
rect 50048 28616 50054 28628
rect 50106 28616 50112 28668
rect 49269 28560 49542 28588
rect 49269 28557 49281 28560
rect 49223 28551 49281 28557
rect 49698 28520 49726 28616
rect 49775 28591 49833 28597
rect 49775 28557 49787 28591
rect 49821 28557 49833 28591
rect 50158 28588 50186 28687
rect 50324 28684 50330 28736
rect 50382 28724 50388 28736
rect 55126 28724 55154 28764
rect 50382 28696 55154 28724
rect 55954 28724 55982 28764
rect 56396 28752 56402 28764
rect 56454 28752 56460 28804
rect 67347 28795 67405 28801
rect 56506 28764 64998 28792
rect 56506 28724 56534 28764
rect 55954 28696 56534 28724
rect 50382 28684 50388 28696
rect 56580 28684 56586 28736
rect 56638 28724 56644 28736
rect 61183 28727 61241 28733
rect 61183 28724 61195 28727
rect 56638 28696 61195 28724
rect 56638 28684 56644 28696
rect 61183 28693 61195 28696
rect 61229 28693 61241 28727
rect 61183 28687 61241 28693
rect 62744 28684 62750 28736
rect 62802 28724 62808 28736
rect 63759 28727 63817 28733
rect 63759 28724 63771 28727
rect 62802 28696 63771 28724
rect 62802 28684 62808 28696
rect 63759 28693 63771 28696
rect 63805 28724 63817 28727
rect 64400 28724 64406 28736
rect 63805 28696 64406 28724
rect 63805 28693 63817 28696
rect 63759 28687 63817 28693
rect 64400 28684 64406 28696
rect 64458 28684 64464 28736
rect 64970 28724 64998 28764
rect 67347 28761 67359 28795
rect 67393 28792 67405 28795
rect 67896 28792 67902 28804
rect 67393 28764 67902 28792
rect 67393 28761 67405 28764
rect 67347 28755 67405 28761
rect 67896 28752 67902 28764
rect 67954 28752 67960 28804
rect 67988 28752 67994 28804
rect 68046 28792 68052 28804
rect 68451 28795 68509 28801
rect 68451 28792 68463 28795
rect 68046 28764 68463 28792
rect 68046 28752 68052 28764
rect 68451 28761 68463 28764
rect 68497 28761 68509 28795
rect 68451 28755 68509 28761
rect 69000 28752 69006 28804
rect 69058 28792 69064 28804
rect 71579 28795 71637 28801
rect 71579 28792 71591 28795
rect 69058 28764 71591 28792
rect 69058 28752 69064 28764
rect 71579 28761 71591 28764
rect 71625 28761 71637 28795
rect 71579 28755 71637 28761
rect 72407 28795 72465 28801
rect 72407 28761 72419 28795
rect 72453 28792 72465 28795
rect 74612 28792 74618 28804
rect 72453 28764 74618 28792
rect 72453 28761 72465 28764
rect 72407 28755 72465 28761
rect 69460 28724 69466 28736
rect 64970 28696 69466 28724
rect 69460 28684 69466 28696
rect 69518 28684 69524 28736
rect 50695 28659 50753 28665
rect 50695 28625 50707 28659
rect 50741 28656 50753 28659
rect 51888 28656 51894 28668
rect 50741 28628 51894 28656
rect 50741 28625 50753 28628
rect 50695 28619 50753 28625
rect 51888 28616 51894 28628
rect 51946 28616 51952 28668
rect 52072 28656 52078 28668
rect 52033 28628 52078 28656
rect 52072 28616 52078 28628
rect 52130 28616 52136 28668
rect 52808 28656 52814 28668
rect 52182 28628 52670 28656
rect 52769 28628 52814 28656
rect 51796 28588 51802 28600
rect 50158 28560 51802 28588
rect 49775 28551 49833 28557
rect 43074 28492 49726 28520
rect 49790 28520 49818 28551
rect 51796 28548 51802 28560
rect 51854 28548 51860 28600
rect 50051 28523 50109 28529
rect 50051 28520 50063 28523
rect 49790 28492 50063 28520
rect 50051 28489 50063 28492
rect 50097 28520 50109 28523
rect 50416 28520 50422 28532
rect 50097 28492 50422 28520
rect 50097 28489 50109 28492
rect 50051 28483 50109 28489
rect 50416 28480 50422 28492
rect 50474 28480 50480 28532
rect 50876 28520 50882 28532
rect 50837 28492 50882 28520
rect 50876 28480 50882 28492
rect 50934 28480 50940 28532
rect 25392 28452 25398 28464
rect 23794 28424 24518 28452
rect 25353 28424 25398 28452
rect 23794 28412 23800 28424
rect 25392 28412 25398 28424
rect 25450 28412 25456 28464
rect 25484 28412 25490 28464
rect 25542 28452 25548 28464
rect 28063 28455 28121 28461
rect 28063 28452 28075 28455
rect 25542 28424 28075 28452
rect 25542 28412 25548 28424
rect 28063 28421 28075 28424
rect 28109 28421 28121 28455
rect 28336 28452 28342 28464
rect 28297 28424 28342 28452
rect 28063 28415 28121 28421
rect 28336 28412 28342 28424
rect 28394 28412 28400 28464
rect 28520 28412 28526 28464
rect 28578 28452 28584 28464
rect 28983 28455 29041 28461
rect 28983 28452 28995 28455
rect 28578 28424 28995 28452
rect 28578 28412 28584 28424
rect 28983 28421 28995 28424
rect 29029 28452 29041 28455
rect 29716 28452 29722 28464
rect 29029 28424 29722 28452
rect 29029 28421 29041 28424
rect 28983 28415 29041 28421
rect 29716 28412 29722 28424
rect 29774 28452 29780 28464
rect 30820 28452 30826 28464
rect 29774 28424 30826 28452
rect 29774 28412 29780 28424
rect 30820 28412 30826 28424
rect 30878 28452 30884 28464
rect 31004 28452 31010 28464
rect 30878 28424 31010 28452
rect 30878 28412 30884 28424
rect 31004 28412 31010 28424
rect 31062 28412 31068 28464
rect 38364 28452 38370 28464
rect 38325 28424 38370 28452
rect 38364 28412 38370 28424
rect 38422 28452 38428 28464
rect 39192 28452 39198 28464
rect 38422 28424 39198 28452
rect 38422 28412 38428 28424
rect 39192 28412 39198 28424
rect 39250 28412 39256 28464
rect 39744 28452 39750 28464
rect 39705 28424 39750 28452
rect 39744 28412 39750 28424
rect 39802 28412 39808 28464
rect 42599 28455 42657 28461
rect 42599 28421 42611 28455
rect 42645 28452 42657 28455
rect 42872 28452 42878 28464
rect 42645 28424 42878 28452
rect 42645 28421 42657 28424
rect 42599 28415 42657 28421
rect 42872 28412 42878 28424
rect 42930 28412 42936 28464
rect 44163 28455 44221 28461
rect 44163 28421 44175 28455
rect 44209 28452 44221 28455
rect 45264 28452 45270 28464
rect 44209 28424 45270 28452
rect 44209 28421 44221 28424
rect 44163 28415 44221 28421
rect 45264 28412 45270 28424
rect 45322 28412 45328 28464
rect 47748 28412 47754 28464
rect 47806 28452 47812 28464
rect 48763 28455 48821 28461
rect 48763 28452 48775 28455
rect 47806 28424 48775 28452
rect 47806 28412 47812 28424
rect 48763 28421 48775 28424
rect 48809 28421 48821 28455
rect 48763 28415 48821 28421
rect 48852 28412 48858 28464
rect 48910 28452 48916 28464
rect 52182 28452 52210 28628
rect 52348 28548 52354 28600
rect 52406 28588 52412 28600
rect 52443 28591 52501 28597
rect 52443 28588 52455 28591
rect 52406 28560 52455 28588
rect 52406 28548 52412 28560
rect 52443 28557 52455 28560
rect 52489 28557 52501 28591
rect 52642 28588 52670 28628
rect 52808 28616 52814 28628
rect 52866 28616 52872 28668
rect 53820 28656 53826 28668
rect 52918 28628 53826 28656
rect 52918 28588 52946 28628
rect 53820 28616 53826 28628
rect 53878 28616 53884 28668
rect 54007 28659 54065 28665
rect 54007 28625 54019 28659
rect 54053 28656 54065 28659
rect 54188 28656 54194 28668
rect 54053 28628 54194 28656
rect 54053 28625 54065 28628
rect 54007 28619 54065 28625
rect 54188 28616 54194 28628
rect 54246 28616 54252 28668
rect 55292 28656 55298 28668
rect 55253 28628 55298 28656
rect 55292 28616 55298 28628
rect 55350 28616 55356 28668
rect 57500 28656 57506 28668
rect 57461 28628 57506 28656
rect 57500 28616 57506 28628
rect 57558 28616 57564 28668
rect 59524 28616 59530 28668
rect 59582 28656 59588 28668
rect 59619 28659 59677 28665
rect 59619 28656 59631 28659
rect 59582 28628 59631 28656
rect 59582 28616 59588 28628
rect 59619 28625 59631 28628
rect 59665 28625 59677 28659
rect 63204 28656 63210 28668
rect 59619 28619 59677 28625
rect 60278 28628 63210 28656
rect 52642 28560 52946 28588
rect 52443 28551 52501 28557
rect 52992 28548 52998 28600
rect 53050 28588 53056 28600
rect 53050 28560 54234 28588
rect 53050 28548 53056 28560
rect 52240 28523 52298 28529
rect 52240 28489 52252 28523
rect 52286 28520 52298 28523
rect 53820 28520 53826 28532
rect 52286 28492 53826 28520
rect 52286 28489 52298 28492
rect 52240 28483 52298 28489
rect 53820 28480 53826 28492
rect 53878 28480 53884 28532
rect 52351 28455 52409 28461
rect 52351 28452 52363 28455
rect 48910 28424 52363 28452
rect 48910 28412 48916 28424
rect 52351 28421 52363 28424
rect 52397 28421 52409 28455
rect 52351 28415 52409 28421
rect 53636 28412 53642 28464
rect 53694 28452 53700 28464
rect 54099 28455 54157 28461
rect 54099 28452 54111 28455
rect 53694 28424 54111 28452
rect 53694 28412 53700 28424
rect 54099 28421 54111 28424
rect 54145 28421 54157 28455
rect 54206 28452 54234 28560
rect 54280 28548 54286 28600
rect 54338 28588 54344 28600
rect 55019 28591 55077 28597
rect 55019 28588 55031 28591
rect 54338 28560 55031 28588
rect 54338 28548 54344 28560
rect 55019 28557 55031 28560
rect 55065 28588 55077 28591
rect 56488 28588 56494 28600
rect 55065 28560 56494 28588
rect 55065 28557 55077 28560
rect 55019 28551 55077 28557
rect 56488 28548 56494 28560
rect 56546 28588 56552 28600
rect 56767 28591 56825 28597
rect 56767 28588 56779 28591
rect 56546 28560 56779 28588
rect 56546 28548 56552 28560
rect 56767 28557 56779 28560
rect 56813 28557 56825 28591
rect 60278 28588 60306 28628
rect 63204 28616 63210 28628
rect 63262 28616 63268 28668
rect 63296 28616 63302 28668
rect 63354 28656 63360 28668
rect 63943 28659 64001 28665
rect 63943 28656 63955 28659
rect 63354 28628 63955 28656
rect 63354 28616 63360 28628
rect 63943 28625 63955 28628
rect 63989 28625 64001 28659
rect 67160 28656 67166 28668
rect 67121 28628 67166 28656
rect 63943 28619 64001 28625
rect 67160 28616 67166 28628
rect 67218 28616 67224 28668
rect 68267 28659 68325 28665
rect 68267 28625 68279 28659
rect 68313 28656 68325 28659
rect 69368 28656 69374 28668
rect 68313 28628 69374 28656
rect 68313 28625 68325 28628
rect 68267 28619 68325 28625
rect 69368 28616 69374 28628
rect 69426 28616 69432 28668
rect 56767 28551 56825 28557
rect 56874 28560 60306 28588
rect 56874 28452 56902 28560
rect 61180 28548 61186 28600
rect 61238 28588 61244 28600
rect 61275 28591 61333 28597
rect 61275 28588 61287 28591
rect 61238 28560 61287 28588
rect 61238 28548 61244 28560
rect 61275 28557 61287 28560
rect 61321 28557 61333 28591
rect 61275 28551 61333 28557
rect 61551 28591 61609 28597
rect 61551 28557 61563 28591
rect 61597 28588 61609 28591
rect 64216 28588 64222 28600
rect 61597 28560 64222 28588
rect 61597 28557 61609 28560
rect 61551 28551 61609 28557
rect 64216 28548 64222 28560
rect 64274 28548 64280 28600
rect 71594 28588 71622 28755
rect 74612 28752 74618 28764
rect 74670 28752 74676 28804
rect 81055 28795 81113 28801
rect 81055 28761 81067 28795
rect 81101 28792 81113 28795
rect 81236 28792 81242 28804
rect 81101 28764 81242 28792
rect 81101 28761 81113 28764
rect 81055 28755 81113 28761
rect 81236 28752 81242 28764
rect 81294 28752 81300 28804
rect 84180 28752 84186 28804
rect 84238 28792 84244 28804
rect 85655 28795 85713 28801
rect 85655 28792 85667 28795
rect 84238 28764 85667 28792
rect 84238 28752 84244 28764
rect 85655 28761 85667 28764
rect 85701 28761 85713 28795
rect 85655 28755 85713 28761
rect 89240 28752 89246 28804
rect 89298 28792 89304 28804
rect 90531 28795 90589 28801
rect 90531 28792 90543 28795
rect 89298 28764 90543 28792
rect 89298 28752 89304 28764
rect 90531 28761 90543 28764
rect 90577 28761 90589 28795
rect 90531 28755 90589 28761
rect 90712 28752 90718 28804
rect 90770 28792 90776 28804
rect 91911 28795 91969 28801
rect 91911 28792 91923 28795
rect 90770 28764 91923 28792
rect 90770 28752 90776 28764
rect 91911 28761 91923 28764
rect 91957 28761 91969 28795
rect 91911 28755 91969 28761
rect 73232 28724 73238 28736
rect 73193 28696 73238 28724
rect 73232 28684 73238 28696
rect 73290 28724 73296 28736
rect 73511 28727 73569 28733
rect 73290 28696 73370 28724
rect 73290 28684 73296 28696
rect 71668 28616 71674 28668
rect 71726 28656 71732 28668
rect 73342 28665 73370 28696
rect 73511 28693 73523 28727
rect 73557 28724 73569 28727
rect 73876 28724 73882 28736
rect 73557 28696 73882 28724
rect 73557 28693 73569 28696
rect 73511 28687 73569 28693
rect 73876 28684 73882 28696
rect 73934 28684 73940 28736
rect 71763 28659 71821 28665
rect 71763 28656 71775 28659
rect 71726 28628 71775 28656
rect 71726 28616 71732 28628
rect 71763 28625 71775 28628
rect 71809 28625 71821 28659
rect 71763 28619 71821 28625
rect 73327 28659 73385 28665
rect 73327 28625 73339 28659
rect 73373 28625 73385 28659
rect 73600 28656 73606 28668
rect 73561 28628 73606 28656
rect 73327 28619 73385 28625
rect 73600 28616 73606 28628
rect 73658 28616 73664 28668
rect 79212 28616 79218 28668
rect 79270 28656 79276 28668
rect 79399 28659 79457 28665
rect 79399 28656 79411 28659
rect 79270 28628 79411 28656
rect 79270 28616 79276 28628
rect 79399 28625 79411 28628
rect 79445 28656 79457 28659
rect 79488 28656 79494 28668
rect 79445 28628 79494 28656
rect 79445 28625 79457 28628
rect 79399 28619 79457 28625
rect 79488 28616 79494 28628
rect 79546 28616 79552 28668
rect 90068 28656 90074 28668
rect 90029 28628 90074 28656
rect 90068 28616 90074 28628
rect 90126 28616 90132 28668
rect 90344 28656 90350 28668
rect 90305 28628 90350 28656
rect 90344 28616 90350 28628
rect 90402 28616 90408 28668
rect 91080 28616 91086 28668
rect 91138 28656 91144 28668
rect 91635 28659 91693 28665
rect 91635 28656 91647 28659
rect 91138 28628 91647 28656
rect 91138 28616 91144 28628
rect 91635 28625 91647 28628
rect 91681 28625 91693 28659
rect 91816 28656 91822 28668
rect 91777 28628 91822 28656
rect 91635 28619 91693 28625
rect 91816 28616 91822 28628
rect 91874 28616 91880 28668
rect 72131 28591 72189 28597
rect 72131 28588 72143 28591
rect 71594 28560 72143 28588
rect 72131 28557 72143 28560
rect 72177 28557 72189 28591
rect 74060 28588 74066 28600
rect 74021 28560 74066 28588
rect 72131 28551 72189 28557
rect 74060 28548 74066 28560
rect 74118 28548 74124 28600
rect 79767 28591 79825 28597
rect 79767 28557 79779 28591
rect 79813 28588 79825 28591
rect 80408 28588 80414 28600
rect 79813 28560 80414 28588
rect 79813 28557 79825 28560
rect 79767 28551 79825 28557
rect 80408 28548 80414 28560
rect 80466 28548 80472 28600
rect 84275 28591 84333 28597
rect 84275 28557 84287 28591
rect 84321 28557 84333 28591
rect 84548 28588 84554 28600
rect 84509 28560 84554 28588
rect 84275 28551 84333 28557
rect 62652 28520 62658 28532
rect 62613 28492 62658 28520
rect 62652 28480 62658 28492
rect 62710 28480 62716 28532
rect 64768 28520 64774 28532
rect 62762 28492 64774 28520
rect 54206 28424 56902 28452
rect 54099 28415 54157 28421
rect 57592 28412 57598 28464
rect 57650 28452 57656 28464
rect 57687 28455 57745 28461
rect 57687 28452 57699 28455
rect 57650 28424 57699 28452
rect 57650 28412 57656 28424
rect 57687 28421 57699 28424
rect 57733 28421 57745 28455
rect 59800 28452 59806 28464
rect 59761 28424 59806 28452
rect 57687 28415 57745 28421
rect 59800 28412 59806 28424
rect 59858 28412 59864 28464
rect 61183 28455 61241 28461
rect 61183 28421 61195 28455
rect 61229 28452 61241 28455
rect 62762 28452 62790 28492
rect 64768 28480 64774 28492
rect 64826 28480 64832 28532
rect 69463 28523 69521 28529
rect 69463 28489 69475 28523
rect 69509 28520 69521 28523
rect 69736 28520 69742 28532
rect 69509 28492 69742 28520
rect 69509 28489 69521 28492
rect 69463 28483 69521 28489
rect 69736 28480 69742 28492
rect 69794 28520 69800 28532
rect 72039 28523 72097 28529
rect 72039 28520 72051 28523
rect 69794 28492 72051 28520
rect 69794 28480 69800 28492
rect 72039 28489 72051 28492
rect 72085 28489 72097 28523
rect 72039 28483 72097 28489
rect 61229 28424 62790 28452
rect 64035 28455 64093 28461
rect 61229 28421 61241 28424
rect 61183 28415 61241 28421
rect 64035 28421 64047 28455
rect 64081 28452 64093 28455
rect 64124 28452 64130 28464
rect 64081 28424 64130 28452
rect 64081 28421 64093 28424
rect 64035 28415 64093 28421
rect 64124 28412 64130 28424
rect 64182 28412 64188 28464
rect 71928 28455 71986 28461
rect 71928 28421 71940 28455
rect 71974 28452 71986 28455
rect 72680 28452 72686 28464
rect 71974 28424 72686 28452
rect 71974 28421 71986 28424
rect 71928 28415 71986 28421
rect 72680 28412 72686 28424
rect 72738 28412 72744 28464
rect 84183 28455 84241 28461
rect 84183 28421 84195 28455
rect 84229 28452 84241 28455
rect 84290 28452 84318 28551
rect 84548 28548 84554 28560
rect 84606 28548 84612 28600
rect 90163 28523 90221 28529
rect 90163 28489 90175 28523
rect 90209 28520 90221 28523
rect 90620 28520 90626 28532
rect 90209 28492 90626 28520
rect 90209 28489 90221 28492
rect 90163 28483 90221 28489
rect 90620 28480 90626 28492
rect 90678 28480 90684 28532
rect 85192 28452 85198 28464
rect 84229 28424 85198 28452
rect 84229 28421 84241 28424
rect 84183 28415 84241 28421
rect 85192 28412 85198 28424
rect 85250 28452 85256 28464
rect 85560 28452 85566 28464
rect 85250 28424 85566 28452
rect 85250 28412 85256 28424
rect 85560 28412 85566 28424
rect 85618 28412 85624 28464
rect 538 28362 93642 28384
rect 538 28310 3680 28362
rect 3732 28310 3744 28362
rect 3796 28310 3808 28362
rect 3860 28310 3872 28362
rect 3924 28310 9008 28362
rect 9060 28310 9072 28362
rect 9124 28310 9136 28362
rect 9188 28310 9200 28362
rect 9252 28310 14336 28362
rect 14388 28310 14400 28362
rect 14452 28310 14464 28362
rect 14516 28310 14528 28362
rect 14580 28310 19664 28362
rect 19716 28310 19728 28362
rect 19780 28310 19792 28362
rect 19844 28310 19856 28362
rect 19908 28310 24992 28362
rect 25044 28310 25056 28362
rect 25108 28310 25120 28362
rect 25172 28310 25184 28362
rect 25236 28310 30320 28362
rect 30372 28310 30384 28362
rect 30436 28310 30448 28362
rect 30500 28310 30512 28362
rect 30564 28310 35648 28362
rect 35700 28310 35712 28362
rect 35764 28310 35776 28362
rect 35828 28310 35840 28362
rect 35892 28310 40976 28362
rect 41028 28310 41040 28362
rect 41092 28310 41104 28362
rect 41156 28310 41168 28362
rect 41220 28310 46304 28362
rect 46356 28310 46368 28362
rect 46420 28310 46432 28362
rect 46484 28310 46496 28362
rect 46548 28310 51632 28362
rect 51684 28310 51696 28362
rect 51748 28310 51760 28362
rect 51812 28310 51824 28362
rect 51876 28310 56960 28362
rect 57012 28310 57024 28362
rect 57076 28310 57088 28362
rect 57140 28310 57152 28362
rect 57204 28310 62288 28362
rect 62340 28310 62352 28362
rect 62404 28310 62416 28362
rect 62468 28310 62480 28362
rect 62532 28310 67616 28362
rect 67668 28310 67680 28362
rect 67732 28310 67744 28362
rect 67796 28310 67808 28362
rect 67860 28310 72944 28362
rect 72996 28310 73008 28362
rect 73060 28310 73072 28362
rect 73124 28310 73136 28362
rect 73188 28310 78272 28362
rect 78324 28310 78336 28362
rect 78388 28310 78400 28362
rect 78452 28310 78464 28362
rect 78516 28310 83600 28362
rect 83652 28310 83664 28362
rect 83716 28310 83728 28362
rect 83780 28310 83792 28362
rect 83844 28310 88928 28362
rect 88980 28310 88992 28362
rect 89044 28310 89056 28362
rect 89108 28310 89120 28362
rect 89172 28310 93642 28362
rect 538 28288 93642 28310
rect 3036 28248 3042 28260
rect 2997 28220 3042 28248
rect 3036 28208 3042 28220
rect 3094 28208 3100 28260
rect 12880 28208 12886 28260
rect 12938 28248 12944 28260
rect 13524 28248 13530 28260
rect 12938 28220 13530 28248
rect 12938 28208 12944 28220
rect 13524 28208 13530 28220
rect 13582 28208 13588 28260
rect 15088 28248 15094 28260
rect 15049 28220 15094 28248
rect 15088 28208 15094 28220
rect 15146 28208 15152 28260
rect 15916 28208 15922 28260
rect 15974 28248 15980 28260
rect 20976 28248 20982 28260
rect 15974 28220 20982 28248
rect 15974 28208 15980 28220
rect 20976 28208 20982 28220
rect 21034 28208 21040 28260
rect 21807 28251 21865 28257
rect 21807 28217 21819 28251
rect 21853 28248 21865 28251
rect 21853 28220 27830 28248
rect 21853 28217 21865 28220
rect 21807 28211 21865 28217
rect 8096 28140 8102 28192
rect 8154 28180 8160 28192
rect 9203 28183 9261 28189
rect 9203 28180 9215 28183
rect 8154 28152 9215 28180
rect 8154 28140 8160 28152
rect 9203 28149 9215 28152
rect 9249 28180 9261 28183
rect 13248 28180 13254 28192
rect 9249 28152 13110 28180
rect 13209 28152 13254 28180
rect 9249 28149 9261 28152
rect 9203 28143 9261 28149
rect 920 28072 926 28124
rect 978 28112 984 28124
rect 1659 28115 1717 28121
rect 1659 28112 1671 28115
rect 978 28084 1671 28112
rect 978 28072 984 28084
rect 1659 28081 1671 28084
rect 1705 28112 1717 28115
rect 2300 28112 2306 28124
rect 1705 28084 2306 28112
rect 1705 28081 1717 28084
rect 1659 28075 1717 28081
rect 2300 28072 2306 28084
rect 2358 28112 2364 28124
rect 3499 28115 3557 28121
rect 3499 28112 3511 28115
rect 2358 28084 3511 28112
rect 2358 28072 2364 28084
rect 3499 28081 3511 28084
rect 3545 28112 3557 28115
rect 6164 28112 6170 28124
rect 3545 28084 6170 28112
rect 3545 28081 3557 28084
rect 3499 28075 3557 28081
rect 6164 28072 6170 28084
rect 6222 28112 6228 28124
rect 6627 28115 6685 28121
rect 6627 28112 6639 28115
rect 6222 28084 6639 28112
rect 6222 28072 6228 28084
rect 6627 28081 6639 28084
rect 6673 28112 6685 28115
rect 8556 28112 8562 28124
rect 6673 28084 8562 28112
rect 6673 28081 6685 28084
rect 6627 28075 6685 28081
rect 8556 28072 8562 28084
rect 8614 28072 8620 28124
rect 11871 28115 11929 28121
rect 11871 28081 11883 28115
rect 11917 28112 11929 28115
rect 11960 28112 11966 28124
rect 11917 28084 11966 28112
rect 11917 28081 11929 28084
rect 11871 28075 11929 28081
rect 11960 28072 11966 28084
rect 12018 28072 12024 28124
rect 1932 28044 1938 28056
rect 1893 28016 1938 28044
rect 1932 28004 1938 28016
rect 1990 28004 1996 28056
rect 6903 28047 6961 28053
rect 6903 28013 6915 28047
rect 6949 28044 6961 28047
rect 7728 28044 7734 28056
rect 6949 28016 7734 28044
rect 6949 28013 6961 28016
rect 6903 28007 6961 28013
rect 7728 28004 7734 28016
rect 7786 28004 7792 28056
rect 8283 28047 8341 28053
rect 8283 28013 8295 28047
rect 8329 28044 8341 28047
rect 9111 28047 9169 28053
rect 9111 28044 9123 28047
rect 8329 28016 9123 28044
rect 8329 28013 8341 28016
rect 8283 28007 8341 28013
rect 9111 28013 9123 28016
rect 9157 28044 9169 28047
rect 9476 28044 9482 28056
rect 9157 28016 9482 28044
rect 9157 28013 9169 28016
rect 9111 28007 9169 28013
rect 9476 28004 9482 28016
rect 9534 28004 9540 28056
rect 10948 28004 10954 28056
rect 11006 28044 11012 28056
rect 12055 28047 12113 28053
rect 12055 28044 12067 28047
rect 11006 28016 12067 28044
rect 11006 28004 11012 28016
rect 12055 28013 12067 28016
rect 12101 28013 12113 28047
rect 12055 28007 12113 28013
rect 12236 28004 12242 28056
rect 12294 28044 12300 28056
rect 12423 28047 12481 28053
rect 12423 28044 12435 28047
rect 12294 28016 12435 28044
rect 12294 28004 12300 28016
rect 12423 28013 12435 28016
rect 12469 28013 12481 28047
rect 12696 28044 12702 28056
rect 12657 28016 12702 28044
rect 12423 28007 12481 28013
rect 12696 28004 12702 28016
rect 12754 28004 12760 28056
rect 12880 28044 12886 28056
rect 12841 28016 12886 28044
rect 12880 28004 12886 28016
rect 12938 28004 12944 28056
rect 11687 27979 11745 27985
rect 11687 27976 11699 27979
rect 7562 27948 11699 27976
rect 4048 27868 4054 27920
rect 4106 27908 4112 27920
rect 7562 27908 7590 27948
rect 11687 27945 11699 27948
rect 11733 27976 11745 27979
rect 12714 27976 12742 28004
rect 11733 27948 12742 27976
rect 13082 27976 13110 28152
rect 13248 28140 13254 28152
rect 13306 28140 13312 28192
rect 15180 28140 15186 28192
rect 15238 28180 15244 28192
rect 15367 28183 15425 28189
rect 15367 28180 15379 28183
rect 15238 28152 15379 28180
rect 15238 28140 15244 28152
rect 15367 28149 15379 28152
rect 15413 28180 15425 28183
rect 17388 28180 17394 28192
rect 15413 28152 17394 28180
rect 15413 28149 15425 28152
rect 15367 28143 15425 28149
rect 15643 28047 15701 28053
rect 15643 28013 15655 28047
rect 15689 28044 15701 28047
rect 15732 28044 15738 28056
rect 15689 28016 15738 28044
rect 15689 28013 15701 28016
rect 15643 28007 15701 28013
rect 15732 28004 15738 28016
rect 15790 28004 15796 28056
rect 15934 28053 15962 28152
rect 17388 28140 17394 28152
rect 17446 28140 17452 28192
rect 21822 28180 21850 28211
rect 21086 28152 21850 28180
rect 16192 28072 16198 28124
rect 16250 28112 16256 28124
rect 16379 28115 16437 28121
rect 16379 28112 16391 28115
rect 16250 28084 16391 28112
rect 16250 28072 16256 28084
rect 16379 28081 16391 28084
rect 16425 28081 16437 28115
rect 16379 28075 16437 28081
rect 16652 28072 16658 28124
rect 16710 28112 16716 28124
rect 17756 28112 17762 28124
rect 16710 28084 17762 28112
rect 16710 28072 16716 28084
rect 17756 28072 17762 28084
rect 17814 28112 17820 28124
rect 17943 28115 18001 28121
rect 17943 28112 17955 28115
rect 17814 28084 17955 28112
rect 17814 28072 17820 28084
rect 17943 28081 17955 28084
rect 17989 28081 18001 28115
rect 18216 28112 18222 28124
rect 18177 28084 18222 28112
rect 17943 28075 18001 28081
rect 18216 28072 18222 28084
rect 18274 28072 18280 28124
rect 19320 28112 19326 28124
rect 19281 28084 19326 28112
rect 19320 28072 19326 28084
rect 19378 28072 19384 28124
rect 21086 28121 21114 28152
rect 23920 28140 23926 28192
rect 23978 28180 23984 28192
rect 24015 28183 24073 28189
rect 24015 28180 24027 28183
rect 23978 28152 24027 28180
rect 23978 28140 23984 28152
rect 24015 28149 24027 28152
rect 24061 28180 24073 28183
rect 27692 28180 27698 28192
rect 24061 28152 24242 28180
rect 27653 28152 27698 28180
rect 24061 28149 24073 28152
rect 24015 28143 24073 28149
rect 24214 28121 24242 28152
rect 27692 28140 27698 28152
rect 27750 28140 27756 28192
rect 27802 28180 27830 28220
rect 28336 28208 28342 28260
rect 28394 28248 28400 28260
rect 35144 28248 35150 28260
rect 28394 28220 35150 28248
rect 28394 28208 28400 28220
rect 35144 28208 35150 28220
rect 35202 28208 35208 28260
rect 35254 28220 35558 28248
rect 30728 28180 30734 28192
rect 27802 28152 30734 28180
rect 30728 28140 30734 28152
rect 30786 28140 30792 28192
rect 31559 28183 31617 28189
rect 31559 28180 31571 28183
rect 30930 28152 31571 28180
rect 21071 28115 21129 28121
rect 21071 28081 21083 28115
rect 21117 28081 21129 28115
rect 21071 28075 21129 28081
rect 24199 28115 24257 28121
rect 24199 28081 24211 28115
rect 24245 28081 24257 28115
rect 24199 28075 24257 28081
rect 24380 28072 24386 28124
rect 24438 28112 24444 28124
rect 30636 28112 30642 28124
rect 24438 28084 30642 28112
rect 24438 28072 24444 28084
rect 30636 28072 30642 28084
rect 30694 28072 30700 28124
rect 30930 28112 30958 28152
rect 31559 28149 31571 28152
rect 31605 28180 31617 28183
rect 35254 28180 35282 28220
rect 35420 28180 35426 28192
rect 31605 28152 35282 28180
rect 35381 28152 35426 28180
rect 31605 28149 31617 28152
rect 31559 28143 31617 28149
rect 35420 28140 35426 28152
rect 35478 28140 35484 28192
rect 35530 28180 35558 28220
rect 36892 28208 36898 28260
rect 36950 28248 36956 28260
rect 40572 28248 40578 28260
rect 36950 28220 40578 28248
rect 36950 28208 36956 28220
rect 40572 28208 40578 28220
rect 40630 28208 40636 28260
rect 46092 28208 46098 28260
rect 46150 28248 46156 28260
rect 46150 28220 49266 28248
rect 46150 28208 46156 28220
rect 38180 28180 38186 28192
rect 35530 28152 38186 28180
rect 38180 28140 38186 28152
rect 38238 28140 38244 28192
rect 39192 28140 39198 28192
rect 39250 28180 39256 28192
rect 40207 28183 40265 28189
rect 40207 28180 40219 28183
rect 39250 28152 40219 28180
rect 39250 28140 39256 28152
rect 40207 28149 40219 28152
rect 40253 28180 40265 28183
rect 41771 28183 41829 28189
rect 40253 28152 40618 28180
rect 40253 28149 40265 28152
rect 40207 28143 40265 28149
rect 31191 28115 31249 28121
rect 31191 28112 31203 28115
rect 30746 28084 30958 28112
rect 31022 28084 31203 28112
rect 15919 28047 15977 28053
rect 15919 28013 15931 28047
rect 15965 28013 15977 28047
rect 15919 28007 15977 28013
rect 16100 28004 16106 28056
rect 16158 28044 16164 28056
rect 16287 28047 16345 28053
rect 16287 28044 16299 28047
rect 16158 28016 16299 28044
rect 16158 28004 16164 28016
rect 16287 28013 16299 28016
rect 16333 28013 16345 28047
rect 18860 28044 18866 28056
rect 16287 28007 16345 28013
rect 17314 28016 18866 28044
rect 17314 27976 17342 28016
rect 18860 28004 18866 28016
rect 18918 28004 18924 28056
rect 20976 28044 20982 28056
rect 20937 28016 20982 28044
rect 20976 28004 20982 28016
rect 21034 28044 21040 28056
rect 21183 28047 21241 28053
rect 21183 28044 21195 28047
rect 21034 28016 21195 28044
rect 21034 28004 21040 28016
rect 21183 28013 21195 28016
rect 21229 28013 21241 28047
rect 21183 28007 21241 28013
rect 21344 28004 21350 28056
rect 21402 28044 21408 28056
rect 21623 28047 21681 28053
rect 21623 28044 21635 28047
rect 21402 28016 21635 28044
rect 21402 28004 21408 28016
rect 21623 28013 21635 28016
rect 21669 28013 21681 28047
rect 21623 28007 21681 28013
rect 23095 28047 23153 28053
rect 23095 28013 23107 28047
rect 23141 28044 23153 28047
rect 23552 28044 23558 28056
rect 23141 28016 23558 28044
rect 23141 28013 23153 28016
rect 23095 28007 23153 28013
rect 23552 28004 23558 28016
rect 23610 28044 23616 28056
rect 24012 28044 24018 28056
rect 23610 28016 24018 28044
rect 23610 28004 23616 28016
rect 24012 28004 24018 28016
rect 24070 28004 24076 28056
rect 24475 28047 24533 28053
rect 24475 28013 24487 28047
rect 24521 28044 24533 28047
rect 24748 28044 24754 28056
rect 24521 28016 24754 28044
rect 24521 28013 24533 28016
rect 24475 28007 24533 28013
rect 24748 28004 24754 28016
rect 24806 28004 24812 28056
rect 25852 28044 25858 28056
rect 25813 28016 25858 28044
rect 25852 28004 25858 28016
rect 25910 28004 25916 28056
rect 27603 28047 27661 28053
rect 27603 28013 27615 28047
rect 27649 28044 27661 28047
rect 29440 28044 29446 28056
rect 27649 28016 29446 28044
rect 27649 28013 27661 28016
rect 27603 28007 27661 28013
rect 29440 28004 29446 28016
rect 29498 28004 29504 28056
rect 29532 28004 29538 28056
rect 29590 28044 29596 28056
rect 29716 28044 29722 28056
rect 29590 28016 29635 28044
rect 29677 28016 29722 28044
rect 29590 28004 29596 28016
rect 29716 28004 29722 28016
rect 29774 28004 29780 28056
rect 29900 28044 29906 28056
rect 29861 28016 29906 28044
rect 29900 28004 29906 28016
rect 29958 28004 29964 28056
rect 29992 28004 29998 28056
rect 30050 28044 30056 28056
rect 30087 28047 30145 28053
rect 30087 28044 30099 28047
rect 30050 28016 30099 28044
rect 30050 28004 30056 28016
rect 30087 28013 30099 28016
rect 30133 28013 30145 28047
rect 30087 28007 30145 28013
rect 30176 28004 30182 28056
rect 30234 28044 30240 28056
rect 30746 28053 30774 28084
rect 30455 28047 30513 28053
rect 30455 28044 30467 28047
rect 30234 28016 30467 28044
rect 30234 28004 30240 28016
rect 30455 28013 30467 28016
rect 30501 28013 30513 28047
rect 30455 28007 30513 28013
rect 30731 28047 30789 28053
rect 30731 28013 30743 28047
rect 30777 28013 30789 28047
rect 30731 28007 30789 28013
rect 30820 28004 30826 28056
rect 30878 28044 30884 28056
rect 30878 28016 30923 28044
rect 30878 28004 30884 28016
rect 13082 27948 17342 27976
rect 11733 27945 11745 27948
rect 11687 27939 11745 27945
rect 19044 27936 19050 27988
rect 19102 27976 19108 27988
rect 19102 27948 21022 27976
rect 19102 27936 19108 27948
rect 4106 27880 7590 27908
rect 8467 27911 8525 27917
rect 4106 27868 4112 27880
rect 8467 27877 8479 27911
rect 8513 27908 8525 27911
rect 8556 27908 8562 27920
rect 8513 27880 8562 27908
rect 8513 27877 8525 27880
rect 8467 27871 8525 27877
rect 8556 27868 8562 27880
rect 8614 27868 8620 27920
rect 9292 27868 9298 27920
rect 9350 27908 9356 27920
rect 14812 27908 14818 27920
rect 9350 27880 14818 27908
rect 9350 27868 9356 27880
rect 14812 27868 14818 27880
rect 14870 27868 14876 27920
rect 15364 27868 15370 27920
rect 15422 27908 15428 27920
rect 17296 27908 17302 27920
rect 15422 27880 17302 27908
rect 15422 27868 15428 27880
rect 17296 27868 17302 27880
rect 17354 27868 17360 27920
rect 17388 27868 17394 27920
rect 17446 27908 17452 27920
rect 20884 27908 20890 27920
rect 17446 27880 20890 27908
rect 17446 27868 17452 27880
rect 20884 27868 20890 27880
rect 20942 27868 20948 27920
rect 20994 27908 21022 27948
rect 21638 27948 23414 27976
rect 21638 27908 21666 27948
rect 23276 27908 23282 27920
rect 20994 27880 21666 27908
rect 23237 27880 23282 27908
rect 23276 27868 23282 27880
rect 23334 27868 23340 27920
rect 23386 27908 23414 27948
rect 23460 27936 23466 27988
rect 23518 27976 23524 27988
rect 24104 27976 24110 27988
rect 23518 27948 24110 27976
rect 23518 27936 23524 27948
rect 24104 27936 24110 27948
rect 24162 27936 24168 27988
rect 31022 27976 31050 28084
rect 31191 28081 31203 28084
rect 31237 28081 31249 28115
rect 34040 28112 34046 28124
rect 31191 28075 31249 28081
rect 31298 28084 34046 28112
rect 31096 28004 31102 28056
rect 31154 28044 31160 28056
rect 31298 28044 31326 28084
rect 34040 28072 34046 28084
rect 34098 28072 34104 28124
rect 34411 28115 34469 28121
rect 34411 28081 34423 28115
rect 34457 28112 34469 28115
rect 34592 28112 34598 28124
rect 34457 28084 34598 28112
rect 34457 28081 34469 28084
rect 34411 28075 34469 28081
rect 34592 28072 34598 28084
rect 34650 28072 34656 28124
rect 40590 28121 40618 28152
rect 41771 28149 41783 28183
rect 41817 28180 41829 28183
rect 44988 28180 44994 28192
rect 41817 28152 44994 28180
rect 41817 28149 41829 28152
rect 41771 28143 41829 28149
rect 44988 28140 44994 28152
rect 45046 28140 45052 28192
rect 49238 28180 49266 28220
rect 49312 28208 49318 28260
rect 49370 28248 49376 28260
rect 49956 28248 49962 28260
rect 49370 28220 49962 28248
rect 49370 28208 49376 28220
rect 49956 28208 49962 28220
rect 50014 28208 50020 28260
rect 50324 28248 50330 28260
rect 50066 28220 50330 28248
rect 50066 28180 50094 28220
rect 50324 28208 50330 28220
rect 50382 28208 50388 28260
rect 50416 28208 50422 28260
rect 50474 28248 50480 28260
rect 50787 28251 50845 28257
rect 50787 28248 50799 28251
rect 50474 28220 50799 28248
rect 50474 28208 50480 28220
rect 50787 28217 50799 28220
rect 50833 28248 50845 28251
rect 52072 28248 52078 28260
rect 50833 28220 52078 28248
rect 50833 28217 50845 28220
rect 50787 28211 50845 28217
rect 52072 28208 52078 28220
rect 52130 28208 52136 28260
rect 53820 28248 53826 28260
rect 53781 28220 53826 28248
rect 53820 28208 53826 28220
rect 53878 28208 53884 28260
rect 53912 28208 53918 28260
rect 53970 28248 53976 28260
rect 59800 28248 59806 28260
rect 53970 28220 59806 28248
rect 53970 28208 53976 28220
rect 59800 28208 59806 28220
rect 59858 28208 59864 28260
rect 63940 28248 63946 28260
rect 63901 28220 63946 28248
rect 63940 28208 63946 28220
rect 63998 28208 64004 28260
rect 64216 28208 64222 28260
rect 64274 28248 64280 28260
rect 64403 28251 64461 28257
rect 64403 28248 64415 28251
rect 64274 28220 64415 28248
rect 64274 28208 64280 28220
rect 64403 28217 64415 28220
rect 64449 28217 64461 28251
rect 64403 28211 64461 28217
rect 74244 28208 74250 28260
rect 74302 28248 74308 28260
rect 75259 28251 75317 28257
rect 75259 28248 75271 28251
rect 74302 28220 75271 28248
rect 74302 28208 74308 28220
rect 75259 28217 75271 28220
rect 75305 28217 75317 28251
rect 80408 28248 80414 28260
rect 80369 28220 80414 28248
rect 75259 28211 75317 28217
rect 80408 28208 80414 28220
rect 80466 28208 80472 28260
rect 89427 28251 89485 28257
rect 89427 28217 89439 28251
rect 89473 28248 89485 28251
rect 90344 28248 90350 28260
rect 89473 28220 90350 28248
rect 89473 28217 89485 28220
rect 89427 28211 89485 28217
rect 90344 28208 90350 28220
rect 90402 28208 90408 28260
rect 49238 28152 50094 28180
rect 40575 28115 40633 28121
rect 40575 28081 40587 28115
rect 40621 28081 40633 28115
rect 40575 28075 40633 28081
rect 42139 28115 42197 28121
rect 42139 28081 42151 28115
rect 42185 28112 42197 28115
rect 42964 28112 42970 28124
rect 42185 28084 42970 28112
rect 42185 28081 42197 28084
rect 42139 28075 42197 28081
rect 31154 28016 31326 28044
rect 31154 28004 31160 28016
rect 31372 28004 31378 28056
rect 31430 28044 31436 28056
rect 33767 28047 33825 28053
rect 33767 28044 33779 28047
rect 31430 28016 33779 28044
rect 31430 28004 31436 28016
rect 33767 28013 33779 28016
rect 33813 28044 33825 28047
rect 33948 28044 33954 28056
rect 33813 28016 33954 28044
rect 33813 28013 33825 28016
rect 33767 28007 33825 28013
rect 33948 28004 33954 28016
rect 34006 28044 34012 28056
rect 34224 28044 34230 28056
rect 34006 28016 34230 28044
rect 34006 28004 34012 28016
rect 34224 28004 34230 28016
rect 34282 28044 34288 28056
rect 34503 28047 34561 28053
rect 34503 28044 34515 28047
rect 34282 28016 34515 28044
rect 34282 28004 34288 28016
rect 34503 28013 34515 28016
rect 34549 28044 34561 28047
rect 35055 28047 35113 28053
rect 35055 28044 35067 28047
rect 34549 28016 35067 28044
rect 34549 28013 34561 28016
rect 34503 28007 34561 28013
rect 35055 28013 35067 28016
rect 35101 28013 35113 28047
rect 35236 28044 35242 28056
rect 35197 28016 35242 28044
rect 35055 28007 35113 28013
rect 35236 28004 35242 28016
rect 35294 28044 35300 28056
rect 35294 28016 35926 28044
rect 35294 28004 35300 28016
rect 25134 27948 31050 27976
rect 25134 27908 25162 27948
rect 31188 27936 31194 27988
rect 31246 27976 31252 27988
rect 35788 27976 35794 27988
rect 31246 27948 35794 27976
rect 31246 27936 31252 27948
rect 35788 27936 35794 27948
rect 35846 27936 35852 27988
rect 35898 27976 35926 28016
rect 36156 28004 36162 28056
rect 36214 28044 36220 28056
rect 36527 28047 36585 28053
rect 36527 28044 36539 28047
rect 36214 28016 36539 28044
rect 36214 28004 36220 28016
rect 36527 28013 36539 28016
rect 36573 28013 36585 28047
rect 38548 28044 38554 28056
rect 36527 28007 36585 28013
rect 36634 28016 38554 28044
rect 36634 27985 36662 28016
rect 38548 28004 38554 28016
rect 38606 28004 38612 28056
rect 40664 28004 40670 28056
rect 40722 28053 40728 28056
rect 40722 28047 40771 28053
rect 40722 28013 40725 28047
rect 40759 28013 40771 28047
rect 40722 28007 40771 28013
rect 41219 28047 41277 28053
rect 41219 28013 41231 28047
rect 41265 28013 41277 28047
rect 41219 28007 41277 28013
rect 41311 28047 41369 28053
rect 41311 28013 41323 28047
rect 41357 28044 41369 28047
rect 41768 28044 41774 28056
rect 41357 28016 41774 28044
rect 41357 28013 41369 28016
rect 41311 28007 41369 28013
rect 40722 28004 40728 28007
rect 36619 27979 36677 27985
rect 36619 27976 36631 27979
rect 35898 27948 36631 27976
rect 36619 27945 36631 27948
rect 36665 27945 36677 27979
rect 36619 27939 36677 27945
rect 36708 27936 36714 27988
rect 36766 27976 36772 27988
rect 38364 27976 38370 27988
rect 36766 27948 38370 27976
rect 36766 27936 36772 27948
rect 38364 27936 38370 27948
rect 38422 27936 38428 27988
rect 38640 27936 38646 27988
rect 38698 27976 38704 27988
rect 40391 27979 40449 27985
rect 40391 27976 40403 27979
rect 38698 27948 40403 27976
rect 38698 27936 38704 27948
rect 40391 27945 40403 27948
rect 40437 27976 40449 27979
rect 41234 27976 41262 28007
rect 41768 28004 41774 28016
rect 41826 28044 41832 28056
rect 42154 28044 42182 28075
rect 42964 28072 42970 28084
rect 43022 28072 43028 28124
rect 44347 28115 44405 28121
rect 44347 28081 44359 28115
rect 44393 28112 44405 28115
rect 45816 28112 45822 28124
rect 44393 28084 45822 28112
rect 44393 28081 44405 28084
rect 44347 28075 44405 28081
rect 45816 28072 45822 28084
rect 45874 28072 45880 28124
rect 48119 28115 48177 28121
rect 48119 28081 48131 28115
rect 48165 28112 48177 28115
rect 48165 28084 48254 28112
rect 48165 28081 48177 28084
rect 48119 28075 48177 28081
rect 43056 28044 43062 28056
rect 41826 28016 42182 28044
rect 43017 28016 43062 28044
rect 41826 28004 41832 28016
rect 43056 28004 43062 28016
rect 43114 28004 43120 28056
rect 43243 28047 43301 28053
rect 43243 28013 43255 28047
rect 43289 28044 43301 28047
rect 43424 28044 43430 28056
rect 43289 28016 43430 28044
rect 43289 28013 43301 28016
rect 43243 28007 43301 28013
rect 43424 28004 43430 28016
rect 43482 28004 43488 28056
rect 43703 28047 43761 28053
rect 43703 28013 43715 28047
rect 43749 28013 43761 28047
rect 43703 28007 43761 28013
rect 42504 27976 42510 27988
rect 40437 27948 42510 27976
rect 40437 27945 40449 27948
rect 40391 27939 40449 27945
rect 42504 27936 42510 27948
rect 42562 27936 42568 27988
rect 43718 27976 43746 28007
rect 43792 28004 43798 28056
rect 43850 28044 43856 28056
rect 43850 28016 43943 28044
rect 43850 28004 43856 28016
rect 44436 28004 44442 28056
rect 44494 28044 44500 28056
rect 44531 28047 44589 28053
rect 44531 28044 44543 28047
rect 44494 28016 44543 28044
rect 44494 28004 44500 28016
rect 44531 28013 44543 28016
rect 44577 28013 44589 28047
rect 47840 28044 47846 28056
rect 44531 28007 44589 28013
rect 44638 28016 47846 28044
rect 42890 27948 43746 27976
rect 43810 27976 43838 28004
rect 44638 27976 44666 28016
rect 47840 28004 47846 28016
rect 47898 28004 47904 28056
rect 48226 28044 48254 28084
rect 48300 28072 48306 28124
rect 48358 28112 48364 28124
rect 48395 28115 48453 28121
rect 48395 28112 48407 28115
rect 48358 28084 48407 28112
rect 48358 28072 48364 28084
rect 48395 28081 48407 28084
rect 48441 28081 48453 28115
rect 50434 28112 50462 28208
rect 51520 28140 51526 28192
rect 51578 28180 51584 28192
rect 56123 28183 56181 28189
rect 56123 28180 56135 28183
rect 51578 28152 56135 28180
rect 51578 28140 51584 28152
rect 56123 28149 56135 28152
rect 56169 28180 56181 28183
rect 56215 28183 56273 28189
rect 56215 28180 56227 28183
rect 56169 28152 56227 28180
rect 56169 28149 56181 28152
rect 56123 28143 56181 28149
rect 56215 28149 56227 28152
rect 56261 28149 56273 28183
rect 56215 28143 56273 28149
rect 57500 28140 57506 28192
rect 57558 28180 57564 28192
rect 58791 28183 58849 28189
rect 58791 28180 58803 28183
rect 57558 28152 58803 28180
rect 57558 28140 57564 28152
rect 58791 28149 58803 28152
rect 58837 28149 58849 28183
rect 65872 28180 65878 28192
rect 58791 28143 58849 28149
rect 62486 28152 65878 28180
rect 52532 28112 52538 28124
rect 48395 28075 48453 28081
rect 49882 28084 50462 28112
rect 51998 28084 52538 28112
rect 49882 28053 49910 28084
rect 49867 28047 49925 28053
rect 48226 28016 49818 28044
rect 43810 27948 44666 27976
rect 46187 27979 46245 27985
rect 42890 27920 42918 27948
rect 46187 27945 46199 27979
rect 46233 27976 46245 27979
rect 46276 27976 46282 27988
rect 46233 27948 46282 27976
rect 46233 27945 46245 27948
rect 46187 27939 46245 27945
rect 46276 27936 46282 27948
rect 46334 27936 46340 27988
rect 23386 27880 25162 27908
rect 25852 27868 25858 27920
rect 25910 27908 25916 27920
rect 31280 27908 31286 27920
rect 25910 27880 31286 27908
rect 25910 27868 25916 27880
rect 31280 27868 31286 27880
rect 31338 27868 31344 27920
rect 31372 27868 31378 27920
rect 31430 27908 31436 27920
rect 38732 27908 38738 27920
rect 31430 27880 38738 27908
rect 31430 27868 31436 27880
rect 38732 27868 38738 27880
rect 38790 27868 38796 27920
rect 42872 27908 42878 27920
rect 42833 27880 42878 27908
rect 42872 27868 42878 27880
rect 42930 27868 42936 27920
rect 43240 27868 43246 27920
rect 43298 27908 43304 27920
rect 47567 27911 47625 27917
rect 47567 27908 47579 27911
rect 43298 27880 47579 27908
rect 43298 27868 43304 27880
rect 47567 27877 47579 27880
rect 47613 27908 47625 27911
rect 48208 27908 48214 27920
rect 47613 27880 48214 27908
rect 47613 27877 47625 27880
rect 47567 27871 47625 27877
rect 48208 27868 48214 27880
rect 48266 27868 48272 27920
rect 48392 27868 48398 27920
rect 48450 27908 48456 27920
rect 49499 27911 49557 27917
rect 49499 27908 49511 27911
rect 48450 27880 49511 27908
rect 48450 27868 48456 27880
rect 49499 27877 49511 27880
rect 49545 27877 49557 27911
rect 49790 27908 49818 28016
rect 49867 28013 49879 28047
rect 49913 28013 49925 28047
rect 50048 28044 50054 28056
rect 50009 28016 50054 28044
rect 49867 28007 49925 28013
rect 50048 28004 50054 28016
rect 50106 28004 50112 28056
rect 50784 28004 50790 28056
rect 50842 28044 50848 28056
rect 51998 28053 52026 28084
rect 52532 28072 52538 28084
rect 52590 28112 52596 28124
rect 52811 28115 52869 28121
rect 52811 28112 52823 28115
rect 52590 28084 52823 28112
rect 52590 28072 52596 28084
rect 52811 28081 52823 28084
rect 52857 28081 52869 28115
rect 52811 28075 52869 28081
rect 52900 28072 52906 28124
rect 52958 28112 52964 28124
rect 57592 28112 57598 28124
rect 52958 28084 57598 28112
rect 52958 28072 52964 28084
rect 57592 28072 57598 28084
rect 57650 28112 57656 28124
rect 57871 28115 57929 28121
rect 57871 28112 57883 28115
rect 57650 28084 57883 28112
rect 57650 28072 57656 28084
rect 57871 28081 57883 28084
rect 57917 28112 57929 28115
rect 57963 28115 58021 28121
rect 57963 28112 57975 28115
rect 57917 28084 57975 28112
rect 57917 28081 57929 28084
rect 57871 28075 57929 28081
rect 57963 28081 57975 28084
rect 58009 28112 58021 28115
rect 58420 28112 58426 28124
rect 58009 28084 58426 28112
rect 58009 28081 58021 28084
rect 57963 28075 58021 28081
rect 58420 28072 58426 28084
rect 58478 28072 58484 28124
rect 51983 28047 52041 28053
rect 51983 28044 51995 28047
rect 50842 28016 51995 28044
rect 50842 28004 50848 28016
rect 51983 28013 51995 28016
rect 52029 28013 52041 28047
rect 51983 28007 52041 28013
rect 52072 28004 52078 28056
rect 52130 28044 52136 28056
rect 52348 28053 52354 28056
rect 52167 28047 52225 28053
rect 52167 28044 52179 28047
rect 52130 28016 52179 28044
rect 52130 28004 52136 28016
rect 52167 28013 52179 28016
rect 52213 28013 52225 28047
rect 52167 28007 52225 28013
rect 52300 28047 52354 28053
rect 52300 28013 52312 28047
rect 52346 28013 52354 28047
rect 52300 28007 52354 28013
rect 52348 28004 52354 28007
rect 52406 28004 52412 28056
rect 53452 28004 53458 28056
rect 53510 28044 53516 28056
rect 53731 28047 53789 28053
rect 53731 28044 53743 28047
rect 53510 28016 53743 28044
rect 53510 28004 53516 28016
rect 53731 28013 53743 28016
rect 53777 28013 53789 28047
rect 53731 28007 53789 28013
rect 56123 28047 56181 28053
rect 56123 28013 56135 28047
rect 56169 28044 56181 28047
rect 56583 28047 56641 28053
rect 56583 28044 56595 28047
rect 56169 28016 56595 28044
rect 56169 28013 56181 28016
rect 56123 28007 56181 28013
rect 56583 28013 56595 28016
rect 56629 28013 56641 28047
rect 57408 28044 57414 28056
rect 57369 28016 57414 28044
rect 56583 28007 56641 28013
rect 57408 28004 57414 28016
rect 57466 28004 57472 28056
rect 57687 28047 57745 28053
rect 57687 28013 57699 28047
rect 57733 28013 57745 28047
rect 57687 28007 57745 28013
rect 50416 27976 50422 27988
rect 50377 27948 50422 27976
rect 50416 27936 50422 27948
rect 50474 27936 50480 27988
rect 52719 27979 52777 27985
rect 52719 27945 52731 27979
rect 52765 27945 52777 27979
rect 52719 27939 52777 27945
rect 53547 27979 53605 27985
rect 53547 27945 53559 27979
rect 53593 27945 53605 27979
rect 56856 27976 56862 27988
rect 56817 27948 56862 27976
rect 53547 27939 53605 27945
rect 50511 27911 50569 27917
rect 50511 27908 50523 27911
rect 49790 27880 50523 27908
rect 49499 27871 49557 27877
rect 50511 27877 50523 27880
rect 50557 27908 50569 27911
rect 51060 27908 51066 27920
rect 50557 27880 51066 27908
rect 50557 27877 50569 27880
rect 50511 27871 50569 27877
rect 51060 27868 51066 27880
rect 51118 27868 51124 27920
rect 51244 27868 51250 27920
rect 51302 27908 51308 27920
rect 52734 27908 52762 27939
rect 53360 27908 53366 27920
rect 51302 27880 52762 27908
rect 53321 27880 53366 27908
rect 51302 27868 51308 27880
rect 53360 27868 53366 27880
rect 53418 27908 53424 27920
rect 53562 27908 53590 27939
rect 56856 27936 56862 27948
rect 56914 27936 56920 27988
rect 56948 27936 56954 27988
rect 57006 27976 57012 27988
rect 57702 27976 57730 28007
rect 58328 28004 58334 28056
rect 58386 28044 58392 28056
rect 58699 28047 58757 28053
rect 58699 28044 58711 28047
rect 58386 28016 58711 28044
rect 58386 28004 58392 28016
rect 58699 28013 58711 28016
rect 58745 28013 58757 28047
rect 58699 28007 58757 28013
rect 62486 27976 62514 28152
rect 65872 28140 65878 28152
rect 65930 28140 65936 28192
rect 71024 28180 71030 28192
rect 65982 28152 71030 28180
rect 62747 28115 62805 28121
rect 62747 28081 62759 28115
rect 62793 28112 62805 28115
rect 62793 28084 64262 28112
rect 62793 28081 62805 28084
rect 62747 28075 62805 28081
rect 62652 28044 62658 28056
rect 62613 28016 62658 28044
rect 62652 28004 62658 28016
rect 62710 28004 62716 28056
rect 62928 28044 62934 28056
rect 62889 28016 62934 28044
rect 62928 28004 62934 28016
rect 62986 28004 62992 28056
rect 64234 28053 64262 28084
rect 64219 28047 64277 28053
rect 64219 28013 64231 28047
rect 64265 28013 64277 28047
rect 64219 28007 64277 28013
rect 64124 27976 64130 27988
rect 57006 27948 57730 27976
rect 57886 27948 62514 27976
rect 64085 27948 64130 27976
rect 57006 27936 57012 27948
rect 53418 27880 53590 27908
rect 56399 27911 56457 27917
rect 53418 27868 53424 27880
rect 56399 27877 56411 27911
rect 56445 27908 56457 27911
rect 57886 27908 57914 27948
rect 64124 27936 64130 27948
rect 64182 27936 64188 27988
rect 56445 27880 57914 27908
rect 56445 27877 56457 27880
rect 56399 27871 56457 27877
rect 58788 27868 58794 27920
rect 58846 27908 58852 27920
rect 65982 27908 66010 28152
rect 71024 28140 71030 28152
rect 71082 28180 71088 28192
rect 73324 28180 73330 28192
rect 71082 28152 73330 28180
rect 71082 28140 71088 28152
rect 73324 28140 73330 28152
rect 73382 28140 73388 28192
rect 79120 28140 79126 28192
rect 79178 28180 79184 28192
rect 81236 28180 81242 28192
rect 79178 28152 81242 28180
rect 79178 28140 79184 28152
rect 81236 28140 81242 28152
rect 81294 28180 81300 28192
rect 81331 28183 81389 28189
rect 81331 28180 81343 28183
rect 81294 28152 81343 28180
rect 81294 28140 81300 28152
rect 81331 28149 81343 28152
rect 81377 28149 81389 28183
rect 83079 28183 83137 28189
rect 83079 28180 83091 28183
rect 81331 28143 81389 28149
rect 81438 28152 83091 28180
rect 67988 28072 67994 28124
rect 68046 28072 68052 28124
rect 72315 28115 72373 28121
rect 72315 28081 72327 28115
rect 72361 28112 72373 28115
rect 73600 28112 73606 28124
rect 72361 28084 73606 28112
rect 72361 28081 72373 28084
rect 72315 28075 72373 28081
rect 73600 28072 73606 28084
rect 73658 28072 73664 28124
rect 74060 28072 74066 28124
rect 74118 28112 74124 28124
rect 74155 28115 74213 28121
rect 74155 28112 74167 28115
rect 74118 28084 74167 28112
rect 74118 28072 74124 28084
rect 74155 28081 74167 28084
rect 74201 28081 74213 28115
rect 74155 28075 74213 28081
rect 79764 28072 79770 28124
rect 79822 28112 79828 28124
rect 79859 28115 79917 28121
rect 79859 28112 79871 28115
rect 79822 28084 79871 28112
rect 79822 28072 79828 28084
rect 79859 28081 79871 28084
rect 79905 28112 79917 28115
rect 79951 28115 80009 28121
rect 79951 28112 79963 28115
rect 79905 28084 79963 28112
rect 79905 28081 79917 28084
rect 79859 28075 79917 28081
rect 79951 28081 79963 28084
rect 79997 28112 80009 28115
rect 81438 28112 81466 28152
rect 83079 28149 83091 28152
rect 83125 28180 83137 28183
rect 83168 28180 83174 28192
rect 83125 28152 83174 28180
rect 83125 28149 83137 28152
rect 83079 28143 83137 28149
rect 83168 28140 83174 28152
rect 83226 28140 83232 28192
rect 83370 28152 85790 28180
rect 79997 28084 81466 28112
rect 79997 28081 80009 28084
rect 79951 28075 80009 28081
rect 68006 28044 68034 28072
rect 68175 28047 68233 28053
rect 68175 28044 68187 28047
rect 68006 28016 68187 28044
rect 68175 28013 68187 28016
rect 68221 28013 68233 28047
rect 69552 28044 69558 28056
rect 69513 28016 69558 28044
rect 68175 28007 68233 28013
rect 69552 28004 69558 28016
rect 69610 28004 69616 28056
rect 69736 28044 69742 28056
rect 69697 28016 69742 28044
rect 69736 28004 69742 28016
rect 69794 28004 69800 28056
rect 72223 28047 72281 28053
rect 72223 28013 72235 28047
rect 72269 28013 72281 28047
rect 72680 28044 72686 28056
rect 72593 28016 72686 28044
rect 72223 28007 72281 28013
rect 67991 27979 68049 27985
rect 67991 27945 68003 27979
rect 68037 27976 68049 27979
rect 68632 27976 68638 27988
rect 68037 27948 68638 27976
rect 68037 27945 68049 27948
rect 67991 27939 68049 27945
rect 68632 27936 68638 27948
rect 68690 27936 68696 27988
rect 70104 27976 70110 27988
rect 70017 27948 70110 27976
rect 70104 27936 70110 27948
rect 70162 27976 70168 27988
rect 72238 27976 72266 28007
rect 72680 28004 72686 28016
rect 72738 28044 72744 28056
rect 73692 28044 73698 28056
rect 72738 28016 73698 28044
rect 72738 28004 72744 28016
rect 73692 28004 73698 28016
rect 73750 28004 73756 28056
rect 73784 28004 73790 28056
rect 73842 28044 73848 28056
rect 73879 28047 73937 28053
rect 73879 28044 73891 28047
rect 73842 28016 73891 28044
rect 73842 28004 73848 28016
rect 73879 28013 73891 28016
rect 73925 28044 73937 28047
rect 75627 28047 75685 28053
rect 75627 28044 75639 28047
rect 73925 28016 75639 28044
rect 73925 28013 73937 28016
rect 73879 28007 73937 28013
rect 75627 28013 75639 28016
rect 75673 28044 75685 28047
rect 77556 28044 77562 28056
rect 75673 28016 77562 28044
rect 75673 28013 75685 28016
rect 75627 28007 75685 28013
rect 77556 28004 77562 28016
rect 77614 28004 77620 28056
rect 80227 28047 80285 28053
rect 80227 28013 80239 28047
rect 80273 28044 80285 28047
rect 81328 28044 81334 28056
rect 80273 28016 81334 28044
rect 80273 28013 80285 28016
rect 80227 28007 80285 28013
rect 81328 28004 81334 28016
rect 81386 28004 81392 28056
rect 83370 28053 83398 28152
rect 83907 28115 83965 28121
rect 83907 28081 83919 28115
rect 83953 28112 83965 28115
rect 84548 28112 84554 28124
rect 83953 28084 84554 28112
rect 83953 28081 83965 28084
rect 83907 28075 83965 28081
rect 84548 28072 84554 28084
rect 84606 28072 84612 28124
rect 85762 28056 85790 28152
rect 90068 28140 90074 28192
rect 90126 28180 90132 28192
rect 90126 28152 91586 28180
rect 90126 28140 90132 28152
rect 87584 28072 87590 28124
rect 87642 28112 87648 28124
rect 90163 28115 90221 28121
rect 90163 28112 90175 28115
rect 87642 28084 90175 28112
rect 87642 28072 87648 28084
rect 90163 28081 90175 28084
rect 90209 28081 90221 28115
rect 90163 28075 90221 28081
rect 81699 28047 81757 28053
rect 81699 28013 81711 28047
rect 81745 28013 81757 28047
rect 81699 28007 81757 28013
rect 83355 28047 83413 28053
rect 83355 28013 83367 28047
rect 83401 28013 83413 28047
rect 83355 28007 83413 28013
rect 83447 28047 83505 28053
rect 83447 28013 83459 28047
rect 83493 28044 83505 28047
rect 84916 28044 84922 28056
rect 83493 28016 84922 28044
rect 83493 28013 83505 28016
rect 83447 28007 83505 28013
rect 73048 27976 73054 27988
rect 70162 27948 73054 27976
rect 70162 27936 70168 27948
rect 73048 27936 73054 27948
rect 73106 27936 73112 27988
rect 80132 27976 80138 27988
rect 80093 27948 80138 27976
rect 80132 27936 80138 27948
rect 80190 27936 80196 27988
rect 81236 27936 81242 27988
rect 81294 27976 81300 27988
rect 81515 27979 81573 27985
rect 81515 27976 81527 27979
rect 81294 27948 81527 27976
rect 81294 27936 81300 27948
rect 81515 27945 81527 27948
rect 81561 27945 81573 27979
rect 81515 27939 81573 27945
rect 68264 27908 68270 27920
rect 58846 27880 66010 27908
rect 68225 27880 68270 27908
rect 58846 27868 58852 27880
rect 68264 27868 68270 27880
rect 68322 27868 68328 27920
rect 79856 27868 79862 27920
rect 79914 27908 79920 27920
rect 81714 27908 81742 28007
rect 84916 28004 84922 28016
rect 84974 28004 84980 28056
rect 85008 28004 85014 28056
rect 85066 28044 85072 28056
rect 85655 28047 85713 28053
rect 85655 28044 85667 28047
rect 85066 28016 85667 28044
rect 85066 28004 85072 28016
rect 85655 28013 85667 28016
rect 85701 28013 85713 28047
rect 85655 28007 85713 28013
rect 85744 28004 85750 28056
rect 85802 28044 85808 28056
rect 85931 28047 85989 28053
rect 85931 28044 85943 28047
rect 85802 28016 85943 28044
rect 85802 28004 85808 28016
rect 85931 28013 85943 28016
rect 85977 28013 85989 28047
rect 86112 28044 86118 28056
rect 86073 28016 86118 28044
rect 85931 28007 85989 28013
rect 86112 28004 86118 28016
rect 86170 28004 86176 28056
rect 89332 28044 89338 28056
rect 89293 28016 89338 28044
rect 89332 28004 89338 28016
rect 89390 28044 89396 28056
rect 89608 28044 89614 28056
rect 89390 28016 89614 28044
rect 89390 28004 89396 28016
rect 89608 28004 89614 28016
rect 89666 28004 89672 28056
rect 90178 28044 90206 28075
rect 90344 28072 90350 28124
rect 90402 28112 90408 28124
rect 91558 28121 91586 28152
rect 91543 28115 91601 28121
rect 90402 28084 91494 28112
rect 90402 28072 90408 28084
rect 91080 28044 91086 28056
rect 90178 28016 90942 28044
rect 91041 28016 91086 28044
rect 82067 27979 82125 27985
rect 82067 27945 82079 27979
rect 82113 27976 82125 27979
rect 83260 27976 83266 27988
rect 82113 27948 83266 27976
rect 82113 27945 82125 27948
rect 82067 27939 82125 27945
rect 83260 27936 83266 27948
rect 83318 27936 83324 27988
rect 85103 27979 85161 27985
rect 85103 27945 85115 27979
rect 85149 27976 85161 27979
rect 86572 27976 86578 27988
rect 85149 27948 86578 27976
rect 85149 27945 85161 27948
rect 85103 27939 85161 27945
rect 86572 27936 86578 27948
rect 86630 27936 86636 27988
rect 89240 27936 89246 27988
rect 89298 27976 89304 27988
rect 90439 27979 90497 27985
rect 90439 27976 90451 27979
rect 89298 27948 90451 27976
rect 89298 27936 89304 27948
rect 90439 27945 90451 27948
rect 90485 27945 90497 27979
rect 90914 27976 90942 28016
rect 91080 28004 91086 28016
rect 91138 28004 91144 28056
rect 91466 28053 91494 28084
rect 91543 28081 91555 28115
rect 91589 28081 91601 28115
rect 91543 28075 91601 28081
rect 91175 28047 91233 28053
rect 91175 28013 91187 28047
rect 91221 28013 91233 28047
rect 91175 28007 91233 28013
rect 91451 28047 91509 28053
rect 91451 28013 91463 28047
rect 91497 28013 91509 28047
rect 91451 28007 91509 28013
rect 91190 27976 91218 28007
rect 90914 27948 91218 27976
rect 90439 27939 90497 27945
rect 79914 27880 81742 27908
rect 79914 27868 79920 27880
rect 538 27818 93642 27840
rect 538 27766 6344 27818
rect 6396 27766 6408 27818
rect 6460 27766 6472 27818
rect 6524 27766 6536 27818
rect 6588 27766 11672 27818
rect 11724 27766 11736 27818
rect 11788 27766 11800 27818
rect 11852 27766 11864 27818
rect 11916 27766 17000 27818
rect 17052 27766 17064 27818
rect 17116 27766 17128 27818
rect 17180 27766 17192 27818
rect 17244 27766 22328 27818
rect 22380 27766 22392 27818
rect 22444 27766 22456 27818
rect 22508 27766 22520 27818
rect 22572 27766 27656 27818
rect 27708 27766 27720 27818
rect 27772 27766 27784 27818
rect 27836 27766 27848 27818
rect 27900 27766 32984 27818
rect 33036 27766 33048 27818
rect 33100 27766 33112 27818
rect 33164 27766 33176 27818
rect 33228 27766 38312 27818
rect 38364 27766 38376 27818
rect 38428 27766 38440 27818
rect 38492 27766 38504 27818
rect 38556 27766 43640 27818
rect 43692 27766 43704 27818
rect 43756 27766 43768 27818
rect 43820 27766 43832 27818
rect 43884 27766 48968 27818
rect 49020 27766 49032 27818
rect 49084 27766 49096 27818
rect 49148 27766 49160 27818
rect 49212 27766 54296 27818
rect 54348 27766 54360 27818
rect 54412 27766 54424 27818
rect 54476 27766 54488 27818
rect 54540 27766 59624 27818
rect 59676 27766 59688 27818
rect 59740 27766 59752 27818
rect 59804 27766 59816 27818
rect 59868 27766 64952 27818
rect 65004 27766 65016 27818
rect 65068 27766 65080 27818
rect 65132 27766 65144 27818
rect 65196 27766 70280 27818
rect 70332 27766 70344 27818
rect 70396 27766 70408 27818
rect 70460 27766 70472 27818
rect 70524 27766 75608 27818
rect 75660 27766 75672 27818
rect 75724 27766 75736 27818
rect 75788 27766 75800 27818
rect 75852 27766 80936 27818
rect 80988 27766 81000 27818
rect 81052 27766 81064 27818
rect 81116 27766 81128 27818
rect 81180 27766 86264 27818
rect 86316 27766 86328 27818
rect 86380 27766 86392 27818
rect 86444 27766 86456 27818
rect 86508 27766 91592 27818
rect 91644 27766 91656 27818
rect 91708 27766 91720 27818
rect 91772 27766 91784 27818
rect 91836 27766 93642 27818
rect 538 27744 93642 27766
rect 1932 27664 1938 27716
rect 1990 27704 1996 27716
rect 2303 27707 2361 27713
rect 2303 27704 2315 27707
rect 1990 27676 2315 27704
rect 1990 27664 1996 27676
rect 2303 27673 2315 27676
rect 2349 27673 2361 27707
rect 7728 27704 7734 27716
rect 7689 27676 7734 27704
rect 2303 27667 2361 27673
rect 7728 27664 7734 27676
rect 7786 27664 7792 27716
rect 8096 27704 8102 27716
rect 8057 27676 8102 27704
rect 8096 27664 8102 27676
rect 8154 27664 8160 27716
rect 8283 27707 8341 27713
rect 8283 27673 8295 27707
rect 8329 27704 8341 27707
rect 8467 27707 8525 27713
rect 8467 27704 8479 27707
rect 8329 27676 8479 27704
rect 8329 27673 8341 27676
rect 8283 27667 8341 27673
rect 8467 27673 8479 27676
rect 8513 27704 8525 27707
rect 15364 27704 15370 27716
rect 8513 27676 15370 27704
rect 8513 27673 8525 27676
rect 8467 27667 8525 27673
rect 8298 27636 8326 27667
rect 15364 27664 15370 27676
rect 15422 27664 15428 27716
rect 15459 27707 15517 27713
rect 15459 27673 15471 27707
rect 15505 27704 15517 27707
rect 15824 27704 15830 27716
rect 15505 27676 15830 27704
rect 15505 27673 15517 27676
rect 15459 27667 15517 27673
rect 7286 27608 8326 27636
rect 920 27568 926 27580
rect 881 27540 926 27568
rect 920 27528 926 27540
rect 978 27528 984 27580
rect 7286 27577 7314 27608
rect 8556 27596 8562 27648
rect 8614 27636 8620 27648
rect 15474 27636 15502 27667
rect 15824 27664 15830 27676
rect 15882 27704 15888 27716
rect 16652 27704 16658 27716
rect 15882 27676 16658 27704
rect 15882 27664 15888 27676
rect 16652 27664 16658 27676
rect 16710 27664 16716 27716
rect 17664 27664 17670 27716
rect 17722 27704 17728 27716
rect 17851 27707 17909 27713
rect 17851 27704 17863 27707
rect 17722 27676 17863 27704
rect 17722 27664 17728 27676
rect 17851 27673 17863 27676
rect 17897 27673 17909 27707
rect 17851 27667 17909 27673
rect 22635 27707 22693 27713
rect 22635 27673 22647 27707
rect 22681 27704 22693 27707
rect 23092 27704 23098 27716
rect 22681 27676 23098 27704
rect 22681 27673 22693 27676
rect 22635 27667 22693 27673
rect 23092 27664 23098 27676
rect 23150 27664 23156 27716
rect 23463 27707 23521 27713
rect 23463 27673 23475 27707
rect 23509 27704 23521 27707
rect 23644 27704 23650 27716
rect 23509 27676 23650 27704
rect 23509 27673 23521 27676
rect 23463 27667 23521 27673
rect 23644 27664 23650 27676
rect 23702 27664 23708 27716
rect 24564 27704 24570 27716
rect 24030 27676 24570 27704
rect 8614 27608 15502 27636
rect 8614 27596 8620 27608
rect 15732 27596 15738 27648
rect 15790 27636 15796 27648
rect 15790 27608 16514 27636
rect 15790 27596 15796 27608
rect 16486 27580 16514 27608
rect 17572 27596 17578 27648
rect 17630 27636 17636 27648
rect 19599 27639 19657 27645
rect 19599 27636 19611 27639
rect 17630 27608 19611 27636
rect 17630 27596 17636 27608
rect 6719 27571 6777 27577
rect 6719 27537 6731 27571
rect 6765 27568 6777 27571
rect 7271 27571 7329 27577
rect 7271 27568 7283 27571
rect 6765 27540 7283 27568
rect 6765 27537 6777 27540
rect 6719 27531 6777 27537
rect 7271 27537 7283 27540
rect 7317 27537 7329 27571
rect 7271 27531 7329 27537
rect 7455 27571 7513 27577
rect 7455 27537 7467 27571
rect 7501 27568 7513 27571
rect 8096 27568 8102 27580
rect 7501 27540 8102 27568
rect 7501 27537 7513 27540
rect 7455 27531 7513 27537
rect 8096 27528 8102 27540
rect 8154 27528 8160 27580
rect 11503 27571 11561 27577
rect 11503 27537 11515 27571
rect 11549 27537 11561 27571
rect 11503 27531 11561 27537
rect 1199 27503 1257 27509
rect 1199 27469 1211 27503
rect 1245 27500 1257 27503
rect 6627 27503 6685 27509
rect 1245 27472 2806 27500
rect 1245 27469 1257 27472
rect 1199 27463 1257 27469
rect 2778 27441 2806 27472
rect 6627 27469 6639 27503
rect 6673 27469 6685 27503
rect 6627 27463 6685 27469
rect 2763 27435 2821 27441
rect 2763 27401 2775 27435
rect 2809 27432 2821 27435
rect 4784 27432 4790 27444
rect 2809 27404 4790 27432
rect 2809 27401 2821 27404
rect 2763 27395 2821 27401
rect 4784 27392 4790 27404
rect 4842 27392 4848 27444
rect 6443 27435 6501 27441
rect 6443 27401 6455 27435
rect 6489 27432 6501 27435
rect 6642 27432 6670 27463
rect 10304 27460 10310 27512
rect 10362 27500 10368 27512
rect 11043 27503 11101 27509
rect 11043 27500 11055 27503
rect 10362 27472 11055 27500
rect 10362 27460 10368 27472
rect 11043 27469 11055 27472
rect 11089 27469 11101 27503
rect 11518 27500 11546 27531
rect 11868 27528 11874 27580
rect 11926 27568 11932 27580
rect 12055 27571 12113 27577
rect 11926 27540 11971 27568
rect 11926 27528 11932 27540
rect 12055 27537 12067 27571
rect 12101 27568 12113 27571
rect 12236 27568 12242 27580
rect 12101 27540 12242 27568
rect 12101 27537 12113 27540
rect 12055 27531 12113 27537
rect 12236 27528 12242 27540
rect 12294 27528 12300 27580
rect 12604 27528 12610 27580
rect 12662 27568 12668 27580
rect 12699 27571 12757 27577
rect 12699 27568 12711 27571
rect 12662 27540 12711 27568
rect 12662 27528 12668 27540
rect 12699 27537 12711 27540
rect 12745 27568 12757 27571
rect 12883 27571 12941 27577
rect 12883 27568 12895 27571
rect 12745 27540 12895 27568
rect 12745 27537 12757 27540
rect 12699 27531 12757 27537
rect 12883 27537 12895 27540
rect 12929 27537 12941 27571
rect 15640 27568 15646 27580
rect 15601 27540 15646 27568
rect 12883 27531 12941 27537
rect 15640 27528 15646 27540
rect 15698 27528 15704 27580
rect 16011 27571 16069 27577
rect 16011 27537 16023 27571
rect 16057 27537 16069 27571
rect 16011 27531 16069 27537
rect 11518 27472 12282 27500
rect 11043 27463 11101 27469
rect 9292 27432 9298 27444
rect 6489 27404 9298 27432
rect 6489 27401 6501 27404
rect 6443 27395 6501 27401
rect 2944 27364 2950 27376
rect 2905 27336 2950 27364
rect 2944 27324 2950 27336
rect 3002 27324 3008 27376
rect 4232 27324 4238 27376
rect 4290 27364 4296 27376
rect 6458 27364 6486 27395
rect 9292 27392 9298 27404
rect 9350 27392 9356 27444
rect 12254 27441 12282 27472
rect 12239 27435 12297 27441
rect 12239 27401 12251 27435
rect 12285 27432 12297 27435
rect 12420 27432 12426 27444
rect 12285 27404 12426 27432
rect 12285 27401 12297 27404
rect 12239 27395 12297 27401
rect 12420 27392 12426 27404
rect 12478 27432 12484 27444
rect 13067 27435 13125 27441
rect 13067 27432 13079 27435
rect 12478 27404 13079 27432
rect 12478 27392 12484 27404
rect 13067 27401 13079 27404
rect 13113 27432 13125 27435
rect 13156 27432 13162 27444
rect 13113 27404 13162 27432
rect 13113 27401 13125 27404
rect 13067 27395 13125 27401
rect 13156 27392 13162 27404
rect 13214 27432 13220 27444
rect 15180 27432 15186 27444
rect 13214 27404 15186 27432
rect 13214 27392 13220 27404
rect 15180 27392 15186 27404
rect 15238 27392 15244 27444
rect 16026 27432 16054 27531
rect 16100 27528 16106 27580
rect 16158 27568 16164 27580
rect 16468 27568 16474 27580
rect 16158 27540 16203 27568
rect 16381 27540 16474 27568
rect 16158 27528 16164 27540
rect 16468 27528 16474 27540
rect 16526 27528 16532 27580
rect 16560 27528 16566 27580
rect 16618 27568 16624 27580
rect 18219 27571 18277 27577
rect 18219 27568 18231 27571
rect 16618 27540 18231 27568
rect 16618 27528 16624 27540
rect 18219 27537 18231 27540
rect 18265 27568 18277 27571
rect 18584 27568 18590 27580
rect 18265 27540 18590 27568
rect 18265 27537 18277 27540
rect 18219 27531 18277 27537
rect 18584 27528 18590 27540
rect 18642 27528 18648 27580
rect 18768 27528 18774 27580
rect 18826 27568 18832 27580
rect 18970 27577 18998 27608
rect 19599 27605 19611 27608
rect 19645 27636 19657 27639
rect 23920 27636 23926 27648
rect 19645 27608 23926 27636
rect 19645 27605 19657 27608
rect 19599 27599 19657 27605
rect 23920 27596 23926 27608
rect 23978 27596 23984 27648
rect 18955 27571 19013 27577
rect 18826 27540 18871 27568
rect 18826 27528 18832 27540
rect 18955 27537 18967 27571
rect 19001 27537 19013 27571
rect 22540 27568 22546 27580
rect 22501 27540 22546 27568
rect 18955 27531 19013 27537
rect 22540 27528 22546 27540
rect 22598 27528 22604 27580
rect 22632 27528 22638 27580
rect 22690 27568 22696 27580
rect 23739 27571 23797 27577
rect 23739 27568 23751 27571
rect 22690 27540 23751 27568
rect 22690 27528 22696 27540
rect 23739 27537 23751 27540
rect 23785 27568 23797 27571
rect 24030 27568 24058 27676
rect 24564 27664 24570 27676
rect 24622 27664 24628 27716
rect 24748 27704 24754 27716
rect 24709 27676 24754 27704
rect 24748 27664 24754 27676
rect 24806 27664 24812 27716
rect 25119 27707 25177 27713
rect 25119 27673 25131 27707
rect 25165 27704 25177 27707
rect 25165 27676 28014 27704
rect 25165 27673 25177 27676
rect 25119 27667 25177 27673
rect 25134 27636 25162 27667
rect 24306 27608 25162 27636
rect 23785 27540 24058 27568
rect 23785 27537 23797 27540
rect 23739 27531 23797 27537
rect 24104 27528 24110 27580
rect 24162 27568 24168 27580
rect 24306 27577 24334 27608
rect 25208 27596 25214 27648
rect 25266 27636 25272 27648
rect 27140 27636 27146 27648
rect 25266 27608 27146 27636
rect 25266 27596 25272 27608
rect 27140 27596 27146 27608
rect 27198 27596 27204 27648
rect 27986 27636 28014 27676
rect 29808 27664 29814 27716
rect 29866 27704 29872 27716
rect 30547 27707 30605 27713
rect 30547 27704 30559 27707
rect 29866 27676 30559 27704
rect 29866 27664 29872 27676
rect 30547 27673 30559 27676
rect 30593 27673 30605 27707
rect 30547 27667 30605 27673
rect 30636 27664 30642 27716
rect 30694 27704 30700 27716
rect 38640 27704 38646 27716
rect 30694 27676 38646 27704
rect 30694 27664 30700 27676
rect 38640 27664 38646 27676
rect 38698 27664 38704 27716
rect 38824 27664 38830 27716
rect 38882 27704 38888 27716
rect 39287 27707 39345 27713
rect 39287 27704 39299 27707
rect 38882 27676 39299 27704
rect 38882 27664 38888 27676
rect 39287 27673 39299 27676
rect 39333 27673 39345 27707
rect 42504 27704 42510 27716
rect 42465 27676 42510 27704
rect 39287 27667 39345 27673
rect 42504 27664 42510 27676
rect 42562 27704 42568 27716
rect 42780 27704 42786 27716
rect 42562 27676 42786 27704
rect 42562 27664 42568 27676
rect 42780 27664 42786 27676
rect 42838 27664 42844 27716
rect 43516 27664 43522 27716
rect 43574 27704 43580 27716
rect 44344 27704 44350 27716
rect 43574 27676 44350 27704
rect 43574 27664 43580 27676
rect 44344 27664 44350 27676
rect 44402 27664 44408 27716
rect 47383 27707 47441 27713
rect 47383 27673 47395 27707
rect 47429 27704 47441 27707
rect 48208 27704 48214 27716
rect 47429 27676 48214 27704
rect 47429 27673 47441 27676
rect 47383 27667 47441 27673
rect 48208 27664 48214 27676
rect 48266 27664 48272 27716
rect 48318 27676 52118 27704
rect 30360 27636 30366 27648
rect 27986 27608 30366 27636
rect 30360 27596 30366 27608
rect 30418 27596 30424 27648
rect 31556 27596 31562 27648
rect 31614 27636 31620 27648
rect 32019 27639 32077 27645
rect 32019 27636 32031 27639
rect 31614 27608 32031 27636
rect 31614 27596 31620 27608
rect 32019 27605 32031 27608
rect 32065 27605 32077 27639
rect 32019 27599 32077 27605
rect 33764 27596 33770 27648
rect 33822 27636 33828 27648
rect 36984 27636 36990 27648
rect 33822 27608 36990 27636
rect 33822 27596 33828 27608
rect 36984 27596 36990 27608
rect 37042 27596 37048 27648
rect 37094 27608 38042 27636
rect 24199 27571 24257 27577
rect 24199 27568 24211 27571
rect 24162 27540 24211 27568
rect 24162 27528 24168 27540
rect 24199 27537 24211 27540
rect 24245 27537 24257 27571
rect 24199 27531 24257 27537
rect 24291 27571 24349 27577
rect 24291 27537 24303 27571
rect 24337 27537 24349 27571
rect 27327 27571 27385 27577
rect 27327 27568 27339 27571
rect 24291 27531 24349 27537
rect 24674 27540 27339 27568
rect 17664 27460 17670 27512
rect 17722 27500 17728 27512
rect 18035 27503 18093 27509
rect 18035 27500 18047 27503
rect 17722 27472 18047 27500
rect 17722 27460 17728 27472
rect 18035 27469 18047 27472
rect 18081 27469 18093 27503
rect 18035 27463 18093 27469
rect 20884 27460 20890 27512
rect 20942 27500 20948 27512
rect 23368 27500 23374 27512
rect 20942 27472 23374 27500
rect 20942 27460 20948 27472
rect 23368 27460 23374 27472
rect 23426 27460 23432 27512
rect 23644 27500 23650 27512
rect 23605 27472 23650 27500
rect 23644 27460 23650 27472
rect 23702 27500 23708 27512
rect 23828 27500 23834 27512
rect 23702 27472 23834 27500
rect 23702 27460 23708 27472
rect 23828 27460 23834 27472
rect 23886 27460 23892 27512
rect 17299 27435 17357 27441
rect 17299 27432 17311 27435
rect 16026 27404 17311 27432
rect 17299 27401 17311 27404
rect 17345 27432 17357 27435
rect 19136 27432 19142 27444
rect 17345 27404 19142 27432
rect 17345 27401 17357 27404
rect 17299 27395 17357 27401
rect 19136 27392 19142 27404
rect 19194 27392 19200 27444
rect 19231 27435 19289 27441
rect 19231 27401 19243 27435
rect 19277 27432 19289 27435
rect 24674 27432 24702 27540
rect 27327 27537 27339 27540
rect 27373 27537 27385 27571
rect 27327 27531 27385 27537
rect 27416 27528 27422 27580
rect 27474 27568 27480 27580
rect 28796 27568 28802 27580
rect 27474 27540 28802 27568
rect 27474 27528 27480 27540
rect 28796 27528 28802 27540
rect 28854 27568 28860 27580
rect 28891 27571 28949 27577
rect 28891 27568 28903 27571
rect 28854 27540 28903 27568
rect 28854 27528 28860 27540
rect 28891 27537 28903 27540
rect 28937 27568 28949 27571
rect 29716 27568 29722 27580
rect 28937 27540 29722 27568
rect 28937 27537 28949 27540
rect 28891 27531 28949 27537
rect 29716 27528 29722 27540
rect 29774 27528 29780 27580
rect 30455 27571 30513 27577
rect 30455 27537 30467 27571
rect 30501 27568 30513 27571
rect 31832 27568 31838 27580
rect 30501 27540 31838 27568
rect 30501 27537 30513 27540
rect 30455 27531 30513 27537
rect 31832 27528 31838 27540
rect 31890 27528 31896 27580
rect 32663 27571 32721 27577
rect 32663 27537 32675 27571
rect 32709 27537 32721 27571
rect 32663 27531 32721 27537
rect 33031 27571 33089 27577
rect 33031 27537 33043 27571
rect 33077 27568 33089 27571
rect 33120 27568 33126 27580
rect 33077 27540 33126 27568
rect 33077 27537 33089 27540
rect 33031 27531 33089 27537
rect 24748 27460 24754 27512
rect 24806 27500 24812 27512
rect 25211 27503 25269 27509
rect 25211 27500 25223 27503
rect 24806 27472 25223 27500
rect 24806 27460 24812 27472
rect 25211 27469 25223 27472
rect 25257 27469 25269 27503
rect 27048 27500 27054 27512
rect 27009 27472 27054 27500
rect 25211 27463 25269 27469
rect 27048 27460 27054 27472
rect 27106 27460 27112 27512
rect 27232 27460 27238 27512
rect 27290 27500 27296 27512
rect 31004 27500 31010 27512
rect 27290 27472 31010 27500
rect 27290 27460 27296 27472
rect 31004 27460 31010 27472
rect 31062 27460 31068 27512
rect 31280 27460 31286 27512
rect 31338 27500 31344 27512
rect 31927 27503 31985 27509
rect 31927 27500 31939 27503
rect 31338 27472 31939 27500
rect 31338 27460 31344 27472
rect 31927 27469 31939 27472
rect 31973 27500 31985 27503
rect 32678 27500 32706 27531
rect 33120 27528 33126 27540
rect 33178 27528 33184 27580
rect 33215 27571 33273 27577
rect 33215 27537 33227 27571
rect 33261 27568 33273 27571
rect 35236 27568 35242 27580
rect 33261 27540 35242 27568
rect 33261 27537 33273 27540
rect 33215 27531 33273 27537
rect 35236 27528 35242 27540
rect 35294 27528 35300 27580
rect 35975 27571 36033 27577
rect 35975 27537 35987 27571
rect 36021 27568 36033 27571
rect 36156 27568 36162 27580
rect 36021 27540 36162 27568
rect 36021 27537 36033 27540
rect 35975 27531 36033 27537
rect 36156 27528 36162 27540
rect 36214 27528 36220 27580
rect 31973 27472 32706 27500
rect 32755 27503 32813 27509
rect 31973 27469 31985 27472
rect 31927 27463 31985 27469
rect 32755 27469 32767 27503
rect 32801 27500 32813 27503
rect 33399 27503 33457 27509
rect 33399 27500 33411 27503
rect 32801 27472 33411 27500
rect 32801 27469 32813 27472
rect 32755 27463 32813 27469
rect 33399 27469 33411 27472
rect 33445 27500 33457 27503
rect 37094 27500 37122 27608
rect 38014 27568 38042 27608
rect 39744 27596 39750 27648
rect 39802 27636 39808 27648
rect 44991 27639 45049 27645
rect 44991 27636 45003 27639
rect 39802 27608 45003 27636
rect 39802 27596 39808 27608
rect 44991 27605 45003 27608
rect 45037 27605 45049 27639
rect 44991 27599 45049 27605
rect 46276 27596 46282 27648
rect 46334 27636 46340 27648
rect 48318 27636 48346 27676
rect 48484 27636 48490 27648
rect 46334 27608 48346 27636
rect 48445 27608 48490 27636
rect 46334 27596 46340 27608
rect 48484 27596 48490 27608
rect 48542 27596 48548 27648
rect 50140 27596 50146 27648
rect 50198 27636 50204 27648
rect 52090 27636 52118 27676
rect 52164 27664 52170 27716
rect 52222 27704 52228 27716
rect 54283 27707 54341 27713
rect 54283 27704 54295 27707
rect 52222 27676 54295 27704
rect 52222 27664 52228 27676
rect 54283 27673 54295 27676
rect 54329 27704 54341 27707
rect 56948 27704 56954 27716
rect 54329 27676 56954 27704
rect 54329 27673 54341 27676
rect 54283 27667 54341 27673
rect 56948 27664 56954 27676
rect 57006 27664 57012 27716
rect 57319 27707 57377 27713
rect 57319 27673 57331 27707
rect 57365 27704 57377 27707
rect 57408 27704 57414 27716
rect 57365 27676 57414 27704
rect 57365 27673 57377 27676
rect 57319 27667 57377 27673
rect 57408 27664 57414 27676
rect 57466 27664 57472 27716
rect 67896 27704 67902 27716
rect 67857 27676 67902 27704
rect 67896 27664 67902 27676
rect 67954 27664 67960 27716
rect 69736 27664 69742 27716
rect 69794 27704 69800 27716
rect 71303 27707 71361 27713
rect 71303 27704 71315 27707
rect 69794 27676 71315 27704
rect 69794 27664 69800 27676
rect 71303 27673 71315 27676
rect 71349 27673 71361 27707
rect 71303 27667 71361 27673
rect 76176 27664 76182 27716
rect 76234 27704 76240 27716
rect 78939 27707 78997 27713
rect 78939 27704 78951 27707
rect 76234 27676 78951 27704
rect 76234 27664 76240 27676
rect 78939 27673 78951 27676
rect 78985 27673 78997 27707
rect 78939 27667 78997 27673
rect 53728 27636 53734 27648
rect 50198 27608 51566 27636
rect 52090 27608 53734 27636
rect 50198 27596 50204 27608
rect 38824 27568 38830 27580
rect 38014 27540 38830 27568
rect 38824 27528 38830 27540
rect 38882 27528 38888 27580
rect 42780 27568 42786 27580
rect 42741 27540 42786 27568
rect 42780 27528 42786 27540
rect 42838 27528 42844 27580
rect 42964 27568 42970 27580
rect 42925 27540 42970 27568
rect 42964 27528 42970 27540
rect 43022 27528 43028 27580
rect 43056 27528 43062 27580
rect 43114 27568 43120 27580
rect 43427 27571 43485 27577
rect 43427 27568 43439 27571
rect 43114 27540 43439 27568
rect 43114 27528 43120 27540
rect 43427 27537 43439 27540
rect 43473 27537 43485 27571
rect 43427 27531 43485 27537
rect 43516 27528 43522 27580
rect 43574 27568 43580 27580
rect 43574 27540 43619 27568
rect 43574 27528 43580 27540
rect 43700 27528 43706 27580
rect 43758 27568 43764 27580
rect 44531 27571 44589 27577
rect 44531 27568 44543 27571
rect 43758 27540 44543 27568
rect 43758 27528 43764 27540
rect 44531 27537 44543 27540
rect 44577 27568 44589 27571
rect 45540 27568 45546 27580
rect 44577 27540 45546 27568
rect 44577 27537 44589 27540
rect 44531 27531 44589 27537
rect 45540 27528 45546 27540
rect 45598 27528 45604 27580
rect 47291 27571 47349 27577
rect 47291 27537 47303 27571
rect 47337 27568 47349 27571
rect 47748 27568 47754 27580
rect 47337 27540 47754 27568
rect 47337 27537 47349 27540
rect 47291 27531 47349 27537
rect 47748 27528 47754 27540
rect 47806 27528 47812 27580
rect 48392 27568 48398 27580
rect 48353 27540 48398 27568
rect 48392 27528 48398 27540
rect 48450 27528 48456 27580
rect 49772 27528 49778 27580
rect 49830 27568 49836 27580
rect 49959 27571 50017 27577
rect 49959 27568 49971 27571
rect 49830 27540 49971 27568
rect 49830 27528 49836 27540
rect 49959 27537 49971 27540
rect 50005 27537 50017 27571
rect 50232 27568 50238 27580
rect 50193 27540 50238 27568
rect 49959 27531 50017 27537
rect 50232 27528 50238 27540
rect 50290 27528 50296 27580
rect 51244 27568 51250 27580
rect 50342 27540 51250 27568
rect 33445 27472 37122 27500
rect 37907 27503 37965 27509
rect 33445 27469 33457 27472
rect 33399 27463 33457 27469
rect 37907 27469 37919 27503
rect 37953 27469 37965 27503
rect 37907 27463 37965 27469
rect 38183 27503 38241 27509
rect 38183 27469 38195 27503
rect 38229 27500 38241 27503
rect 38229 27472 39790 27500
rect 38229 27469 38241 27472
rect 38183 27463 38241 27469
rect 19277 27404 24702 27432
rect 19277 27401 19289 27404
rect 19231 27395 19289 27401
rect 24840 27392 24846 27444
rect 24898 27432 24904 27444
rect 26956 27432 26962 27444
rect 24898 27404 26962 27432
rect 24898 27392 24904 27404
rect 26956 27392 26962 27404
rect 27014 27392 27020 27444
rect 28612 27432 28618 27444
rect 28525 27404 28618 27432
rect 28612 27392 28618 27404
rect 28670 27432 28676 27444
rect 31372 27432 31378 27444
rect 28670 27404 31378 27432
rect 28670 27392 28676 27404
rect 31372 27392 31378 27404
rect 31430 27392 31436 27444
rect 35236 27432 35242 27444
rect 31574 27404 35242 27432
rect 4290 27336 6486 27364
rect 4290 27324 4296 27336
rect 7544 27324 7550 27376
rect 7602 27364 7608 27376
rect 10580 27364 10586 27376
rect 7602 27336 10586 27364
rect 7602 27324 7608 27336
rect 10580 27324 10586 27336
rect 10638 27324 10644 27376
rect 10859 27367 10917 27373
rect 10859 27333 10871 27367
rect 10905 27364 10917 27367
rect 11868 27364 11874 27376
rect 10905 27336 11874 27364
rect 10905 27333 10917 27336
rect 10859 27327 10917 27333
rect 11868 27324 11874 27336
rect 11926 27364 11932 27376
rect 12144 27364 12150 27376
rect 11926 27336 12150 27364
rect 11926 27324 11932 27336
rect 12144 27324 12150 27336
rect 12202 27324 12208 27376
rect 15272 27324 15278 27376
rect 15330 27364 15336 27376
rect 15367 27367 15425 27373
rect 15367 27364 15379 27367
rect 15330 27336 15379 27364
rect 15330 27324 15336 27336
rect 15367 27333 15379 27336
rect 15413 27364 15425 27367
rect 16008 27364 16014 27376
rect 15413 27336 16014 27364
rect 15413 27333 15425 27336
rect 15367 27327 15425 27333
rect 16008 27324 16014 27336
rect 16066 27324 16072 27376
rect 17020 27364 17026 27376
rect 16981 27336 17026 27364
rect 17020 27324 17026 27336
rect 17078 27324 17084 27376
rect 17112 27324 17118 27376
rect 17170 27364 17176 27376
rect 22908 27364 22914 27376
rect 17170 27336 22914 27364
rect 17170 27324 17176 27336
rect 22908 27324 22914 27336
rect 22966 27324 22972 27376
rect 23368 27324 23374 27376
rect 23426 27364 23432 27376
rect 31574 27364 31602 27404
rect 35236 27392 35242 27404
rect 35294 27392 35300 27444
rect 35788 27432 35794 27444
rect 35749 27404 35794 27432
rect 35788 27392 35794 27404
rect 35846 27392 35852 27444
rect 37723 27435 37781 27441
rect 37723 27432 37735 27435
rect 35990 27404 37735 27432
rect 31740 27364 31746 27376
rect 23426 27336 31602 27364
rect 31653 27336 31746 27364
rect 23426 27324 23432 27336
rect 31740 27324 31746 27336
rect 31798 27364 31804 27376
rect 33120 27364 33126 27376
rect 31798 27336 33126 27364
rect 31798 27324 31804 27336
rect 33120 27324 33126 27336
rect 33178 27324 33184 27376
rect 34408 27324 34414 27376
rect 34466 27364 34472 27376
rect 35990 27364 36018 27404
rect 37723 27401 37735 27404
rect 37769 27432 37781 27435
rect 37922 27432 37950 27463
rect 39762 27441 39790 27472
rect 42228 27460 42234 27512
rect 42286 27500 42292 27512
rect 43074 27500 43102 27528
rect 42286 27472 43102 27500
rect 44071 27503 44129 27509
rect 42286 27460 42292 27472
rect 44071 27469 44083 27503
rect 44117 27500 44129 27503
rect 45138 27503 45196 27509
rect 45138 27500 45150 27503
rect 44117 27472 45150 27500
rect 44117 27469 44129 27472
rect 44071 27463 44129 27469
rect 45138 27469 45150 27472
rect 45184 27469 45196 27503
rect 45356 27500 45362 27512
rect 45317 27472 45362 27500
rect 45138 27463 45196 27469
rect 45356 27460 45362 27472
rect 45414 27460 45420 27512
rect 50342 27500 50370 27540
rect 51244 27528 51250 27540
rect 51302 27528 51308 27580
rect 51538 27577 51566 27608
rect 53728 27596 53734 27608
rect 53786 27596 53792 27648
rect 53820 27596 53826 27648
rect 53878 27636 53884 27648
rect 58607 27639 58665 27645
rect 58607 27636 58619 27639
rect 53878 27608 54234 27636
rect 53878 27596 53884 27608
rect 51523 27571 51581 27577
rect 51523 27537 51535 27571
rect 51569 27537 51581 27571
rect 51523 27531 51581 27537
rect 51612 27528 51618 27580
rect 51670 27568 51676 27580
rect 52075 27571 52133 27577
rect 52075 27568 52087 27571
rect 51670 27540 52087 27568
rect 51670 27528 51676 27540
rect 52075 27537 52087 27540
rect 52121 27568 52133 27571
rect 53360 27568 53366 27580
rect 52121 27540 53366 27568
rect 52121 27537 52133 27540
rect 52075 27531 52133 27537
rect 53360 27528 53366 27540
rect 53418 27528 53424 27580
rect 54004 27568 54010 27580
rect 53965 27540 54010 27568
rect 54004 27528 54010 27540
rect 54062 27528 54068 27580
rect 54206 27577 54234 27608
rect 57426 27608 58619 27636
rect 57426 27577 57454 27608
rect 58607 27605 58619 27608
rect 58653 27636 58665 27639
rect 58788 27636 58794 27648
rect 58653 27608 58794 27636
rect 58653 27605 58665 27608
rect 58607 27599 58665 27605
rect 58788 27596 58794 27608
rect 58846 27596 58852 27648
rect 61919 27639 61977 27645
rect 61919 27605 61931 27639
rect 61965 27636 61977 27639
rect 62100 27636 62106 27648
rect 61965 27608 62106 27636
rect 61965 27605 61977 27608
rect 61919 27599 61977 27605
rect 62100 27596 62106 27608
rect 62158 27636 62164 27648
rect 62158 27608 63526 27636
rect 62158 27596 62164 27608
rect 54191 27571 54249 27577
rect 54191 27537 54203 27571
rect 54237 27537 54249 27571
rect 54191 27531 54249 27537
rect 57411 27571 57469 27577
rect 57411 27537 57423 27571
rect 57457 27537 57469 27571
rect 57411 27531 57469 27537
rect 57684 27528 57690 27580
rect 57742 27568 57748 27580
rect 57779 27571 57837 27577
rect 57779 27568 57791 27571
rect 57742 27540 57791 27568
rect 57742 27528 57748 27540
rect 57779 27537 57791 27540
rect 57825 27537 57837 27571
rect 61827 27571 61885 27577
rect 61827 27568 61839 27571
rect 57779 27531 57837 27537
rect 57978 27540 61839 27568
rect 45466 27472 50370 27500
rect 50695 27503 50753 27509
rect 37769 27404 37950 27432
rect 39747 27435 39805 27441
rect 37769 27401 37781 27404
rect 37723 27395 37781 27401
rect 39747 27401 39759 27435
rect 39793 27432 39805 27435
rect 44344 27432 44350 27444
rect 39793 27404 43838 27432
rect 44305 27404 44350 27432
rect 39793 27401 39805 27404
rect 39747 27395 39805 27401
rect 36156 27364 36162 27376
rect 34466 27336 36018 27364
rect 36117 27336 36162 27364
rect 34466 27324 34472 27336
rect 36156 27324 36162 27336
rect 36214 27324 36220 27376
rect 42964 27324 42970 27376
rect 43022 27364 43028 27376
rect 43700 27364 43706 27376
rect 43022 27336 43706 27364
rect 43022 27324 43028 27336
rect 43700 27324 43706 27336
rect 43758 27324 43764 27376
rect 43810 27364 43838 27404
rect 44344 27392 44350 27404
rect 44402 27392 44408 27444
rect 45264 27432 45270 27444
rect 45225 27404 45270 27432
rect 45264 27392 45270 27404
rect 45322 27392 45328 27444
rect 45466 27364 45494 27472
rect 50695 27469 50707 27503
rect 50741 27500 50753 27503
rect 51428 27500 51434 27512
rect 50741 27472 51434 27500
rect 50741 27469 50753 27472
rect 50695 27463 50753 27469
rect 51428 27460 51434 27472
rect 51486 27460 51492 27512
rect 51891 27503 51949 27509
rect 51891 27469 51903 27503
rect 51937 27500 51949 27503
rect 52348 27500 52354 27512
rect 51937 27472 52354 27500
rect 51937 27469 51949 27472
rect 51891 27463 51949 27469
rect 52348 27460 52354 27472
rect 52406 27460 52412 27512
rect 55292 27460 55298 27512
rect 55350 27500 55356 27512
rect 57978 27500 58006 27540
rect 61827 27537 61839 27540
rect 61873 27568 61885 27571
rect 62195 27571 62253 27577
rect 62195 27568 62207 27571
rect 61873 27540 62207 27568
rect 61873 27537 61885 27540
rect 61827 27531 61885 27537
rect 62195 27537 62207 27540
rect 62241 27568 62253 27571
rect 63296 27568 63302 27580
rect 62241 27540 63302 27568
rect 62241 27537 62253 27540
rect 62195 27531 62253 27537
rect 63296 27528 63302 27540
rect 63354 27528 63360 27580
rect 55350 27472 58006 27500
rect 58055 27503 58113 27509
rect 55350 27460 55356 27472
rect 58055 27469 58067 27503
rect 58101 27469 58113 27503
rect 58420 27500 58426 27512
rect 58381 27472 58426 27500
rect 58055 27463 58113 27469
rect 45635 27435 45693 27441
rect 45635 27401 45647 27435
rect 45681 27432 45693 27435
rect 45681 27404 51842 27432
rect 45681 27401 45693 27404
rect 45635 27395 45693 27401
rect 43810 27336 45494 27364
rect 45540 27324 45546 27376
rect 45598 27364 45604 27376
rect 48668 27364 48674 27376
rect 45598 27336 48674 27364
rect 45598 27324 45604 27336
rect 48668 27324 48674 27336
rect 48726 27324 48732 27376
rect 49772 27324 49778 27376
rect 49830 27364 49836 27376
rect 50784 27364 50790 27376
rect 49830 27336 50790 27364
rect 49830 27324 49836 27336
rect 50784 27324 50790 27336
rect 50842 27324 50848 27376
rect 51152 27324 51158 27376
rect 51210 27364 51216 27376
rect 51339 27367 51397 27373
rect 51339 27364 51351 27367
rect 51210 27336 51351 27364
rect 51210 27324 51216 27336
rect 51339 27333 51351 27336
rect 51385 27364 51397 27367
rect 51520 27364 51526 27376
rect 51385 27336 51526 27364
rect 51385 27333 51397 27336
rect 51339 27327 51397 27333
rect 51520 27324 51526 27336
rect 51578 27324 51584 27376
rect 51814 27364 51842 27404
rect 56948 27392 56954 27444
rect 57006 27432 57012 27444
rect 58070 27432 58098 27463
rect 58420 27460 58426 27472
rect 58478 27460 58484 27512
rect 62652 27460 62658 27512
rect 62710 27500 62716 27512
rect 62839 27503 62897 27509
rect 62839 27500 62851 27503
rect 62710 27472 62851 27500
rect 62710 27460 62716 27472
rect 62839 27469 62851 27472
rect 62885 27469 62897 27503
rect 63388 27500 63394 27512
rect 63349 27472 63394 27500
rect 62839 27463 62897 27469
rect 63388 27460 63394 27472
rect 63446 27460 63452 27512
rect 63498 27500 63526 27608
rect 63667 27571 63725 27577
rect 63667 27537 63679 27571
rect 63713 27568 63725 27571
rect 64124 27568 64130 27580
rect 63713 27540 64130 27568
rect 63713 27537 63725 27540
rect 63667 27531 63725 27537
rect 64124 27528 64130 27540
rect 64182 27528 64188 27580
rect 67914 27568 67942 27664
rect 68175 27639 68233 27645
rect 68175 27605 68187 27639
rect 68221 27636 68233 27639
rect 70104 27636 70110 27648
rect 68221 27608 70110 27636
rect 68221 27605 68233 27608
rect 68175 27599 68233 27605
rect 70104 27596 70110 27608
rect 70162 27596 70168 27648
rect 73048 27596 73054 27648
rect 73106 27636 73112 27648
rect 74523 27639 74581 27645
rect 74523 27636 74535 27639
rect 73106 27608 74535 27636
rect 73106 27596 73112 27608
rect 74523 27605 74535 27608
rect 74569 27605 74581 27639
rect 74523 27599 74581 27605
rect 68083 27571 68141 27577
rect 68083 27568 68095 27571
rect 67914 27540 68095 27568
rect 68083 27537 68095 27540
rect 68129 27537 68141 27571
rect 68264 27568 68270 27580
rect 68225 27540 68270 27568
rect 68083 27531 68141 27537
rect 68264 27528 68270 27540
rect 68322 27528 68328 27580
rect 70935 27571 70993 27577
rect 70935 27537 70947 27571
rect 70981 27568 70993 27571
rect 71668 27568 71674 27580
rect 70981 27540 71674 27568
rect 70981 27537 70993 27540
rect 70935 27531 70993 27537
rect 71668 27528 71674 27540
rect 71726 27568 71732 27580
rect 71726 27540 72450 27568
rect 71726 27528 71732 27540
rect 63851 27503 63909 27509
rect 63851 27500 63863 27503
rect 63498 27472 63863 27500
rect 63851 27469 63863 27472
rect 63897 27500 63909 27503
rect 65412 27500 65418 27512
rect 63897 27472 65418 27500
rect 63897 27469 63909 27472
rect 63851 27463 63909 27469
rect 65412 27460 65418 27472
rect 65470 27460 65476 27512
rect 67068 27500 67074 27512
rect 65522 27472 67074 27500
rect 65522 27432 65550 27472
rect 67068 27460 67074 27472
rect 67126 27460 67132 27512
rect 67988 27460 67994 27512
rect 68046 27500 68052 27512
rect 69831 27503 69889 27509
rect 69831 27500 69843 27503
rect 68046 27472 69843 27500
rect 68046 27460 68052 27472
rect 69831 27469 69843 27472
rect 69877 27500 69889 27503
rect 72039 27503 72097 27509
rect 72039 27500 72051 27503
rect 69877 27472 72051 27500
rect 69877 27469 69889 27472
rect 69831 27463 69889 27469
rect 72039 27469 72051 27472
rect 72085 27469 72097 27503
rect 72312 27500 72318 27512
rect 72273 27472 72318 27500
rect 72039 27463 72097 27469
rect 57006 27404 58098 27432
rect 62118 27404 65550 27432
rect 57006 27392 57012 27404
rect 62118 27364 62146 27404
rect 66148 27392 66154 27444
rect 66206 27432 66212 27444
rect 70012 27432 70018 27444
rect 66206 27404 70018 27432
rect 66206 27392 66212 27404
rect 70012 27392 70018 27404
rect 70070 27392 70076 27444
rect 51814 27336 62146 27364
rect 68264 27324 68270 27376
rect 68322 27364 68328 27376
rect 68451 27367 68509 27373
rect 68451 27364 68463 27367
rect 68322 27336 68463 27364
rect 68322 27324 68328 27336
rect 68451 27333 68463 27336
rect 68497 27333 68509 27367
rect 68451 27327 68509 27333
rect 68724 27324 68730 27376
rect 68782 27364 68788 27376
rect 71119 27367 71177 27373
rect 71119 27364 71131 27367
rect 68782 27336 71131 27364
rect 68782 27324 68788 27336
rect 71119 27333 71131 27336
rect 71165 27364 71177 27367
rect 71487 27367 71545 27373
rect 71487 27364 71499 27367
rect 71165 27336 71499 27364
rect 71165 27333 71177 27336
rect 71119 27327 71177 27333
rect 71487 27333 71499 27336
rect 71533 27364 71545 27367
rect 71944 27364 71950 27376
rect 71533 27336 71950 27364
rect 71533 27333 71545 27336
rect 71487 27327 71545 27333
rect 71944 27324 71950 27336
rect 72002 27324 72008 27376
rect 72054 27364 72082 27463
rect 72312 27460 72318 27472
rect 72370 27460 72376 27512
rect 72422 27500 72450 27540
rect 73692 27528 73698 27580
rect 73750 27568 73756 27580
rect 74707 27571 74765 27577
rect 74707 27568 74719 27571
rect 73750 27540 74719 27568
rect 73750 27528 73756 27540
rect 74707 27537 74719 27540
rect 74753 27537 74765 27571
rect 74707 27531 74765 27537
rect 78111 27571 78169 27577
rect 78111 27537 78123 27571
rect 78157 27568 78169 27571
rect 78660 27568 78666 27580
rect 78157 27540 78666 27568
rect 78157 27537 78169 27540
rect 78111 27531 78169 27537
rect 78660 27528 78666 27540
rect 78718 27528 78724 27580
rect 75624 27500 75630 27512
rect 72422 27472 75630 27500
rect 75624 27460 75630 27472
rect 75682 27460 75688 27512
rect 78954 27500 78982 27667
rect 80132 27664 80138 27716
rect 80190 27704 80196 27716
rect 80592 27704 80598 27716
rect 80190 27676 80598 27704
rect 80190 27664 80196 27676
rect 80592 27664 80598 27676
rect 80650 27704 80656 27716
rect 83815 27707 83873 27713
rect 80650 27676 82294 27704
rect 80650 27664 80656 27676
rect 81420 27636 81426 27648
rect 79782 27608 81426 27636
rect 79782 27577 79810 27608
rect 81420 27596 81426 27608
rect 81478 27636 81484 27648
rect 82159 27639 82217 27645
rect 82159 27636 82171 27639
rect 81478 27608 82171 27636
rect 81478 27596 81484 27608
rect 82159 27605 82171 27608
rect 82205 27605 82217 27639
rect 82266 27636 82294 27676
rect 83815 27673 83827 27707
rect 83861 27704 83873 27707
rect 90068 27704 90074 27716
rect 83861 27676 90074 27704
rect 83861 27673 83873 27676
rect 83815 27667 83873 27673
rect 90068 27664 90074 27676
rect 90126 27704 90132 27716
rect 90528 27704 90534 27716
rect 90126 27676 90298 27704
rect 90489 27676 90534 27704
rect 90126 27664 90132 27676
rect 84824 27636 84830 27648
rect 82266 27608 84830 27636
rect 82159 27599 82217 27605
rect 84824 27596 84830 27608
rect 84882 27596 84888 27648
rect 89792 27636 89798 27648
rect 87694 27608 89798 27636
rect 87694 27580 87722 27608
rect 89792 27596 89798 27608
rect 89850 27596 89856 27648
rect 90270 27645 90298 27676
rect 90528 27664 90534 27676
rect 90586 27664 90592 27716
rect 91080 27664 91086 27716
rect 91138 27704 91144 27716
rect 91727 27707 91785 27713
rect 91727 27704 91739 27707
rect 91138 27676 91739 27704
rect 91138 27664 91144 27676
rect 91727 27673 91739 27676
rect 91773 27673 91785 27707
rect 91727 27667 91785 27673
rect 90255 27639 90313 27645
rect 90255 27605 90267 27639
rect 90301 27605 90313 27639
rect 90255 27599 90313 27605
rect 79767 27571 79825 27577
rect 79767 27537 79779 27571
rect 79813 27537 79825 27571
rect 79767 27531 79825 27537
rect 79948 27528 79954 27580
rect 80006 27568 80012 27580
rect 80135 27571 80193 27577
rect 80135 27568 80147 27571
rect 80006 27540 80147 27568
rect 80006 27528 80012 27540
rect 80135 27537 80147 27540
rect 80181 27537 80193 27571
rect 80135 27531 80193 27537
rect 80316 27528 80322 27580
rect 80374 27568 80380 27580
rect 82067 27571 82125 27577
rect 82067 27568 82079 27571
rect 80374 27540 82079 27568
rect 80374 27528 80380 27540
rect 82067 27537 82079 27540
rect 82113 27537 82125 27571
rect 82067 27531 82125 27537
rect 83171 27571 83229 27577
rect 83171 27537 83183 27571
rect 83217 27537 83229 27571
rect 83171 27531 83229 27537
rect 79859 27503 79917 27509
rect 79859 27500 79871 27503
rect 78954 27472 79871 27500
rect 79859 27469 79871 27472
rect 79905 27469 79917 27503
rect 79859 27463 79917 27469
rect 73603 27435 73661 27441
rect 73603 27401 73615 27435
rect 73649 27432 73661 27435
rect 75532 27432 75538 27444
rect 73649 27404 75538 27432
rect 73649 27401 73661 27404
rect 73603 27395 73661 27401
rect 75532 27392 75538 27404
rect 75590 27392 75596 27444
rect 78203 27435 78261 27441
rect 78203 27401 78215 27435
rect 78249 27432 78261 27435
rect 79764 27432 79770 27444
rect 78249 27404 79770 27432
rect 78249 27401 78261 27404
rect 78203 27395 78261 27401
rect 79764 27392 79770 27404
rect 79822 27392 79828 27444
rect 73784 27364 73790 27376
rect 72054 27336 73790 27364
rect 73784 27324 73790 27336
rect 73842 27324 73848 27376
rect 73876 27324 73882 27376
rect 73934 27364 73940 27376
rect 74799 27367 74857 27373
rect 74799 27364 74811 27367
rect 73934 27336 74811 27364
rect 73934 27324 73940 27336
rect 74799 27333 74811 27336
rect 74845 27333 74857 27367
rect 74799 27327 74857 27333
rect 79028 27324 79034 27376
rect 79086 27364 79092 27376
rect 79215 27367 79273 27373
rect 79215 27364 79227 27367
rect 79086 27336 79227 27364
rect 79086 27324 79092 27336
rect 79215 27333 79227 27336
rect 79261 27333 79273 27367
rect 79874 27364 79902 27463
rect 80224 27460 80230 27512
rect 80282 27500 80288 27512
rect 83186 27500 83214 27531
rect 83260 27528 83266 27580
rect 83318 27577 83324 27580
rect 83318 27571 83376 27577
rect 83318 27537 83330 27571
rect 83364 27537 83376 27571
rect 84551 27571 84609 27577
rect 84551 27568 84563 27571
rect 83318 27531 83376 27537
rect 83462 27540 84563 27568
rect 83318 27528 83324 27531
rect 83462 27500 83490 27540
rect 84551 27537 84563 27540
rect 84597 27568 84609 27571
rect 84735 27571 84793 27577
rect 84735 27568 84747 27571
rect 84597 27540 84747 27568
rect 84597 27537 84609 27540
rect 84551 27531 84609 27537
rect 84735 27537 84747 27540
rect 84781 27537 84793 27571
rect 85287 27571 85345 27577
rect 85287 27568 85299 27571
rect 84735 27531 84793 27537
rect 84842 27540 85299 27568
rect 80282 27472 83214 27500
rect 83278 27472 83490 27500
rect 83539 27503 83597 27509
rect 80282 27460 80288 27472
rect 80500 27392 80506 27444
rect 80558 27432 80564 27444
rect 83278 27432 83306 27472
rect 83539 27469 83551 27503
rect 83585 27500 83597 27503
rect 84088 27500 84094 27512
rect 83585 27472 84094 27500
rect 83585 27469 83597 27472
rect 83539 27463 83597 27469
rect 84088 27460 84094 27472
rect 84146 27460 84152 27512
rect 80558 27404 83306 27432
rect 83447 27435 83505 27441
rect 80558 27392 80564 27404
rect 83447 27401 83459 27435
rect 83493 27432 83505 27435
rect 84842 27432 84870 27540
rect 85287 27537 85299 27540
rect 85333 27568 85345 27571
rect 86112 27568 86118 27580
rect 85333 27540 86118 27568
rect 85333 27537 85345 27540
rect 85287 27531 85345 27537
rect 86112 27528 86118 27540
rect 86170 27528 86176 27580
rect 87676 27568 87682 27580
rect 87589 27540 87682 27568
rect 87676 27528 87682 27540
rect 87734 27528 87740 27580
rect 89240 27568 89246 27580
rect 89201 27540 89246 27568
rect 89240 27528 89246 27540
rect 89298 27528 89304 27580
rect 90344 27528 90350 27580
rect 90402 27568 90408 27580
rect 90439 27571 90497 27577
rect 90439 27568 90451 27571
rect 90402 27540 90451 27568
rect 90402 27528 90408 27540
rect 90439 27537 90451 27540
rect 90485 27537 90497 27571
rect 90546 27568 90574 27664
rect 91635 27571 91693 27577
rect 91635 27568 91647 27571
rect 90546 27540 91647 27568
rect 90439 27531 90497 27537
rect 91635 27537 91647 27540
rect 91681 27537 91693 27571
rect 91635 27531 91693 27537
rect 85744 27500 85750 27512
rect 85705 27472 85750 27500
rect 85744 27460 85750 27472
rect 85802 27460 85808 27512
rect 86130 27500 86158 27528
rect 87771 27503 87829 27509
rect 87771 27500 87783 27503
rect 86130 27472 87783 27500
rect 87771 27469 87783 27472
rect 87817 27469 87829 27503
rect 87771 27463 87829 27469
rect 85008 27432 85014 27444
rect 83493 27404 84870 27432
rect 84969 27404 85014 27432
rect 83493 27401 83505 27404
rect 83447 27395 83505 27401
rect 85008 27392 85014 27404
rect 85066 27392 85072 27444
rect 87584 27364 87590 27376
rect 79874 27336 87590 27364
rect 79215 27327 79273 27333
rect 87584 27324 87590 27336
rect 87642 27324 87648 27376
rect 89332 27364 89338 27376
rect 89293 27336 89338 27364
rect 89332 27324 89338 27336
rect 89390 27324 89396 27376
rect 538 27274 93642 27296
rect 538 27222 3680 27274
rect 3732 27222 3744 27274
rect 3796 27222 3808 27274
rect 3860 27222 3872 27274
rect 3924 27222 9008 27274
rect 9060 27222 9072 27274
rect 9124 27222 9136 27274
rect 9188 27222 9200 27274
rect 9252 27222 14336 27274
rect 14388 27222 14400 27274
rect 14452 27222 14464 27274
rect 14516 27222 14528 27274
rect 14580 27222 19664 27274
rect 19716 27222 19728 27274
rect 19780 27222 19792 27274
rect 19844 27222 19856 27274
rect 19908 27222 24992 27274
rect 25044 27222 25056 27274
rect 25108 27222 25120 27274
rect 25172 27222 25184 27274
rect 25236 27222 30320 27274
rect 30372 27222 30384 27274
rect 30436 27222 30448 27274
rect 30500 27222 30512 27274
rect 30564 27222 35648 27274
rect 35700 27222 35712 27274
rect 35764 27222 35776 27274
rect 35828 27222 35840 27274
rect 35892 27222 40976 27274
rect 41028 27222 41040 27274
rect 41092 27222 41104 27274
rect 41156 27222 41168 27274
rect 41220 27222 46304 27274
rect 46356 27222 46368 27274
rect 46420 27222 46432 27274
rect 46484 27222 46496 27274
rect 46548 27222 51632 27274
rect 51684 27222 51696 27274
rect 51748 27222 51760 27274
rect 51812 27222 51824 27274
rect 51876 27222 56960 27274
rect 57012 27222 57024 27274
rect 57076 27222 57088 27274
rect 57140 27222 57152 27274
rect 57204 27222 62288 27274
rect 62340 27222 62352 27274
rect 62404 27222 62416 27274
rect 62468 27222 62480 27274
rect 62532 27222 67616 27274
rect 67668 27222 67680 27274
rect 67732 27222 67744 27274
rect 67796 27222 67808 27274
rect 67860 27222 72944 27274
rect 72996 27222 73008 27274
rect 73060 27222 73072 27274
rect 73124 27222 73136 27274
rect 73188 27222 78272 27274
rect 78324 27222 78336 27274
rect 78388 27222 78400 27274
rect 78452 27222 78464 27274
rect 78516 27222 83600 27274
rect 83652 27222 83664 27274
rect 83716 27222 83728 27274
rect 83780 27222 83792 27274
rect 83844 27222 88928 27274
rect 88980 27222 88992 27274
rect 89044 27222 89056 27274
rect 89108 27222 89120 27274
rect 89172 27222 93642 27274
rect 538 27200 93642 27222
rect 3867 27163 3925 27169
rect 3867 27129 3879 27163
rect 3913 27160 3925 27163
rect 4048 27160 4054 27172
rect 3913 27132 4054 27160
rect 3913 27129 3925 27132
rect 3867 27123 3925 27129
rect 4048 27120 4054 27132
rect 4106 27120 4112 27172
rect 9292 27160 9298 27172
rect 9253 27132 9298 27160
rect 9292 27120 9298 27132
rect 9350 27120 9356 27172
rect 11687 27163 11745 27169
rect 11687 27129 11699 27163
rect 11733 27160 11745 27163
rect 12144 27160 12150 27172
rect 11733 27132 12150 27160
rect 11733 27129 11745 27132
rect 11687 27123 11745 27129
rect 12144 27120 12150 27132
rect 12202 27160 12208 27172
rect 12696 27160 12702 27172
rect 12202 27132 12702 27160
rect 12202 27120 12208 27132
rect 12696 27120 12702 27132
rect 12754 27120 12760 27172
rect 13156 27160 13162 27172
rect 13117 27132 13162 27160
rect 13156 27120 13162 27132
rect 13214 27120 13220 27172
rect 16468 27160 16474 27172
rect 15106 27132 16330 27160
rect 16429 27132 16474 27160
rect 4600 27052 4606 27104
rect 4658 27092 4664 27104
rect 4658 27064 10534 27092
rect 4658 27052 4664 27064
rect 2303 27027 2361 27033
rect 2303 26993 2315 27027
rect 2349 27024 2361 27027
rect 2944 27024 2950 27036
rect 2349 26996 2950 27024
rect 2349 26993 2361 26996
rect 2303 26987 2361 26993
rect 2944 26984 2950 26996
rect 3002 27024 3008 27036
rect 10506 27024 10534 27064
rect 10580 27052 10586 27104
rect 10638 27092 10644 27104
rect 14999 27095 15057 27101
rect 14999 27092 15011 27095
rect 10638 27064 15011 27092
rect 10638 27052 10644 27064
rect 14999 27061 15011 27064
rect 15045 27061 15057 27095
rect 14999 27055 15057 27061
rect 3002 26996 4186 27024
rect 10506 26996 11914 27024
rect 3002 26984 3008 26996
rect 2579 26959 2637 26965
rect 2579 26925 2591 26959
rect 2625 26956 2637 26959
rect 4048 26956 4054 26968
rect 2625 26928 4054 26956
rect 2625 26925 2637 26928
rect 2579 26919 2637 26925
rect 4048 26916 4054 26928
rect 4106 26916 4112 26968
rect 4158 26897 4186 26996
rect 4416 26916 4422 26968
rect 4474 26956 4480 26968
rect 4692 26956 4698 26968
rect 4474 26928 4698 26956
rect 4474 26916 4480 26928
rect 4692 26916 4698 26928
rect 4750 26956 4756 26968
rect 4787 26959 4845 26965
rect 4787 26956 4799 26959
rect 4750 26928 4799 26956
rect 4750 26916 4756 26928
rect 4787 26925 4799 26928
rect 4833 26925 4845 26959
rect 4787 26919 4845 26925
rect 9292 26916 9298 26968
rect 9350 26956 9356 26968
rect 9387 26959 9445 26965
rect 9387 26956 9399 26959
rect 9350 26928 9399 26956
rect 9350 26916 9356 26928
rect 9387 26925 9399 26928
rect 9433 26925 9445 26959
rect 9387 26919 9445 26925
rect 9571 26959 9629 26965
rect 9571 26925 9583 26959
rect 9617 26956 9629 26959
rect 10120 26956 10126 26968
rect 9617 26928 10126 26956
rect 9617 26925 9629 26928
rect 9571 26919 9629 26925
rect 10120 26916 10126 26928
rect 10178 26916 10184 26968
rect 10304 26916 10310 26968
rect 10362 26956 10368 26968
rect 10362 26928 10455 26956
rect 10362 26916 10368 26928
rect 4143 26891 4201 26897
rect 4143 26857 4155 26891
rect 4189 26888 4201 26891
rect 5520 26888 5526 26900
rect 4189 26860 5526 26888
rect 4189 26857 4201 26860
rect 4143 26851 4201 26857
rect 5520 26848 5526 26860
rect 5578 26848 5584 26900
rect 9016 26848 9022 26900
rect 9074 26888 9080 26900
rect 10322 26888 10350 26916
rect 10672 26888 10678 26900
rect 9074 26860 9522 26888
rect 9074 26848 9080 26860
rect 4784 26780 4790 26832
rect 4842 26820 4848 26832
rect 4971 26823 5029 26829
rect 4971 26820 4983 26823
rect 4842 26792 4983 26820
rect 4842 26780 4848 26792
rect 4971 26789 4983 26792
rect 5017 26789 5029 26823
rect 9494 26820 9522 26860
rect 10230 26860 10350 26888
rect 10633 26860 10678 26888
rect 10230 26820 10258 26860
rect 10672 26848 10678 26860
rect 10730 26848 10736 26900
rect 9494 26792 10258 26820
rect 11886 26820 11914 26996
rect 12052 26984 12058 27036
rect 12110 27024 12116 27036
rect 12791 27027 12849 27033
rect 12791 27024 12803 27027
rect 12110 26996 12803 27024
rect 12110 26984 12116 26996
rect 12791 26993 12803 26996
rect 12837 26993 12849 27027
rect 12791 26987 12849 26993
rect 11963 26959 12021 26965
rect 11963 26925 11975 26959
rect 12009 26925 12021 26959
rect 12420 26956 12426 26968
rect 12381 26928 12426 26956
rect 11963 26919 12021 26925
rect 11978 26888 12006 26919
rect 12420 26916 12426 26928
rect 12478 26916 12484 26968
rect 12696 26956 12702 26968
rect 12657 26928 12702 26956
rect 12696 26916 12702 26928
rect 12754 26916 12760 26968
rect 13251 26959 13309 26965
rect 13251 26956 13263 26959
rect 12898 26928 13263 26956
rect 12898 26888 12926 26928
rect 13251 26925 13263 26928
rect 13297 26956 13309 26959
rect 15106 26956 15134 27132
rect 16103 27095 16161 27101
rect 16103 27061 16115 27095
rect 16149 27061 16161 27095
rect 16302 27092 16330 27132
rect 16468 27120 16474 27132
rect 16526 27120 16532 27172
rect 16560 27120 16566 27172
rect 16618 27160 16624 27172
rect 16747 27163 16805 27169
rect 16747 27160 16759 27163
rect 16618 27132 16759 27160
rect 16618 27120 16624 27132
rect 16747 27129 16759 27132
rect 16793 27160 16805 27163
rect 19599 27163 19657 27169
rect 19599 27160 19611 27163
rect 16793 27132 19611 27160
rect 16793 27129 16805 27132
rect 16747 27123 16805 27129
rect 19599 27129 19611 27132
rect 19645 27160 19657 27163
rect 19645 27132 24610 27160
rect 19645 27129 19657 27132
rect 19599 27123 19657 27129
rect 17572 27092 17578 27104
rect 16302 27064 17578 27092
rect 16103 27055 16161 27061
rect 15640 27024 15646 27036
rect 15198 26996 15646 27024
rect 15198 26965 15226 26996
rect 15640 26984 15646 26996
rect 15698 27024 15704 27036
rect 16118 27024 16146 27055
rect 17572 27052 17578 27064
rect 17630 27052 17636 27104
rect 17756 27052 17762 27104
rect 17814 27092 17820 27104
rect 17851 27095 17909 27101
rect 17851 27092 17863 27095
rect 17814 27064 17863 27092
rect 17814 27052 17820 27064
rect 17851 27061 17863 27064
rect 17897 27061 17909 27095
rect 23736 27092 23742 27104
rect 17851 27055 17909 27061
rect 20902 27064 23742 27092
rect 15698 26996 16146 27024
rect 16210 26996 16698 27024
rect 15698 26984 15704 26996
rect 13297 26928 15134 26956
rect 15183 26959 15241 26965
rect 13297 26925 13309 26928
rect 13251 26919 13309 26925
rect 15183 26925 15195 26959
rect 15229 26925 15241 26959
rect 15183 26919 15241 26925
rect 16210 26888 16238 26996
rect 16287 26959 16345 26965
rect 16287 26925 16299 26959
rect 16333 26925 16345 26959
rect 16287 26919 16345 26925
rect 16379 26959 16437 26965
rect 16379 26925 16391 26959
rect 16425 26956 16437 26959
rect 16560 26956 16566 26968
rect 16425 26928 16566 26956
rect 16425 26925 16437 26928
rect 16379 26919 16437 26925
rect 11978 26860 12926 26888
rect 12990 26860 16238 26888
rect 16302 26888 16330 26919
rect 16560 26916 16566 26928
rect 16618 26916 16624 26968
rect 16670 26956 16698 26996
rect 17020 26984 17026 27036
rect 17078 27024 17084 27036
rect 18311 27027 18369 27033
rect 18311 27024 18323 27027
rect 17078 26996 18323 27024
rect 17078 26984 17084 26996
rect 18311 26993 18323 26996
rect 18357 26993 18369 27027
rect 18311 26987 18369 26993
rect 17664 26956 17670 26968
rect 16670 26928 17670 26956
rect 17664 26916 17670 26928
rect 17722 26916 17728 26968
rect 17756 26916 17762 26968
rect 17814 26956 17820 26968
rect 18035 26959 18093 26965
rect 18035 26956 18047 26959
rect 17814 26928 18047 26956
rect 17814 26916 17820 26928
rect 18035 26925 18047 26928
rect 18081 26925 18093 26959
rect 18035 26919 18093 26925
rect 18142 26928 18998 26956
rect 16931 26891 16989 26897
rect 16931 26888 16943 26891
rect 16302 26860 16943 26888
rect 12990 26820 13018 26860
rect 16931 26857 16943 26860
rect 16977 26888 16989 26891
rect 18142 26888 18170 26928
rect 16977 26860 18170 26888
rect 18970 26888 18998 26928
rect 19136 26916 19142 26968
rect 19194 26956 19200 26968
rect 20902 26965 20930 27064
rect 23736 27052 23742 27064
rect 23794 27052 23800 27104
rect 24472 27092 24478 27104
rect 23938 27064 24478 27092
rect 22540 26984 22546 27036
rect 22598 27024 22604 27036
rect 23938 27033 23966 27064
rect 24472 27052 24478 27064
rect 24530 27052 24536 27104
rect 24582 27092 24610 27132
rect 24656 27120 24662 27172
rect 24714 27160 24720 27172
rect 24714 27132 29946 27160
rect 24714 27120 24720 27132
rect 25579 27095 25637 27101
rect 24582 27064 25438 27092
rect 23187 27027 23245 27033
rect 23187 27024 23199 27027
rect 22598 26996 23199 27024
rect 22598 26984 22604 26996
rect 23187 26993 23199 26996
rect 23233 26993 23245 27027
rect 23187 26987 23245 26993
rect 23923 27027 23981 27033
rect 23923 26993 23935 27027
rect 23969 26993 23981 27027
rect 24104 27024 24110 27036
rect 24065 26996 24110 27024
rect 23923 26987 23981 26993
rect 24104 26984 24110 26996
rect 24162 27024 24168 27036
rect 25303 27027 25361 27033
rect 25303 27024 25315 27027
rect 24162 26996 25315 27024
rect 24162 26984 24168 26996
rect 25303 26993 25315 26996
rect 25349 26993 25361 27027
rect 25410 27024 25438 27064
rect 25579 27061 25591 27095
rect 25625 27092 25637 27095
rect 25852 27092 25858 27104
rect 25625 27064 25858 27092
rect 25625 27061 25637 27064
rect 25579 27055 25637 27061
rect 25852 27052 25858 27064
rect 25910 27052 25916 27104
rect 26956 27052 26962 27104
rect 27014 27092 27020 27104
rect 27014 27064 27922 27092
rect 27014 27052 27020 27064
rect 25410 26996 27830 27024
rect 25303 26987 25361 26993
rect 20519 26959 20577 26965
rect 20519 26956 20531 26959
rect 19194 26928 20531 26956
rect 19194 26916 19200 26928
rect 20519 26925 20531 26928
rect 20565 26956 20577 26959
rect 20887 26959 20945 26965
rect 20887 26956 20899 26959
rect 20565 26928 20899 26956
rect 20565 26925 20577 26928
rect 20519 26919 20577 26925
rect 20887 26925 20899 26928
rect 20933 26925 20945 26959
rect 22908 26956 22914 26968
rect 22869 26928 22914 26956
rect 20887 26919 20945 26925
rect 22908 26916 22914 26928
rect 22966 26956 22972 26968
rect 23831 26959 23889 26965
rect 23831 26956 23843 26959
rect 22966 26928 23843 26956
rect 22966 26916 22972 26928
rect 23831 26925 23843 26928
rect 23877 26925 23889 26959
rect 23831 26919 23889 26925
rect 23644 26888 23650 26900
rect 18970 26860 23650 26888
rect 16977 26857 16989 26860
rect 16931 26851 16989 26857
rect 23644 26848 23650 26860
rect 23702 26848 23708 26900
rect 11886 26792 13018 26820
rect 4971 26783 5029 26789
rect 18768 26780 18774 26832
rect 18826 26820 18832 26832
rect 20703 26823 20761 26829
rect 20703 26820 20715 26823
rect 18826 26792 20715 26820
rect 18826 26780 18832 26792
rect 20703 26789 20715 26792
rect 20749 26789 20761 26823
rect 23846 26820 23874 26919
rect 24012 26916 24018 26968
rect 24070 26956 24076 26968
rect 24199 26959 24257 26965
rect 24199 26956 24211 26959
rect 24070 26928 24211 26956
rect 24070 26916 24076 26928
rect 24199 26925 24211 26928
rect 24245 26925 24257 26959
rect 24199 26919 24257 26925
rect 24567 26959 24625 26965
rect 24567 26925 24579 26959
rect 24613 26956 24625 26959
rect 24656 26956 24662 26968
rect 24613 26928 24662 26956
rect 24613 26925 24625 26928
rect 24567 26919 24625 26925
rect 24656 26916 24662 26928
rect 24714 26916 24720 26968
rect 25211 26959 25269 26965
rect 25211 26925 25223 26959
rect 25257 26956 25269 26959
rect 25852 26956 25858 26968
rect 25257 26928 25858 26956
rect 25257 26925 25269 26928
rect 25211 26919 25269 26925
rect 25852 26916 25858 26928
rect 25910 26916 25916 26968
rect 27600 26956 27606 26968
rect 27561 26928 27606 26956
rect 27600 26916 27606 26928
rect 27658 26916 27664 26968
rect 23920 26848 23926 26900
rect 23978 26888 23984 26900
rect 27695 26891 27753 26897
rect 27695 26888 27707 26891
rect 23978 26860 27707 26888
rect 23978 26848 23984 26860
rect 27695 26857 27707 26860
rect 27741 26857 27753 26891
rect 27802 26888 27830 26996
rect 27894 26956 27922 27064
rect 27968 27052 27974 27104
rect 28026 27092 28032 27104
rect 28612 27092 28618 27104
rect 28026 27064 28618 27092
rect 28026 27052 28032 27064
rect 28612 27052 28618 27064
rect 28670 27052 28676 27104
rect 29167 27095 29225 27101
rect 29167 27061 29179 27095
rect 29213 27092 29225 27095
rect 29918 27092 29946 27132
rect 30728 27120 30734 27172
rect 30786 27160 30792 27172
rect 33764 27160 33770 27172
rect 30786 27132 33770 27160
rect 30786 27120 30792 27132
rect 33764 27120 33770 27132
rect 33822 27120 33828 27172
rect 33948 27160 33954 27172
rect 33909 27132 33954 27160
rect 33948 27120 33954 27132
rect 34006 27160 34012 27172
rect 34043 27163 34101 27169
rect 34043 27160 34055 27163
rect 34006 27132 34055 27160
rect 34006 27120 34012 27132
rect 34043 27129 34055 27132
rect 34089 27129 34101 27163
rect 34043 27123 34101 27129
rect 34132 27120 34138 27172
rect 34190 27160 34196 27172
rect 34319 27163 34377 27169
rect 34319 27160 34331 27163
rect 34190 27132 34331 27160
rect 34190 27120 34196 27132
rect 34319 27129 34331 27132
rect 34365 27129 34377 27163
rect 34319 27123 34377 27129
rect 35236 27120 35242 27172
rect 35294 27160 35300 27172
rect 35699 27163 35757 27169
rect 35699 27160 35711 27163
rect 35294 27132 35711 27160
rect 35294 27120 35300 27132
rect 35699 27129 35711 27132
rect 35745 27160 35757 27163
rect 43240 27160 43246 27172
rect 35745 27132 36110 27160
rect 35745 27129 35757 27132
rect 35699 27123 35757 27129
rect 30820 27092 30826 27104
rect 29213 27064 29854 27092
rect 29918 27064 30826 27092
rect 29213 27061 29225 27064
rect 29167 27055 29225 27061
rect 29182 26956 29210 27055
rect 29440 27024 29446 27036
rect 29401 26996 29446 27024
rect 29440 26984 29446 26996
rect 29498 26984 29504 27036
rect 29826 27024 29854 27064
rect 30820 27052 30826 27064
rect 30878 27052 30884 27104
rect 31464 27052 31470 27104
rect 31522 27092 31528 27104
rect 31559 27095 31617 27101
rect 31559 27092 31571 27095
rect 31522 27064 31571 27092
rect 31522 27052 31528 27064
rect 31559 27061 31571 27064
rect 31605 27061 31617 27095
rect 31559 27055 31617 27061
rect 31648 27052 31654 27104
rect 31706 27092 31712 27104
rect 32939 27095 32997 27101
rect 32939 27092 32951 27095
rect 31706 27064 32951 27092
rect 31706 27052 31712 27064
rect 32939 27061 32951 27064
rect 32985 27092 32997 27095
rect 33031 27095 33089 27101
rect 33031 27092 33043 27095
rect 32985 27064 33043 27092
rect 32985 27061 32997 27064
rect 32939 27055 32997 27061
rect 33031 27061 33043 27064
rect 33077 27061 33089 27095
rect 33031 27055 33089 27061
rect 33120 27052 33126 27104
rect 33178 27092 33184 27104
rect 35604 27092 35610 27104
rect 33178 27064 35610 27092
rect 33178 27052 33184 27064
rect 35604 27052 35610 27064
rect 35662 27052 35668 27104
rect 31280 27024 31286 27036
rect 29826 26996 30314 27024
rect 30286 26968 30314 26996
rect 30930 26996 31286 27024
rect 27894 26928 29210 26956
rect 29808 26916 29814 26968
rect 29866 26956 29872 26968
rect 29903 26959 29961 26965
rect 29903 26956 29915 26959
rect 29866 26928 29915 26956
rect 29866 26916 29872 26928
rect 29903 26925 29915 26928
rect 29949 26925 29961 26959
rect 30087 26959 30145 26965
rect 30087 26956 30099 26959
rect 29903 26919 29961 26925
rect 30010 26928 30099 26956
rect 29348 26888 29354 26900
rect 27802 26860 29354 26888
rect 27695 26851 27753 26857
rect 29348 26848 29354 26860
rect 29406 26848 29412 26900
rect 29259 26823 29317 26829
rect 29259 26820 29271 26823
rect 23846 26792 29271 26820
rect 20703 26783 20761 26789
rect 29259 26789 29271 26792
rect 29305 26820 29317 26823
rect 30010 26820 30038 26928
rect 30087 26925 30099 26928
rect 30133 26925 30145 26959
rect 30087 26919 30145 26925
rect 30268 26916 30274 26968
rect 30326 26956 30332 26968
rect 30455 26959 30513 26965
rect 30455 26956 30467 26959
rect 30326 26928 30467 26956
rect 30326 26916 30332 26928
rect 30455 26925 30467 26928
rect 30501 26925 30513 26959
rect 30455 26919 30513 26925
rect 30639 26959 30697 26965
rect 30639 26925 30651 26959
rect 30685 26956 30697 26959
rect 30728 26956 30734 26968
rect 30685 26928 30734 26956
rect 30685 26925 30697 26928
rect 30639 26919 30697 26925
rect 30728 26916 30734 26928
rect 30786 26916 30792 26968
rect 30930 26820 30958 26996
rect 31280 26984 31286 26996
rect 31338 26984 31344 27036
rect 35883 27027 35941 27033
rect 35883 27024 35895 27027
rect 31482 26996 35895 27024
rect 31188 26956 31194 26968
rect 29305 26792 30958 26820
rect 31022 26928 31194 26956
rect 31022 26820 31050 26928
rect 31188 26916 31194 26928
rect 31246 26916 31252 26968
rect 31482 26965 31510 26996
rect 35883 26993 35895 26996
rect 35929 26993 35941 27027
rect 36082 27024 36110 27132
rect 42522 27132 43246 27160
rect 36156 27052 36162 27104
rect 36214 27092 36220 27104
rect 42522 27092 42550 27132
rect 43240 27120 43246 27132
rect 43298 27120 43304 27172
rect 43427 27163 43485 27169
rect 43427 27129 43439 27163
rect 43473 27160 43485 27163
rect 45356 27160 45362 27172
rect 43473 27132 45362 27160
rect 43473 27129 43485 27132
rect 43427 27123 43485 27129
rect 45356 27120 45362 27132
rect 45414 27120 45420 27172
rect 48668 27120 48674 27172
rect 48726 27160 48732 27172
rect 55292 27160 55298 27172
rect 48726 27132 55298 27160
rect 48726 27120 48732 27132
rect 55292 27120 55298 27132
rect 55350 27120 55356 27172
rect 56488 27160 56494 27172
rect 56449 27132 56494 27160
rect 56488 27120 56494 27132
rect 56546 27120 56552 27172
rect 58328 27160 58334 27172
rect 56598 27132 58190 27160
rect 58289 27132 58334 27160
rect 51152 27092 51158 27104
rect 36214 27064 42550 27092
rect 42614 27064 51158 27092
rect 36214 27052 36220 27064
rect 36082 26996 36570 27024
rect 35883 26987 35941 26993
rect 36542 26968 36570 26996
rect 39008 26984 39014 27036
rect 39066 27024 39072 27036
rect 42614 27024 42642 27064
rect 51152 27052 51158 27064
rect 51210 27052 51216 27104
rect 52900 27092 52906 27104
rect 52861 27064 52906 27092
rect 52900 27052 52906 27064
rect 52958 27052 52964 27104
rect 53728 27052 53734 27104
rect 53786 27092 53792 27104
rect 56598 27092 56626 27132
rect 53786 27064 56626 27092
rect 58162 27092 58190 27132
rect 58328 27120 58334 27132
rect 58386 27120 58392 27172
rect 91172 27160 91178 27172
rect 58438 27132 91178 27160
rect 58438 27092 58466 27132
rect 91172 27120 91178 27132
rect 91230 27120 91236 27172
rect 58162 27064 58466 27092
rect 53786 27052 53792 27064
rect 63388 27052 63394 27104
rect 63446 27092 63452 27104
rect 64955 27095 65013 27101
rect 64955 27092 64967 27095
rect 63446 27064 64967 27092
rect 63446 27052 63452 27064
rect 64955 27061 64967 27064
rect 65001 27061 65013 27095
rect 66148 27092 66154 27104
rect 66109 27064 66154 27092
rect 64955 27055 65013 27061
rect 66148 27052 66154 27064
rect 66206 27052 66212 27104
rect 69368 27092 69374 27104
rect 69329 27064 69374 27092
rect 69368 27052 69374 27064
rect 69426 27052 69432 27104
rect 70751 27095 70809 27101
rect 70751 27061 70763 27095
rect 70797 27092 70809 27095
rect 71116 27092 71122 27104
rect 70797 27064 71122 27092
rect 70797 27061 70809 27064
rect 70751 27055 70809 27061
rect 71116 27052 71122 27064
rect 71174 27052 71180 27104
rect 73695 27095 73753 27101
rect 73695 27092 73707 27095
rect 72422 27064 73707 27092
rect 39066 26996 42642 27024
rect 43795 27027 43853 27033
rect 39066 26984 39072 26996
rect 43795 26993 43807 27027
rect 43841 27024 43853 27027
rect 43979 27027 44037 27033
rect 43979 27024 43991 27027
rect 43841 26996 43991 27024
rect 43841 26993 43853 26996
rect 43795 26987 43853 26993
rect 43979 26993 43991 26996
rect 44025 27024 44037 27027
rect 44160 27024 44166 27036
rect 44025 26996 44166 27024
rect 44025 26993 44037 26996
rect 43979 26987 44037 26993
rect 31467 26959 31525 26965
rect 31467 26925 31479 26959
rect 31513 26925 31525 26959
rect 31467 26919 31525 26925
rect 33215 26959 33273 26965
rect 33215 26925 33227 26959
rect 33261 26956 33273 26959
rect 35144 26956 35150 26968
rect 33261 26928 35150 26956
rect 33261 26925 33273 26928
rect 33215 26919 33273 26925
rect 35144 26916 35150 26928
rect 35202 26916 35208 26968
rect 36340 26956 36346 26968
rect 36301 26928 36346 26956
rect 36340 26916 36346 26928
rect 36398 26916 36404 26968
rect 36524 26956 36530 26968
rect 36437 26928 36530 26956
rect 36524 26916 36530 26928
rect 36582 26916 36588 26968
rect 36708 26916 36714 26968
rect 36766 26956 36772 26968
rect 36895 26959 36953 26965
rect 36895 26956 36907 26959
rect 36766 26928 36907 26956
rect 36766 26916 36772 26928
rect 36895 26925 36907 26928
rect 36941 26925 36953 26959
rect 36895 26919 36953 26925
rect 37079 26959 37137 26965
rect 37079 26925 37091 26959
rect 37125 26956 37137 26959
rect 39284 26956 39290 26968
rect 37125 26928 39290 26956
rect 37125 26925 37137 26928
rect 37079 26919 37137 26925
rect 39284 26916 39290 26928
rect 39342 26916 39348 26968
rect 42415 26959 42473 26965
rect 42415 26925 42427 26959
rect 42461 26925 42473 26959
rect 42415 26919 42473 26925
rect 34960 26888 34966 26900
rect 31574 26860 34966 26888
rect 31574 26820 31602 26860
rect 34960 26848 34966 26860
rect 35018 26848 35024 26900
rect 35604 26888 35610 26900
rect 35517 26860 35610 26888
rect 35604 26848 35610 26860
rect 35662 26888 35668 26900
rect 36726 26888 36754 26916
rect 35662 26860 36754 26888
rect 42430 26888 42458 26919
rect 42504 26916 42510 26968
rect 42562 26956 42568 26968
rect 42875 26959 42933 26965
rect 42875 26956 42887 26959
rect 42562 26928 42887 26956
rect 42562 26916 42568 26928
rect 42875 26925 42887 26928
rect 42921 26925 42933 26959
rect 42875 26919 42933 26925
rect 42967 26959 43025 26965
rect 42967 26925 42979 26959
rect 43013 26956 43025 26959
rect 43810 26956 43838 26987
rect 44160 26984 44166 26996
rect 44218 26984 44224 27036
rect 44344 26984 44350 27036
rect 44402 27024 44408 27036
rect 48392 27024 48398 27036
rect 44402 26996 48398 27024
rect 44402 26984 44408 26996
rect 48392 26984 48398 26996
rect 48450 26984 48456 27036
rect 48855 27027 48913 27033
rect 48855 26993 48867 27027
rect 48901 27024 48913 27027
rect 50140 27024 50146 27036
rect 48901 26996 50002 27024
rect 50101 26996 50146 27024
rect 48901 26993 48913 26996
rect 48855 26987 48913 26993
rect 43013 26928 43838 26956
rect 48487 26959 48545 26965
rect 43013 26925 43025 26928
rect 42967 26919 43025 26925
rect 48487 26925 48499 26959
rect 48533 26956 48545 26959
rect 48576 26956 48582 26968
rect 48533 26928 48582 26956
rect 48533 26925 48545 26928
rect 48487 26919 48545 26925
rect 42982 26888 43010 26919
rect 48576 26916 48582 26928
rect 48634 26916 48640 26968
rect 49867 26959 49925 26965
rect 49867 26925 49879 26959
rect 49913 26925 49925 26959
rect 49974 26956 50002 26996
rect 50140 26984 50146 26996
rect 50198 26984 50204 27036
rect 51428 27024 51434 27036
rect 50342 26996 51290 27024
rect 51389 26996 51434 27024
rect 50232 26956 50238 26968
rect 49974 26928 50238 26956
rect 49867 26919 49925 26925
rect 42430 26860 43010 26888
rect 48303 26891 48361 26897
rect 35662 26848 35668 26860
rect 48303 26857 48315 26891
rect 48349 26888 48361 26891
rect 49312 26888 49318 26900
rect 48349 26860 49318 26888
rect 48349 26857 48361 26860
rect 48303 26851 48361 26857
rect 49312 26848 49318 26860
rect 49370 26848 49376 26900
rect 49683 26891 49741 26897
rect 49683 26857 49695 26891
rect 49729 26888 49741 26891
rect 49882 26888 49910 26919
rect 50232 26916 50238 26928
rect 50290 26916 50296 26968
rect 50342 26888 50370 26996
rect 50416 26916 50422 26968
rect 50474 26916 50480 26968
rect 51060 26916 51066 26968
rect 51118 26956 51124 26968
rect 51155 26959 51213 26965
rect 51155 26956 51167 26959
rect 51118 26928 51167 26956
rect 51118 26916 51124 26928
rect 51155 26925 51167 26928
rect 51201 26925 51213 26959
rect 51262 26956 51290 26996
rect 51428 26984 51434 26996
rect 51486 26984 51492 27036
rect 52164 26984 52170 27036
rect 52222 27024 52228 27036
rect 52535 27027 52593 27033
rect 52535 27024 52547 27027
rect 52222 26996 52547 27024
rect 52222 26984 52228 26996
rect 52535 26993 52547 26996
rect 52581 26993 52593 27027
rect 52535 26987 52593 26993
rect 52550 26956 52578 26987
rect 56488 26984 56494 27036
rect 56546 27024 56552 27036
rect 56767 27027 56825 27033
rect 56767 27024 56779 27027
rect 56546 26996 56779 27024
rect 56546 26984 56552 26996
rect 56767 26993 56779 26996
rect 56813 26993 56825 27027
rect 56767 26987 56825 26993
rect 61180 26984 61186 27036
rect 61238 27024 61244 27036
rect 62379 27027 62437 27033
rect 62379 27024 62391 27027
rect 61238 26996 62391 27024
rect 61238 26984 61244 26996
rect 62379 26993 62391 26996
rect 62425 26993 62437 27027
rect 62652 27024 62658 27036
rect 62613 26996 62658 27024
rect 62379 26987 62437 26993
rect 62652 26984 62658 26996
rect 62710 26984 62716 27036
rect 63296 26984 63302 27036
rect 63354 27024 63360 27036
rect 63759 27027 63817 27033
rect 63759 27024 63771 27027
rect 63354 26996 63771 27024
rect 63354 26984 63360 26996
rect 63759 26993 63771 26996
rect 63805 26993 63817 27027
rect 63759 26987 63817 26993
rect 64124 26984 64130 27036
rect 64182 27024 64188 27036
rect 65691 27027 65749 27033
rect 65691 27024 65703 27027
rect 64182 26996 65703 27024
rect 64182 26984 64188 26996
rect 65691 26993 65703 26996
rect 65737 26993 65749 27027
rect 65691 26987 65749 26993
rect 53639 26959 53697 26965
rect 53639 26956 53651 26959
rect 51262 26928 52486 26956
rect 52550 26928 53651 26956
rect 51155 26919 51213 26925
rect 49729 26860 49818 26888
rect 49882 26860 50370 26888
rect 49729 26857 49741 26860
rect 49683 26851 49741 26857
rect 31022 26792 31602 26820
rect 32939 26823 32997 26829
rect 29305 26789 29317 26792
rect 29259 26783 29317 26789
rect 32939 26789 32951 26823
rect 32985 26820 32997 26823
rect 34408 26820 34414 26832
rect 32985 26792 34414 26820
rect 32985 26789 32997 26792
rect 32939 26783 32997 26789
rect 34408 26780 34414 26792
rect 34466 26780 34472 26832
rect 49790 26820 49818 26860
rect 50434 26832 50462 26916
rect 52458 26888 52486 26928
rect 53639 26925 53651 26928
rect 53685 26925 53697 26959
rect 53639 26919 53697 26925
rect 56856 26916 56862 26968
rect 56914 26956 56920 26968
rect 57043 26959 57101 26965
rect 57043 26956 57055 26959
rect 56914 26928 57055 26956
rect 56914 26916 56920 26928
rect 57043 26925 57055 26928
rect 57089 26925 57101 26959
rect 57043 26919 57101 26925
rect 65047 26959 65105 26965
rect 65047 26925 65059 26959
rect 65093 26925 65105 26959
rect 65412 26956 65418 26968
rect 65373 26928 65418 26956
rect 65047 26919 65105 26925
rect 53452 26888 53458 26900
rect 52458 26860 53458 26888
rect 53452 26848 53458 26860
rect 53510 26888 53516 26900
rect 53731 26891 53789 26897
rect 53731 26888 53743 26891
rect 53510 26860 53743 26888
rect 53510 26848 53516 26860
rect 53731 26857 53743 26860
rect 53777 26857 53789 26891
rect 65062 26888 65090 26919
rect 65412 26916 65418 26928
rect 65470 26916 65476 26968
rect 66166 26888 66194 27052
rect 67988 27024 67994 27036
rect 67949 26996 67994 27024
rect 67988 26984 67994 26996
rect 68046 26984 68052 27036
rect 68264 27024 68270 27036
rect 68225 26996 68270 27024
rect 68264 26984 68270 26996
rect 68322 26984 68328 27036
rect 68448 26984 68454 27036
rect 68506 27024 68512 27036
rect 69739 27027 69797 27033
rect 69739 27024 69751 27027
rect 68506 26996 69751 27024
rect 68506 26984 68512 26996
rect 69739 26993 69751 26996
rect 69785 26993 69797 27027
rect 70104 27024 70110 27036
rect 70065 26996 70110 27024
rect 69739 26987 69797 26993
rect 70104 26984 70110 26996
rect 70162 26984 70168 27036
rect 71671 27027 71729 27033
rect 71671 26993 71683 27027
rect 71717 27024 71729 27027
rect 72312 27024 72318 27036
rect 71717 26996 72318 27024
rect 71717 26993 71729 26996
rect 71671 26987 71729 26993
rect 72312 26984 72318 26996
rect 72370 26984 72376 27036
rect 68356 26916 68362 26968
rect 68414 26956 68420 26968
rect 70659 26959 70717 26965
rect 70659 26956 70671 26959
rect 68414 26928 70671 26956
rect 68414 26916 68420 26928
rect 70659 26925 70671 26928
rect 70705 26925 70717 26959
rect 70659 26919 70717 26925
rect 72223 26959 72281 26965
rect 72223 26925 72235 26959
rect 72269 26956 72281 26959
rect 72422 26956 72450 27064
rect 73695 27061 73707 27064
rect 73741 27061 73753 27095
rect 75624 27092 75630 27104
rect 73695 27055 73753 27061
rect 73802 27064 74566 27092
rect 75585 27064 75630 27092
rect 73600 27024 73606 27036
rect 72514 26996 73606 27024
rect 72514 26965 72542 26996
rect 73600 26984 73606 26996
rect 73658 26984 73664 27036
rect 72269 26928 72450 26956
rect 72499 26959 72557 26965
rect 72269 26925 72281 26928
rect 72223 26919 72281 26925
rect 72499 26925 72511 26959
rect 72545 26925 72557 26959
rect 72499 26919 72557 26925
rect 72683 26959 72741 26965
rect 72683 26925 72695 26959
rect 72729 26956 72741 26959
rect 73051 26959 73109 26965
rect 73051 26956 73063 26959
rect 72729 26928 73063 26956
rect 72729 26925 72741 26928
rect 72683 26919 72741 26925
rect 73051 26925 73063 26928
rect 73097 26925 73109 26959
rect 73324 26956 73330 26968
rect 73237 26928 73330 26956
rect 73051 26919 73109 26925
rect 65062 26860 66194 26888
rect 53731 26851 53789 26857
rect 70012 26848 70018 26900
rect 70070 26888 70076 26900
rect 70291 26891 70349 26897
rect 70291 26888 70303 26891
rect 70070 26860 70303 26888
rect 70070 26848 70076 26860
rect 70291 26857 70303 26860
rect 70337 26857 70349 26891
rect 70291 26851 70349 26857
rect 70567 26891 70625 26897
rect 70567 26857 70579 26891
rect 70613 26888 70625 26891
rect 70840 26888 70846 26900
rect 70613 26860 70846 26888
rect 70613 26857 70625 26860
rect 70567 26851 70625 26857
rect 70840 26848 70846 26860
rect 70898 26848 70904 26900
rect 70932 26848 70938 26900
rect 70990 26888 70996 26900
rect 71208 26888 71214 26900
rect 70990 26860 71035 26888
rect 71169 26860 71214 26888
rect 70990 26848 70996 26860
rect 71208 26848 71214 26860
rect 71266 26848 71272 26900
rect 71300 26848 71306 26900
rect 71358 26888 71364 26900
rect 71484 26888 71490 26900
rect 71358 26860 71403 26888
rect 71445 26860 71490 26888
rect 71358 26848 71364 26860
rect 71484 26848 71490 26860
rect 71542 26848 71548 26900
rect 71944 26848 71950 26900
rect 72002 26888 72008 26900
rect 72698 26888 72726 26919
rect 72002 26860 72726 26888
rect 73066 26888 73094 26919
rect 73324 26916 73330 26928
rect 73382 26956 73388 26968
rect 73802 26965 73830 27064
rect 74431 27027 74489 27033
rect 74431 27024 74443 27027
rect 73986 26996 74443 27024
rect 73787 26959 73845 26965
rect 73787 26956 73799 26959
rect 73382 26928 73799 26956
rect 73382 26916 73388 26928
rect 73787 26925 73799 26928
rect 73833 26925 73845 26959
rect 73787 26919 73845 26925
rect 73876 26916 73882 26968
rect 73934 26956 73940 26968
rect 73986 26956 74014 26996
rect 74431 26993 74443 26996
rect 74477 26993 74489 27027
rect 74431 26987 74489 26993
rect 73934 26928 74014 26956
rect 74155 26959 74213 26965
rect 73934 26916 73940 26928
rect 74155 26925 74167 26959
rect 74201 26925 74213 26959
rect 74155 26919 74213 26925
rect 74170 26888 74198 26919
rect 73066 26860 74198 26888
rect 74538 26888 74566 27064
rect 75624 27052 75630 27064
rect 75682 27052 75688 27104
rect 79031 27095 79089 27101
rect 79031 27061 79043 27095
rect 79077 27092 79089 27095
rect 79212 27092 79218 27104
rect 79077 27064 79218 27092
rect 79077 27061 79089 27064
rect 79031 27055 79089 27061
rect 79212 27052 79218 27064
rect 79270 27052 79276 27104
rect 87676 27092 87682 27104
rect 87637 27064 87682 27092
rect 87676 27052 87682 27064
rect 87734 27052 87740 27104
rect 78203 27027 78261 27033
rect 78203 26993 78215 27027
rect 78249 27024 78261 27027
rect 79491 27027 79549 27033
rect 79491 27024 79503 27027
rect 78249 26996 79503 27024
rect 78249 26993 78261 26996
rect 78203 26987 78261 26993
rect 79491 26993 79503 26996
rect 79537 26993 79549 27027
rect 79491 26987 79549 26993
rect 80595 27027 80653 27033
rect 80595 26993 80607 27027
rect 80641 26993 80653 27027
rect 80595 26987 80653 26993
rect 85379 27027 85437 27033
rect 85379 26993 85391 27027
rect 85425 27024 85437 27027
rect 85744 27024 85750 27036
rect 85425 26996 85750 27024
rect 85425 26993 85437 26996
rect 85379 26987 85437 26993
rect 75532 26956 75538 26968
rect 75493 26928 75538 26956
rect 75532 26916 75538 26928
rect 75590 26916 75596 26968
rect 78111 26959 78169 26965
rect 78111 26925 78123 26959
rect 78157 26956 78169 26959
rect 79028 26956 79034 26968
rect 78157 26928 79034 26956
rect 78157 26925 78169 26928
rect 78111 26919 78169 26925
rect 79028 26916 79034 26928
rect 79086 26916 79092 26968
rect 79212 26956 79218 26968
rect 79173 26928 79218 26956
rect 79212 26916 79218 26928
rect 79270 26916 79276 26968
rect 80610 26956 80638 26987
rect 85744 26984 85750 26996
rect 85802 26984 85808 27036
rect 86572 27024 86578 27036
rect 86533 26996 86578 27024
rect 86572 26984 86578 26996
rect 86630 26984 86636 27036
rect 89332 26984 89338 27036
rect 89390 27024 89396 27036
rect 90715 27027 90773 27033
rect 90715 27024 90727 27027
rect 89390 26996 90727 27024
rect 89390 26984 89396 26996
rect 90715 26993 90727 26996
rect 90761 26993 90773 27027
rect 90715 26987 90773 26993
rect 79322 26928 80638 26956
rect 74538 26860 78522 26888
rect 72002 26848 72008 26860
rect 50324 26820 50330 26832
rect 49790 26792 50330 26820
rect 50324 26780 50330 26792
rect 50382 26780 50388 26832
rect 50416 26780 50422 26832
rect 50474 26780 50480 26832
rect 69920 26820 69926 26832
rect 69881 26792 69926 26820
rect 69920 26780 69926 26792
rect 69978 26780 69984 26832
rect 78494 26820 78522 26860
rect 78660 26848 78666 26900
rect 78718 26888 78724 26900
rect 79322 26888 79350 26928
rect 84088 26916 84094 26968
rect 84146 26956 84152 26968
rect 85011 26959 85069 26965
rect 85011 26956 85023 26959
rect 84146 26928 85023 26956
rect 84146 26916 84152 26928
rect 85011 26925 85023 26928
rect 85057 26956 85069 26959
rect 85471 26959 85529 26965
rect 85471 26956 85483 26959
rect 85057 26928 85483 26956
rect 85057 26925 85069 26928
rect 85011 26919 85069 26925
rect 85471 26925 85483 26928
rect 85517 26925 85529 26959
rect 85471 26919 85529 26925
rect 85560 26916 85566 26968
rect 85618 26956 85624 26968
rect 86207 26959 86265 26965
rect 86207 26956 86219 26959
rect 85618 26928 86219 26956
rect 85618 26916 85624 26928
rect 86207 26925 86219 26928
rect 86253 26956 86265 26959
rect 86299 26959 86357 26965
rect 86299 26956 86311 26959
rect 86253 26928 86311 26956
rect 86253 26925 86265 26928
rect 86207 26919 86265 26925
rect 86299 26925 86311 26928
rect 86345 26956 86357 26959
rect 90255 26959 90313 26965
rect 90255 26956 90267 26959
rect 86345 26928 90267 26956
rect 86345 26925 86357 26928
rect 86299 26919 86357 26925
rect 90255 26925 90267 26928
rect 90301 26956 90313 26959
rect 90436 26956 90442 26968
rect 90301 26928 90442 26956
rect 90301 26925 90313 26928
rect 90255 26919 90313 26925
rect 90436 26916 90442 26928
rect 90494 26916 90500 26968
rect 92095 26959 92153 26965
rect 92095 26956 92107 26959
rect 90546 26928 92107 26956
rect 80500 26888 80506 26900
rect 78718 26860 79350 26888
rect 80150 26860 80506 26888
rect 78718 26848 78724 26860
rect 80150 26820 80178 26860
rect 80500 26848 80506 26860
rect 80558 26848 80564 26900
rect 84824 26888 84830 26900
rect 84785 26860 84830 26888
rect 84824 26848 84830 26860
rect 84882 26848 84888 26900
rect 89608 26848 89614 26900
rect 89666 26888 89672 26900
rect 90546 26888 90574 26928
rect 92095 26925 92107 26928
rect 92141 26925 92153 26959
rect 92095 26919 92153 26925
rect 89666 26860 90574 26888
rect 89666 26848 89672 26860
rect 78494 26792 80178 26820
rect 538 26730 93642 26752
rect 538 26678 6344 26730
rect 6396 26678 6408 26730
rect 6460 26678 6472 26730
rect 6524 26678 6536 26730
rect 6588 26678 11672 26730
rect 11724 26678 11736 26730
rect 11788 26678 11800 26730
rect 11852 26678 11864 26730
rect 11916 26678 17000 26730
rect 17052 26678 17064 26730
rect 17116 26678 17128 26730
rect 17180 26678 17192 26730
rect 17244 26678 22328 26730
rect 22380 26678 22392 26730
rect 22444 26678 22456 26730
rect 22508 26678 22520 26730
rect 22572 26678 27656 26730
rect 27708 26678 27720 26730
rect 27772 26678 27784 26730
rect 27836 26678 27848 26730
rect 27900 26678 32984 26730
rect 33036 26678 33048 26730
rect 33100 26678 33112 26730
rect 33164 26678 33176 26730
rect 33228 26678 38312 26730
rect 38364 26678 38376 26730
rect 38428 26678 38440 26730
rect 38492 26678 38504 26730
rect 38556 26678 43640 26730
rect 43692 26678 43704 26730
rect 43756 26678 43768 26730
rect 43820 26678 43832 26730
rect 43884 26678 48968 26730
rect 49020 26678 49032 26730
rect 49084 26678 49096 26730
rect 49148 26678 49160 26730
rect 49212 26678 54296 26730
rect 54348 26678 54360 26730
rect 54412 26678 54424 26730
rect 54476 26678 54488 26730
rect 54540 26678 59624 26730
rect 59676 26678 59688 26730
rect 59740 26678 59752 26730
rect 59804 26678 59816 26730
rect 59868 26678 64952 26730
rect 65004 26678 65016 26730
rect 65068 26678 65080 26730
rect 65132 26678 65144 26730
rect 65196 26678 70280 26730
rect 70332 26678 70344 26730
rect 70396 26678 70408 26730
rect 70460 26678 70472 26730
rect 70524 26678 75608 26730
rect 75660 26678 75672 26730
rect 75724 26678 75736 26730
rect 75788 26678 75800 26730
rect 75852 26678 80936 26730
rect 80988 26678 81000 26730
rect 81052 26678 81064 26730
rect 81116 26678 81128 26730
rect 81180 26678 86264 26730
rect 86316 26678 86328 26730
rect 86380 26678 86392 26730
rect 86444 26678 86456 26730
rect 86508 26678 91592 26730
rect 91644 26678 91656 26730
rect 91708 26678 91720 26730
rect 91772 26678 91784 26730
rect 91836 26678 93642 26730
rect 538 26656 93642 26678
rect 3956 26616 3962 26628
rect 3917 26588 3962 26616
rect 3956 26576 3962 26588
rect 4014 26576 4020 26628
rect 5520 26616 5526 26628
rect 5433 26588 5526 26616
rect 5520 26576 5526 26588
rect 5578 26616 5584 26628
rect 6164 26616 6170 26628
rect 5578 26588 6170 26616
rect 5578 26576 5584 26588
rect 6164 26576 6170 26588
rect 6222 26616 6228 26628
rect 7271 26619 7329 26625
rect 7271 26616 7283 26619
rect 6222 26588 7283 26616
rect 6222 26576 6228 26588
rect 7271 26585 7283 26588
rect 7317 26585 7329 26619
rect 7271 26579 7329 26585
rect 23644 26576 23650 26628
rect 23702 26616 23708 26628
rect 25392 26616 25398 26628
rect 23702 26588 25398 26616
rect 23702 26576 23708 26588
rect 25392 26576 25398 26588
rect 25450 26576 25456 26628
rect 38088 26616 38094 26628
rect 38049 26588 38094 26616
rect 38088 26576 38094 26588
rect 38146 26616 38152 26628
rect 38275 26619 38333 26625
rect 38275 26616 38287 26619
rect 38146 26588 38287 26616
rect 38146 26576 38152 26588
rect 38275 26585 38287 26588
rect 38321 26616 38333 26619
rect 39376 26616 39382 26628
rect 38321 26588 39382 26616
rect 38321 26585 38333 26588
rect 38275 26579 38333 26585
rect 39376 26576 39382 26588
rect 39434 26576 39440 26628
rect 3683 26483 3741 26489
rect 3683 26449 3695 26483
rect 3729 26480 3741 26483
rect 3974 26480 4002 26576
rect 5538 26489 5566 26576
rect 31372 26508 31378 26560
rect 31430 26548 31436 26560
rect 37171 26551 37229 26557
rect 37171 26548 37183 26551
rect 31430 26520 35374 26548
rect 31430 26508 31436 26520
rect 3729 26452 4002 26480
rect 5523 26483 5581 26489
rect 3729 26449 3741 26452
rect 3683 26443 3741 26449
rect 5523 26449 5535 26483
rect 5569 26449 5581 26483
rect 5523 26443 5581 26449
rect 34132 26440 34138 26492
rect 34190 26480 34196 26492
rect 35346 26489 35374 26520
rect 35898 26520 37183 26548
rect 35898 26489 35926 26520
rect 37171 26517 37183 26520
rect 37217 26548 37229 26551
rect 42872 26548 42878 26560
rect 37217 26520 42878 26548
rect 37217 26517 37229 26520
rect 37171 26511 37229 26517
rect 42872 26508 42878 26520
rect 42930 26508 42936 26560
rect 34411 26483 34469 26489
rect 34411 26480 34423 26483
rect 34190 26452 34423 26480
rect 34190 26440 34196 26452
rect 34411 26449 34423 26452
rect 34457 26449 34469 26483
rect 34411 26443 34469 26449
rect 34595 26483 34653 26489
rect 34595 26449 34607 26483
rect 34641 26480 34653 26483
rect 35147 26483 35205 26489
rect 35147 26480 35159 26483
rect 34641 26452 35159 26480
rect 34641 26449 34653 26452
rect 34595 26443 34653 26449
rect 35147 26449 35159 26452
rect 35193 26449 35205 26483
rect 35147 26443 35205 26449
rect 35331 26483 35389 26489
rect 35331 26449 35343 26483
rect 35377 26480 35389 26483
rect 35883 26483 35941 26489
rect 35883 26480 35895 26483
rect 35377 26452 35895 26480
rect 35377 26449 35389 26452
rect 35331 26443 35389 26449
rect 35883 26449 35895 26452
rect 35929 26449 35941 26483
rect 35883 26443 35941 26449
rect 5796 26412 5802 26424
rect 5757 26384 5802 26412
rect 5796 26372 5802 26384
rect 5854 26372 5860 26424
rect 33948 26372 33954 26424
rect 34006 26412 34012 26424
rect 34610 26412 34638 26443
rect 35972 26440 35978 26492
rect 36030 26480 36036 26492
rect 37079 26483 37137 26489
rect 37079 26480 37091 26483
rect 36030 26452 37091 26480
rect 36030 26440 36036 26452
rect 37079 26449 37091 26452
rect 37125 26449 37137 26483
rect 37079 26443 37137 26449
rect 38088 26440 38094 26492
rect 38146 26480 38152 26492
rect 38827 26483 38885 26489
rect 38827 26480 38839 26483
rect 38146 26452 38839 26480
rect 38146 26440 38152 26452
rect 38827 26449 38839 26452
rect 38873 26449 38885 26483
rect 39284 26480 39290 26492
rect 39245 26452 39290 26480
rect 38827 26443 38885 26449
rect 39284 26440 39290 26452
rect 39342 26440 39348 26492
rect 39376 26440 39382 26492
rect 39434 26480 39440 26492
rect 39434 26452 39479 26480
rect 39434 26440 39440 26452
rect 38548 26412 38554 26424
rect 34006 26384 34638 26412
rect 38461 26384 38554 26412
rect 34006 26372 34012 26384
rect 38548 26372 38554 26384
rect 38606 26412 38612 26424
rect 38643 26415 38701 26421
rect 38643 26412 38655 26415
rect 38606 26384 38655 26412
rect 38606 26372 38612 26384
rect 38643 26381 38655 26384
rect 38689 26381 38701 26415
rect 38643 26375 38701 26381
rect 6624 26304 6630 26356
rect 6682 26344 6688 26356
rect 7087 26347 7145 26353
rect 7087 26344 7099 26347
rect 6682 26316 7099 26344
rect 6682 26304 6688 26316
rect 7087 26313 7099 26316
rect 7133 26344 7145 26347
rect 11500 26344 11506 26356
rect 7133 26316 11506 26344
rect 7133 26313 7145 26316
rect 7087 26307 7145 26313
rect 11500 26304 11506 26316
rect 11558 26344 11564 26356
rect 11558 26316 67114 26344
rect 11558 26304 11564 26316
rect 67086 26288 67114 26316
rect 3496 26236 3502 26288
rect 3554 26276 3560 26288
rect 3775 26279 3833 26285
rect 3775 26276 3787 26279
rect 3554 26248 3787 26276
rect 3554 26236 3560 26248
rect 3775 26245 3787 26248
rect 3821 26245 3833 26279
rect 3775 26239 3833 26245
rect 34684 26236 34690 26288
rect 34742 26276 34748 26288
rect 35607 26279 35665 26285
rect 35607 26276 35619 26279
rect 34742 26248 35619 26276
rect 34742 26236 34748 26248
rect 35607 26245 35619 26248
rect 35653 26245 35665 26279
rect 35607 26239 35665 26245
rect 36800 26236 36806 26288
rect 36858 26276 36864 26288
rect 37720 26276 37726 26288
rect 36858 26248 37726 26276
rect 36858 26236 36864 26248
rect 37720 26236 37726 26248
rect 37778 26276 37784 26288
rect 38548 26276 38554 26288
rect 37778 26248 38554 26276
rect 37778 26236 37784 26248
rect 38548 26236 38554 26248
rect 38606 26236 38612 26288
rect 39839 26279 39897 26285
rect 39839 26245 39851 26279
rect 39885 26276 39897 26279
rect 40848 26276 40854 26288
rect 39885 26248 40854 26276
rect 39885 26245 39897 26248
rect 39839 26239 39897 26245
rect 40848 26236 40854 26248
rect 40906 26236 40912 26288
rect 67068 26236 67074 26288
rect 67126 26276 67132 26288
rect 69920 26276 69926 26288
rect 67126 26248 69926 26276
rect 67126 26236 67132 26248
rect 69920 26236 69926 26248
rect 69978 26236 69984 26288
rect 538 26186 8450 26208
rect 538 26134 3680 26186
rect 3732 26134 3744 26186
rect 3796 26134 3808 26186
rect 3860 26134 3872 26186
rect 3924 26134 8450 26186
rect 538 26112 8450 26134
rect 34118 26186 43410 26208
rect 34118 26134 35648 26186
rect 35700 26134 35712 26186
rect 35764 26134 35776 26186
rect 35828 26134 35840 26186
rect 35892 26134 40976 26186
rect 41028 26134 41040 26186
rect 41092 26134 41104 26186
rect 41156 26134 41168 26186
rect 41220 26134 43410 26186
rect 34118 26112 43410 26134
rect 3867 26075 3925 26081
rect 3867 26041 3879 26075
rect 3913 26072 3925 26075
rect 4048 26072 4054 26084
rect 3913 26044 4054 26072
rect 3913 26041 3925 26044
rect 3867 26035 3925 26041
rect 4048 26032 4054 26044
rect 4106 26032 4112 26084
rect 6624 26072 6630 26084
rect 6585 26044 6630 26072
rect 6624 26032 6630 26044
rect 6682 26032 6688 26084
rect 35972 26072 35978 26084
rect 35933 26044 35978 26072
rect 35972 26032 35978 26044
rect 36030 26032 36036 26084
rect 36524 26032 36530 26084
rect 36582 26072 36588 26084
rect 36711 26075 36769 26081
rect 36711 26072 36723 26075
rect 36582 26044 36723 26072
rect 36582 26032 36588 26044
rect 36711 26041 36723 26044
rect 36757 26041 36769 26075
rect 36711 26035 36769 26041
rect 4232 26004 4238 26016
rect 2962 25976 4238 26004
rect 2579 25939 2637 25945
rect 2579 25905 2591 25939
rect 2625 25936 2637 25939
rect 2962 25936 2990 25976
rect 4232 25964 4238 25976
rect 4290 26004 4296 26016
rect 4508 26004 4514 26016
rect 4290 25976 4514 26004
rect 4290 25964 4296 25976
rect 4508 25964 4514 25976
rect 4566 25964 4572 26016
rect 2625 25908 2990 25936
rect 2625 25905 2637 25908
rect 2579 25899 2637 25905
rect 2760 25828 2766 25880
rect 2818 25868 2824 25880
rect 2962 25877 2990 25908
rect 2855 25871 2913 25877
rect 2855 25868 2867 25871
rect 2818 25840 2867 25868
rect 2818 25828 2824 25840
rect 2855 25837 2867 25840
rect 2901 25837 2913 25871
rect 2855 25831 2913 25837
rect 2947 25871 3005 25877
rect 2947 25837 2959 25871
rect 2993 25837 3005 25871
rect 2947 25831 3005 25837
rect 3407 25871 3465 25877
rect 3407 25837 3419 25871
rect 3453 25837 3465 25871
rect 3407 25831 3465 25837
rect 2870 25800 2898 25831
rect 3422 25800 3450 25831
rect 3496 25828 3502 25880
rect 3554 25868 3560 25880
rect 3591 25871 3649 25877
rect 3591 25868 3603 25871
rect 3554 25840 3603 25868
rect 3554 25828 3560 25840
rect 3591 25837 3603 25840
rect 3637 25837 3649 25871
rect 3591 25831 3649 25837
rect 6259 25871 6317 25877
rect 6259 25837 6271 25871
rect 6305 25868 6317 25871
rect 6642 25868 6670 26032
rect 36726 26004 36754 26035
rect 39284 26032 39290 26084
rect 39342 26072 39348 26084
rect 42047 26075 42105 26081
rect 42047 26072 42059 26075
rect 39342 26044 42059 26072
rect 39342 26032 39348 26044
rect 42047 26041 42059 26044
rect 42093 26041 42105 26075
rect 42047 26035 42105 26041
rect 36726 25976 37950 26004
rect 31832 25896 31838 25948
rect 31890 25936 31896 25948
rect 34684 25936 34690 25948
rect 31890 25908 34546 25936
rect 34645 25908 34690 25936
rect 31890 25896 31896 25908
rect 34408 25868 34414 25880
rect 6305 25840 6670 25868
rect 34369 25840 34414 25868
rect 6305 25837 6317 25840
rect 6259 25831 6317 25837
rect 34408 25828 34414 25840
rect 34466 25828 34472 25880
rect 34518 25868 34546 25908
rect 34684 25896 34690 25908
rect 34742 25896 34748 25948
rect 36619 25939 36677 25945
rect 36619 25905 36631 25939
rect 36665 25936 36677 25939
rect 36708 25936 36714 25948
rect 36665 25908 36714 25936
rect 36665 25905 36677 25908
rect 36619 25899 36677 25905
rect 36708 25896 36714 25908
rect 36766 25936 36772 25948
rect 36766 25908 37582 25936
rect 36766 25896 36772 25908
rect 37554 25877 37582 25908
rect 37922 25877 37950 25976
rect 42504 25936 42510 25948
rect 40958 25908 42510 25936
rect 40958 25877 40986 25908
rect 42504 25896 42510 25908
rect 42562 25896 42568 25948
rect 36895 25871 36953 25877
rect 36895 25868 36907 25871
rect 34518 25840 36907 25868
rect 36895 25837 36907 25840
rect 36941 25837 36953 25871
rect 37355 25871 37413 25877
rect 37355 25868 37367 25871
rect 36895 25831 36953 25837
rect 37094 25840 37367 25868
rect 2870 25772 3450 25800
rect 6351 25803 6409 25809
rect 6351 25769 6363 25803
rect 6397 25800 6409 25803
rect 6624 25800 6630 25812
rect 6397 25772 6630 25800
rect 6397 25769 6409 25772
rect 6351 25763 6409 25769
rect 6624 25760 6630 25772
rect 6682 25760 6688 25812
rect 37094 25732 37122 25840
rect 37355 25837 37367 25840
rect 37401 25837 37413 25871
rect 37355 25831 37413 25837
rect 37539 25871 37597 25877
rect 37539 25837 37551 25871
rect 37585 25837 37597 25871
rect 37539 25831 37597 25837
rect 37907 25871 37965 25877
rect 37907 25837 37919 25871
rect 37953 25837 37965 25871
rect 37907 25831 37965 25837
rect 37999 25871 38057 25877
rect 37999 25837 38011 25871
rect 38045 25837 38057 25871
rect 37999 25831 38057 25837
rect 40943 25871 41001 25877
rect 40943 25837 40955 25871
rect 40989 25837 41001 25871
rect 40943 25831 41001 25837
rect 41955 25871 42013 25877
rect 41955 25837 41967 25871
rect 42001 25868 42013 25871
rect 42228 25868 42234 25880
rect 42001 25840 42234 25868
rect 42001 25837 42013 25840
rect 41955 25831 42013 25837
rect 37168 25760 37174 25812
rect 37226 25800 37232 25812
rect 38014 25800 38042 25831
rect 42228 25828 42234 25840
rect 42286 25828 42292 25880
rect 37226 25772 38042 25800
rect 37226 25760 37232 25772
rect 38824 25732 38830 25744
rect 37094 25704 38830 25732
rect 38824 25692 38830 25704
rect 38882 25732 38888 25744
rect 41035 25735 41093 25741
rect 41035 25732 41047 25735
rect 38882 25704 41047 25732
rect 38882 25692 38888 25704
rect 41035 25701 41047 25704
rect 41081 25701 41093 25735
rect 41035 25695 41093 25701
rect 538 25642 8450 25664
rect 538 25590 6344 25642
rect 6396 25590 6408 25642
rect 6460 25590 6472 25642
rect 6524 25590 6536 25642
rect 6588 25590 8450 25642
rect 538 25568 8450 25590
rect 34118 25642 43410 25664
rect 34118 25590 38312 25642
rect 38364 25590 38376 25642
rect 38428 25590 38440 25642
rect 38492 25590 38504 25642
rect 38556 25590 43410 25642
rect 34118 25568 43410 25590
rect 16744 25488 16750 25540
rect 16802 25528 16808 25540
rect 70196 25528 70202 25540
rect 16802 25500 70202 25528
rect 16802 25488 16808 25500
rect 70196 25488 70202 25500
rect 70254 25488 70260 25540
rect 2760 25420 2766 25472
rect 2818 25460 2824 25472
rect 4232 25460 4238 25472
rect 2818 25432 4238 25460
rect 2818 25420 2824 25432
rect 4232 25420 4238 25432
rect 4290 25460 4296 25472
rect 5796 25460 5802 25472
rect 4290 25432 4738 25460
rect 5757 25432 5802 25460
rect 4290 25420 4296 25432
rect 4710 25401 4738 25432
rect 5796 25420 5802 25432
rect 5854 25420 5860 25472
rect 34408 25460 34414 25472
rect 34369 25432 34414 25460
rect 34408 25420 34414 25432
rect 34466 25460 34472 25472
rect 36800 25460 36806 25472
rect 34466 25432 36806 25460
rect 34466 25420 34472 25432
rect 36800 25420 36806 25432
rect 36858 25460 36864 25472
rect 39931 25463 39989 25469
rect 39931 25460 39943 25463
rect 36858 25432 39943 25460
rect 36858 25420 36864 25432
rect 39931 25429 39943 25432
rect 39977 25460 39989 25463
rect 41771 25463 41829 25469
rect 39977 25432 40158 25460
rect 39977 25429 39989 25432
rect 39931 25423 39989 25429
rect 3499 25395 3557 25401
rect 3499 25361 3511 25395
rect 3545 25361 3557 25395
rect 3499 25355 3557 25361
rect 4695 25395 4753 25401
rect 4695 25361 4707 25395
rect 4741 25392 4753 25395
rect 5247 25395 5305 25401
rect 5247 25392 5259 25395
rect 4741 25364 5259 25392
rect 4741 25361 4753 25364
rect 4695 25355 4753 25361
rect 5247 25361 5259 25364
rect 5293 25361 5305 25395
rect 5247 25355 5305 25361
rect 5431 25395 5489 25401
rect 5431 25361 5443 25395
rect 5477 25392 5489 25395
rect 6624 25392 6630 25404
rect 5477 25364 6630 25392
rect 5477 25361 5489 25364
rect 5431 25355 5489 25361
rect 3514 25188 3542 25355
rect 6624 25352 6630 25364
rect 6682 25352 6688 25404
rect 37447 25395 37505 25401
rect 37447 25361 37459 25395
rect 37493 25392 37505 25395
rect 37631 25395 37689 25401
rect 37631 25392 37643 25395
rect 37493 25364 37643 25392
rect 37493 25361 37505 25364
rect 37447 25355 37505 25361
rect 37631 25361 37643 25364
rect 37677 25392 37689 25395
rect 38088 25392 38094 25404
rect 37677 25364 38094 25392
rect 37677 25361 37689 25364
rect 37631 25355 37689 25361
rect 38088 25352 38094 25364
rect 38146 25392 38152 25404
rect 38643 25395 38701 25401
rect 38643 25392 38655 25395
rect 38146 25364 38655 25392
rect 38146 25352 38152 25364
rect 38643 25361 38655 25364
rect 38689 25361 38701 25395
rect 38824 25392 38830 25404
rect 38785 25364 38830 25392
rect 38643 25355 38701 25361
rect 38824 25352 38830 25364
rect 38882 25352 38888 25404
rect 40130 25401 40158 25432
rect 41771 25429 41783 25463
rect 41817 25460 41829 25463
rect 42504 25460 42510 25472
rect 41817 25432 42510 25460
rect 41817 25429 41829 25432
rect 41771 25423 41829 25429
rect 42504 25420 42510 25432
rect 42562 25420 42568 25472
rect 40115 25395 40173 25401
rect 40115 25361 40127 25395
rect 40161 25361 40173 25395
rect 40115 25355 40173 25361
rect 4419 25327 4477 25333
rect 4419 25293 4431 25327
rect 4465 25324 4477 25327
rect 4600 25324 4606 25336
rect 4465 25296 4606 25324
rect 4465 25293 4477 25296
rect 4419 25287 4477 25293
rect 4600 25284 4606 25296
rect 4658 25284 4664 25336
rect 37536 25284 37542 25336
rect 37594 25324 37600 25336
rect 37723 25327 37781 25333
rect 37723 25324 37735 25327
rect 37594 25296 37735 25324
rect 37594 25284 37600 25296
rect 37723 25293 37735 25296
rect 37769 25324 37781 25327
rect 37907 25327 37965 25333
rect 37907 25324 37919 25327
rect 37769 25296 37919 25324
rect 37769 25293 37781 25296
rect 37723 25287 37781 25293
rect 37907 25293 37919 25296
rect 37953 25293 37965 25327
rect 37907 25287 37965 25293
rect 39195 25327 39253 25333
rect 39195 25293 39207 25327
rect 39241 25324 39253 25327
rect 40391 25327 40449 25333
rect 40391 25324 40403 25327
rect 39241 25296 40403 25324
rect 39241 25293 39253 25296
rect 39195 25287 39253 25293
rect 40391 25293 40403 25296
rect 40437 25293 40449 25327
rect 40391 25287 40449 25293
rect 3591 25259 3649 25265
rect 3591 25225 3603 25259
rect 3637 25256 3649 25259
rect 4140 25256 4146 25268
rect 3637 25228 4146 25256
rect 3637 25225 3649 25228
rect 3591 25219 3649 25225
rect 4140 25216 4146 25228
rect 4198 25216 4204 25268
rect 3867 25191 3925 25197
rect 3867 25188 3879 25191
rect 3514 25160 3879 25188
rect 3867 25157 3879 25160
rect 3913 25188 3925 25191
rect 4048 25188 4054 25200
rect 3913 25160 4054 25188
rect 3913 25157 3925 25160
rect 3867 25151 3925 25157
rect 4048 25148 4054 25160
rect 4106 25148 4112 25200
rect 23828 25148 23834 25200
rect 23886 25188 23892 25200
rect 39284 25188 39290 25200
rect 23886 25160 39290 25188
rect 23886 25148 23892 25160
rect 39284 25148 39290 25160
rect 39342 25148 39348 25200
rect 538 25098 8450 25120
rect 538 25046 3680 25098
rect 3732 25046 3744 25098
rect 3796 25046 3808 25098
rect 3860 25046 3872 25098
rect 3924 25046 8450 25098
rect 538 25024 8450 25046
rect 34118 25098 43410 25120
rect 34118 25046 35648 25098
rect 35700 25046 35712 25098
rect 35764 25046 35776 25098
rect 35828 25046 35840 25098
rect 35892 25046 40976 25098
rect 41028 25046 41040 25098
rect 41092 25046 41104 25098
rect 41156 25046 41168 25098
rect 41220 25046 43410 25098
rect 34118 25024 43410 25046
rect 1843 24987 1901 24993
rect 1843 24953 1855 24987
rect 1889 24984 1901 24987
rect 2760 24984 2766 24996
rect 1889 24956 2766 24984
rect 1889 24953 1901 24956
rect 1843 24947 1901 24953
rect 2760 24944 2766 24956
rect 2818 24944 2824 24996
rect 7084 24944 7090 24996
rect 7142 24984 7148 24996
rect 35144 24984 35150 24996
rect 7142 24956 7590 24984
rect 35105 24956 35150 24984
rect 7142 24944 7148 24956
rect 7562 24925 7590 24956
rect 35144 24944 35150 24956
rect 35202 24944 35208 24996
rect 42228 24984 42234 24996
rect 42189 24956 42234 24984
rect 42228 24944 42234 24956
rect 42286 24944 42292 24996
rect 7271 24919 7329 24925
rect 7271 24885 7283 24919
rect 7317 24885 7329 24919
rect 7271 24879 7329 24885
rect 7547 24919 7605 24925
rect 7547 24885 7559 24919
rect 7593 24916 7605 24919
rect 9019 24919 9077 24925
rect 9019 24916 9031 24919
rect 7593 24888 9031 24916
rect 7593 24885 7605 24888
rect 7547 24879 7605 24885
rect 9019 24885 9031 24888
rect 9065 24885 9077 24919
rect 9019 24879 9077 24885
rect 2763 24851 2821 24857
rect 2763 24817 2775 24851
rect 2809 24848 2821 24851
rect 3404 24848 3410 24860
rect 2809 24820 3410 24848
rect 2809 24817 2821 24820
rect 2763 24811 2821 24817
rect 3404 24808 3410 24820
rect 3462 24808 3468 24860
rect 5060 24808 5066 24860
rect 5118 24848 5124 24860
rect 7286 24848 7314 24879
rect 34868 24876 34874 24928
rect 34926 24916 34932 24928
rect 35975 24919 36033 24925
rect 35975 24916 35987 24919
rect 34926 24888 35987 24916
rect 34926 24876 34932 24888
rect 35975 24885 35987 24888
rect 36021 24916 36033 24919
rect 36021 24888 36202 24916
rect 36021 24885 36033 24888
rect 35975 24879 36033 24885
rect 36174 24857 36202 24888
rect 35607 24851 35665 24857
rect 35607 24848 35619 24851
rect 5118 24820 35619 24848
rect 5118 24808 5124 24820
rect 35607 24817 35619 24820
rect 35653 24848 35665 24851
rect 35791 24851 35849 24857
rect 35791 24848 35803 24851
rect 35653 24820 35803 24848
rect 35653 24817 35665 24820
rect 35607 24811 35665 24817
rect 35791 24817 35803 24820
rect 35837 24817 35849 24851
rect 35791 24811 35849 24817
rect 36159 24851 36217 24857
rect 36159 24817 36171 24851
rect 36205 24817 36217 24851
rect 36159 24811 36217 24817
rect 1659 24783 1717 24789
rect 1659 24749 1671 24783
rect 1705 24780 1717 24783
rect 3039 24783 3097 24789
rect 1705 24752 2162 24780
rect 1705 24749 1717 24752
rect 1659 24743 1717 24749
rect 2134 24653 2162 24752
rect 3039 24749 3051 24783
rect 3085 24780 3097 24783
rect 4692 24780 4698 24792
rect 3085 24752 4698 24780
rect 3085 24749 3097 24752
rect 3039 24743 3097 24749
rect 4692 24740 4698 24752
rect 4750 24740 4756 24792
rect 7084 24780 7090 24792
rect 7045 24752 7090 24780
rect 7084 24740 7090 24752
rect 7142 24740 7148 24792
rect 34408 24780 34414 24792
rect 21638 24752 34414 24780
rect 4048 24672 4054 24724
rect 4106 24712 4112 24724
rect 4419 24715 4477 24721
rect 4419 24712 4431 24715
rect 4106 24684 4431 24712
rect 4106 24672 4112 24684
rect 4419 24681 4431 24684
rect 4465 24712 4477 24715
rect 16744 24712 16750 24724
rect 4465 24684 16750 24712
rect 4465 24681 4477 24684
rect 4419 24675 4477 24681
rect 16744 24672 16750 24684
rect 16802 24672 16808 24724
rect 21531 24715 21589 24721
rect 21531 24681 21543 24715
rect 21577 24712 21589 24715
rect 21638 24712 21666 24752
rect 34408 24740 34414 24752
rect 34466 24740 34472 24792
rect 35331 24783 35389 24789
rect 35331 24749 35343 24783
rect 35377 24749 35389 24783
rect 35806 24780 35834 24811
rect 38180 24808 38186 24860
rect 38238 24848 38244 24860
rect 38824 24848 38830 24860
rect 38238 24820 38830 24848
rect 38238 24808 38244 24820
rect 38824 24808 38830 24820
rect 38882 24808 38888 24860
rect 40848 24808 40854 24860
rect 40906 24848 40912 24860
rect 40943 24851 41001 24857
rect 40943 24848 40955 24851
rect 40906 24820 40955 24848
rect 40906 24808 40912 24820
rect 40943 24817 40955 24820
rect 40989 24817 41001 24851
rect 40943 24811 41001 24817
rect 36343 24783 36401 24789
rect 36343 24780 36355 24783
rect 35806 24752 36355 24780
rect 35331 24743 35389 24749
rect 36343 24749 36355 24752
rect 36389 24780 36401 24783
rect 36892 24780 36898 24792
rect 36389 24752 36898 24780
rect 36389 24749 36401 24752
rect 36343 24743 36401 24749
rect 21577 24684 21666 24712
rect 21577 24681 21589 24684
rect 21531 24675 21589 24681
rect 25392 24672 25398 24724
rect 25450 24712 25456 24724
rect 34963 24715 35021 24721
rect 34963 24712 34975 24715
rect 25450 24684 34975 24712
rect 25450 24672 25456 24684
rect 34963 24681 34975 24684
rect 35009 24712 35021 24715
rect 35346 24712 35374 24743
rect 36892 24740 36898 24752
rect 36950 24740 36956 24792
rect 37076 24780 37082 24792
rect 37037 24752 37082 24780
rect 37076 24740 37082 24752
rect 37134 24740 37140 24792
rect 40667 24783 40725 24789
rect 40667 24780 40679 24783
rect 40498 24752 40679 24780
rect 35009 24684 35374 24712
rect 37447 24715 37505 24721
rect 35009 24681 35021 24684
rect 34963 24675 35021 24681
rect 37447 24681 37459 24715
rect 37493 24712 37505 24715
rect 38180 24712 38186 24724
rect 37493 24684 38186 24712
rect 37493 24681 37505 24684
rect 37447 24675 37505 24681
rect 38180 24672 38186 24684
rect 38238 24672 38244 24724
rect 2119 24647 2177 24653
rect 2119 24613 2131 24647
rect 2165 24644 2177 24647
rect 3680 24644 3686 24656
rect 2165 24616 3686 24644
rect 2165 24613 2177 24616
rect 2119 24607 2177 24613
rect 3680 24604 3686 24616
rect 3738 24604 3744 24656
rect 4603 24647 4661 24653
rect 4603 24613 4615 24647
rect 4649 24644 4661 24647
rect 6716 24644 6722 24656
rect 4649 24616 6722 24644
rect 4649 24613 4661 24616
rect 4603 24607 4661 24613
rect 6716 24604 6722 24616
rect 6774 24604 6780 24656
rect 9019 24647 9077 24653
rect 9019 24613 9031 24647
rect 9065 24644 9077 24647
rect 9844 24644 9850 24656
rect 9065 24616 9850 24644
rect 9065 24613 9077 24616
rect 9019 24607 9077 24613
rect 9844 24604 9850 24616
rect 9902 24644 9908 24656
rect 21439 24647 21497 24653
rect 21439 24644 21451 24647
rect 9902 24616 21451 24644
rect 9902 24604 9908 24616
rect 21439 24613 21451 24616
rect 21485 24613 21497 24647
rect 21439 24607 21497 24613
rect 36708 24604 36714 24656
rect 36766 24644 36772 24656
rect 40498 24653 40526 24752
rect 40667 24749 40679 24752
rect 40713 24749 40725 24783
rect 40667 24743 40725 24749
rect 40483 24647 40541 24653
rect 40483 24644 40495 24647
rect 36766 24616 40495 24644
rect 36766 24604 36772 24616
rect 40483 24613 40495 24616
rect 40529 24613 40541 24647
rect 40483 24607 40541 24613
rect 538 24554 8450 24576
rect 538 24502 6344 24554
rect 6396 24502 6408 24554
rect 6460 24502 6472 24554
rect 6524 24502 6536 24554
rect 6588 24502 8450 24554
rect 538 24480 8450 24502
rect 34118 24554 43410 24576
rect 34118 24502 38312 24554
rect 38364 24502 38376 24554
rect 38428 24502 38440 24554
rect 38492 24502 38504 24554
rect 38556 24502 43410 24554
rect 34118 24480 43410 24502
rect 4692 24440 4698 24452
rect 4653 24412 4698 24440
rect 4692 24400 4698 24412
rect 4750 24400 4756 24452
rect 4894 24412 7682 24440
rect 2484 24332 2490 24384
rect 2542 24372 2548 24384
rect 3315 24375 3373 24381
rect 3315 24372 3327 24375
rect 2542 24344 3327 24372
rect 2542 24332 2548 24344
rect 3315 24341 3327 24344
rect 3361 24372 3373 24375
rect 4894 24372 4922 24412
rect 5060 24372 5066 24384
rect 3361 24344 4922 24372
rect 5021 24344 5066 24372
rect 3361 24341 3373 24344
rect 3315 24335 3373 24341
rect 3680 24304 3686 24316
rect 3593 24276 3686 24304
rect 3680 24264 3686 24276
rect 3738 24264 3744 24316
rect 3790 24313 3818 24344
rect 5060 24332 5066 24344
rect 5118 24332 5124 24384
rect 7544 24372 7550 24384
rect 7505 24344 7550 24372
rect 7544 24332 7550 24344
rect 7602 24332 7608 24384
rect 7654 24372 7682 24412
rect 37076 24400 37082 24452
rect 37134 24440 37140 24452
rect 37171 24443 37229 24449
rect 37171 24440 37183 24443
rect 37134 24412 37183 24440
rect 37134 24400 37140 24412
rect 37171 24409 37183 24412
rect 37217 24409 37229 24443
rect 37171 24403 37229 24409
rect 15272 24372 15278 24384
rect 7654 24344 15278 24372
rect 15272 24332 15278 24344
rect 15330 24332 15336 24384
rect 3775 24307 3833 24313
rect 3775 24273 3787 24307
rect 3821 24273 3833 24307
rect 4140 24304 4146 24316
rect 4101 24276 4146 24304
rect 3775 24267 3833 24273
rect 4140 24264 4146 24276
rect 4198 24264 4204 24316
rect 4232 24264 4238 24316
rect 4290 24304 4296 24316
rect 4290 24276 4335 24304
rect 4290 24264 4296 24276
rect 3698 24168 3726 24264
rect 5078 24168 5106 24332
rect 5983 24307 6041 24313
rect 5983 24273 5995 24307
rect 6029 24304 6041 24307
rect 10672 24304 10678 24316
rect 6029 24276 10678 24304
rect 6029 24273 6041 24276
rect 5983 24267 6041 24273
rect 10672 24264 10678 24276
rect 10730 24264 10736 24316
rect 35144 24264 35150 24316
rect 35202 24304 35208 24316
rect 35331 24307 35389 24313
rect 35331 24304 35343 24307
rect 35202 24276 35343 24304
rect 35202 24264 35208 24276
rect 35331 24273 35343 24276
rect 35377 24273 35389 24307
rect 35331 24267 35389 24273
rect 36984 24264 36990 24316
rect 37042 24304 37048 24316
rect 37079 24307 37137 24313
rect 37079 24304 37091 24307
rect 37042 24276 37091 24304
rect 37042 24264 37048 24276
rect 37079 24273 37091 24276
rect 37125 24304 37137 24307
rect 37355 24307 37413 24313
rect 37355 24304 37367 24307
rect 37125 24276 37367 24304
rect 37125 24273 37137 24276
rect 37079 24267 37137 24273
rect 37355 24273 37367 24276
rect 37401 24304 37413 24307
rect 39468 24304 39474 24316
rect 37401 24276 39474 24304
rect 37401 24273 37413 24276
rect 37355 24267 37413 24273
rect 39468 24264 39474 24276
rect 39526 24264 39532 24316
rect 5707 24239 5765 24245
rect 5707 24205 5719 24239
rect 5753 24236 5765 24239
rect 6716 24236 6722 24248
rect 5753 24208 6722 24236
rect 5753 24205 5765 24208
rect 5707 24199 5765 24205
rect 6716 24196 6722 24208
rect 6774 24236 6780 24248
rect 7544 24236 7550 24248
rect 6774 24208 7550 24236
rect 6774 24196 6780 24208
rect 7544 24196 7550 24208
rect 7602 24196 7608 24248
rect 3698 24140 5106 24168
rect 35147 24171 35205 24177
rect 35147 24137 35159 24171
rect 35193 24168 35205 24171
rect 36708 24168 36714 24180
rect 35193 24140 36714 24168
rect 35193 24137 35205 24140
rect 35147 24131 35205 24137
rect 36708 24128 36714 24140
rect 36766 24128 36772 24180
rect 39468 24128 39474 24180
rect 39526 24168 39532 24180
rect 70012 24168 70018 24180
rect 39526 24140 70018 24168
rect 39526 24128 39532 24140
rect 70012 24128 70018 24140
rect 70070 24128 70076 24180
rect 7268 24100 7274 24112
rect 7229 24072 7274 24100
rect 7268 24060 7274 24072
rect 7326 24060 7332 24112
rect 30268 24100 30274 24112
rect 8482 24072 30274 24100
rect 538 24010 8450 24032
rect 538 23958 3680 24010
rect 3732 23958 3744 24010
rect 3796 23958 3808 24010
rect 3860 23958 3872 24010
rect 3924 23958 8450 24010
rect 538 23936 8450 23958
rect 7268 23856 7274 23908
rect 7326 23896 7332 23908
rect 7547 23899 7605 23905
rect 7547 23896 7559 23899
rect 7326 23868 7559 23896
rect 7326 23856 7332 23868
rect 7547 23865 7559 23868
rect 7593 23896 7605 23899
rect 8482 23896 8510 24072
rect 30268 24060 30274 24072
rect 30326 24060 30332 24112
rect 34118 24010 43410 24032
rect 34118 23958 35648 24010
rect 35700 23958 35712 24010
rect 35764 23958 35776 24010
rect 35828 23958 35840 24010
rect 35892 23958 40976 24010
rect 41028 23958 41040 24010
rect 41092 23958 41104 24010
rect 41156 23958 41168 24010
rect 41220 23958 43410 24010
rect 34118 23936 43410 23958
rect 33948 23896 33954 23908
rect 7593 23868 8510 23896
rect 8574 23868 33954 23896
rect 7593 23865 7605 23868
rect 7547 23859 7605 23865
rect 6900 23788 6906 23840
rect 6958 23828 6964 23840
rect 8574 23828 8602 23868
rect 33948 23856 33954 23868
rect 34006 23856 34012 23908
rect 34040 23856 34046 23908
rect 34098 23896 34104 23908
rect 34503 23899 34561 23905
rect 34503 23896 34515 23899
rect 34098 23868 34515 23896
rect 34098 23856 34104 23868
rect 34503 23865 34515 23868
rect 34549 23896 34561 23899
rect 34687 23899 34745 23905
rect 34687 23896 34699 23899
rect 34549 23868 34699 23896
rect 34549 23865 34561 23868
rect 34503 23859 34561 23865
rect 34687 23865 34699 23868
rect 34733 23865 34745 23899
rect 34868 23896 34874 23908
rect 34829 23868 34874 23896
rect 34687 23859 34745 23865
rect 6958 23800 8602 23828
rect 6958 23788 6964 23800
rect 2027 23763 2085 23769
rect 2027 23729 2039 23763
rect 2073 23760 2085 23763
rect 2073 23732 2438 23760
rect 2073 23729 2085 23732
rect 2027 23723 2085 23729
rect 2410 23701 2438 23732
rect 6624 23720 6630 23772
rect 6682 23760 6688 23772
rect 31372 23760 31378 23772
rect 6682 23732 31378 23760
rect 6682 23720 6688 23732
rect 31372 23720 31378 23732
rect 31430 23760 31436 23772
rect 33951 23763 34009 23769
rect 33951 23760 33963 23763
rect 31430 23732 33963 23760
rect 31430 23720 31436 23732
rect 33951 23729 33963 23732
rect 33997 23729 34009 23763
rect 33951 23723 34009 23729
rect 2303 23695 2361 23701
rect 2303 23661 2315 23695
rect 2349 23661 2361 23695
rect 2303 23655 2361 23661
rect 2395 23695 2453 23701
rect 2395 23661 2407 23695
rect 2441 23692 2453 23695
rect 2484 23692 2490 23704
rect 2441 23664 2490 23692
rect 2441 23661 2453 23664
rect 2395 23655 2453 23661
rect 2318 23624 2346 23655
rect 2484 23652 2490 23664
rect 2542 23652 2548 23704
rect 2668 23652 2674 23704
rect 2726 23692 2732 23704
rect 2855 23695 2913 23701
rect 2855 23692 2867 23695
rect 2726 23664 2867 23692
rect 2726 23652 2732 23664
rect 2855 23661 2867 23664
rect 2901 23661 2913 23695
rect 2855 23655 2913 23661
rect 3039 23695 3097 23701
rect 3039 23661 3051 23695
rect 3085 23692 3097 23695
rect 3588 23692 3594 23704
rect 3085 23664 3594 23692
rect 3085 23661 3097 23664
rect 3039 23655 3097 23661
rect 3588 23652 3594 23664
rect 3646 23652 3652 23704
rect 7179 23695 7237 23701
rect 7179 23661 7191 23695
rect 7225 23692 7237 23695
rect 7268 23692 7274 23704
rect 7225 23664 7274 23692
rect 7225 23661 7237 23664
rect 7179 23655 7237 23661
rect 7268 23652 7274 23664
rect 7326 23652 7332 23704
rect 34592 23652 34598 23704
rect 34650 23692 34656 23704
rect 34702 23692 34730 23859
rect 34868 23856 34874 23868
rect 34926 23856 34932 23908
rect 36800 23856 36806 23908
rect 36858 23896 36864 23908
rect 37079 23899 37137 23905
rect 37079 23896 37091 23899
rect 36858 23868 37091 23896
rect 36858 23856 36864 23868
rect 37079 23865 37091 23868
rect 37125 23865 37137 23899
rect 37079 23859 37137 23865
rect 34886 23760 34914 23856
rect 35254 23800 36202 23828
rect 35055 23763 35113 23769
rect 35055 23760 35067 23763
rect 34886 23732 35067 23760
rect 35055 23729 35067 23732
rect 35101 23729 35113 23763
rect 35055 23723 35113 23729
rect 35254 23701 35282 23800
rect 35239 23695 35297 23701
rect 35239 23692 35251 23695
rect 34650 23664 35251 23692
rect 34650 23652 34656 23664
rect 35239 23661 35251 23664
rect 35285 23661 35297 23695
rect 35239 23655 35297 23661
rect 35604 23652 35610 23704
rect 35662 23692 35668 23704
rect 35699 23695 35757 23701
rect 35699 23692 35711 23695
rect 35662 23664 35711 23692
rect 35662 23652 35668 23664
rect 35699 23661 35711 23664
rect 35745 23661 35757 23695
rect 35699 23655 35757 23661
rect 35791 23695 35849 23701
rect 35791 23661 35803 23695
rect 35837 23692 35849 23695
rect 36174 23692 36202 23800
rect 36343 23763 36401 23769
rect 36343 23729 36355 23763
rect 36389 23760 36401 23763
rect 37539 23763 37597 23769
rect 37539 23760 37551 23763
rect 36389 23732 37551 23760
rect 36389 23729 36401 23732
rect 36343 23723 36401 23729
rect 37539 23729 37551 23732
rect 37585 23729 37597 23763
rect 37539 23723 37597 23729
rect 42320 23720 42326 23772
rect 42378 23760 42384 23772
rect 68264 23760 68270 23772
rect 42378 23732 68270 23760
rect 42378 23720 42384 23732
rect 68264 23720 68270 23732
rect 68322 23760 68328 23772
rect 70932 23760 70938 23772
rect 68322 23732 70938 23760
rect 68322 23720 68328 23732
rect 70932 23720 70938 23732
rect 70990 23720 70996 23772
rect 35837 23664 36202 23692
rect 35837 23661 35849 23664
rect 35791 23655 35849 23661
rect 2686 23624 2714 23652
rect 2318 23596 2714 23624
rect 35714 23624 35742 23655
rect 36800 23652 36806 23704
rect 36858 23692 36864 23704
rect 37263 23695 37321 23701
rect 37263 23692 37275 23695
rect 36858 23664 37275 23692
rect 36858 23652 36864 23664
rect 37263 23661 37275 23664
rect 37309 23661 37321 23695
rect 37263 23655 37321 23661
rect 36524 23624 36530 23636
rect 35714 23596 36530 23624
rect 36524 23584 36530 23596
rect 36582 23584 36588 23636
rect 3312 23556 3318 23568
rect 3273 23528 3318 23556
rect 3312 23516 3318 23528
rect 3370 23516 3376 23568
rect 7271 23559 7329 23565
rect 7271 23525 7283 23559
rect 7317 23556 7329 23559
rect 9016 23556 9022 23568
rect 7317 23528 9022 23556
rect 7317 23525 7329 23528
rect 7271 23519 7329 23525
rect 9016 23516 9022 23528
rect 9074 23516 9080 23568
rect 38640 23516 38646 23568
rect 38698 23556 38704 23568
rect 38827 23559 38885 23565
rect 38827 23556 38839 23559
rect 38698 23528 38839 23556
rect 38698 23516 38704 23528
rect 38827 23525 38839 23528
rect 38873 23556 38885 23559
rect 43516 23556 43522 23568
rect 38873 23528 43522 23556
rect 38873 23525 38885 23528
rect 38827 23519 38885 23525
rect 43516 23516 43522 23528
rect 43574 23516 43580 23568
rect 538 23466 8450 23488
rect 538 23414 6344 23466
rect 6396 23414 6408 23466
rect 6460 23414 6472 23466
rect 6524 23414 6536 23466
rect 6588 23414 8450 23466
rect 538 23392 8450 23414
rect 34118 23466 43410 23488
rect 34118 23414 38312 23466
rect 38364 23414 38376 23466
rect 38428 23414 38440 23466
rect 38492 23414 38504 23466
rect 38556 23414 43410 23466
rect 34118 23392 43410 23414
rect 3588 23352 3594 23364
rect 3549 23324 3594 23352
rect 3588 23312 3594 23324
rect 3646 23312 3652 23364
rect 6535 23355 6593 23361
rect 6535 23352 6547 23355
rect 4802 23324 6547 23352
rect 3404 23244 3410 23296
rect 3462 23284 3468 23296
rect 4802 23284 4830 23324
rect 6535 23321 6547 23324
rect 6581 23352 6593 23355
rect 6716 23352 6722 23364
rect 6581 23324 6722 23352
rect 6581 23321 6593 23324
rect 6535 23315 6593 23321
rect 6716 23312 6722 23324
rect 6774 23312 6780 23364
rect 33951 23355 34009 23361
rect 33951 23321 33963 23355
rect 33997 23352 34009 23355
rect 34779 23355 34837 23361
rect 34779 23352 34791 23355
rect 33997 23324 34791 23352
rect 33997 23321 34009 23324
rect 33951 23315 34009 23321
rect 34779 23321 34791 23324
rect 34825 23321 34837 23355
rect 39468 23352 39474 23364
rect 39429 23324 39474 23352
rect 34779 23315 34837 23321
rect 39468 23312 39474 23324
rect 39526 23312 39532 23364
rect 3462 23256 4830 23284
rect 3462 23244 3468 23256
rect 3496 23216 3502 23228
rect 3457 23188 3502 23216
rect 3496 23176 3502 23188
rect 3554 23176 3560 23228
rect 4802 23225 4830 23256
rect 6443 23287 6501 23293
rect 6443 23253 6455 23287
rect 6489 23284 6501 23287
rect 6624 23284 6630 23296
rect 6489 23256 6630 23284
rect 6489 23253 6501 23256
rect 6443 23247 6501 23253
rect 6624 23244 6630 23256
rect 6682 23244 6688 23296
rect 39560 23244 39566 23296
rect 39618 23284 39624 23296
rect 39618 23256 40894 23284
rect 39618 23244 39624 23256
rect 4787 23219 4845 23225
rect 4787 23185 4799 23219
rect 4833 23185 4845 23219
rect 34408 23216 34414 23228
rect 34369 23188 34414 23216
rect 4787 23179 4845 23185
rect 34408 23176 34414 23188
rect 34466 23216 34472 23228
rect 34963 23219 35021 23225
rect 34963 23216 34975 23219
rect 34466 23188 34975 23216
rect 34466 23176 34472 23188
rect 34963 23185 34975 23188
rect 35009 23185 35021 23219
rect 38180 23216 38186 23228
rect 38141 23188 38186 23216
rect 34963 23179 35021 23185
rect 38180 23176 38186 23188
rect 38238 23176 38244 23228
rect 40498 23225 40526 23256
rect 40483 23219 40541 23225
rect 40483 23185 40495 23219
rect 40529 23216 40541 23219
rect 40529 23188 40563 23216
rect 40529 23185 40541 23188
rect 40483 23179 40541 23185
rect 5063 23151 5121 23157
rect 5063 23117 5075 23151
rect 5109 23148 5121 23151
rect 7176 23148 7182 23160
rect 5109 23120 7182 23148
rect 5109 23117 5121 23120
rect 5063 23111 5121 23117
rect 7176 23108 7182 23120
rect 7234 23108 7240 23160
rect 40866 23157 40894 23256
rect 37907 23151 37965 23157
rect 37907 23148 37919 23151
rect 37738 23120 37919 23148
rect 3496 22972 3502 23024
rect 3554 23012 3560 23024
rect 3775 23015 3833 23021
rect 3775 23012 3787 23015
rect 3554 22984 3787 23012
rect 3554 22972 3560 22984
rect 3775 22981 3787 22984
rect 3821 22981 3833 23015
rect 3775 22975 3833 22981
rect 34595 23015 34653 23021
rect 34595 22981 34607 23015
rect 34641 23012 34653 23015
rect 35328 23012 35334 23024
rect 34641 22984 35334 23012
rect 34641 22981 34653 22984
rect 34595 22975 34653 22981
rect 35328 22972 35334 22984
rect 35386 22972 35392 23024
rect 36708 22972 36714 23024
rect 36766 23012 36772 23024
rect 37738 23021 37766 23120
rect 37907 23117 37919 23120
rect 37953 23117 37965 23151
rect 37907 23111 37965 23117
rect 40851 23151 40909 23157
rect 40851 23117 40863 23151
rect 40897 23148 40909 23151
rect 42320 23148 42326 23160
rect 40897 23120 42326 23148
rect 40897 23117 40909 23120
rect 40851 23111 40909 23117
rect 42320 23108 42326 23120
rect 42378 23108 42384 23160
rect 37723 23015 37781 23021
rect 37723 23012 37735 23015
rect 36766 22984 37735 23012
rect 36766 22972 36772 22984
rect 37723 22981 37735 22984
rect 37769 22981 37781 23015
rect 37723 22975 37781 22981
rect 40575 23015 40633 23021
rect 40575 22981 40587 23015
rect 40621 23012 40633 23015
rect 40664 23012 40670 23024
rect 40621 22984 40670 23012
rect 40621 22981 40633 22984
rect 40575 22975 40633 22981
rect 40664 22972 40670 22984
rect 40722 22972 40728 23024
rect 538 22922 8450 22944
rect 538 22870 3680 22922
rect 3732 22870 3744 22922
rect 3796 22870 3808 22922
rect 3860 22870 3872 22922
rect 3924 22870 8450 22922
rect 538 22848 8450 22870
rect 34118 22922 43410 22944
rect 34118 22870 35648 22922
rect 35700 22870 35712 22922
rect 35764 22870 35776 22922
rect 35828 22870 35840 22922
rect 35892 22870 40976 22922
rect 41028 22870 41040 22922
rect 41092 22870 41104 22922
rect 41156 22870 41168 22922
rect 41220 22870 43410 22922
rect 34118 22848 43410 22870
rect 6624 22808 6630 22820
rect 6585 22780 6630 22808
rect 6624 22768 6630 22780
rect 6682 22768 6688 22820
rect 34592 22808 34598 22820
rect 34553 22780 34598 22808
rect 34592 22768 34598 22780
rect 34650 22768 34656 22820
rect 3223 22743 3281 22749
rect 3223 22709 3235 22743
rect 3269 22740 3281 22743
rect 3496 22740 3502 22752
rect 3269 22712 3502 22740
rect 3269 22709 3281 22712
rect 3223 22703 3281 22709
rect 3496 22700 3502 22712
rect 3554 22700 3560 22752
rect 1935 22675 1993 22681
rect 1935 22641 1947 22675
rect 1981 22672 1993 22675
rect 3312 22672 3318 22684
rect 1981 22644 3318 22672
rect 1981 22641 1993 22644
rect 1935 22635 1993 22641
rect 3312 22632 3318 22644
rect 3370 22632 3376 22684
rect 3404 22632 3410 22684
rect 3462 22672 3468 22684
rect 3462 22644 3507 22672
rect 3462 22632 3468 22644
rect 1659 22607 1717 22613
rect 1659 22573 1671 22607
rect 1705 22604 1717 22607
rect 3422 22604 3450 22632
rect 1705 22576 3450 22604
rect 1705 22573 1717 22576
rect 1659 22567 1717 22573
rect 3588 22564 3594 22616
rect 3646 22604 3652 22616
rect 4235 22607 4293 22613
rect 4235 22604 4247 22607
rect 3646 22576 4247 22604
rect 3646 22564 3652 22576
rect 4235 22573 4247 22576
rect 4281 22604 4293 22607
rect 4416 22604 4422 22616
rect 4281 22576 4422 22604
rect 4281 22573 4293 22576
rect 4235 22567 4293 22573
rect 4416 22564 4422 22576
rect 4474 22564 4480 22616
rect 6259 22607 6317 22613
rect 6259 22573 6271 22607
rect 6305 22604 6317 22607
rect 6642 22604 6670 22768
rect 30360 22632 30366 22684
rect 30418 22672 30424 22684
rect 42320 22672 42326 22684
rect 30418 22644 40802 22672
rect 42281 22644 42326 22672
rect 30418 22632 30424 22644
rect 6305 22576 6670 22604
rect 6305 22573 6317 22576
rect 6259 22567 6317 22573
rect 30912 22564 30918 22616
rect 30970 22604 30976 22616
rect 33951 22607 34009 22613
rect 33951 22604 33963 22607
rect 30970 22576 33963 22604
rect 30970 22564 30976 22576
rect 33951 22573 33963 22576
rect 33997 22604 34009 22607
rect 34411 22607 34469 22613
rect 34411 22604 34423 22607
rect 33997 22576 34423 22604
rect 33997 22573 34009 22576
rect 33951 22567 34009 22573
rect 34411 22573 34423 22576
rect 34457 22604 34469 22607
rect 34963 22607 35021 22613
rect 34963 22604 34975 22607
rect 34457 22576 34975 22604
rect 34457 22573 34469 22576
rect 34411 22567 34469 22573
rect 34963 22573 34975 22576
rect 35009 22573 35021 22607
rect 34963 22567 35021 22573
rect 36892 22564 36898 22616
rect 36950 22604 36956 22616
rect 37355 22607 37413 22613
rect 37355 22604 37367 22607
rect 36950 22576 37367 22604
rect 36950 22564 36956 22576
rect 37355 22573 37367 22576
rect 37401 22604 37413 22607
rect 37539 22607 37597 22613
rect 37539 22604 37551 22607
rect 37401 22576 37551 22604
rect 37401 22573 37413 22576
rect 37355 22567 37413 22573
rect 37539 22573 37551 22576
rect 37585 22573 37597 22607
rect 38640 22604 38646 22616
rect 38601 22576 38646 22604
rect 37539 22567 37597 22573
rect 38640 22564 38646 22576
rect 38698 22564 38704 22616
rect 40667 22607 40725 22613
rect 40667 22604 40679 22607
rect 40498 22576 40679 22604
rect 6351 22539 6409 22545
rect 6351 22505 6363 22539
rect 6397 22536 6409 22539
rect 6624 22536 6630 22548
rect 6397 22508 6630 22536
rect 6397 22505 6409 22508
rect 6351 22499 6409 22505
rect 6624 22496 6630 22508
rect 6682 22496 6688 22548
rect 36524 22496 36530 22548
rect 36582 22536 36588 22548
rect 38735 22539 38793 22545
rect 38735 22536 38747 22539
rect 36582 22508 38747 22536
rect 36582 22496 36588 22508
rect 38735 22505 38747 22508
rect 38781 22505 38793 22539
rect 38735 22499 38793 22505
rect 4416 22468 4422 22480
rect 4377 22440 4422 22468
rect 4416 22428 4422 22440
rect 4474 22428 4480 22480
rect 34776 22468 34782 22480
rect 34737 22440 34782 22468
rect 34776 22428 34782 22440
rect 34834 22428 34840 22480
rect 37723 22471 37781 22477
rect 37723 22437 37735 22471
rect 37769 22468 37781 22471
rect 38088 22468 38094 22480
rect 37769 22440 38094 22468
rect 37769 22437 37781 22440
rect 37723 22431 37781 22437
rect 38088 22428 38094 22440
rect 38146 22428 38152 22480
rect 39652 22428 39658 22480
rect 39710 22468 39716 22480
rect 40498 22477 40526 22576
rect 40667 22573 40679 22576
rect 40713 22573 40725 22607
rect 40667 22567 40725 22573
rect 40483 22471 40541 22477
rect 40483 22468 40495 22471
rect 39710 22440 40495 22468
rect 39710 22428 39716 22440
rect 40483 22437 40495 22440
rect 40529 22437 40541 22471
rect 40774 22468 40802 22644
rect 42320 22632 42326 22644
rect 42378 22632 42384 22684
rect 40940 22604 40946 22616
rect 40901 22576 40946 22604
rect 40940 22564 40946 22576
rect 40998 22564 41004 22616
rect 41970 22508 43102 22536
rect 41970 22468 41998 22508
rect 43074 22480 43102 22508
rect 43056 22468 43062 22480
rect 40774 22440 41998 22468
rect 43017 22440 43062 22468
rect 40483 22431 40541 22437
rect 43056 22428 43062 22440
rect 43114 22428 43120 22480
rect 538 22378 8450 22400
rect 538 22326 6344 22378
rect 6396 22326 6408 22378
rect 6460 22326 6472 22378
rect 6524 22326 6536 22378
rect 6588 22326 8450 22378
rect 538 22304 8450 22326
rect 34118 22378 43410 22400
rect 34118 22326 38312 22378
rect 38364 22326 38376 22378
rect 38428 22326 38440 22378
rect 38492 22326 38504 22378
rect 38556 22326 43410 22378
rect 34118 22304 43410 22326
rect 3683 22267 3741 22273
rect 3683 22233 3695 22267
rect 3729 22264 3741 22267
rect 3864 22264 3870 22276
rect 3729 22236 3870 22264
rect 3729 22233 3741 22236
rect 3683 22227 3741 22233
rect 3864 22224 3870 22236
rect 3922 22264 3928 22276
rect 4600 22264 4606 22276
rect 3922 22236 4606 22264
rect 3922 22224 3928 22236
rect 4600 22224 4606 22236
rect 4658 22224 4664 22276
rect 7176 22264 7182 22276
rect 7137 22236 7182 22264
rect 7176 22224 7182 22236
rect 7234 22224 7240 22276
rect 39284 22224 39290 22276
rect 39342 22264 39348 22276
rect 39563 22267 39621 22273
rect 39563 22264 39575 22267
rect 39342 22236 39575 22264
rect 39342 22224 39348 22236
rect 39563 22233 39575 22236
rect 39609 22233 39621 22267
rect 40940 22264 40946 22276
rect 40901 22236 40946 22264
rect 39563 22227 39621 22233
rect 40940 22224 40946 22236
rect 40998 22224 41004 22276
rect 2668 22156 2674 22208
rect 2726 22196 2732 22208
rect 4416 22196 4422 22208
rect 2726 22168 4422 22196
rect 2726 22156 2732 22168
rect 4416 22156 4422 22168
rect 4474 22196 4480 22208
rect 4474 22168 6762 22196
rect 4474 22156 4480 22168
rect 2303 22131 2361 22137
rect 2303 22097 2315 22131
rect 2349 22097 2361 22131
rect 2303 22091 2361 22097
rect 2318 22060 2346 22091
rect 2760 22088 2766 22140
rect 2818 22128 2824 22140
rect 3959 22131 4017 22137
rect 3959 22128 3971 22131
rect 2818 22100 3971 22128
rect 2818 22088 2824 22100
rect 3959 22097 3971 22100
rect 4005 22128 4017 22131
rect 4511 22131 4569 22137
rect 4511 22128 4523 22131
rect 4005 22100 4523 22128
rect 4005 22097 4017 22100
rect 3959 22091 4017 22097
rect 4511 22097 4523 22100
rect 4557 22097 4569 22131
rect 4511 22091 4569 22097
rect 4695 22131 4753 22137
rect 4695 22097 4707 22131
rect 4741 22128 4753 22131
rect 6072 22128 6078 22140
rect 4741 22100 6078 22128
rect 4741 22097 4753 22100
rect 4695 22091 4753 22097
rect 6072 22088 6078 22100
rect 6130 22088 6136 22140
rect 6182 22137 6210 22168
rect 6167 22131 6225 22137
rect 6167 22097 6179 22131
rect 6213 22097 6225 22131
rect 6167 22091 6225 22097
rect 6259 22131 6317 22137
rect 6259 22097 6271 22131
rect 6305 22128 6317 22131
rect 6624 22128 6630 22140
rect 6305 22100 6394 22128
rect 6585 22100 6630 22128
rect 6305 22097 6317 22100
rect 6259 22091 6317 22097
rect 3588 22060 3594 22072
rect 2318 22032 3594 22060
rect 3588 22020 3594 22032
rect 3646 22020 3652 22072
rect 3864 22060 3870 22072
rect 3825 22032 3870 22060
rect 3864 22020 3870 22032
rect 3922 22020 3928 22072
rect 5891 22063 5949 22069
rect 5891 22029 5903 22063
rect 5937 22060 5949 22063
rect 6366 22060 6394 22100
rect 6624 22088 6630 22100
rect 6682 22088 6688 22140
rect 6734 22137 6762 22168
rect 6719 22131 6777 22137
rect 6719 22097 6731 22131
rect 6765 22097 6777 22131
rect 6719 22091 6777 22097
rect 35331 22131 35389 22137
rect 35331 22097 35343 22131
rect 35377 22128 35389 22131
rect 35420 22128 35426 22140
rect 35377 22100 35426 22128
rect 35377 22097 35389 22100
rect 35331 22091 35389 22097
rect 35420 22088 35426 22100
rect 35478 22128 35484 22140
rect 35607 22131 35665 22137
rect 35607 22128 35619 22131
rect 35478 22100 35619 22128
rect 35478 22088 35484 22100
rect 35607 22097 35619 22100
rect 35653 22128 35665 22131
rect 36524 22128 36530 22140
rect 35653 22100 36530 22128
rect 35653 22097 35665 22100
rect 35607 22091 35665 22097
rect 36524 22088 36530 22100
rect 36582 22088 36588 22140
rect 36616 22088 36622 22140
rect 36674 22128 36680 22140
rect 39931 22131 39989 22137
rect 39931 22128 39943 22131
rect 36674 22100 39943 22128
rect 36674 22088 36680 22100
rect 39931 22097 39943 22100
rect 39977 22128 39989 22131
rect 40483 22131 40541 22137
rect 40483 22128 40495 22131
rect 39977 22100 40495 22128
rect 39977 22097 39989 22100
rect 39931 22091 39989 22097
rect 40483 22097 40495 22100
rect 40529 22097 40541 22131
rect 40664 22128 40670 22140
rect 40625 22100 40670 22128
rect 40483 22091 40541 22097
rect 40664 22088 40670 22100
rect 40722 22088 40728 22140
rect 5937 22032 6394 22060
rect 5937 22029 5949 22032
rect 5891 22023 5949 22029
rect 6366 21992 6394 22032
rect 39284 22020 39290 22072
rect 39342 22060 39348 22072
rect 39747 22063 39805 22069
rect 39747 22060 39759 22063
rect 39342 22032 39759 22060
rect 39342 22020 39348 22032
rect 39747 22029 39759 22032
rect 39793 22029 39805 22063
rect 39747 22023 39805 22029
rect 8372 21992 8378 22004
rect 6366 21964 8378 21992
rect 8372 21952 8378 21964
rect 8430 21952 8436 22004
rect 2487 21927 2545 21933
rect 2487 21893 2499 21927
rect 2533 21924 2545 21927
rect 2760 21924 2766 21936
rect 2533 21896 2766 21924
rect 2533 21893 2545 21896
rect 2487 21887 2545 21893
rect 2760 21884 2766 21896
rect 2818 21884 2824 21936
rect 4968 21924 4974 21936
rect 4929 21896 4974 21924
rect 4968 21884 4974 21896
rect 5026 21884 5032 21936
rect 35420 21924 35426 21936
rect 35381 21896 35426 21924
rect 35420 21884 35426 21896
rect 35478 21884 35484 21936
rect 538 21834 8450 21856
rect 538 21782 3680 21834
rect 3732 21782 3744 21834
rect 3796 21782 3808 21834
rect 3860 21782 3872 21834
rect 3924 21782 8450 21834
rect 538 21760 8450 21782
rect 34118 21834 43410 21856
rect 34118 21782 35648 21834
rect 35700 21782 35712 21834
rect 35764 21782 35776 21834
rect 35828 21782 35840 21834
rect 35892 21782 40976 21834
rect 41028 21782 41040 21834
rect 41092 21782 41104 21834
rect 41156 21782 41168 21834
rect 41220 21782 43410 21834
rect 34118 21760 43410 21782
rect 67068 21748 67074 21800
rect 67126 21788 67132 21800
rect 71208 21788 71214 21800
rect 67126 21760 71214 21788
rect 67126 21748 67132 21760
rect 71208 21748 71214 21760
rect 71266 21748 71272 21800
rect 3683 21723 3741 21729
rect 3683 21689 3695 21723
rect 3729 21720 3741 21723
rect 4508 21720 4514 21732
rect 3729 21692 4514 21720
rect 3729 21689 3741 21692
rect 3683 21683 3741 21689
rect 3882 21593 3910 21692
rect 4508 21680 4514 21692
rect 4566 21680 4572 21732
rect 33951 21723 34009 21729
rect 33951 21689 33963 21723
rect 33997 21720 34009 21723
rect 34963 21723 35021 21729
rect 34963 21720 34975 21723
rect 33997 21692 34975 21720
rect 33997 21689 34009 21692
rect 33951 21683 34009 21689
rect 3867 21587 3925 21593
rect 3867 21553 3879 21587
rect 3913 21553 3925 21587
rect 3867 21547 3925 21553
rect 2668 21516 2674 21528
rect 2629 21488 2674 21516
rect 2668 21476 2674 21488
rect 2726 21476 2732 21528
rect 2760 21476 2766 21528
rect 2818 21516 2824 21528
rect 3959 21519 4017 21525
rect 3959 21516 3971 21519
rect 2818 21488 3971 21516
rect 2818 21476 2824 21488
rect 3959 21485 3971 21488
rect 4005 21485 4017 21519
rect 3959 21479 4017 21485
rect 4511 21519 4569 21525
rect 4511 21485 4523 21519
rect 4557 21485 4569 21519
rect 4511 21479 4569 21485
rect 4695 21519 4753 21525
rect 4695 21485 4707 21519
rect 4741 21516 4753 21519
rect 6164 21516 6170 21528
rect 4741 21488 6170 21516
rect 4741 21485 4753 21488
rect 4695 21479 4753 21485
rect 3974 21448 4002 21479
rect 4526 21448 4554 21479
rect 6164 21476 6170 21488
rect 6222 21476 6228 21528
rect 34426 21525 34454 21692
rect 34963 21689 34975 21692
rect 35009 21689 35021 21723
rect 34963 21683 35021 21689
rect 35515 21723 35573 21729
rect 35515 21689 35527 21723
rect 35561 21720 35573 21723
rect 36708 21720 36714 21732
rect 35561 21692 36714 21720
rect 35561 21689 35573 21692
rect 35515 21683 35573 21689
rect 35622 21593 35650 21692
rect 36708 21680 36714 21692
rect 36766 21720 36772 21732
rect 39652 21720 39658 21732
rect 36766 21692 39658 21720
rect 36766 21680 36772 21692
rect 39652 21680 39658 21692
rect 39710 21680 39716 21732
rect 38732 21612 38738 21664
rect 38790 21652 38796 21664
rect 43056 21652 43062 21664
rect 38790 21624 43062 21652
rect 38790 21612 38796 21624
rect 43056 21612 43062 21624
rect 43114 21612 43120 21664
rect 35607 21587 35665 21593
rect 35607 21553 35619 21587
rect 35653 21553 35665 21587
rect 35607 21547 35665 21553
rect 36524 21544 36530 21596
rect 36582 21584 36588 21596
rect 36984 21584 36990 21596
rect 36582 21556 36990 21584
rect 36582 21544 36588 21556
rect 36984 21544 36990 21556
rect 37042 21544 37048 21596
rect 34411 21519 34469 21525
rect 34411 21485 34423 21519
rect 34457 21485 34469 21519
rect 35880 21516 35886 21528
rect 35841 21488 35886 21516
rect 34411 21479 34469 21485
rect 35880 21476 35886 21488
rect 35938 21476 35944 21528
rect 39836 21516 39842 21528
rect 39797 21488 39842 21516
rect 39836 21476 39842 21488
rect 39894 21516 39900 21528
rect 40115 21519 40173 21525
rect 40115 21516 40127 21519
rect 39894 21488 40127 21516
rect 39894 21476 39900 21488
rect 40115 21485 40127 21488
rect 40161 21516 40173 21519
rect 41492 21516 41498 21528
rect 40161 21488 41498 21516
rect 40161 21485 40173 21488
rect 40115 21479 40173 21485
rect 41492 21476 41498 21488
rect 41550 21476 41556 21528
rect 5060 21448 5066 21460
rect 3974 21420 4554 21448
rect 5021 21420 5066 21448
rect 5060 21408 5066 21420
rect 5118 21408 5124 21460
rect 2855 21383 2913 21389
rect 2855 21349 2867 21383
rect 2901 21380 2913 21383
rect 3312 21380 3318 21392
rect 2901 21352 3318 21380
rect 2901 21349 2913 21352
rect 2855 21343 2913 21349
rect 3312 21340 3318 21352
rect 3370 21340 3376 21392
rect 34592 21380 34598 21392
rect 34553 21352 34598 21380
rect 34592 21340 34598 21352
rect 34650 21340 34656 21392
rect 34776 21380 34782 21392
rect 34737 21352 34782 21380
rect 34776 21340 34782 21352
rect 34834 21340 34840 21392
rect 39468 21340 39474 21392
rect 39526 21380 39532 21392
rect 39931 21383 39989 21389
rect 39931 21380 39943 21383
rect 39526 21352 39943 21380
rect 39526 21340 39532 21352
rect 39931 21349 39943 21352
rect 39977 21349 39989 21383
rect 43056 21380 43062 21392
rect 43017 21352 43062 21380
rect 39931 21343 39989 21349
rect 43056 21340 43062 21352
rect 43114 21340 43120 21392
rect 538 21290 8450 21312
rect 538 21238 6344 21290
rect 6396 21238 6408 21290
rect 6460 21238 6472 21290
rect 6524 21238 6536 21290
rect 6588 21238 8450 21290
rect 538 21216 8450 21238
rect 34118 21290 43410 21312
rect 34118 21238 38312 21290
rect 38364 21238 38376 21290
rect 38428 21238 38440 21290
rect 38492 21238 38504 21290
rect 38556 21238 43410 21290
rect 34118 21216 43410 21238
rect 6072 21136 6078 21188
rect 6130 21176 6136 21188
rect 7087 21179 7145 21185
rect 7087 21176 7099 21179
rect 6130 21148 7099 21176
rect 6130 21136 6136 21148
rect 7087 21145 7099 21148
rect 7133 21145 7145 21179
rect 7087 21139 7145 21145
rect 34132 21136 34138 21188
rect 34190 21176 34196 21188
rect 34411 21179 34469 21185
rect 34411 21176 34423 21179
rect 34190 21148 34423 21176
rect 34190 21136 34196 21148
rect 34411 21145 34423 21148
rect 34457 21145 34469 21179
rect 35328 21176 35334 21188
rect 34411 21139 34469 21145
rect 34794 21148 35334 21176
rect 6167 21111 6225 21117
rect 6167 21077 6179 21111
rect 6213 21108 6225 21111
rect 6900 21108 6906 21120
rect 6213 21080 6906 21108
rect 6213 21077 6225 21080
rect 6167 21071 6225 21077
rect 6900 21068 6906 21080
rect 6958 21108 6964 21120
rect 6958 21080 7038 21108
rect 6958 21068 6964 21080
rect 3404 21000 3410 21052
rect 3462 21040 3468 21052
rect 4511 21043 4569 21049
rect 4511 21040 4523 21043
rect 3462 21012 4523 21040
rect 3462 21000 3468 21012
rect 4511 21009 4523 21012
rect 4557 21009 4569 21043
rect 4511 21003 4569 21009
rect 6351 21043 6409 21049
rect 6351 21009 6363 21043
rect 6397 21040 6409 21043
rect 6716 21040 6722 21052
rect 6397 21012 6722 21040
rect 6397 21009 6409 21012
rect 6351 21003 6409 21009
rect 6716 21000 6722 21012
rect 6774 21000 6780 21052
rect 7010 21049 7038 21080
rect 6995 21043 7053 21049
rect 6995 21009 7007 21043
rect 7041 21009 7053 21043
rect 34426 21040 34454 21139
rect 34500 21040 34506 21052
rect 34413 21012 34506 21040
rect 6995 21003 7053 21009
rect 34500 21000 34506 21012
rect 34558 21040 34564 21052
rect 34794 21049 34822 21148
rect 35328 21136 35334 21148
rect 35386 21136 35392 21188
rect 37444 21136 37450 21188
rect 37502 21176 37508 21188
rect 37539 21179 37597 21185
rect 37539 21176 37551 21179
rect 37502 21148 37551 21176
rect 37502 21136 37508 21148
rect 37539 21145 37551 21148
rect 37585 21145 37597 21179
rect 37539 21139 37597 21145
rect 39652 21136 39658 21188
rect 39710 21176 39716 21188
rect 39747 21179 39805 21185
rect 39747 21176 39759 21179
rect 39710 21148 39759 21176
rect 39710 21136 39716 21148
rect 39747 21145 39759 21148
rect 39793 21145 39805 21179
rect 39747 21139 39805 21145
rect 35420 21108 35426 21120
rect 35254 21080 35426 21108
rect 35254 21049 35282 21080
rect 35420 21068 35426 21080
rect 35478 21068 35484 21120
rect 35880 21108 35886 21120
rect 35841 21080 35886 21108
rect 35880 21068 35886 21080
rect 35938 21068 35944 21120
rect 39011 21111 39069 21117
rect 39011 21077 39023 21111
rect 39057 21108 39069 21111
rect 39057 21080 39606 21108
rect 39057 21077 39069 21080
rect 39011 21071 39069 21077
rect 34595 21043 34653 21049
rect 34595 21040 34607 21043
rect 34558 21012 34607 21040
rect 34558 21000 34564 21012
rect 34595 21009 34607 21012
rect 34641 21009 34653 21043
rect 34595 21003 34653 21009
rect 34779 21043 34837 21049
rect 34779 21009 34791 21043
rect 34825 21009 34837 21043
rect 34779 21003 34837 21009
rect 35239 21043 35297 21049
rect 35239 21009 35251 21043
rect 35285 21009 35297 21043
rect 35239 21003 35297 21009
rect 35328 21000 35334 21052
rect 35386 21040 35392 21052
rect 36616 21040 36622 21052
rect 35386 21012 36622 21040
rect 35386 21000 35392 21012
rect 36616 21000 36622 21012
rect 36674 21040 36680 21052
rect 37907 21043 37965 21049
rect 37907 21040 37919 21043
rect 36674 21012 37919 21040
rect 36674 21000 36680 21012
rect 37907 21009 37919 21012
rect 37953 21009 37965 21043
rect 37907 21003 37965 21009
rect 38088 21000 38094 21052
rect 38146 21040 38152 21052
rect 38459 21043 38517 21049
rect 38459 21040 38471 21043
rect 38146 21012 38471 21040
rect 38146 21000 38152 21012
rect 38459 21009 38471 21012
rect 38505 21009 38517 21043
rect 38459 21003 38517 21009
rect 38643 21043 38701 21049
rect 38643 21009 38655 21043
rect 38689 21040 38701 21043
rect 39468 21040 39474 21052
rect 38689 21012 39474 21040
rect 38689 21009 38701 21012
rect 38643 21003 38701 21009
rect 39468 21000 39474 21012
rect 39526 21000 39532 21052
rect 39578 21040 39606 21080
rect 40207 21043 40265 21049
rect 40207 21040 40219 21043
rect 39578 21012 40219 21040
rect 40207 21009 40219 21012
rect 40253 21009 40265 21043
rect 40207 21003 40265 21009
rect 4787 20975 4845 20981
rect 4787 20941 4799 20975
rect 4833 20972 4845 20975
rect 4968 20972 4974 20984
rect 4833 20944 4974 20972
rect 4833 20941 4845 20944
rect 4787 20935 4845 20941
rect 4968 20932 4974 20944
rect 5026 20932 5032 20984
rect 37444 20932 37450 20984
rect 37502 20972 37508 20984
rect 37723 20975 37781 20981
rect 37723 20972 37735 20975
rect 37502 20944 37735 20972
rect 37502 20932 37508 20944
rect 37723 20941 37735 20944
rect 37769 20941 37781 20975
rect 37723 20935 37781 20941
rect 39652 20932 39658 20984
rect 39710 20972 39716 20984
rect 39931 20975 39989 20981
rect 39931 20972 39943 20975
rect 39710 20944 39943 20972
rect 39710 20932 39716 20944
rect 39931 20941 39943 20944
rect 39977 20941 39989 20975
rect 39931 20935 39989 20941
rect 41492 20836 41498 20848
rect 41453 20808 41498 20836
rect 41492 20796 41498 20808
rect 41550 20796 41556 20848
rect 538 20746 8450 20768
rect 538 20694 3680 20746
rect 3732 20694 3744 20746
rect 3796 20694 3808 20746
rect 3860 20694 3872 20746
rect 3924 20694 8450 20746
rect 538 20672 8450 20694
rect 34118 20746 43410 20768
rect 34118 20694 35648 20746
rect 35700 20694 35712 20746
rect 35764 20694 35776 20746
rect 35828 20694 35840 20746
rect 35892 20694 40976 20746
rect 41028 20694 41040 20746
rect 41092 20694 41104 20746
rect 41156 20694 41168 20746
rect 41220 20694 43410 20746
rect 34118 20672 43410 20694
rect 2392 20632 2398 20644
rect 2353 20604 2398 20632
rect 2392 20592 2398 20604
rect 2450 20592 2456 20644
rect 6164 20592 6170 20644
rect 6222 20632 6228 20644
rect 6351 20635 6409 20641
rect 6351 20632 6363 20635
rect 6222 20604 6363 20632
rect 6222 20592 6228 20604
rect 6351 20601 6363 20604
rect 6397 20601 6409 20635
rect 6351 20595 6409 20601
rect 34684 20592 34690 20644
rect 34742 20632 34748 20644
rect 36067 20635 36125 20641
rect 36067 20632 36079 20635
rect 34742 20604 36079 20632
rect 34742 20592 34748 20604
rect 36067 20601 36079 20604
rect 36113 20601 36125 20635
rect 36067 20595 36125 20601
rect 2410 20496 2438 20592
rect 2579 20499 2637 20505
rect 2579 20496 2591 20499
rect 2410 20468 2591 20496
rect 2579 20465 2591 20468
rect 2625 20465 2637 20499
rect 2579 20459 2637 20465
rect 2760 20428 2766 20440
rect 2721 20400 2766 20428
rect 2760 20388 2766 20400
rect 2818 20388 2824 20440
rect 3312 20428 3318 20440
rect 3273 20400 3318 20428
rect 3312 20388 3318 20400
rect 3370 20388 3376 20440
rect 3499 20431 3557 20437
rect 3499 20397 3511 20431
rect 3545 20428 3557 20431
rect 4232 20428 4238 20440
rect 3545 20400 4238 20428
rect 3545 20397 3557 20400
rect 3499 20391 3557 20397
rect 4232 20388 4238 20400
rect 4290 20388 4296 20440
rect 6259 20431 6317 20437
rect 6259 20397 6271 20431
rect 6305 20428 6317 20431
rect 36082 20428 36110 20595
rect 39652 20592 39658 20644
rect 39710 20632 39716 20644
rect 40391 20635 40449 20641
rect 40391 20632 40403 20635
rect 39710 20604 40403 20632
rect 39710 20592 39716 20604
rect 40391 20601 40403 20604
rect 40437 20632 40449 20635
rect 40483 20635 40541 20641
rect 40483 20632 40495 20635
rect 40437 20604 40495 20632
rect 40437 20601 40449 20604
rect 40391 20595 40449 20601
rect 40483 20601 40495 20604
rect 40529 20601 40541 20635
rect 40483 20595 40541 20601
rect 43056 20496 43062 20508
rect 36358 20468 43062 20496
rect 36251 20431 36309 20437
rect 36251 20428 36263 20431
rect 6305 20400 6670 20428
rect 36082 20400 36263 20428
rect 6305 20397 6317 20400
rect 6259 20391 6317 20397
rect 3330 20360 3358 20388
rect 3588 20360 3594 20372
rect 3330 20332 3594 20360
rect 3588 20320 3594 20332
rect 3646 20320 3652 20372
rect 3867 20363 3925 20369
rect 3867 20329 3879 20363
rect 3913 20360 3925 20363
rect 4048 20360 4054 20372
rect 3913 20332 4054 20360
rect 3913 20329 3925 20332
rect 3867 20323 3925 20329
rect 4048 20320 4054 20332
rect 4106 20320 4112 20372
rect 6642 20301 6670 20400
rect 36251 20397 36263 20400
rect 36297 20397 36309 20431
rect 36251 20391 36309 20397
rect 30268 20320 30274 20372
rect 30326 20360 30332 20372
rect 36358 20360 36386 20468
rect 43056 20456 43062 20468
rect 43114 20456 43120 20508
rect 40391 20431 40449 20437
rect 40391 20397 40403 20431
rect 40437 20428 40449 20431
rect 40667 20431 40725 20437
rect 40667 20428 40679 20431
rect 40437 20400 40679 20428
rect 40437 20397 40449 20400
rect 40391 20391 40449 20397
rect 40667 20397 40679 20400
rect 40713 20397 40725 20431
rect 40940 20428 40946 20440
rect 40901 20400 40946 20428
rect 40667 20391 40725 20397
rect 40940 20388 40946 20400
rect 40998 20388 41004 20440
rect 42320 20360 42326 20372
rect 30326 20332 36386 20360
rect 42281 20332 42326 20360
rect 30326 20320 30332 20332
rect 42320 20320 42326 20332
rect 42378 20320 42384 20372
rect 6627 20295 6685 20301
rect 6627 20261 6639 20295
rect 6673 20292 6685 20295
rect 6808 20292 6814 20304
rect 6673 20264 6814 20292
rect 6673 20261 6685 20264
rect 6627 20255 6685 20261
rect 6808 20252 6814 20264
rect 6866 20252 6872 20304
rect 34408 20292 34414 20304
rect 34369 20264 34414 20292
rect 34408 20252 34414 20264
rect 34466 20252 34472 20304
rect 36432 20292 36438 20304
rect 36393 20264 36438 20292
rect 36432 20252 36438 20264
rect 36490 20252 36496 20304
rect 43056 20292 43062 20304
rect 43017 20264 43062 20292
rect 43056 20252 43062 20264
rect 43114 20252 43120 20304
rect 538 20202 8450 20224
rect 538 20150 6344 20202
rect 6396 20150 6408 20202
rect 6460 20150 6472 20202
rect 6524 20150 6536 20202
rect 6588 20150 8450 20202
rect 538 20128 8450 20150
rect 34118 20202 43410 20224
rect 34118 20150 38312 20202
rect 38364 20150 38376 20202
rect 38428 20150 38440 20202
rect 38492 20150 38504 20202
rect 38556 20150 43410 20202
rect 34118 20128 43410 20150
rect 39103 20091 39161 20097
rect 39103 20057 39115 20091
rect 39149 20088 39161 20091
rect 39284 20088 39290 20100
rect 39149 20060 39290 20088
rect 39149 20057 39161 20060
rect 39103 20051 39161 20057
rect 39284 20048 39290 20060
rect 39342 20048 39348 20100
rect 6808 20020 6814 20032
rect 6769 19992 6814 20020
rect 6808 19980 6814 19992
rect 6866 19980 6872 20032
rect 39394 19992 39974 20020
rect 5060 19912 5066 19964
rect 5118 19952 5124 19964
rect 5431 19955 5489 19961
rect 5431 19952 5443 19955
rect 5118 19924 5443 19952
rect 5118 19912 5124 19924
rect 5431 19921 5443 19924
rect 5477 19921 5489 19955
rect 5431 19915 5489 19921
rect 37628 19912 37634 19964
rect 37686 19952 37692 19964
rect 39394 19961 39422 19992
rect 39946 19961 39974 19992
rect 67160 19980 67166 20032
rect 67218 20020 67224 20032
rect 70472 20020 70478 20032
rect 67218 19992 70478 20020
rect 67218 19980 67224 19992
rect 70472 19980 70478 19992
rect 70530 20020 70536 20032
rect 71300 20020 71306 20032
rect 70530 19992 71306 20020
rect 70530 19980 70536 19992
rect 71300 19980 71306 19992
rect 71358 19980 71364 20032
rect 39379 19955 39437 19961
rect 39379 19952 39391 19955
rect 37686 19924 39391 19952
rect 37686 19912 37692 19924
rect 39379 19921 39391 19924
rect 39425 19921 39437 19955
rect 39839 19955 39897 19961
rect 39839 19952 39851 19955
rect 39379 19915 39437 19921
rect 39578 19924 39851 19952
rect 5155 19887 5213 19893
rect 5155 19853 5167 19887
rect 5201 19884 5213 19887
rect 6716 19884 6722 19896
rect 5201 19856 6722 19884
rect 5201 19853 5213 19856
rect 5155 19847 5213 19853
rect 6716 19844 6722 19856
rect 6774 19844 6780 19896
rect 39192 19884 39198 19896
rect 39153 19856 39198 19884
rect 39192 19844 39198 19856
rect 39250 19844 39256 19896
rect 30820 19776 30826 19828
rect 30878 19816 30884 19828
rect 39578 19816 39606 19924
rect 39839 19921 39851 19924
rect 39885 19921 39897 19955
rect 39839 19915 39897 19921
rect 39931 19955 39989 19961
rect 39931 19921 39943 19955
rect 39977 19952 39989 19955
rect 41587 19955 41645 19961
rect 39977 19924 40011 19952
rect 39977 19921 39989 19924
rect 39931 19915 39989 19921
rect 41587 19921 41599 19955
rect 41633 19952 41645 19955
rect 42320 19952 42326 19964
rect 41633 19924 42326 19952
rect 41633 19921 41645 19924
rect 41587 19915 41645 19921
rect 42320 19912 42326 19924
rect 42378 19912 42384 19964
rect 40483 19887 40541 19893
rect 40483 19853 40495 19887
rect 40529 19884 40541 19887
rect 40940 19884 40946 19896
rect 40529 19856 40946 19884
rect 40529 19853 40541 19856
rect 40483 19847 40541 19853
rect 40940 19844 40946 19856
rect 40998 19844 41004 19896
rect 40667 19819 40725 19825
rect 40667 19816 40679 19819
rect 30878 19788 40679 19816
rect 30878 19776 30884 19788
rect 40667 19785 40679 19788
rect 40713 19816 40725 19819
rect 41679 19819 41737 19825
rect 41679 19816 41691 19819
rect 40713 19788 41691 19816
rect 40713 19785 40725 19788
rect 40667 19779 40725 19785
rect 41679 19785 41691 19788
rect 41725 19785 41737 19819
rect 41679 19779 41737 19785
rect 6716 19708 6722 19760
rect 6774 19748 6780 19760
rect 6992 19748 6998 19760
rect 6774 19720 6998 19748
rect 6774 19708 6780 19720
rect 6992 19708 6998 19720
rect 7050 19708 7056 19760
rect 538 19658 8450 19680
rect 538 19606 3680 19658
rect 3732 19606 3744 19658
rect 3796 19606 3808 19658
rect 3860 19606 3872 19658
rect 3924 19606 8450 19658
rect 538 19584 8450 19606
rect 34118 19658 43410 19680
rect 34118 19606 35648 19658
rect 35700 19606 35712 19658
rect 35764 19606 35776 19658
rect 35828 19606 35840 19658
rect 35892 19606 40976 19658
rect 41028 19606 41040 19658
rect 41092 19606 41104 19658
rect 41156 19606 41168 19658
rect 41220 19606 43410 19658
rect 34118 19584 43410 19606
rect 4232 19544 4238 19556
rect 4193 19516 4238 19544
rect 4232 19504 4238 19516
rect 4290 19504 4296 19556
rect 34500 19504 34506 19556
rect 34558 19544 34564 19556
rect 34595 19547 34653 19553
rect 34595 19544 34607 19547
rect 34558 19516 34607 19544
rect 34558 19504 34564 19516
rect 34595 19513 34607 19516
rect 34641 19513 34653 19547
rect 34595 19507 34653 19513
rect 34960 19504 34966 19556
rect 35018 19544 35024 19556
rect 35515 19547 35573 19553
rect 35515 19544 35527 19547
rect 35018 19516 35527 19544
rect 35018 19504 35024 19516
rect 35515 19513 35527 19516
rect 35561 19513 35573 19547
rect 35515 19507 35573 19513
rect 37355 19547 37413 19553
rect 37355 19513 37367 19547
rect 37401 19544 37413 19547
rect 37444 19544 37450 19556
rect 37401 19516 37450 19544
rect 37401 19513 37413 19516
rect 37355 19507 37413 19513
rect 37444 19504 37450 19516
rect 37502 19504 37508 19556
rect 1935 19411 1993 19417
rect 1935 19377 1947 19411
rect 1981 19408 1993 19411
rect 4048 19408 4054 19420
rect 1981 19380 4054 19408
rect 1981 19377 1993 19380
rect 1935 19371 1993 19377
rect 4048 19368 4054 19380
rect 4106 19368 4112 19420
rect 37462 19417 37490 19504
rect 37447 19411 37505 19417
rect 37447 19377 37459 19411
rect 37493 19377 37505 19411
rect 37447 19371 37505 19377
rect 39011 19411 39069 19417
rect 39011 19377 39023 19411
rect 39057 19408 39069 19411
rect 39931 19411 39989 19417
rect 39931 19408 39943 19411
rect 39057 19380 39943 19408
rect 39057 19377 39069 19380
rect 39011 19371 39069 19377
rect 39931 19377 39943 19380
rect 39977 19377 39989 19411
rect 39931 19371 39989 19377
rect 1659 19343 1717 19349
rect 1659 19309 1671 19343
rect 1705 19340 1717 19343
rect 3315 19343 3373 19349
rect 1705 19312 2622 19340
rect 1705 19309 1717 19312
rect 1659 19303 1717 19309
rect 2594 19204 2622 19312
rect 3315 19309 3327 19343
rect 3361 19340 3373 19343
rect 3959 19343 4017 19349
rect 3959 19340 3971 19343
rect 3361 19312 3971 19340
rect 3361 19309 3373 19312
rect 3315 19303 3373 19309
rect 3959 19309 3971 19312
rect 4005 19340 4017 19343
rect 4140 19340 4146 19352
rect 4005 19312 4146 19340
rect 4005 19309 4017 19312
rect 3959 19303 4017 19309
rect 4140 19300 4146 19312
rect 4198 19300 4204 19352
rect 35420 19340 35426 19352
rect 35381 19312 35426 19340
rect 35420 19300 35426 19312
rect 35478 19300 35484 19352
rect 37628 19340 37634 19352
rect 37589 19312 37634 19340
rect 37628 19300 37634 19312
rect 37686 19300 37692 19352
rect 38183 19343 38241 19349
rect 38183 19309 38195 19343
rect 38229 19309 38241 19343
rect 38183 19303 38241 19309
rect 38367 19343 38425 19349
rect 38367 19309 38379 19343
rect 38413 19340 38425 19343
rect 38916 19340 38922 19352
rect 38413 19312 38922 19340
rect 38413 19309 38425 19312
rect 38367 19303 38425 19309
rect 36432 19232 36438 19284
rect 36490 19272 36496 19284
rect 38198 19272 38226 19303
rect 38916 19300 38922 19312
rect 38974 19340 38980 19352
rect 39026 19340 39054 19371
rect 38974 19312 39054 19340
rect 39839 19343 39897 19349
rect 38974 19300 38980 19312
rect 39839 19309 39851 19343
rect 39885 19340 39897 19343
rect 40572 19340 40578 19352
rect 39885 19312 40578 19340
rect 39885 19309 39897 19312
rect 39839 19303 39897 19309
rect 40572 19300 40578 19312
rect 40630 19300 40636 19352
rect 36490 19244 38226 19272
rect 38735 19275 38793 19281
rect 36490 19232 36496 19244
rect 38735 19241 38747 19275
rect 38781 19272 38793 19275
rect 39376 19272 39382 19284
rect 38781 19244 39382 19272
rect 38781 19241 38793 19244
rect 38735 19235 38793 19241
rect 39376 19232 39382 19244
rect 39434 19232 39440 19284
rect 3496 19204 3502 19216
rect 2594 19176 3502 19204
rect 3496 19164 3502 19176
rect 3554 19164 3560 19216
rect 34408 19204 34414 19216
rect 34369 19176 34414 19204
rect 34408 19164 34414 19176
rect 34466 19164 34472 19216
rect 538 19114 8450 19136
rect 538 19062 6344 19114
rect 6396 19062 6408 19114
rect 6460 19062 6472 19114
rect 6524 19062 6536 19114
rect 6588 19062 8450 19114
rect 538 19040 8450 19062
rect 34118 19114 43410 19136
rect 34118 19062 38312 19114
rect 38364 19062 38376 19114
rect 38428 19062 38440 19114
rect 38492 19062 38504 19114
rect 38556 19062 43410 19114
rect 34118 19040 43410 19062
rect 5891 19003 5949 19009
rect 5891 18969 5903 19003
rect 5937 19000 5949 19003
rect 5980 19000 5986 19012
rect 5937 18972 5986 19000
rect 5937 18969 5949 18972
rect 5891 18963 5949 18969
rect 5980 18960 5986 18972
rect 6038 18960 6044 19012
rect 39011 19003 39069 19009
rect 39011 18969 39023 19003
rect 39057 19000 39069 19003
rect 39652 19000 39658 19012
rect 39057 18972 39658 19000
rect 39057 18969 39069 18972
rect 39011 18963 39069 18969
rect 3315 18935 3373 18941
rect 3315 18901 3327 18935
rect 3361 18932 3373 18935
rect 4324 18932 4330 18944
rect 3361 18904 4330 18932
rect 3361 18901 3373 18904
rect 3315 18895 3373 18901
rect 3588 18824 3594 18876
rect 3646 18864 3652 18876
rect 3790 18873 3818 18904
rect 4324 18892 4330 18904
rect 4382 18892 4388 18944
rect 3683 18867 3741 18873
rect 3683 18864 3695 18867
rect 3646 18836 3695 18864
rect 3646 18824 3652 18836
rect 3683 18833 3695 18836
rect 3729 18833 3741 18867
rect 3683 18827 3741 18833
rect 3775 18867 3833 18873
rect 3775 18833 3787 18867
rect 3821 18833 3833 18867
rect 4235 18867 4293 18873
rect 4235 18864 4247 18867
rect 3775 18827 3833 18833
rect 3882 18836 4247 18864
rect 3698 18796 3726 18827
rect 3882 18796 3910 18836
rect 4235 18833 4247 18836
rect 4281 18833 4293 18867
rect 4416 18864 4422 18876
rect 4377 18836 4422 18864
rect 4235 18827 4293 18833
rect 4416 18824 4422 18836
rect 4474 18824 4480 18876
rect 5998 18873 6026 18960
rect 34886 18904 35190 18932
rect 5983 18867 6041 18873
rect 5983 18833 5995 18867
rect 6029 18833 6041 18867
rect 5983 18827 6041 18833
rect 6167 18867 6225 18873
rect 6167 18833 6179 18867
rect 6213 18864 6225 18867
rect 6719 18867 6777 18873
rect 6719 18864 6731 18867
rect 6213 18836 6731 18864
rect 6213 18833 6225 18836
rect 6167 18827 6225 18833
rect 6719 18833 6731 18836
rect 6765 18833 6777 18867
rect 6900 18864 6906 18876
rect 6861 18836 6906 18864
rect 6719 18827 6777 18833
rect 3698 18768 3910 18796
rect 3882 18660 3910 18768
rect 4600 18728 4606 18740
rect 4561 18700 4606 18728
rect 4600 18688 4606 18700
rect 4658 18688 4664 18740
rect 6182 18660 6210 18827
rect 6900 18824 6906 18836
rect 6958 18824 6964 18876
rect 34408 18864 34414 18876
rect 34369 18836 34414 18864
rect 34408 18824 34414 18836
rect 34466 18824 34472 18876
rect 34592 18873 34598 18876
rect 34580 18867 34598 18873
rect 34580 18833 34592 18867
rect 34650 18864 34656 18876
rect 34886 18864 34914 18904
rect 34650 18836 34914 18864
rect 34580 18827 34598 18833
rect 34592 18824 34598 18827
rect 34650 18824 34656 18836
rect 34960 18824 34966 18876
rect 35018 18864 35024 18876
rect 35162 18873 35190 18904
rect 35055 18867 35113 18873
rect 35055 18864 35067 18867
rect 35018 18836 35067 18864
rect 35018 18824 35024 18836
rect 35055 18833 35067 18836
rect 35101 18833 35113 18867
rect 35055 18827 35113 18833
rect 35147 18867 35205 18873
rect 35147 18833 35159 18867
rect 35193 18864 35205 18867
rect 37628 18864 37634 18876
rect 35193 18836 37634 18864
rect 35193 18833 35205 18836
rect 35147 18827 35205 18833
rect 37628 18824 37634 18836
rect 37686 18824 37692 18876
rect 39118 18873 39146 18972
rect 39652 18960 39658 18972
rect 39710 18960 39716 19012
rect 40572 18960 40578 19012
rect 40630 19000 40636 19012
rect 40667 19003 40725 19009
rect 40667 19000 40679 19003
rect 40630 18972 40679 19000
rect 40630 18960 40636 18972
rect 40667 18969 40679 18972
rect 40713 18969 40725 19003
rect 40667 18963 40725 18969
rect 39103 18867 39161 18873
rect 39103 18833 39115 18867
rect 39149 18833 39161 18867
rect 39376 18864 39382 18876
rect 39337 18836 39382 18864
rect 39103 18827 39161 18833
rect 39376 18824 39382 18836
rect 39434 18824 39440 18876
rect 7084 18728 7090 18740
rect 7045 18700 7090 18728
rect 7084 18688 7090 18700
rect 7142 18688 7148 18740
rect 35512 18728 35518 18740
rect 35473 18700 35518 18728
rect 35512 18688 35518 18700
rect 35570 18688 35576 18740
rect 3882 18632 6210 18660
rect 40682 18660 40710 18963
rect 70380 18824 70386 18876
rect 70438 18864 70444 18876
rect 70840 18864 70846 18876
rect 70438 18836 70846 18864
rect 70438 18824 70444 18836
rect 70840 18824 70846 18836
rect 70898 18824 70904 18876
rect 43332 18660 43338 18672
rect 40682 18632 43338 18660
rect 43332 18620 43338 18632
rect 43390 18620 43396 18672
rect 538 18570 8450 18592
rect 538 18518 3680 18570
rect 3732 18518 3744 18570
rect 3796 18518 3808 18570
rect 3860 18518 3872 18570
rect 3924 18518 8450 18570
rect 538 18496 8450 18518
rect 34118 18570 43410 18592
rect 34118 18518 35648 18570
rect 35700 18518 35712 18570
rect 35764 18518 35776 18570
rect 35828 18518 35840 18570
rect 35892 18518 40976 18570
rect 41028 18518 41040 18570
rect 41092 18518 41104 18570
rect 41156 18518 41168 18570
rect 41220 18518 43410 18570
rect 34118 18496 43410 18518
rect 6900 18416 6906 18468
rect 6958 18456 6964 18468
rect 7271 18459 7329 18465
rect 7271 18456 7283 18459
rect 6958 18428 7283 18456
rect 6958 18416 6964 18428
rect 7271 18425 7283 18428
rect 7317 18425 7329 18459
rect 36619 18459 36677 18465
rect 36619 18456 36631 18459
rect 7271 18419 7329 18425
rect 34794 18428 36631 18456
rect 3959 18323 4017 18329
rect 3959 18289 3971 18323
rect 4005 18320 4017 18323
rect 4600 18320 4606 18332
rect 4005 18292 4606 18320
rect 4005 18289 4017 18292
rect 3959 18283 4017 18289
rect 4600 18280 4606 18292
rect 4658 18280 4664 18332
rect 34794 18329 34822 18428
rect 36619 18425 36631 18428
rect 36665 18456 36677 18459
rect 36708 18456 36714 18468
rect 36665 18428 36714 18456
rect 36665 18425 36677 18428
rect 36619 18419 36677 18425
rect 36708 18416 36714 18428
rect 36766 18416 36772 18468
rect 39652 18416 39658 18468
rect 39710 18456 39716 18468
rect 40299 18459 40357 18465
rect 40299 18456 40311 18459
rect 39710 18428 40311 18456
rect 39710 18416 39716 18428
rect 40299 18425 40311 18428
rect 40345 18425 40357 18459
rect 40299 18419 40357 18425
rect 34779 18323 34837 18329
rect 34779 18289 34791 18323
rect 34825 18289 34837 18323
rect 34779 18283 34837 18289
rect 35055 18323 35113 18329
rect 35055 18289 35067 18323
rect 35101 18320 35113 18323
rect 35512 18320 35518 18332
rect 35101 18292 35518 18320
rect 35101 18289 35113 18292
rect 35055 18283 35113 18289
rect 35512 18280 35518 18292
rect 35570 18280 35576 18332
rect 40314 18320 40342 18419
rect 40483 18323 40541 18329
rect 40483 18320 40495 18323
rect 40314 18292 40495 18320
rect 40483 18289 40495 18292
rect 40529 18289 40541 18323
rect 43516 18320 43522 18332
rect 40483 18283 40541 18289
rect 40590 18292 43522 18320
rect 3496 18212 3502 18264
rect 3554 18252 3560 18264
rect 3683 18255 3741 18261
rect 3683 18252 3695 18255
rect 3554 18224 3695 18252
rect 3554 18212 3560 18224
rect 3683 18221 3695 18224
rect 3729 18252 3741 18255
rect 7179 18255 7237 18261
rect 3729 18224 5566 18252
rect 3729 18221 3741 18224
rect 3683 18215 3741 18221
rect 5538 18128 5566 18224
rect 7179 18221 7191 18255
rect 7225 18252 7237 18255
rect 7225 18224 7314 18252
rect 7225 18221 7237 18224
rect 7179 18215 7237 18221
rect 7286 18128 7314 18224
rect 35420 18212 35426 18264
rect 35478 18252 35484 18264
rect 35478 18224 36478 18252
rect 35478 18212 35484 18224
rect 36450 18193 36478 18224
rect 36435 18187 36493 18193
rect 36435 18153 36447 18187
rect 36481 18184 36493 18187
rect 40590 18184 40618 18292
rect 43516 18280 43522 18292
rect 43574 18280 43580 18332
rect 40756 18252 40762 18264
rect 40717 18224 40762 18252
rect 40756 18212 40762 18224
rect 40814 18212 40820 18264
rect 36481 18156 40618 18184
rect 36481 18153 36493 18156
rect 36435 18147 36493 18153
rect 5060 18116 5066 18128
rect 5021 18088 5066 18116
rect 5060 18076 5066 18088
rect 5118 18076 5124 18128
rect 5520 18116 5526 18128
rect 5481 18088 5526 18116
rect 5520 18076 5526 18088
rect 5578 18076 5584 18128
rect 7268 18076 7274 18128
rect 7326 18116 7332 18128
rect 7455 18119 7513 18125
rect 7455 18116 7467 18119
rect 7326 18088 7467 18116
rect 7326 18076 7332 18088
rect 7455 18085 7467 18088
rect 7501 18085 7513 18119
rect 34408 18116 34414 18128
rect 34369 18088 34414 18116
rect 7455 18079 7513 18085
rect 34408 18076 34414 18088
rect 34466 18076 34472 18128
rect 42044 18116 42050 18128
rect 42005 18088 42050 18116
rect 42044 18076 42050 18088
rect 42102 18076 42108 18128
rect 538 18026 8450 18048
rect 538 17974 6344 18026
rect 6396 17974 6408 18026
rect 6460 17974 6472 18026
rect 6524 17974 6536 18026
rect 6588 17974 8450 18026
rect 538 17952 8450 17974
rect 34118 18026 43410 18048
rect 34118 17974 38312 18026
rect 38364 17974 38376 18026
rect 38428 17974 38440 18026
rect 38492 17974 38504 18026
rect 38556 17974 43410 18026
rect 34118 17952 43410 17974
rect 4416 17872 4422 17924
rect 4474 17912 4480 17924
rect 4787 17915 4845 17921
rect 4787 17912 4799 17915
rect 4474 17884 4799 17912
rect 4474 17872 4480 17884
rect 4787 17881 4799 17884
rect 4833 17881 4845 17915
rect 4787 17875 4845 17881
rect 41035 17915 41093 17921
rect 41035 17881 41047 17915
rect 41081 17912 41093 17915
rect 42044 17912 42050 17924
rect 41081 17884 42050 17912
rect 41081 17881 41093 17884
rect 41035 17875 41093 17881
rect 40759 17847 40817 17853
rect 40759 17844 40771 17847
rect 39394 17816 40771 17844
rect 4695 17779 4753 17785
rect 4695 17745 4707 17779
rect 4741 17776 4753 17779
rect 5060 17776 5066 17788
rect 4741 17748 5066 17776
rect 4741 17745 4753 17748
rect 4695 17739 4753 17745
rect 5060 17736 5066 17748
rect 5118 17736 5124 17788
rect 5983 17779 6041 17785
rect 5983 17745 5995 17779
rect 6029 17776 6041 17779
rect 7084 17776 7090 17788
rect 6029 17748 7090 17776
rect 6029 17745 6041 17748
rect 5983 17739 6041 17745
rect 7084 17736 7090 17748
rect 7142 17736 7148 17788
rect 38088 17736 38094 17788
rect 38146 17776 38152 17788
rect 38643 17779 38701 17785
rect 38643 17776 38655 17779
rect 38146 17748 38655 17776
rect 38146 17736 38152 17748
rect 38643 17745 38655 17748
rect 38689 17776 38701 17779
rect 39192 17776 39198 17788
rect 38689 17748 39198 17776
rect 38689 17745 38701 17748
rect 38643 17739 38701 17745
rect 39192 17736 39198 17748
rect 39250 17736 39256 17788
rect 39394 17785 39422 17816
rect 40759 17813 40771 17816
rect 40805 17813 40817 17847
rect 40759 17807 40817 17813
rect 39379 17779 39437 17785
rect 39379 17745 39391 17779
rect 39425 17745 39437 17779
rect 40664 17776 40670 17788
rect 40577 17748 40670 17776
rect 39379 17739 39437 17745
rect 40664 17736 40670 17748
rect 40722 17776 40728 17788
rect 41050 17776 41078 17875
rect 42044 17872 42050 17884
rect 42102 17872 42108 17924
rect 40722 17748 41078 17776
rect 40722 17736 40728 17748
rect 5520 17668 5526 17720
rect 5578 17708 5584 17720
rect 5707 17711 5765 17717
rect 5707 17708 5719 17711
rect 5578 17680 5719 17708
rect 5578 17668 5584 17680
rect 5707 17677 5719 17680
rect 5753 17708 5765 17711
rect 6072 17708 6078 17720
rect 5753 17680 6078 17708
rect 5753 17677 5765 17680
rect 5707 17671 5765 17677
rect 6072 17668 6078 17680
rect 6130 17708 6136 17720
rect 6992 17708 6998 17720
rect 6130 17680 6998 17708
rect 6130 17668 6136 17680
rect 6992 17668 6998 17680
rect 7050 17708 7056 17720
rect 7455 17711 7513 17717
rect 7455 17708 7467 17711
rect 7050 17680 7467 17708
rect 7050 17668 7056 17680
rect 7455 17677 7467 17680
rect 7501 17677 7513 17711
rect 38459 17711 38517 17717
rect 38459 17708 38471 17711
rect 7455 17671 7513 17677
rect 38290 17680 38471 17708
rect 5060 17572 5066 17584
rect 5021 17544 5066 17572
rect 5060 17532 5066 17544
rect 5118 17532 5124 17584
rect 7268 17572 7274 17584
rect 7229 17544 7274 17572
rect 7268 17532 7274 17544
rect 7326 17532 7332 17584
rect 37536 17532 37542 17584
rect 37594 17572 37600 17584
rect 37996 17572 38002 17584
rect 37594 17544 38002 17572
rect 37594 17532 37600 17544
rect 37996 17532 38002 17544
rect 38054 17572 38060 17584
rect 38290 17581 38318 17680
rect 38459 17677 38471 17680
rect 38505 17677 38517 17711
rect 38459 17671 38517 17677
rect 39747 17711 39805 17717
rect 39747 17677 39759 17711
rect 39793 17708 39805 17711
rect 40756 17708 40762 17720
rect 39793 17680 40762 17708
rect 39793 17677 39805 17680
rect 39747 17671 39805 17677
rect 40756 17668 40762 17680
rect 40814 17668 40820 17720
rect 38275 17575 38333 17581
rect 38275 17572 38287 17575
rect 38054 17544 38287 17572
rect 38054 17532 38060 17544
rect 38275 17541 38287 17544
rect 38321 17541 38333 17575
rect 38275 17535 38333 17541
rect 538 17482 8450 17504
rect 538 17430 3680 17482
rect 3732 17430 3744 17482
rect 3796 17430 3808 17482
rect 3860 17430 3872 17482
rect 3924 17430 8450 17482
rect 538 17408 8450 17430
rect 34118 17482 43410 17504
rect 34118 17430 35648 17482
rect 35700 17430 35712 17482
rect 35764 17430 35776 17482
rect 35828 17430 35840 17482
rect 35892 17430 40976 17482
rect 41028 17430 41040 17482
rect 41092 17430 41104 17482
rect 41156 17430 41168 17482
rect 41220 17430 43410 17482
rect 34118 17408 43410 17430
rect 36708 17260 36714 17312
rect 36766 17300 36772 17312
rect 39744 17300 39750 17312
rect 36766 17272 39750 17300
rect 36766 17260 36772 17272
rect 39744 17260 39750 17272
rect 39802 17260 39808 17312
rect 37263 17235 37321 17241
rect 37263 17201 37275 17235
rect 37309 17232 37321 17235
rect 37352 17232 37358 17244
rect 37309 17204 37358 17232
rect 37309 17201 37321 17204
rect 37263 17195 37321 17201
rect 37352 17192 37358 17204
rect 37410 17192 37416 17244
rect 39192 17192 39198 17244
rect 39250 17232 39256 17244
rect 39250 17204 39974 17232
rect 39250 17192 39256 17204
rect 35975 17167 36033 17173
rect 35975 17133 35987 17167
rect 36021 17133 36033 17167
rect 35975 17127 36033 17133
rect 36159 17167 36217 17173
rect 36159 17133 36171 17167
rect 36205 17133 36217 17167
rect 36159 17127 36217 17133
rect 34408 17028 34414 17040
rect 34369 17000 34414 17028
rect 34408 16988 34414 17000
rect 34466 16988 34472 17040
rect 35883 17031 35941 17037
rect 35883 16997 35895 17031
rect 35929 17028 35941 17031
rect 35990 17028 36018 17127
rect 36174 17096 36202 17127
rect 36340 17124 36346 17176
rect 36398 17164 36404 17176
rect 36619 17167 36677 17173
rect 36619 17164 36631 17167
rect 36398 17136 36631 17164
rect 36398 17124 36404 17136
rect 36619 17133 36631 17136
rect 36665 17133 36677 17167
rect 36619 17127 36677 17133
rect 36711 17167 36769 17173
rect 36711 17133 36723 17167
rect 36757 17133 36769 17167
rect 38732 17164 38738 17176
rect 38693 17136 38738 17164
rect 36711 17127 36769 17133
rect 36432 17096 36438 17108
rect 36174 17068 36438 17096
rect 36432 17056 36438 17068
rect 36490 17096 36496 17108
rect 36726 17096 36754 17127
rect 38732 17124 38738 17136
rect 38790 17164 38796 17176
rect 39011 17167 39069 17173
rect 39011 17164 39023 17167
rect 38790 17136 39023 17164
rect 38790 17124 38796 17136
rect 39011 17133 39023 17136
rect 39057 17133 39069 17167
rect 39836 17164 39842 17176
rect 39797 17136 39842 17164
rect 39011 17127 39069 17133
rect 39836 17124 39842 17136
rect 39894 17124 39900 17176
rect 39946 17164 39974 17204
rect 40023 17167 40081 17173
rect 40023 17164 40035 17167
rect 39946 17136 40035 17164
rect 40023 17133 40035 17136
rect 40069 17164 40081 17167
rect 40575 17167 40633 17173
rect 40575 17164 40587 17167
rect 40069 17136 40587 17164
rect 40069 17133 40081 17136
rect 40023 17127 40081 17133
rect 40575 17133 40587 17136
rect 40621 17133 40633 17167
rect 40756 17164 40762 17176
rect 40717 17136 40762 17164
rect 40575 17127 40633 17133
rect 40756 17124 40762 17136
rect 40814 17124 40820 17176
rect 38824 17096 38830 17108
rect 36490 17068 36754 17096
rect 38785 17068 38830 17096
rect 36490 17056 36496 17068
rect 38824 17056 38830 17068
rect 38882 17056 38888 17108
rect 37720 17028 37726 17040
rect 35929 17000 37726 17028
rect 35929 16997 35941 17000
rect 35883 16991 35941 16997
rect 37720 16988 37726 17000
rect 37778 17028 37784 17040
rect 39563 17031 39621 17037
rect 39563 17028 39575 17031
rect 37778 17000 39575 17028
rect 37778 16988 37784 17000
rect 39563 16997 39575 17000
rect 39609 17028 39621 17031
rect 39836 17028 39842 17040
rect 39609 17000 39842 17028
rect 39609 16997 39621 17000
rect 39563 16991 39621 16997
rect 39836 16988 39842 17000
rect 39894 16988 39900 17040
rect 41032 17028 41038 17040
rect 40993 17000 41038 17028
rect 41032 16988 41038 17000
rect 41090 16988 41096 17040
rect 538 16938 8450 16960
rect 538 16886 6344 16938
rect 6396 16886 6408 16938
rect 6460 16886 6472 16938
rect 6524 16886 6536 16938
rect 6588 16886 8450 16938
rect 538 16864 8450 16886
rect 34118 16938 43410 16960
rect 34118 16886 38312 16938
rect 38364 16886 38376 16938
rect 38428 16886 38440 16938
rect 38492 16886 38504 16938
rect 38556 16886 43410 16938
rect 34118 16864 43410 16886
rect 4692 16784 4698 16836
rect 4750 16824 4756 16836
rect 5063 16827 5121 16833
rect 5063 16824 5075 16827
rect 4750 16796 5075 16824
rect 4750 16784 4756 16796
rect 5063 16793 5075 16796
rect 5109 16824 5121 16827
rect 5247 16827 5305 16833
rect 5247 16824 5259 16827
rect 5109 16796 5259 16824
rect 5109 16793 5121 16796
rect 5063 16787 5121 16793
rect 5247 16793 5259 16796
rect 5293 16824 5305 16827
rect 5293 16796 6394 16824
rect 5293 16793 5305 16796
rect 5247 16787 5305 16793
rect 5814 16697 5842 16796
rect 6366 16697 6394 16796
rect 36340 16784 36346 16836
rect 36398 16824 36404 16836
rect 37631 16827 37689 16833
rect 37631 16824 37643 16827
rect 36398 16796 37643 16824
rect 36398 16784 36404 16796
rect 37631 16793 37643 16796
rect 37677 16793 37689 16827
rect 37631 16787 37689 16793
rect 39744 16784 39750 16836
rect 39802 16824 39808 16836
rect 39839 16827 39897 16833
rect 39839 16824 39851 16827
rect 39802 16796 39851 16824
rect 39802 16784 39808 16796
rect 39839 16793 39851 16796
rect 39885 16793 39897 16827
rect 39839 16787 39897 16793
rect 5799 16691 5857 16697
rect 5799 16657 5811 16691
rect 5845 16657 5857 16691
rect 5799 16651 5857 16657
rect 6351 16691 6409 16697
rect 6351 16657 6363 16691
rect 6397 16657 6409 16691
rect 6351 16651 6409 16657
rect 6535 16691 6593 16697
rect 6535 16657 6547 16691
rect 6581 16688 6593 16691
rect 7176 16688 7182 16700
rect 6581 16660 7182 16688
rect 6581 16657 6593 16660
rect 6535 16651 6593 16657
rect 7176 16648 7182 16660
rect 7234 16648 7240 16700
rect 37539 16691 37597 16697
rect 37539 16657 37551 16691
rect 37585 16688 37597 16691
rect 38640 16688 38646 16700
rect 37585 16660 38646 16688
rect 37585 16657 37597 16660
rect 37539 16651 37597 16657
rect 38640 16648 38646 16660
rect 38698 16648 38704 16700
rect 38732 16648 38738 16700
rect 38790 16688 38796 16700
rect 40299 16691 40357 16697
rect 38790 16660 40158 16688
rect 38790 16648 38796 16660
rect 5523 16623 5581 16629
rect 5523 16589 5535 16623
rect 5569 16620 5581 16623
rect 5704 16620 5710 16632
rect 5569 16592 5710 16620
rect 5569 16589 5581 16592
rect 5523 16583 5581 16589
rect 5704 16580 5710 16592
rect 5762 16580 5768 16632
rect 39744 16580 39750 16632
rect 39802 16620 39808 16632
rect 40023 16623 40081 16629
rect 40023 16620 40035 16623
rect 39802 16592 40035 16620
rect 39802 16580 39808 16592
rect 40023 16589 40035 16592
rect 40069 16589 40081 16623
rect 40130 16620 40158 16660
rect 40299 16657 40311 16691
rect 40345 16688 40357 16691
rect 41032 16688 41038 16700
rect 40345 16660 41038 16688
rect 40345 16657 40357 16660
rect 40299 16651 40357 16657
rect 41032 16648 41038 16660
rect 41090 16648 41096 16700
rect 41676 16620 41682 16632
rect 40130 16592 41682 16620
rect 40023 16583 40081 16589
rect 41676 16580 41682 16592
rect 41734 16580 41740 16632
rect 6716 16552 6722 16564
rect 6677 16524 6722 16552
rect 6716 16512 6722 16524
rect 6774 16512 6780 16564
rect 538 16394 8450 16416
rect 538 16342 3680 16394
rect 3732 16342 3744 16394
rect 3796 16342 3808 16394
rect 3860 16342 3872 16394
rect 3924 16342 8450 16394
rect 538 16320 8450 16342
rect 34118 16394 43410 16416
rect 34118 16342 35648 16394
rect 35700 16342 35712 16394
rect 35764 16342 35776 16394
rect 35828 16342 35840 16394
rect 35892 16342 40976 16394
rect 41028 16342 41040 16394
rect 41092 16342 41104 16394
rect 41156 16342 41168 16394
rect 41220 16342 43410 16394
rect 34118 16320 43410 16342
rect 4692 16240 4698 16292
rect 4750 16280 4756 16292
rect 5431 16283 5489 16289
rect 5431 16280 5443 16283
rect 4750 16252 5443 16280
rect 4750 16240 4756 16252
rect 5431 16249 5443 16252
rect 5477 16280 5489 16283
rect 5615 16283 5673 16289
rect 5615 16280 5627 16283
rect 5477 16252 5627 16280
rect 5477 16249 5489 16252
rect 5431 16243 5489 16249
rect 5615 16249 5627 16252
rect 5661 16249 5673 16283
rect 36340 16280 36346 16292
rect 36301 16252 36346 16280
rect 5615 16243 5673 16249
rect 36340 16240 36346 16252
rect 36398 16280 36404 16292
rect 37996 16280 38002 16292
rect 36398 16252 38002 16280
rect 36398 16240 36404 16252
rect 3867 16215 3925 16221
rect 3867 16181 3879 16215
rect 3913 16212 3925 16215
rect 4876 16212 4882 16224
rect 3913 16184 4882 16212
rect 3913 16181 3925 16184
rect 3867 16175 3925 16181
rect 4066 16153 4094 16184
rect 4876 16172 4882 16184
rect 4934 16172 4940 16224
rect 36542 16153 36570 16252
rect 37996 16240 38002 16252
rect 38054 16240 38060 16292
rect 36726 16184 37674 16212
rect 4051 16147 4109 16153
rect 4051 16113 4063 16147
rect 4097 16113 4109 16147
rect 6535 16147 6593 16153
rect 6535 16144 6547 16147
rect 4051 16107 4109 16113
rect 5538 16116 6547 16144
rect 4143 16079 4201 16085
rect 4143 16045 4155 16079
rect 4189 16076 4201 16079
rect 4692 16076 4698 16088
rect 4189 16048 4698 16076
rect 4189 16045 4201 16048
rect 4143 16039 4201 16045
rect 4692 16036 4698 16048
rect 4750 16036 4756 16088
rect 4879 16079 4937 16085
rect 4879 16045 4891 16079
rect 4925 16076 4937 16079
rect 5538 16076 5566 16116
rect 6535 16113 6547 16116
rect 6581 16113 6593 16147
rect 6535 16107 6593 16113
rect 36527 16147 36585 16153
rect 36527 16113 36539 16147
rect 36573 16113 36585 16147
rect 36527 16107 36585 16113
rect 4925 16048 5566 16076
rect 6443 16079 6501 16085
rect 4925 16045 4937 16048
rect 4879 16039 4937 16045
rect 6443 16045 6455 16079
rect 6489 16076 6501 16079
rect 6489 16048 6854 16076
rect 6489 16045 6501 16048
rect 6443 16039 6501 16045
rect 5244 16008 5250 16020
rect 5205 15980 5250 16008
rect 5244 15968 5250 15980
rect 5302 15968 5308 16020
rect 6826 15949 6854 16048
rect 36432 16036 36438 16088
rect 36490 16076 36496 16088
rect 36726 16085 36754 16184
rect 36711 16079 36769 16085
rect 36711 16076 36723 16079
rect 36490 16048 36723 16076
rect 36490 16036 36496 16048
rect 36711 16045 36723 16048
rect 36757 16045 36769 16079
rect 37168 16076 37174 16088
rect 37129 16048 37174 16076
rect 36711 16039 36769 16045
rect 37168 16036 37174 16048
rect 37226 16036 37232 16088
rect 37263 16079 37321 16085
rect 37263 16045 37275 16079
rect 37309 16076 37321 16079
rect 37646 16076 37674 16184
rect 37309 16048 37674 16076
rect 38735 16079 38793 16085
rect 37309 16045 37321 16048
rect 37263 16039 37321 16045
rect 38735 16045 38747 16079
rect 38781 16076 38793 16079
rect 38916 16076 38922 16088
rect 38781 16048 38922 16076
rect 38781 16045 38793 16048
rect 38735 16039 38793 16045
rect 38916 16036 38922 16048
rect 38974 16036 38980 16088
rect 37186 16008 37214 16036
rect 38827 16011 38885 16017
rect 38827 16008 38839 16011
rect 37186 15980 38839 16008
rect 38827 15977 38839 15980
rect 38873 15977 38885 16011
rect 38827 15971 38885 15977
rect 6811 15943 6869 15949
rect 6811 15909 6823 15943
rect 6857 15940 6869 15943
rect 6992 15940 6998 15952
rect 6857 15912 6998 15940
rect 6857 15909 6869 15912
rect 6811 15903 6869 15909
rect 6992 15900 6998 15912
rect 7050 15900 7056 15952
rect 37720 15940 37726 15952
rect 37681 15912 37726 15940
rect 37720 15900 37726 15912
rect 37778 15900 37784 15952
rect 538 15850 8450 15872
rect 538 15798 6344 15850
rect 6396 15798 6408 15850
rect 6460 15798 6472 15850
rect 6524 15798 6536 15850
rect 6588 15798 8450 15850
rect 538 15776 8450 15798
rect 34118 15850 43410 15872
rect 34118 15798 38312 15850
rect 38364 15798 38376 15850
rect 38428 15798 38440 15850
rect 38492 15798 38504 15850
rect 38556 15798 43410 15850
rect 68356 15832 68362 15884
rect 68414 15872 68420 15884
rect 70472 15872 70478 15884
rect 68414 15844 70478 15872
rect 68414 15832 68420 15844
rect 70472 15832 70478 15844
rect 70530 15872 70536 15884
rect 71484 15872 71490 15884
rect 70530 15844 71490 15872
rect 70530 15832 70536 15844
rect 71484 15832 71490 15844
rect 71542 15832 71548 15884
rect 34118 15776 43410 15798
rect 36708 15696 36714 15748
rect 36766 15736 36772 15748
rect 36803 15739 36861 15745
rect 36803 15736 36815 15739
rect 36766 15708 36815 15736
rect 36766 15696 36772 15708
rect 36803 15705 36815 15708
rect 36849 15705 36861 15739
rect 36803 15699 36861 15705
rect 5244 15560 5250 15612
rect 5302 15600 5308 15612
rect 5707 15603 5765 15609
rect 5707 15600 5719 15603
rect 5302 15572 5719 15600
rect 5302 15560 5308 15572
rect 5707 15569 5719 15572
rect 5753 15569 5765 15603
rect 36818 15600 36846 15699
rect 37076 15600 37082 15612
rect 36818 15572 37082 15600
rect 5707 15563 5765 15569
rect 37076 15560 37082 15572
rect 37134 15560 37140 15612
rect 37352 15600 37358 15612
rect 37313 15572 37358 15600
rect 37352 15560 37358 15572
rect 37410 15560 37416 15612
rect 5431 15535 5489 15541
rect 5431 15501 5443 15535
rect 5477 15532 5489 15535
rect 6072 15532 6078 15544
rect 5477 15504 6078 15532
rect 5477 15501 5489 15504
rect 5431 15495 5489 15501
rect 6072 15492 6078 15504
rect 6130 15532 6136 15544
rect 7179 15535 7237 15541
rect 7179 15532 7191 15535
rect 6130 15504 7191 15532
rect 6130 15492 6136 15504
rect 7179 15501 7191 15504
rect 7225 15501 7237 15535
rect 7179 15495 7237 15501
rect 6992 15396 6998 15408
rect 6953 15368 6998 15396
rect 6992 15356 6998 15368
rect 7050 15356 7056 15408
rect 38640 15396 38646 15408
rect 38553 15368 38646 15396
rect 38640 15356 38646 15368
rect 38698 15396 38704 15408
rect 43516 15396 43522 15408
rect 38698 15368 43522 15396
rect 38698 15356 38704 15368
rect 43516 15356 43522 15368
rect 43574 15356 43580 15408
rect 538 15306 8450 15328
rect 538 15254 3680 15306
rect 3732 15254 3744 15306
rect 3796 15254 3808 15306
rect 3860 15254 3872 15306
rect 3924 15254 8450 15306
rect 538 15232 8450 15254
rect 34118 15306 43410 15328
rect 34118 15254 35648 15306
rect 35700 15254 35712 15306
rect 35764 15254 35776 15306
rect 35828 15254 35840 15306
rect 35892 15254 40976 15306
rect 41028 15254 41040 15306
rect 41092 15254 41104 15306
rect 41156 15254 41168 15306
rect 41220 15254 43410 15306
rect 34118 15232 43410 15254
rect 7176 15192 7182 15204
rect 7137 15164 7182 15192
rect 7176 15152 7182 15164
rect 7234 15152 7240 15204
rect 37076 15192 37082 15204
rect 37037 15164 37082 15192
rect 37076 15152 37082 15164
rect 37134 15152 37140 15204
rect 37094 15056 37122 15152
rect 37263 15059 37321 15065
rect 37263 15056 37275 15059
rect 37094 15028 37275 15056
rect 37263 15025 37275 15028
rect 37309 15025 37321 15059
rect 37263 15019 37321 15025
rect 37539 15059 37597 15065
rect 37539 15025 37551 15059
rect 37585 15056 37597 15059
rect 37720 15056 37726 15068
rect 37585 15028 37726 15056
rect 37585 15025 37597 15028
rect 37539 15019 37597 15025
rect 37720 15016 37726 15028
rect 37778 15016 37784 15068
rect 7087 14991 7145 14997
rect 7087 14957 7099 14991
rect 7133 14988 7145 14991
rect 7133 14960 7406 14988
rect 7133 14957 7145 14960
rect 7087 14951 7145 14957
rect 7378 14864 7406 14960
rect 38916 14920 38922 14932
rect 38877 14892 38922 14920
rect 38916 14880 38922 14892
rect 38974 14880 38980 14932
rect 7360 14852 7366 14864
rect 7321 14824 7366 14852
rect 7360 14812 7366 14824
rect 7418 14812 7424 14864
rect 34408 14852 34414 14864
rect 34369 14824 34414 14852
rect 34408 14812 34414 14824
rect 34466 14812 34472 14864
rect 538 14762 8450 14784
rect 538 14710 6344 14762
rect 6396 14710 6408 14762
rect 6460 14710 6472 14762
rect 6524 14710 6536 14762
rect 6588 14710 8450 14762
rect 538 14688 8450 14710
rect 34118 14762 43410 14784
rect 34118 14710 38312 14762
rect 38364 14710 38376 14762
rect 38428 14710 38440 14762
rect 38492 14710 38504 14762
rect 38556 14710 43410 14762
rect 34118 14688 43410 14710
rect 6072 14648 6078 14660
rect 5722 14620 6078 14648
rect 5722 14521 5750 14620
rect 6072 14608 6078 14620
rect 6130 14648 6136 14660
rect 7455 14651 7513 14657
rect 7455 14648 7467 14651
rect 6130 14620 7467 14648
rect 6130 14608 6136 14620
rect 7455 14617 7467 14620
rect 7501 14617 7513 14651
rect 7455 14611 7513 14617
rect 5707 14515 5765 14521
rect 5707 14481 5719 14515
rect 5753 14481 5765 14515
rect 5707 14475 5765 14481
rect 5983 14515 6041 14521
rect 5983 14481 5995 14515
rect 6029 14512 6041 14515
rect 6716 14512 6722 14524
rect 6029 14484 6722 14512
rect 6029 14481 6041 14484
rect 5983 14475 6041 14481
rect 6716 14472 6722 14484
rect 6774 14472 6780 14524
rect 7360 14512 7366 14524
rect 7321 14484 7366 14512
rect 7360 14472 7366 14484
rect 7418 14472 7424 14524
rect 538 14218 8450 14240
rect 538 14166 3680 14218
rect 3732 14166 3744 14218
rect 3796 14166 3808 14218
rect 3860 14166 3872 14218
rect 3924 14166 8450 14218
rect 538 14144 8450 14166
rect 34118 14218 43410 14240
rect 34118 14166 35648 14218
rect 35700 14166 35712 14218
rect 35764 14166 35776 14218
rect 35828 14166 35840 14218
rect 35892 14166 40976 14218
rect 41028 14166 41040 14218
rect 41092 14166 41104 14218
rect 41156 14166 41168 14218
rect 41220 14166 43410 14218
rect 34118 14144 43410 14166
rect 538 13674 8450 13696
rect 538 13622 6344 13674
rect 6396 13622 6408 13674
rect 6460 13622 6472 13674
rect 6524 13622 6536 13674
rect 6588 13622 8450 13674
rect 538 13600 8450 13622
rect 34118 13674 43410 13696
rect 34118 13622 38312 13674
rect 38364 13622 38376 13674
rect 38428 13622 38440 13674
rect 38492 13622 38504 13674
rect 38556 13622 43410 13674
rect 34118 13600 43410 13622
rect 538 13130 8450 13152
rect 538 13078 3680 13130
rect 3732 13078 3744 13130
rect 3796 13078 3808 13130
rect 3860 13078 3872 13130
rect 3924 13078 8450 13130
rect 538 13056 8450 13078
rect 34118 13130 43410 13152
rect 34118 13078 35648 13130
rect 35700 13078 35712 13130
rect 35764 13078 35776 13130
rect 35828 13078 35840 13130
rect 35892 13078 40976 13130
rect 41028 13078 41040 13130
rect 41092 13078 41104 13130
rect 41156 13078 41168 13130
rect 41220 13078 43410 13130
rect 34118 13056 43410 13078
rect 538 12586 8450 12608
rect 538 12534 6344 12586
rect 6396 12534 6408 12586
rect 6460 12534 6472 12586
rect 6524 12534 6536 12586
rect 6588 12534 8450 12586
rect 538 12512 8450 12534
rect 34118 12586 43410 12608
rect 34118 12534 38312 12586
rect 38364 12534 38376 12586
rect 38428 12534 38440 12586
rect 38492 12534 38504 12586
rect 38556 12534 43410 12586
rect 34118 12512 43410 12534
rect 538 12042 8450 12064
rect 538 11990 3680 12042
rect 3732 11990 3744 12042
rect 3796 11990 3808 12042
rect 3860 11990 3872 12042
rect 3924 11990 8450 12042
rect 538 11968 8450 11990
rect 34118 12042 43410 12064
rect 34118 11990 35648 12042
rect 35700 11990 35712 12042
rect 35764 11990 35776 12042
rect 35828 11990 35840 12042
rect 35892 11990 40976 12042
rect 41028 11990 41040 12042
rect 41092 11990 41104 12042
rect 41156 11990 41168 12042
rect 41220 11990 43410 12042
rect 34118 11968 43410 11990
rect 38916 11616 38922 11668
rect 38974 11656 38980 11668
rect 43516 11656 43522 11668
rect 38974 11628 43522 11656
rect 38974 11616 38980 11628
rect 43516 11616 43522 11628
rect 43574 11616 43580 11668
rect 538 11498 8450 11520
rect 538 11446 6344 11498
rect 6396 11446 6408 11498
rect 6460 11446 6472 11498
rect 6524 11446 6536 11498
rect 6588 11446 8450 11498
rect 538 11424 8450 11446
rect 34118 11498 43410 11520
rect 34118 11446 38312 11498
rect 38364 11446 38376 11498
rect 38428 11446 38440 11498
rect 38492 11446 38504 11498
rect 38556 11446 43410 11498
rect 34118 11424 43410 11446
rect 538 10954 8450 10976
rect 538 10902 3680 10954
rect 3732 10902 3744 10954
rect 3796 10902 3808 10954
rect 3860 10902 3872 10954
rect 3924 10902 8450 10954
rect 538 10880 8450 10902
rect 34118 10954 43410 10976
rect 34118 10902 35648 10954
rect 35700 10902 35712 10954
rect 35764 10902 35776 10954
rect 35828 10902 35840 10954
rect 35892 10902 40976 10954
rect 41028 10902 41040 10954
rect 41092 10902 41104 10954
rect 41156 10902 41168 10954
rect 41220 10902 43410 10954
rect 34118 10880 43410 10902
rect 34408 10500 34414 10512
rect 34369 10472 34414 10500
rect 34408 10460 34414 10472
rect 34466 10460 34472 10512
rect 538 10410 8450 10432
rect 538 10358 6344 10410
rect 6396 10358 6408 10410
rect 6460 10358 6472 10410
rect 6524 10358 6536 10410
rect 6588 10358 8450 10410
rect 538 10336 8450 10358
rect 34118 10410 43410 10432
rect 34118 10358 38312 10410
rect 38364 10358 38376 10410
rect 38428 10358 38440 10410
rect 38492 10358 38504 10410
rect 38556 10358 43410 10410
rect 34118 10336 43410 10358
rect 7547 10231 7605 10237
rect 7547 10197 7559 10231
rect 7593 10228 7605 10231
rect 11132 10228 11138 10240
rect 7593 10200 11138 10228
rect 7593 10197 7605 10200
rect 7547 10191 7605 10197
rect 5707 10163 5765 10169
rect 5707 10129 5719 10163
rect 5753 10160 5765 10163
rect 6072 10160 6078 10172
rect 5753 10132 6078 10160
rect 5753 10129 5765 10132
rect 5707 10123 5765 10129
rect 6072 10120 6078 10132
rect 6130 10160 6136 10172
rect 7639 10163 7697 10169
rect 7639 10160 7651 10163
rect 6130 10132 7651 10160
rect 6130 10120 6136 10132
rect 7639 10129 7651 10132
rect 7685 10129 7697 10163
rect 7639 10123 7697 10129
rect 5983 10095 6041 10101
rect 5983 10061 5995 10095
rect 6029 10092 6041 10095
rect 7746 10092 7774 10200
rect 11132 10188 11138 10200
rect 11190 10188 11196 10240
rect 6029 10064 7774 10092
rect 6029 10061 6041 10064
rect 5983 10055 6041 10061
rect 7084 9956 7090 9968
rect 7045 9928 7090 9956
rect 7084 9916 7090 9928
rect 7142 9916 7148 9968
rect 538 9866 8450 9888
rect 538 9814 3680 9866
rect 3732 9814 3744 9866
rect 3796 9814 3808 9866
rect 3860 9814 3872 9866
rect 3924 9814 8450 9866
rect 538 9792 8450 9814
rect 34118 9866 43410 9888
rect 34118 9814 35648 9866
rect 35700 9814 35712 9866
rect 35764 9814 35776 9866
rect 35828 9814 35840 9866
rect 35892 9814 40976 9866
rect 41028 9814 41040 9866
rect 41092 9814 41104 9866
rect 41156 9814 41168 9866
rect 41220 9814 43410 9866
rect 34118 9792 43410 9814
rect 538 9322 8450 9344
rect 538 9270 6344 9322
rect 6396 9270 6408 9322
rect 6460 9270 6472 9322
rect 6524 9270 6536 9322
rect 6588 9270 8450 9322
rect 538 9248 8450 9270
rect 34118 9322 43410 9344
rect 34118 9270 38312 9322
rect 38364 9270 38376 9322
rect 38428 9270 38440 9322
rect 38492 9270 38504 9322
rect 38556 9270 43410 9322
rect 34118 9248 43410 9270
rect 538 8778 8450 8800
rect 538 8726 3680 8778
rect 3732 8726 3744 8778
rect 3796 8726 3808 8778
rect 3860 8726 3872 8778
rect 3924 8726 8450 8778
rect 538 8704 8450 8726
rect 34118 8778 43410 8800
rect 34118 8726 35648 8778
rect 35700 8726 35712 8778
rect 35764 8726 35776 8778
rect 35828 8726 35840 8778
rect 35892 8726 40976 8778
rect 41028 8726 41040 8778
rect 41092 8726 41104 8778
rect 41156 8726 41168 8778
rect 41220 8726 43410 8778
rect 34118 8704 43410 8726
rect 538 8234 8450 8256
rect 538 8182 6344 8234
rect 6396 8182 6408 8234
rect 6460 8182 6472 8234
rect 6524 8182 6536 8234
rect 6588 8182 8450 8234
rect 538 8160 8450 8182
rect 34118 8234 43410 8256
rect 34118 8182 38312 8234
rect 38364 8182 38376 8234
rect 38428 8182 38440 8234
rect 38492 8182 38504 8234
rect 38556 8182 43410 8234
rect 34118 8160 43410 8182
rect 538 7690 8450 7712
rect 538 7638 3680 7690
rect 3732 7638 3744 7690
rect 3796 7638 3808 7690
rect 3860 7638 3872 7690
rect 3924 7638 8450 7690
rect 538 7616 8450 7638
rect 34118 7690 43410 7712
rect 34118 7638 35648 7690
rect 35700 7638 35712 7690
rect 35764 7638 35776 7690
rect 35828 7638 35840 7690
rect 35892 7638 40976 7690
rect 41028 7638 41040 7690
rect 41092 7638 41104 7690
rect 41156 7638 41168 7690
rect 41220 7638 43410 7690
rect 34118 7616 43410 7638
rect 538 7146 8450 7168
rect 538 7094 6344 7146
rect 6396 7094 6408 7146
rect 6460 7094 6472 7146
rect 6524 7094 6536 7146
rect 6588 7094 8450 7146
rect 538 7072 8450 7094
rect 34118 7146 43410 7168
rect 34118 7094 38312 7146
rect 38364 7094 38376 7146
rect 38428 7094 38440 7146
rect 38492 7094 38504 7146
rect 38556 7094 43410 7146
rect 34118 7072 43410 7094
rect 538 6602 8450 6624
rect 538 6550 3680 6602
rect 3732 6550 3744 6602
rect 3796 6550 3808 6602
rect 3860 6550 3872 6602
rect 3924 6550 8450 6602
rect 538 6528 8450 6550
rect 34118 6602 43410 6624
rect 34118 6550 35648 6602
rect 35700 6550 35712 6602
rect 35764 6550 35776 6602
rect 35828 6550 35840 6602
rect 35892 6550 40976 6602
rect 41028 6550 41040 6602
rect 41092 6550 41104 6602
rect 41156 6550 41168 6602
rect 41220 6550 43410 6602
rect 34118 6528 43410 6550
rect 538 6058 8450 6080
rect 538 6006 6344 6058
rect 6396 6006 6408 6058
rect 6460 6006 6472 6058
rect 6524 6006 6536 6058
rect 6588 6006 8450 6058
rect 538 5984 8450 6006
rect 34118 6058 43410 6080
rect 34118 6006 38312 6058
rect 38364 6006 38376 6058
rect 38428 6006 38440 6058
rect 38492 6006 38504 6058
rect 38556 6006 43410 6058
rect 34118 5984 43410 6006
rect 538 5514 8450 5536
rect 538 5462 3680 5514
rect 3732 5462 3744 5514
rect 3796 5462 3808 5514
rect 3860 5462 3872 5514
rect 3924 5462 8450 5514
rect 538 5440 8450 5462
rect 34118 5514 43410 5536
rect 34118 5462 35648 5514
rect 35700 5462 35712 5514
rect 35764 5462 35776 5514
rect 35828 5462 35840 5514
rect 35892 5462 40976 5514
rect 41028 5462 41040 5514
rect 41092 5462 41104 5514
rect 41156 5462 41168 5514
rect 41220 5462 43410 5514
rect 34118 5440 43410 5462
rect 538 4970 8450 4992
rect 538 4918 6344 4970
rect 6396 4918 6408 4970
rect 6460 4918 6472 4970
rect 6524 4918 6536 4970
rect 6588 4918 8450 4970
rect 538 4896 8450 4918
rect 34118 4970 43410 4992
rect 34118 4918 38312 4970
rect 38364 4918 38376 4970
rect 38428 4918 38440 4970
rect 38492 4918 38504 4970
rect 38556 4918 43410 4970
rect 34118 4896 43410 4918
rect 538 4426 8450 4448
rect 538 4374 3680 4426
rect 3732 4374 3744 4426
rect 3796 4374 3808 4426
rect 3860 4374 3872 4426
rect 3924 4374 8450 4426
rect 538 4352 8450 4374
rect 34118 4426 43410 4448
rect 34118 4374 35648 4426
rect 35700 4374 35712 4426
rect 35764 4374 35776 4426
rect 35828 4374 35840 4426
rect 35892 4374 40976 4426
rect 41028 4374 41040 4426
rect 41092 4374 41104 4426
rect 41156 4374 41168 4426
rect 41220 4374 43410 4426
rect 34118 4352 43410 4374
rect 538 3882 8450 3904
rect 538 3830 6344 3882
rect 6396 3830 6408 3882
rect 6460 3830 6472 3882
rect 6524 3830 6536 3882
rect 6588 3830 8450 3882
rect 538 3808 8450 3830
rect 34118 3882 43410 3904
rect 34118 3830 38312 3882
rect 38364 3830 38376 3882
rect 38428 3830 38440 3882
rect 38492 3830 38504 3882
rect 38556 3830 43410 3882
rect 34118 3808 43410 3830
rect 538 3338 8450 3360
rect 538 3286 3680 3338
rect 3732 3286 3744 3338
rect 3796 3286 3808 3338
rect 3860 3286 3872 3338
rect 3924 3286 8450 3338
rect 538 3264 8450 3286
rect 34118 3338 43410 3360
rect 34118 3286 35648 3338
rect 35700 3286 35712 3338
rect 35764 3286 35776 3338
rect 35828 3286 35840 3338
rect 35892 3286 40976 3338
rect 41028 3286 41040 3338
rect 41092 3286 41104 3338
rect 41156 3286 41168 3338
rect 41220 3286 43410 3338
rect 34118 3264 43410 3286
rect 538 2794 8450 2816
rect 538 2742 6344 2794
rect 6396 2742 6408 2794
rect 6460 2742 6472 2794
rect 6524 2742 6536 2794
rect 6588 2742 8450 2794
rect 538 2720 8450 2742
rect 34118 2794 43410 2816
rect 34118 2742 38312 2794
rect 38364 2742 38376 2794
rect 38428 2742 38440 2794
rect 38492 2742 38504 2794
rect 38556 2742 43410 2794
rect 34118 2720 43410 2742
rect 43059 2683 43117 2689
rect 43059 2649 43071 2683
rect 43105 2680 43117 2683
rect 43240 2680 43246 2692
rect 43105 2652 43246 2680
rect 43105 2649 43117 2652
rect 43059 2643 43117 2649
rect 43240 2640 43246 2652
rect 43298 2640 43304 2692
rect 31372 2300 31378 2352
rect 31430 2340 31436 2352
rect 34411 2343 34469 2349
rect 34411 2340 34423 2343
rect 31430 2312 34423 2340
rect 31430 2300 31436 2312
rect 34411 2309 34423 2312
rect 34457 2309 34469 2343
rect 34411 2303 34469 2309
rect 538 2250 8450 2272
rect 538 2198 3680 2250
rect 3732 2198 3744 2250
rect 3796 2198 3808 2250
rect 3860 2198 3872 2250
rect 3924 2198 8450 2250
rect 538 2176 8450 2198
rect 34118 2250 43410 2272
rect 34118 2198 35648 2250
rect 35700 2198 35712 2250
rect 35764 2198 35776 2250
rect 35828 2198 35840 2250
rect 35892 2198 40976 2250
rect 41028 2198 41040 2250
rect 41092 2198 41104 2250
rect 41156 2198 41168 2250
rect 41220 2198 43410 2250
rect 34118 2176 43410 2198
rect 7084 2096 7090 2148
rect 7142 2136 7148 2148
rect 31372 2136 31378 2148
rect 7142 2108 31378 2136
rect 7142 2096 7148 2108
rect 31372 2096 31378 2108
rect 31430 2096 31436 2148
rect 538 1706 8450 1728
rect 538 1654 6344 1706
rect 6396 1654 6408 1706
rect 6460 1654 6472 1706
rect 6524 1654 6536 1706
rect 6588 1654 8450 1706
rect 538 1632 8450 1654
rect 34118 1706 43410 1728
rect 34118 1654 38312 1706
rect 38364 1654 38376 1706
rect 38428 1654 38440 1706
rect 38492 1654 38504 1706
rect 38556 1654 43410 1706
rect 34118 1632 43410 1654
rect 538 1162 8450 1184
rect 538 1110 3680 1162
rect 3732 1110 3744 1162
rect 3796 1110 3808 1162
rect 3860 1110 3872 1162
rect 3924 1110 8450 1162
rect 538 1088 8450 1110
rect 34118 1162 43410 1184
rect 34118 1110 35648 1162
rect 35700 1110 35712 1162
rect 35764 1110 35776 1162
rect 35828 1110 35840 1162
rect 35892 1110 40976 1162
rect 41028 1110 41040 1162
rect 41092 1110 41104 1162
rect 41156 1110 41168 1162
rect 41220 1110 43410 1162
rect 34118 1088 43410 1110
rect 538 618 8450 640
rect 538 566 6344 618
rect 6396 566 6408 618
rect 6460 566 6472 618
rect 6524 566 6536 618
rect 6588 566 8450 618
rect 538 544 8450 566
rect 34118 618 43410 640
rect 34118 566 38312 618
rect 38364 566 38376 618
rect 38428 566 38440 618
rect 38492 566 38504 618
rect 38556 566 43410 618
rect 34118 544 43410 566
rect 538 74 8450 96
rect 538 22 3680 74
rect 3732 22 3744 74
rect 3796 22 3808 74
rect 3860 22 3872 74
rect 3924 22 8450 74
rect 538 0 8450 22
rect 34118 74 43410 96
rect 34118 22 35648 74
rect 35700 22 35712 74
rect 35764 22 35776 74
rect 35828 22 35840 74
rect 35892 22 40976 74
rect 41028 22 41040 74
rect 41092 22 41104 74
rect 41156 22 41168 74
rect 41220 22 43410 74
rect 34118 0 43410 22
<< via1 >>
rect 6344 41910 6396 41962
rect 6408 41910 6460 41962
rect 6472 41910 6524 41962
rect 6536 41910 6588 41962
rect 11672 41910 11724 41962
rect 11736 41910 11788 41962
rect 11800 41910 11852 41962
rect 11864 41910 11916 41962
rect 17000 41910 17052 41962
rect 17064 41910 17116 41962
rect 17128 41910 17180 41962
rect 17192 41910 17244 41962
rect 22328 41910 22380 41962
rect 22392 41910 22444 41962
rect 22456 41910 22508 41962
rect 22520 41910 22572 41962
rect 27656 41910 27708 41962
rect 27720 41910 27772 41962
rect 27784 41910 27836 41962
rect 27848 41910 27900 41962
rect 32984 41910 33036 41962
rect 33048 41910 33100 41962
rect 33112 41910 33164 41962
rect 33176 41910 33228 41962
rect 38312 41910 38364 41962
rect 38376 41910 38428 41962
rect 38440 41910 38492 41962
rect 38504 41910 38556 41962
rect 43640 41910 43692 41962
rect 43704 41910 43756 41962
rect 43768 41910 43820 41962
rect 43832 41910 43884 41962
rect 48968 41910 49020 41962
rect 49032 41910 49084 41962
rect 49096 41910 49148 41962
rect 49160 41910 49212 41962
rect 54296 41910 54348 41962
rect 54360 41910 54412 41962
rect 54424 41910 54476 41962
rect 54488 41910 54540 41962
rect 59624 41910 59676 41962
rect 59688 41910 59740 41962
rect 59752 41910 59804 41962
rect 59816 41910 59868 41962
rect 64952 41910 65004 41962
rect 65016 41910 65068 41962
rect 65080 41910 65132 41962
rect 65144 41910 65196 41962
rect 70280 41910 70332 41962
rect 70344 41910 70396 41962
rect 70408 41910 70460 41962
rect 70472 41910 70524 41962
rect 75608 41910 75660 41962
rect 75672 41910 75724 41962
rect 75736 41910 75788 41962
rect 75800 41910 75852 41962
rect 80936 41910 80988 41962
rect 81000 41910 81052 41962
rect 81064 41910 81116 41962
rect 81128 41910 81180 41962
rect 86264 41910 86316 41962
rect 86328 41910 86380 41962
rect 86392 41910 86444 41962
rect 86456 41910 86508 41962
rect 91592 41910 91644 41962
rect 91656 41910 91708 41962
rect 91720 41910 91772 41962
rect 91784 41910 91836 41962
rect 65326 41604 65378 41656
rect 68546 41604 68598 41656
rect 88142 41604 88194 41656
rect 89338 41647 89390 41656
rect 89338 41613 89347 41647
rect 89347 41613 89381 41647
rect 89381 41613 89390 41647
rect 89338 41604 89390 41613
rect 3502 41468 3554 41520
rect 20614 41468 20666 41520
rect 67442 41468 67494 41520
rect 73238 41468 73290 41520
rect 3680 41366 3732 41418
rect 3744 41366 3796 41418
rect 3808 41366 3860 41418
rect 3872 41366 3924 41418
rect 9008 41366 9060 41418
rect 9072 41366 9124 41418
rect 9136 41366 9188 41418
rect 9200 41366 9252 41418
rect 14336 41366 14388 41418
rect 14400 41366 14452 41418
rect 14464 41366 14516 41418
rect 14528 41366 14580 41418
rect 19664 41366 19716 41418
rect 19728 41366 19780 41418
rect 19792 41366 19844 41418
rect 19856 41366 19908 41418
rect 24992 41366 25044 41418
rect 25056 41366 25108 41418
rect 25120 41366 25172 41418
rect 25184 41366 25236 41418
rect 30320 41366 30372 41418
rect 30384 41366 30436 41418
rect 30448 41366 30500 41418
rect 30512 41366 30564 41418
rect 35648 41366 35700 41418
rect 35712 41366 35764 41418
rect 35776 41366 35828 41418
rect 35840 41366 35892 41418
rect 40976 41366 41028 41418
rect 41040 41366 41092 41418
rect 41104 41366 41156 41418
rect 41168 41366 41220 41418
rect 46304 41366 46356 41418
rect 46368 41366 46420 41418
rect 46432 41366 46484 41418
rect 46496 41366 46548 41418
rect 51632 41366 51684 41418
rect 51696 41366 51748 41418
rect 51760 41366 51812 41418
rect 51824 41366 51876 41418
rect 56960 41366 57012 41418
rect 57024 41366 57076 41418
rect 57088 41366 57140 41418
rect 57152 41366 57204 41418
rect 62288 41366 62340 41418
rect 62352 41366 62404 41418
rect 62416 41366 62468 41418
rect 62480 41366 62532 41418
rect 67616 41366 67668 41418
rect 67680 41366 67732 41418
rect 67744 41366 67796 41418
rect 67808 41366 67860 41418
rect 72944 41366 72996 41418
rect 73008 41366 73060 41418
rect 73072 41366 73124 41418
rect 73136 41366 73188 41418
rect 78272 41366 78324 41418
rect 78336 41366 78388 41418
rect 78400 41366 78452 41418
rect 78464 41366 78516 41418
rect 83600 41366 83652 41418
rect 83664 41366 83716 41418
rect 83728 41366 83780 41418
rect 83792 41366 83844 41418
rect 88928 41366 88980 41418
rect 88992 41366 89044 41418
rect 89056 41366 89108 41418
rect 89120 41366 89172 41418
rect 2398 41264 2450 41316
rect 3502 41307 3554 41316
rect 3502 41273 3511 41307
rect 3511 41273 3545 41307
rect 3545 41273 3554 41307
rect 3502 41264 3554 41273
rect 17394 41264 17446 41316
rect 24386 41264 24438 41316
rect 27054 41264 27106 41316
rect 31746 41264 31798 41316
rect 48858 41264 48910 41316
rect 53734 41264 53786 41316
rect 3502 41060 3554 41112
rect 4606 41103 4658 41112
rect 4606 41069 4615 41103
rect 4615 41069 4649 41103
rect 4649 41069 4658 41103
rect 4606 41060 4658 41069
rect 6170 41060 6222 41112
rect 12334 41103 12386 41112
rect 12334 41069 12343 41103
rect 12343 41069 12377 41103
rect 12377 41069 12386 41103
rect 12334 41060 12386 41069
rect 37082 41128 37134 41180
rect 13070 40992 13122 41044
rect 7826 40967 7878 40976
rect 7826 40933 7835 40967
rect 7835 40933 7869 40967
rect 7869 40933 7878 40967
rect 7826 40924 7878 40933
rect 8010 40967 8062 40976
rect 8010 40933 8019 40967
rect 8019 40933 8053 40967
rect 8053 40933 8062 40967
rect 8010 40924 8062 40933
rect 13438 40967 13490 40976
rect 13438 40933 13447 40967
rect 13447 40933 13481 40967
rect 13481 40933 13490 40967
rect 13438 40924 13490 40933
rect 17762 41103 17814 41112
rect 17762 41069 17771 41103
rect 17771 41069 17805 41103
rect 17805 41069 17814 41103
rect 17762 41060 17814 41069
rect 14910 40924 14962 40976
rect 17394 40924 17446 40976
rect 20890 40924 20942 40976
rect 25674 41060 25726 41112
rect 28434 41060 28486 41112
rect 28802 41060 28854 41112
rect 32758 41060 32810 41112
rect 36346 41103 36398 41112
rect 36346 41069 36355 41103
rect 36355 41069 36389 41103
rect 36389 41069 36398 41103
rect 36346 41060 36398 41069
rect 26778 40924 26830 40976
rect 28526 40924 28578 40976
rect 29354 40924 29406 40976
rect 30458 40967 30510 40976
rect 30458 40933 30467 40967
rect 30467 40933 30501 40967
rect 30501 40933 30510 40967
rect 30458 40924 30510 40933
rect 31562 40924 31614 40976
rect 32758 40924 32810 40976
rect 40854 41060 40906 41112
rect 50790 41128 50842 41180
rect 52538 41128 52590 41180
rect 61094 41264 61146 41316
rect 83082 41264 83134 41316
rect 47110 41103 47162 41112
rect 37542 40967 37594 40976
rect 37542 40933 37551 40967
rect 37551 40933 37585 40967
rect 37585 40933 37594 40967
rect 37542 40924 37594 40933
rect 47110 41069 47119 41103
rect 47119 41069 47153 41103
rect 47153 41069 47162 41103
rect 47110 41060 47162 41069
rect 47386 41103 47438 41112
rect 47386 41069 47395 41103
rect 47395 41069 47429 41103
rect 47429 41069 47438 41103
rect 47386 41060 47438 41069
rect 51066 41060 51118 41112
rect 51434 41103 51486 41112
rect 44074 40992 44126 41044
rect 46742 40924 46794 40976
rect 47110 40924 47162 40976
rect 49502 40924 49554 40976
rect 51434 41069 51443 41103
rect 51443 41069 51477 41103
rect 51477 41069 51486 41103
rect 51434 41060 51486 41069
rect 54654 41103 54706 41112
rect 54654 41069 54663 41103
rect 54663 41069 54697 41103
rect 54697 41069 54706 41103
rect 54654 41060 54706 41069
rect 56034 41060 56086 41112
rect 56770 41103 56822 41112
rect 56770 41069 56779 41103
rect 56779 41069 56813 41103
rect 56813 41069 56822 41103
rect 56770 41060 56822 41069
rect 60266 41103 60318 41112
rect 60266 41069 60275 41103
rect 60275 41069 60309 41103
rect 60309 41069 60318 41103
rect 60266 41060 60318 41069
rect 55574 40924 55626 40976
rect 55850 40924 55902 40976
rect 56678 40924 56730 40976
rect 58058 40924 58110 40976
rect 58702 40924 58754 40976
rect 61738 41060 61790 41112
rect 65326 41060 65378 41112
rect 73698 41060 73750 41112
rect 73882 41103 73934 41112
rect 73882 41069 73891 41103
rect 73891 41069 73925 41103
rect 73925 41069 73934 41103
rect 73882 41060 73934 41069
rect 79494 41060 79546 41112
rect 81150 41060 81202 41112
rect 83634 41128 83686 41180
rect 81426 41060 81478 41112
rect 85658 41103 85710 41112
rect 61738 40924 61790 40976
rect 63578 40924 63630 40976
rect 75998 40924 76050 40976
rect 85014 40924 85066 40976
rect 85658 41069 85667 41103
rect 85667 41069 85701 41103
rect 85701 41069 85710 41103
rect 85658 41060 85710 41069
rect 88142 40924 88194 40976
rect 6344 40822 6396 40874
rect 6408 40822 6460 40874
rect 6472 40822 6524 40874
rect 6536 40822 6588 40874
rect 11672 40822 11724 40874
rect 11736 40822 11788 40874
rect 11800 40822 11852 40874
rect 11864 40822 11916 40874
rect 17000 40822 17052 40874
rect 17064 40822 17116 40874
rect 17128 40822 17180 40874
rect 17192 40822 17244 40874
rect 22328 40822 22380 40874
rect 22392 40822 22444 40874
rect 22456 40822 22508 40874
rect 22520 40822 22572 40874
rect 27656 40822 27708 40874
rect 27720 40822 27772 40874
rect 27784 40822 27836 40874
rect 27848 40822 27900 40874
rect 32984 40822 33036 40874
rect 33048 40822 33100 40874
rect 33112 40822 33164 40874
rect 33176 40822 33228 40874
rect 38312 40822 38364 40874
rect 38376 40822 38428 40874
rect 38440 40822 38492 40874
rect 38504 40822 38556 40874
rect 43640 40822 43692 40874
rect 43704 40822 43756 40874
rect 43768 40822 43820 40874
rect 43832 40822 43884 40874
rect 48968 40822 49020 40874
rect 49032 40822 49084 40874
rect 49096 40822 49148 40874
rect 49160 40822 49212 40874
rect 54296 40822 54348 40874
rect 54360 40822 54412 40874
rect 54424 40822 54476 40874
rect 54488 40822 54540 40874
rect 59624 40822 59676 40874
rect 59688 40822 59740 40874
rect 59752 40822 59804 40874
rect 59816 40822 59868 40874
rect 64952 40822 65004 40874
rect 65016 40822 65068 40874
rect 65080 40822 65132 40874
rect 65144 40822 65196 40874
rect 70280 40822 70332 40874
rect 70344 40822 70396 40874
rect 70408 40822 70460 40874
rect 70472 40822 70524 40874
rect 75608 40822 75660 40874
rect 75672 40822 75724 40874
rect 75736 40822 75788 40874
rect 75800 40822 75852 40874
rect 80936 40822 80988 40874
rect 81000 40822 81052 40874
rect 81064 40822 81116 40874
rect 81128 40822 81180 40874
rect 86264 40822 86316 40874
rect 86328 40822 86380 40874
rect 86392 40822 86444 40874
rect 86456 40822 86508 40874
rect 91592 40822 91644 40874
rect 91656 40822 91708 40874
rect 91720 40822 91772 40874
rect 91784 40822 91836 40874
rect 3502 40720 3554 40772
rect 6170 40720 6222 40772
rect 14910 40720 14962 40772
rect 29262 40720 29314 40772
rect 17394 40652 17446 40704
rect 28526 40695 28578 40704
rect 28526 40661 28535 40695
rect 28535 40661 28569 40695
rect 28569 40661 28578 40695
rect 28526 40652 28578 40661
rect 6 40584 58 40636
rect 3502 40627 3554 40636
rect 3502 40593 3511 40627
rect 3511 40593 3545 40627
rect 3545 40593 3554 40627
rect 3502 40584 3554 40593
rect 4054 40584 4106 40636
rect 5066 40584 5118 40636
rect 2490 40423 2542 40432
rect 2490 40389 2499 40423
rect 2499 40389 2533 40423
rect 2533 40389 2542 40423
rect 2490 40380 2542 40389
rect 4882 40516 4934 40568
rect 4606 40448 4658 40500
rect 6170 40516 6222 40568
rect 8010 40584 8062 40636
rect 9758 40584 9810 40636
rect 13438 40584 13490 40636
rect 14634 40584 14686 40636
rect 7366 40516 7418 40568
rect 11046 40559 11098 40568
rect 11046 40525 11055 40559
rect 11055 40525 11089 40559
rect 11089 40525 11098 40559
rect 11046 40516 11098 40525
rect 14174 40516 14226 40568
rect 14910 40559 14962 40568
rect 14910 40525 14919 40559
rect 14919 40525 14953 40559
rect 14953 40525 14962 40559
rect 14910 40516 14962 40525
rect 5342 40423 5394 40432
rect 5342 40389 5351 40423
rect 5351 40389 5385 40423
rect 5385 40389 5394 40423
rect 5342 40380 5394 40389
rect 8010 40423 8062 40432
rect 8010 40389 8019 40423
rect 8019 40389 8053 40423
rect 8053 40389 8062 40423
rect 8010 40380 8062 40389
rect 12150 40448 12202 40500
rect 13070 40380 13122 40432
rect 17394 40559 17446 40568
rect 17394 40525 17403 40559
rect 17403 40525 17437 40559
rect 17437 40525 17446 40559
rect 17394 40516 17446 40525
rect 17670 40559 17722 40568
rect 17670 40525 17679 40559
rect 17679 40525 17713 40559
rect 17713 40525 17722 40559
rect 17670 40516 17722 40525
rect 25674 40584 25726 40636
rect 26778 40627 26830 40636
rect 26778 40593 26787 40627
rect 26787 40593 26821 40627
rect 26821 40593 26830 40627
rect 26778 40584 26830 40593
rect 30458 40584 30510 40636
rect 21258 40559 21310 40568
rect 21258 40525 21267 40559
rect 21267 40525 21301 40559
rect 21301 40525 21310 40559
rect 21258 40516 21310 40525
rect 21994 40516 22046 40568
rect 27054 40559 27106 40568
rect 27054 40525 27063 40559
rect 27063 40525 27097 40559
rect 27097 40525 27106 40559
rect 27054 40516 27106 40525
rect 32298 40516 32350 40568
rect 34138 40584 34190 40636
rect 36622 40584 36674 40636
rect 37542 40584 37594 40636
rect 39106 40584 39158 40636
rect 41498 40584 41550 40636
rect 44074 40584 44126 40636
rect 47110 40720 47162 40772
rect 51066 40652 51118 40704
rect 56770 40652 56822 40704
rect 49502 40627 49554 40636
rect 49502 40593 49511 40627
rect 49511 40593 49545 40627
rect 49545 40593 49554 40627
rect 49502 40584 49554 40593
rect 51250 40584 51302 40636
rect 55574 40627 55626 40636
rect 55574 40593 55583 40627
rect 55583 40593 55617 40627
rect 55617 40593 55626 40627
rect 55574 40584 55626 40593
rect 56126 40584 56178 40636
rect 57322 40584 57374 40636
rect 58058 40627 58110 40636
rect 58058 40593 58067 40627
rect 58067 40593 58101 40627
rect 58101 40593 58110 40627
rect 58058 40584 58110 40593
rect 58702 40584 58754 40636
rect 61646 40584 61698 40636
rect 62658 40584 62710 40636
rect 62934 40584 62986 40636
rect 63578 40627 63630 40636
rect 63578 40593 63587 40627
rect 63587 40593 63621 40627
rect 63621 40593 63630 40627
rect 63578 40584 63630 40593
rect 34598 40559 34650 40568
rect 17854 40380 17906 40432
rect 20890 40423 20942 40432
rect 20890 40389 20899 40423
rect 20899 40389 20933 40423
rect 20933 40389 20942 40423
rect 20890 40380 20942 40389
rect 34598 40525 34607 40559
rect 34607 40525 34641 40559
rect 34641 40525 34650 40559
rect 34598 40516 34650 40525
rect 34690 40380 34742 40432
rect 39658 40559 39710 40568
rect 39658 40525 39667 40559
rect 39667 40525 39701 40559
rect 39701 40525 39710 40559
rect 39658 40516 39710 40525
rect 39934 40559 39986 40568
rect 39934 40525 39943 40559
rect 39943 40525 39977 40559
rect 39977 40525 39986 40559
rect 39934 40516 39986 40525
rect 41590 40516 41642 40568
rect 43982 40516 44034 40568
rect 45730 40559 45782 40568
rect 45730 40525 45739 40559
rect 45739 40525 45773 40559
rect 45773 40525 45782 40559
rect 45730 40516 45782 40525
rect 46650 40516 46702 40568
rect 49778 40559 49830 40568
rect 49778 40525 49787 40559
rect 49787 40525 49821 40559
rect 49821 40525 49830 40559
rect 49778 40516 49830 40525
rect 55850 40559 55902 40568
rect 55850 40525 55859 40559
rect 55859 40525 55893 40559
rect 55893 40525 55902 40559
rect 55850 40516 55902 40525
rect 56678 40516 56730 40568
rect 61370 40559 61422 40568
rect 61370 40525 61379 40559
rect 61379 40525 61413 40559
rect 61413 40525 61422 40559
rect 61370 40516 61422 40525
rect 61738 40516 61790 40568
rect 62750 40516 62802 40568
rect 68178 40516 68230 40568
rect 68362 40584 68414 40636
rect 70754 40584 70806 40636
rect 71122 40720 71174 40772
rect 71214 40584 71266 40636
rect 69926 40516 69978 40568
rect 41406 40448 41458 40500
rect 42694 40448 42746 40500
rect 51342 40380 51394 40432
rect 59530 40448 59582 40500
rect 56862 40380 56914 40432
rect 62658 40423 62710 40432
rect 62658 40389 62667 40423
rect 62667 40389 62701 40423
rect 62701 40389 62710 40423
rect 62658 40380 62710 40389
rect 64038 40380 64090 40432
rect 72226 40423 72278 40432
rect 72226 40389 72235 40423
rect 72235 40389 72269 40423
rect 72269 40389 72278 40423
rect 72226 40380 72278 40389
rect 73606 40559 73658 40568
rect 73606 40525 73615 40559
rect 73615 40525 73649 40559
rect 73649 40525 73658 40559
rect 73606 40516 73658 40525
rect 73698 40516 73750 40568
rect 73698 40380 73750 40432
rect 74710 40423 74762 40432
rect 74710 40389 74719 40423
rect 74719 40389 74753 40423
rect 74753 40389 74762 40423
rect 74710 40380 74762 40389
rect 78114 40584 78166 40636
rect 78574 40584 78626 40636
rect 75998 40516 76050 40568
rect 76366 40516 76418 40568
rect 79494 40652 79546 40704
rect 82346 40763 82398 40772
rect 80598 40584 80650 40636
rect 80874 40627 80926 40636
rect 80874 40593 80883 40627
rect 80883 40593 80917 40627
rect 80917 40593 80926 40627
rect 80874 40584 80926 40593
rect 82346 40729 82355 40763
rect 82355 40729 82389 40763
rect 82389 40729 82398 40763
rect 82346 40720 82398 40729
rect 88142 40763 88194 40772
rect 88142 40729 88151 40763
rect 88151 40729 88185 40763
rect 88185 40729 88194 40763
rect 88142 40720 88194 40729
rect 81150 40652 81202 40704
rect 82070 40627 82122 40636
rect 82070 40593 82079 40627
rect 82079 40593 82113 40627
rect 82113 40593 82122 40627
rect 82070 40584 82122 40593
rect 82530 40627 82582 40636
rect 82530 40593 82539 40627
rect 82539 40593 82573 40627
rect 82573 40593 82582 40627
rect 82530 40584 82582 40593
rect 85014 40584 85066 40636
rect 85474 40584 85526 40636
rect 83634 40516 83686 40568
rect 84186 40559 84238 40568
rect 84186 40525 84195 40559
rect 84195 40525 84229 40559
rect 84229 40525 84238 40559
rect 84186 40516 84238 40525
rect 88142 40516 88194 40568
rect 88510 40559 88562 40568
rect 88510 40525 88519 40559
rect 88519 40525 88553 40559
rect 88553 40525 88562 40559
rect 88510 40516 88562 40525
rect 75998 40380 76050 40432
rect 78114 40423 78166 40432
rect 78114 40389 78123 40423
rect 78123 40389 78157 40423
rect 78157 40389 78166 40423
rect 78114 40380 78166 40389
rect 79218 40380 79270 40432
rect 80874 40380 80926 40432
rect 88142 40380 88194 40432
rect 90166 40380 90218 40432
rect 90994 40559 91046 40568
rect 90994 40525 91003 40559
rect 91003 40525 91037 40559
rect 91037 40525 91046 40559
rect 90994 40516 91046 40525
rect 90534 40423 90586 40432
rect 90534 40389 90543 40423
rect 90543 40389 90577 40423
rect 90577 40389 90586 40423
rect 90534 40380 90586 40389
rect 90994 40380 91046 40432
rect 92834 40380 92886 40432
rect 3680 40278 3732 40330
rect 3744 40278 3796 40330
rect 3808 40278 3860 40330
rect 3872 40278 3924 40330
rect 9008 40278 9060 40330
rect 9072 40278 9124 40330
rect 9136 40278 9188 40330
rect 9200 40278 9252 40330
rect 14336 40278 14388 40330
rect 14400 40278 14452 40330
rect 14464 40278 14516 40330
rect 14528 40278 14580 40330
rect 19664 40278 19716 40330
rect 19728 40278 19780 40330
rect 19792 40278 19844 40330
rect 19856 40278 19908 40330
rect 24992 40278 25044 40330
rect 25056 40278 25108 40330
rect 25120 40278 25172 40330
rect 25184 40278 25236 40330
rect 30320 40278 30372 40330
rect 30384 40278 30436 40330
rect 30448 40278 30500 40330
rect 30512 40278 30564 40330
rect 35648 40278 35700 40330
rect 35712 40278 35764 40330
rect 35776 40278 35828 40330
rect 35840 40278 35892 40330
rect 40976 40278 41028 40330
rect 41040 40278 41092 40330
rect 41104 40278 41156 40330
rect 41168 40278 41220 40330
rect 46304 40278 46356 40330
rect 46368 40278 46420 40330
rect 46432 40278 46484 40330
rect 46496 40278 46548 40330
rect 51632 40278 51684 40330
rect 51696 40278 51748 40330
rect 51760 40278 51812 40330
rect 51824 40278 51876 40330
rect 56960 40278 57012 40330
rect 57024 40278 57076 40330
rect 57088 40278 57140 40330
rect 57152 40278 57204 40330
rect 62288 40278 62340 40330
rect 62352 40278 62404 40330
rect 62416 40278 62468 40330
rect 62480 40278 62532 40330
rect 67616 40278 67668 40330
rect 67680 40278 67732 40330
rect 67744 40278 67796 40330
rect 67808 40278 67860 40330
rect 72944 40278 72996 40330
rect 73008 40278 73060 40330
rect 73072 40278 73124 40330
rect 73136 40278 73188 40330
rect 78272 40278 78324 40330
rect 78336 40278 78388 40330
rect 78400 40278 78452 40330
rect 78464 40278 78516 40330
rect 83600 40278 83652 40330
rect 83664 40278 83716 40330
rect 83728 40278 83780 40330
rect 83792 40278 83844 40330
rect 88928 40278 88980 40330
rect 88992 40278 89044 40330
rect 89056 40278 89108 40330
rect 89120 40278 89172 40330
rect 2490 40176 2542 40228
rect 11966 40176 12018 40228
rect 12334 40176 12386 40228
rect 14174 40219 14226 40228
rect 14174 40185 14183 40219
rect 14183 40185 14217 40219
rect 14217 40185 14226 40219
rect 14174 40176 14226 40185
rect 19510 40176 19562 40228
rect 39658 40176 39710 40228
rect 41590 40219 41642 40228
rect 41590 40185 41599 40219
rect 41599 40185 41633 40219
rect 41633 40185 41642 40219
rect 41590 40176 41642 40185
rect 46742 40176 46794 40228
rect 8102 40151 8154 40160
rect 8102 40117 8111 40151
rect 8111 40117 8145 40151
rect 8145 40117 8154 40151
rect 8102 40108 8154 40117
rect 11046 40108 11098 40160
rect 13070 40108 13122 40160
rect 13530 40108 13582 40160
rect 16658 40108 16710 40160
rect 6170 40040 6222 40092
rect 7826 40040 7878 40092
rect 8010 40040 8062 40092
rect 17394 40040 17446 40092
rect 20890 40040 20942 40092
rect 8102 39972 8154 40024
rect 11046 39972 11098 40024
rect 13254 39972 13306 40024
rect 13898 40015 13950 40024
rect 13898 39981 13907 40015
rect 13907 39981 13941 40015
rect 13941 39981 13950 40015
rect 13898 39972 13950 39981
rect 19050 40015 19102 40024
rect 8010 39947 8062 39956
rect 8010 39913 8019 39947
rect 8019 39913 8053 39947
rect 8053 39913 8062 39947
rect 8010 39904 8062 39913
rect 12242 39904 12294 39956
rect 12978 39904 13030 39956
rect 19050 39981 19059 40015
rect 19059 39981 19093 40015
rect 19093 39981 19102 40015
rect 19050 39972 19102 39981
rect 32758 40108 32810 40160
rect 27054 40040 27106 40092
rect 28802 40040 28854 40092
rect 34598 40040 34650 40092
rect 27146 39972 27198 40024
rect 27422 40015 27474 40024
rect 27422 39981 27431 40015
rect 27431 39981 27465 40015
rect 27465 39981 27474 40015
rect 27422 39972 27474 39981
rect 31378 39972 31430 40024
rect 32114 40015 32166 40024
rect 31562 39904 31614 39956
rect 32114 39981 32123 40015
rect 32123 39981 32157 40015
rect 32157 39981 32166 40015
rect 32114 39972 32166 39981
rect 38094 40040 38146 40092
rect 45730 40040 45782 40092
rect 39198 39972 39250 40024
rect 41958 40015 42010 40024
rect 41958 39981 41967 40015
rect 41967 39981 42001 40015
rect 42001 39981 42010 40015
rect 41958 39972 42010 39981
rect 46742 40015 46794 40024
rect 46742 39981 46751 40015
rect 46751 39981 46785 40015
rect 46785 39981 46794 40015
rect 46742 39972 46794 39981
rect 55850 40176 55902 40228
rect 61370 40176 61422 40228
rect 63486 40176 63538 40228
rect 67442 40176 67494 40228
rect 50054 40108 50106 40160
rect 51434 40040 51486 40092
rect 49502 40015 49554 40024
rect 34230 39904 34282 39956
rect 35426 39904 35478 39956
rect 20246 39836 20298 39888
rect 25582 39836 25634 39888
rect 27146 39836 27198 39888
rect 28434 39836 28486 39888
rect 33310 39836 33362 39888
rect 40302 39904 40354 39956
rect 49502 39981 49511 40015
rect 49511 39981 49545 40015
rect 49545 39981 49554 40015
rect 49502 39972 49554 39981
rect 51158 39972 51210 40024
rect 54654 40015 54706 40024
rect 54654 39981 54663 40015
rect 54663 39981 54697 40015
rect 54697 39981 54706 40015
rect 54654 39972 54706 39981
rect 57322 40108 57374 40160
rect 64038 40108 64090 40160
rect 62106 40040 62158 40092
rect 49870 39904 49922 39956
rect 37082 39879 37134 39888
rect 37082 39845 37091 39879
rect 37091 39845 37125 39879
rect 37125 39845 37134 39879
rect 37082 39836 37134 39845
rect 38094 39836 38146 39888
rect 43062 39879 43114 39888
rect 43062 39845 43071 39879
rect 43071 39845 43105 39879
rect 43105 39845 43114 39879
rect 43062 39836 43114 39845
rect 55206 40015 55258 40024
rect 55206 39981 55215 40015
rect 55215 39981 55249 40015
rect 55249 39981 55258 40015
rect 55390 40015 55442 40024
rect 55206 39972 55258 39981
rect 55390 39981 55399 40015
rect 55399 39981 55433 40015
rect 55433 39981 55442 40015
rect 55390 39972 55442 39981
rect 56862 39972 56914 40024
rect 60266 39972 60318 40024
rect 59990 39904 60042 39956
rect 62658 39972 62710 40024
rect 65970 40040 66022 40092
rect 72226 40176 72278 40228
rect 75906 40176 75958 40228
rect 74710 40108 74762 40160
rect 83726 40108 83778 40160
rect 90534 40108 90586 40160
rect 68546 40083 68598 40092
rect 68546 40049 68555 40083
rect 68555 40049 68589 40083
rect 68589 40049 68598 40083
rect 68546 40040 68598 40049
rect 68454 40015 68506 40024
rect 63118 39904 63170 39956
rect 67994 39904 68046 39956
rect 68454 39981 68463 40015
rect 68463 39981 68497 40015
rect 68497 39981 68506 40015
rect 68454 39972 68506 39981
rect 71214 39972 71266 40024
rect 71582 40015 71634 40024
rect 71582 39981 71591 40015
rect 71591 39981 71625 40015
rect 71625 39981 71634 40015
rect 71582 39972 71634 39981
rect 72042 40040 72094 40092
rect 73330 40040 73382 40092
rect 75446 40040 75498 40092
rect 72870 39972 72922 40024
rect 74066 40015 74118 40024
rect 74066 39981 74075 40015
rect 74075 39981 74109 40015
rect 74109 39981 74118 40015
rect 74066 39972 74118 39981
rect 75262 39972 75314 40024
rect 55022 39836 55074 39888
rect 55390 39836 55442 39888
rect 55850 39836 55902 39888
rect 67166 39836 67218 39888
rect 72778 39904 72830 39956
rect 74526 39904 74578 39956
rect 71122 39879 71174 39888
rect 71122 39845 71131 39879
rect 71131 39845 71165 39879
rect 71165 39845 71174 39879
rect 71122 39836 71174 39845
rect 73606 39836 73658 39888
rect 74158 39836 74210 39888
rect 75262 39836 75314 39888
rect 75446 39836 75498 39888
rect 76274 39904 76326 39956
rect 77102 39972 77154 40024
rect 77654 39904 77706 39956
rect 79862 39972 79914 40024
rect 81150 40015 81202 40024
rect 81150 39981 81159 40015
rect 81159 39981 81193 40015
rect 81193 39981 81202 40015
rect 81150 39972 81202 39981
rect 82346 40040 82398 40092
rect 88418 40040 88470 40092
rect 89338 40083 89390 40092
rect 89338 40049 89347 40083
rect 89347 40049 89381 40083
rect 89381 40049 89390 40083
rect 89338 40040 89390 40049
rect 83910 39972 83962 40024
rect 85842 40015 85894 40024
rect 85842 39981 85851 40015
rect 85851 39981 85885 40015
rect 85885 39981 85894 40015
rect 85842 39972 85894 39981
rect 88786 39972 88838 40024
rect 88694 39904 88746 39956
rect 82806 39836 82858 39888
rect 85658 39879 85710 39888
rect 85658 39845 85667 39879
rect 85667 39845 85701 39879
rect 85701 39845 85710 39879
rect 85658 39836 85710 39845
rect 6344 39734 6396 39786
rect 6408 39734 6460 39786
rect 6472 39734 6524 39786
rect 6536 39734 6588 39786
rect 11672 39734 11724 39786
rect 11736 39734 11788 39786
rect 11800 39734 11852 39786
rect 11864 39734 11916 39786
rect 17000 39734 17052 39786
rect 17064 39734 17116 39786
rect 17128 39734 17180 39786
rect 17192 39734 17244 39786
rect 22328 39734 22380 39786
rect 22392 39734 22444 39786
rect 22456 39734 22508 39786
rect 22520 39734 22572 39786
rect 27656 39734 27708 39786
rect 27720 39734 27772 39786
rect 27784 39734 27836 39786
rect 27848 39734 27900 39786
rect 32984 39734 33036 39786
rect 33048 39734 33100 39786
rect 33112 39734 33164 39786
rect 33176 39734 33228 39786
rect 38312 39734 38364 39786
rect 38376 39734 38428 39786
rect 38440 39734 38492 39786
rect 38504 39734 38556 39786
rect 43640 39734 43692 39786
rect 43704 39734 43756 39786
rect 43768 39734 43820 39786
rect 43832 39734 43884 39786
rect 48968 39734 49020 39786
rect 49032 39734 49084 39786
rect 49096 39734 49148 39786
rect 49160 39734 49212 39786
rect 54296 39734 54348 39786
rect 54360 39734 54412 39786
rect 54424 39734 54476 39786
rect 54488 39734 54540 39786
rect 59624 39734 59676 39786
rect 59688 39734 59740 39786
rect 59752 39734 59804 39786
rect 59816 39734 59868 39786
rect 64952 39734 65004 39786
rect 65016 39734 65068 39786
rect 65080 39734 65132 39786
rect 65144 39734 65196 39786
rect 70280 39734 70332 39786
rect 70344 39734 70396 39786
rect 70408 39734 70460 39786
rect 70472 39734 70524 39786
rect 75608 39734 75660 39786
rect 75672 39734 75724 39786
rect 75736 39734 75788 39786
rect 75800 39734 75852 39786
rect 80936 39734 80988 39786
rect 81000 39734 81052 39786
rect 81064 39734 81116 39786
rect 81128 39734 81180 39786
rect 86264 39734 86316 39786
rect 86328 39734 86380 39786
rect 86392 39734 86444 39786
rect 86456 39734 86508 39786
rect 91592 39734 91644 39786
rect 91656 39734 91708 39786
rect 91720 39734 91772 39786
rect 91784 39734 91836 39786
rect 4606 39632 4658 39684
rect 10954 39632 11006 39684
rect 15922 39632 15974 39684
rect 38094 39632 38146 39684
rect 39474 39632 39526 39684
rect 41958 39632 42010 39684
rect 42878 39632 42930 39684
rect 47662 39632 47714 39684
rect 49502 39675 49554 39684
rect 49502 39641 49511 39675
rect 49511 39641 49545 39675
rect 49545 39641 49554 39675
rect 49502 39632 49554 39641
rect 49778 39675 49830 39684
rect 49778 39641 49787 39675
rect 49787 39641 49821 39675
rect 49821 39641 49830 39675
rect 49778 39632 49830 39641
rect 49870 39632 49922 39684
rect 5342 39496 5394 39548
rect 13622 39564 13674 39616
rect 13898 39564 13950 39616
rect 3502 39471 3554 39480
rect 3502 39437 3511 39471
rect 3511 39437 3545 39471
rect 3545 39437 3554 39471
rect 3502 39428 3554 39437
rect 11506 39428 11558 39480
rect 12242 39496 12294 39548
rect 18774 39564 18826 39616
rect 21258 39564 21310 39616
rect 32298 39607 32350 39616
rect 17486 39539 17538 39548
rect 17486 39505 17495 39539
rect 17495 39505 17529 39539
rect 17529 39505 17538 39539
rect 17486 39496 17538 39505
rect 12334 39428 12386 39480
rect 17394 39360 17446 39412
rect 12242 39292 12294 39344
rect 17762 39335 17814 39344
rect 17762 39301 17771 39335
rect 17771 39301 17805 39335
rect 17805 39301 17814 39335
rect 17762 39292 17814 39301
rect 21074 39471 21126 39480
rect 21074 39437 21083 39471
rect 21083 39437 21117 39471
rect 21117 39437 21126 39471
rect 21074 39428 21126 39437
rect 27974 39496 28026 39548
rect 31562 39539 31614 39548
rect 31562 39505 31571 39539
rect 31571 39505 31605 39539
rect 31605 39505 31614 39539
rect 31562 39496 31614 39505
rect 32022 39539 32074 39548
rect 32022 39505 32031 39539
rect 32031 39505 32065 39539
rect 32065 39505 32074 39539
rect 32022 39496 32074 39505
rect 32298 39573 32307 39607
rect 32307 39573 32341 39607
rect 32341 39573 32350 39607
rect 32298 39564 32350 39573
rect 32758 39564 32810 39616
rect 55298 39632 55350 39684
rect 56678 39632 56730 39684
rect 57322 39632 57374 39684
rect 58610 39632 58662 39684
rect 62106 39632 62158 39684
rect 70754 39564 70806 39616
rect 34046 39539 34098 39548
rect 34046 39505 34055 39539
rect 34055 39505 34089 39539
rect 34089 39505 34098 39539
rect 34046 39496 34098 39505
rect 34874 39496 34926 39548
rect 36346 39496 36398 39548
rect 40394 39496 40446 39548
rect 41314 39496 41366 39548
rect 24202 39360 24254 39412
rect 27054 39403 27106 39412
rect 27054 39369 27063 39403
rect 27063 39369 27097 39403
rect 27097 39369 27106 39403
rect 31930 39428 31982 39480
rect 33310 39471 33362 39480
rect 33310 39437 33319 39471
rect 33319 39437 33353 39471
rect 33353 39437 33362 39471
rect 33310 39428 33362 39437
rect 28250 39403 28302 39412
rect 27054 39360 27106 39369
rect 18314 39292 18366 39344
rect 28250 39369 28259 39403
rect 28259 39369 28293 39403
rect 28293 39369 28302 39403
rect 28250 39360 28302 39369
rect 37818 39360 37870 39412
rect 43062 39496 43114 39548
rect 49502 39496 49554 39548
rect 53918 39496 53970 39548
rect 55390 39539 55442 39548
rect 55390 39505 55399 39539
rect 55399 39505 55433 39539
rect 55433 39505 55442 39539
rect 55390 39496 55442 39505
rect 56862 39496 56914 39548
rect 64682 39496 64734 39548
rect 67810 39496 67862 39548
rect 67994 39539 68046 39548
rect 67994 39505 68003 39539
rect 68003 39505 68037 39539
rect 68037 39505 68046 39539
rect 67994 39496 68046 39505
rect 68270 39539 68322 39548
rect 68270 39505 68279 39539
rect 68279 39505 68313 39539
rect 68313 39505 68322 39539
rect 68270 39496 68322 39505
rect 70846 39539 70898 39548
rect 70846 39505 70855 39539
rect 70855 39505 70889 39539
rect 70889 39505 70898 39539
rect 70846 39496 70898 39505
rect 72870 39539 72922 39548
rect 72870 39505 72879 39539
rect 72879 39505 72913 39539
rect 72913 39505 72922 39539
rect 72870 39496 72922 39505
rect 54654 39428 54706 39480
rect 55206 39428 55258 39480
rect 30642 39292 30694 39344
rect 31838 39292 31890 39344
rect 34506 39335 34558 39344
rect 34506 39301 34515 39335
rect 34515 39301 34549 39335
rect 34549 39301 34558 39335
rect 34506 39292 34558 39301
rect 34874 39335 34926 39344
rect 34874 39301 34883 39335
rect 34883 39301 34917 39335
rect 34917 39301 34926 39335
rect 34874 39292 34926 39301
rect 56586 39360 56638 39412
rect 56770 39360 56822 39412
rect 43062 39292 43114 39344
rect 45178 39292 45230 39344
rect 54194 39335 54246 39344
rect 54194 39301 54203 39335
rect 54203 39301 54237 39335
rect 54237 39301 54246 39335
rect 54194 39292 54246 39301
rect 65234 39471 65286 39480
rect 65234 39437 65243 39471
rect 65243 39437 65277 39471
rect 65277 39437 65286 39471
rect 65234 39428 65286 39437
rect 65510 39471 65562 39480
rect 65510 39437 65519 39471
rect 65519 39437 65553 39471
rect 65553 39437 65562 39471
rect 65510 39428 65562 39437
rect 68178 39471 68230 39480
rect 68178 39437 68187 39471
rect 68187 39437 68221 39471
rect 68221 39437 68230 39471
rect 68178 39428 68230 39437
rect 71214 39428 71266 39480
rect 73882 39564 73934 39616
rect 73422 39496 73474 39548
rect 77194 39496 77246 39548
rect 77470 39564 77522 39616
rect 79402 39632 79454 39684
rect 84186 39675 84238 39684
rect 83726 39564 83778 39616
rect 84186 39641 84195 39675
rect 84195 39641 84229 39675
rect 84229 39641 84238 39675
rect 84186 39632 84238 39641
rect 88510 39632 88562 39684
rect 88234 39564 88286 39616
rect 88326 39564 88378 39616
rect 90166 39564 90218 39616
rect 77654 39539 77706 39548
rect 77654 39505 77663 39539
rect 77663 39505 77697 39539
rect 77697 39505 77706 39539
rect 77654 39496 77706 39505
rect 82070 39496 82122 39548
rect 83910 39539 83962 39548
rect 83910 39505 83919 39539
rect 83919 39505 83953 39539
rect 83953 39505 83962 39539
rect 83910 39496 83962 39505
rect 84462 39539 84514 39548
rect 84462 39505 84471 39539
rect 84471 39505 84505 39539
rect 84505 39505 84514 39539
rect 84462 39496 84514 39505
rect 88694 39539 88746 39548
rect 88694 39505 88703 39539
rect 88703 39505 88737 39539
rect 88737 39505 88746 39539
rect 88694 39496 88746 39505
rect 77562 39428 77614 39480
rect 88142 39428 88194 39480
rect 88602 39428 88654 39480
rect 62750 39292 62802 39344
rect 66798 39335 66850 39344
rect 66798 39301 66807 39335
rect 66807 39301 66841 39335
rect 66841 39301 66850 39335
rect 66798 39292 66850 39301
rect 67994 39292 68046 39344
rect 69926 39292 69978 39344
rect 71306 39335 71358 39344
rect 71306 39301 71315 39335
rect 71315 39301 71349 39335
rect 71349 39301 71358 39335
rect 79218 39360 79270 39412
rect 71306 39292 71358 39301
rect 79862 39292 79914 39344
rect 3680 39190 3732 39242
rect 3744 39190 3796 39242
rect 3808 39190 3860 39242
rect 3872 39190 3924 39242
rect 9008 39190 9060 39242
rect 9072 39190 9124 39242
rect 9136 39190 9188 39242
rect 9200 39190 9252 39242
rect 14336 39190 14388 39242
rect 14400 39190 14452 39242
rect 14464 39190 14516 39242
rect 14528 39190 14580 39242
rect 19664 39190 19716 39242
rect 19728 39190 19780 39242
rect 19792 39190 19844 39242
rect 19856 39190 19908 39242
rect 24992 39190 25044 39242
rect 25056 39190 25108 39242
rect 25120 39190 25172 39242
rect 25184 39190 25236 39242
rect 30320 39190 30372 39242
rect 30384 39190 30436 39242
rect 30448 39190 30500 39242
rect 30512 39190 30564 39242
rect 35648 39190 35700 39242
rect 35712 39190 35764 39242
rect 35776 39190 35828 39242
rect 35840 39190 35892 39242
rect 40976 39190 41028 39242
rect 41040 39190 41092 39242
rect 41104 39190 41156 39242
rect 41168 39190 41220 39242
rect 46304 39190 46356 39242
rect 46368 39190 46420 39242
rect 46432 39190 46484 39242
rect 46496 39190 46548 39242
rect 51632 39190 51684 39242
rect 51696 39190 51748 39242
rect 51760 39190 51812 39242
rect 51824 39190 51876 39242
rect 56960 39190 57012 39242
rect 57024 39190 57076 39242
rect 57088 39190 57140 39242
rect 57152 39190 57204 39242
rect 62288 39190 62340 39242
rect 62352 39190 62404 39242
rect 62416 39190 62468 39242
rect 62480 39190 62532 39242
rect 67616 39190 67668 39242
rect 67680 39190 67732 39242
rect 67744 39190 67796 39242
rect 67808 39190 67860 39242
rect 72944 39190 72996 39242
rect 73008 39190 73060 39242
rect 73072 39190 73124 39242
rect 73136 39190 73188 39242
rect 78272 39190 78324 39242
rect 78336 39190 78388 39242
rect 78400 39190 78452 39242
rect 78464 39190 78516 39242
rect 83600 39190 83652 39242
rect 83664 39190 83716 39242
rect 83728 39190 83780 39242
rect 83792 39190 83844 39242
rect 88928 39190 88980 39242
rect 88992 39190 89044 39242
rect 89056 39190 89108 39242
rect 89120 39190 89172 39242
rect 19050 39088 19102 39140
rect 18774 39020 18826 39072
rect 21074 39088 21126 39140
rect 27422 39088 27474 39140
rect 32022 39088 32074 39140
rect 34690 39131 34742 39140
rect 34690 39097 34699 39131
rect 34699 39097 34733 39131
rect 34733 39097 34742 39131
rect 34690 39088 34742 39097
rect 41774 39088 41826 39140
rect 44810 39088 44862 39140
rect 2490 38995 2542 39004
rect 2490 38961 2499 38995
rect 2499 38961 2533 38995
rect 2533 38961 2542 38995
rect 2490 38952 2542 38961
rect 3502 38952 3554 39004
rect 8010 38952 8062 39004
rect 8654 38952 8706 39004
rect 12242 38995 12294 39004
rect 12242 38961 12251 38995
rect 12251 38961 12285 38995
rect 12285 38961 12294 38995
rect 12242 38952 12294 38961
rect 17486 38952 17538 39004
rect 2214 38927 2266 38936
rect 2214 38893 2223 38927
rect 2223 38893 2257 38927
rect 2257 38893 2266 38927
rect 2214 38884 2266 38893
rect 3410 38884 3462 38936
rect 9114 38927 9166 38936
rect 4330 38816 4382 38868
rect 8102 38859 8154 38868
rect 8102 38825 8111 38859
rect 8111 38825 8145 38859
rect 8145 38825 8154 38859
rect 8102 38816 8154 38825
rect 9114 38893 9123 38927
rect 9123 38893 9157 38927
rect 9157 38893 9166 38927
rect 9114 38884 9166 38893
rect 13622 38927 13674 38936
rect 9758 38816 9810 38868
rect 3410 38748 3462 38800
rect 4054 38791 4106 38800
rect 4054 38757 4063 38791
rect 4063 38757 4097 38791
rect 4097 38757 4106 38791
rect 4054 38748 4106 38757
rect 9114 38748 9166 38800
rect 9482 38748 9534 38800
rect 13622 38893 13631 38927
rect 13631 38893 13665 38927
rect 13665 38893 13674 38927
rect 13622 38884 13674 38893
rect 19050 38884 19102 38936
rect 20246 38927 20298 38936
rect 20246 38893 20255 38927
rect 20255 38893 20289 38927
rect 20289 38893 20298 38927
rect 20246 38884 20298 38893
rect 25674 38884 25726 38936
rect 27422 38884 27474 38936
rect 27514 38884 27566 38936
rect 27974 38884 28026 38936
rect 16014 38859 16066 38868
rect 16014 38825 16023 38859
rect 16023 38825 16057 38859
rect 16057 38825 16066 38859
rect 16014 38816 16066 38825
rect 16750 38816 16802 38868
rect 32758 38884 32810 38936
rect 32666 38816 32718 38868
rect 34874 39020 34926 39072
rect 39474 39020 39526 39072
rect 47202 39063 47254 39072
rect 47202 39029 47211 39063
rect 47211 39029 47245 39063
rect 47245 39029 47254 39063
rect 50330 39088 50382 39140
rect 50514 39088 50566 39140
rect 52170 39088 52222 39140
rect 54194 39088 54246 39140
rect 55114 39088 55166 39140
rect 55850 39088 55902 39140
rect 65510 39088 65562 39140
rect 68270 39131 68322 39140
rect 68270 39097 68279 39131
rect 68279 39097 68313 39131
rect 68313 39097 68322 39131
rect 68270 39088 68322 39097
rect 74066 39131 74118 39140
rect 74066 39097 74075 39131
rect 74075 39097 74109 39131
rect 74109 39097 74118 39131
rect 74066 39088 74118 39097
rect 75446 39088 75498 39140
rect 90166 39131 90218 39140
rect 47202 39020 47254 39029
rect 34506 38952 34558 39004
rect 40854 38995 40906 39004
rect 40854 38961 40863 38995
rect 40863 38961 40897 38995
rect 40897 38961 40906 38995
rect 41314 38995 41366 39004
rect 40854 38952 40906 38961
rect 41314 38961 41323 38995
rect 41323 38961 41357 38995
rect 41357 38961 41366 38995
rect 41314 38952 41366 38961
rect 43062 38995 43114 39004
rect 43062 38961 43071 38995
rect 43071 38961 43105 38995
rect 43105 38961 43114 38995
rect 43062 38952 43114 38961
rect 34690 38884 34742 38936
rect 41774 38927 41826 38936
rect 41314 38816 41366 38868
rect 14082 38748 14134 38800
rect 33402 38791 33454 38800
rect 33402 38757 33411 38791
rect 33411 38757 33445 38791
rect 33445 38757 33454 38791
rect 33402 38748 33454 38757
rect 41774 38893 41783 38927
rect 41783 38893 41817 38927
rect 41817 38893 41826 38927
rect 41774 38884 41826 38893
rect 43154 38927 43206 38936
rect 43154 38893 43163 38927
rect 43163 38893 43197 38927
rect 43197 38893 43206 38927
rect 43154 38884 43206 38893
rect 47478 38952 47530 39004
rect 51158 38995 51210 39004
rect 51158 38961 51167 38995
rect 51167 38961 51201 38995
rect 51201 38961 51210 38995
rect 51158 38952 51210 38961
rect 53918 38995 53970 39004
rect 46006 38884 46058 38936
rect 47294 38927 47346 38936
rect 47294 38893 47303 38927
rect 47303 38893 47337 38927
rect 47337 38893 47346 38927
rect 47294 38884 47346 38893
rect 48030 38927 48082 38936
rect 48030 38893 48039 38927
rect 48039 38893 48073 38927
rect 48073 38893 48082 38927
rect 48030 38884 48082 38893
rect 44718 38816 44770 38868
rect 44810 38816 44862 38868
rect 50422 38884 50474 38936
rect 42326 38791 42378 38800
rect 42326 38757 42335 38791
rect 42335 38757 42369 38791
rect 42369 38757 42378 38791
rect 42326 38748 42378 38757
rect 47386 38791 47438 38800
rect 47386 38757 47395 38791
rect 47395 38757 47429 38791
rect 47429 38757 47438 38791
rect 47386 38748 47438 38757
rect 47570 38748 47622 38800
rect 51710 38884 51762 38936
rect 53918 38961 53927 38995
rect 53927 38961 53961 38995
rect 53961 38961 53970 38995
rect 53918 38952 53970 38961
rect 52170 38927 52222 38936
rect 52170 38893 52179 38927
rect 52179 38893 52213 38927
rect 52213 38893 52222 38927
rect 52170 38884 52222 38893
rect 52262 38927 52314 38936
rect 52262 38893 52271 38927
rect 52271 38893 52305 38927
rect 52305 38893 52314 38927
rect 55114 38952 55166 39004
rect 52262 38884 52314 38893
rect 55390 39020 55442 39072
rect 55482 39020 55534 39072
rect 70846 39020 70898 39072
rect 59990 38952 60042 39004
rect 63026 38952 63078 39004
rect 60358 38927 60410 38936
rect 60358 38893 60367 38927
rect 60367 38893 60401 38927
rect 60401 38893 60410 38927
rect 60358 38884 60410 38893
rect 61370 38884 61422 38936
rect 62934 38884 62986 38936
rect 64130 38927 64182 38936
rect 64130 38893 64139 38927
rect 64139 38893 64173 38927
rect 64173 38893 64182 38927
rect 64130 38884 64182 38893
rect 64774 38927 64826 38936
rect 50790 38816 50842 38868
rect 63670 38816 63722 38868
rect 64774 38893 64783 38927
rect 64783 38893 64817 38927
rect 64817 38893 64826 38927
rect 64774 38884 64826 38893
rect 73974 38952 74026 39004
rect 74158 38952 74210 39004
rect 90166 39097 90175 39131
rect 90175 39097 90209 39131
rect 90209 39097 90218 39131
rect 90166 39088 90218 39097
rect 66798 38927 66850 38936
rect 66798 38893 66807 38927
rect 66807 38893 66841 38927
rect 66841 38893 66850 38927
rect 66798 38884 66850 38893
rect 60266 38748 60318 38800
rect 64774 38748 64826 38800
rect 68638 38927 68690 38936
rect 68638 38893 68647 38927
rect 68647 38893 68681 38927
rect 68681 38893 68690 38927
rect 68638 38884 68690 38893
rect 69006 38927 69058 38936
rect 69006 38893 69015 38927
rect 69015 38893 69049 38927
rect 69049 38893 69058 38927
rect 69006 38884 69058 38893
rect 68362 38748 68414 38800
rect 73698 38884 73750 38936
rect 90166 38952 90218 39004
rect 73790 38816 73842 38868
rect 76274 38884 76326 38936
rect 76458 38884 76510 38936
rect 77102 38927 77154 38936
rect 77102 38893 77111 38927
rect 77111 38893 77145 38927
rect 77145 38893 77154 38927
rect 77102 38884 77154 38893
rect 77470 38748 77522 38800
rect 90718 38927 90770 38936
rect 90718 38893 90727 38927
rect 90727 38893 90761 38927
rect 90761 38893 90770 38927
rect 90718 38884 90770 38893
rect 80414 38748 80466 38800
rect 91454 38748 91506 38800
rect 6344 38646 6396 38698
rect 6408 38646 6460 38698
rect 6472 38646 6524 38698
rect 6536 38646 6588 38698
rect 11672 38646 11724 38698
rect 11736 38646 11788 38698
rect 11800 38646 11852 38698
rect 11864 38646 11916 38698
rect 17000 38646 17052 38698
rect 17064 38646 17116 38698
rect 17128 38646 17180 38698
rect 17192 38646 17244 38698
rect 22328 38646 22380 38698
rect 22392 38646 22444 38698
rect 22456 38646 22508 38698
rect 22520 38646 22572 38698
rect 27656 38646 27708 38698
rect 27720 38646 27772 38698
rect 27784 38646 27836 38698
rect 27848 38646 27900 38698
rect 32984 38646 33036 38698
rect 33048 38646 33100 38698
rect 33112 38646 33164 38698
rect 33176 38646 33228 38698
rect 38312 38646 38364 38698
rect 38376 38646 38428 38698
rect 38440 38646 38492 38698
rect 38504 38646 38556 38698
rect 43640 38646 43692 38698
rect 43704 38646 43756 38698
rect 43768 38646 43820 38698
rect 43832 38646 43884 38698
rect 48968 38646 49020 38698
rect 49032 38646 49084 38698
rect 49096 38646 49148 38698
rect 49160 38646 49212 38698
rect 54296 38646 54348 38698
rect 54360 38646 54412 38698
rect 54424 38646 54476 38698
rect 54488 38646 54540 38698
rect 59624 38646 59676 38698
rect 59688 38646 59740 38698
rect 59752 38646 59804 38698
rect 59816 38646 59868 38698
rect 64952 38646 65004 38698
rect 65016 38646 65068 38698
rect 65080 38646 65132 38698
rect 65144 38646 65196 38698
rect 70280 38646 70332 38698
rect 70344 38646 70396 38698
rect 70408 38646 70460 38698
rect 70472 38646 70524 38698
rect 75608 38646 75660 38698
rect 75672 38646 75724 38698
rect 75736 38646 75788 38698
rect 75800 38646 75852 38698
rect 80936 38646 80988 38698
rect 81000 38646 81052 38698
rect 81064 38646 81116 38698
rect 81128 38646 81180 38698
rect 86264 38646 86316 38698
rect 86328 38646 86380 38698
rect 86392 38646 86444 38698
rect 86456 38646 86508 38698
rect 91592 38646 91644 38698
rect 91656 38646 91708 38698
rect 91720 38646 91772 38698
rect 91784 38646 91836 38698
rect 2490 38587 2542 38596
rect 2490 38553 2499 38587
rect 2499 38553 2533 38587
rect 2533 38553 2542 38587
rect 2490 38544 2542 38553
rect 4330 38451 4382 38460
rect 4330 38417 4339 38451
rect 4339 38417 4373 38451
rect 4373 38417 4382 38451
rect 4330 38408 4382 38417
rect 9298 38408 9350 38460
rect 13070 38544 13122 38596
rect 29354 38587 29406 38596
rect 16750 38519 16802 38528
rect 16750 38485 16759 38519
rect 16759 38485 16793 38519
rect 16793 38485 16802 38519
rect 16750 38476 16802 38485
rect 16014 38408 16066 38460
rect 16382 38451 16434 38460
rect 16382 38417 16391 38451
rect 16391 38417 16425 38451
rect 16425 38417 16434 38451
rect 16382 38408 16434 38417
rect 17762 38451 17814 38460
rect 17762 38417 17771 38451
rect 17771 38417 17805 38451
rect 17805 38417 17814 38451
rect 17762 38408 17814 38417
rect 27054 38476 27106 38528
rect 2398 38340 2450 38392
rect 4054 38383 4106 38392
rect 4054 38349 4063 38383
rect 4063 38349 4097 38383
rect 4097 38349 4106 38383
rect 4054 38340 4106 38349
rect 7642 38340 7694 38392
rect 10310 38383 10362 38392
rect 10310 38349 10319 38383
rect 10319 38349 10353 38383
rect 10353 38349 10362 38383
rect 10310 38340 10362 38349
rect 5894 38247 5946 38256
rect 5894 38213 5903 38247
rect 5903 38213 5937 38247
rect 5937 38213 5946 38247
rect 5894 38204 5946 38213
rect 10770 38204 10822 38256
rect 11966 38204 12018 38256
rect 15738 38204 15790 38256
rect 15922 38204 15974 38256
rect 17578 38247 17630 38256
rect 17578 38213 17587 38247
rect 17587 38213 17621 38247
rect 17621 38213 17630 38247
rect 17578 38204 17630 38213
rect 17670 38204 17722 38256
rect 25674 38408 25726 38460
rect 29354 38553 29363 38587
rect 29363 38553 29397 38587
rect 29397 38553 29406 38587
rect 29354 38544 29406 38553
rect 28250 38408 28302 38460
rect 34690 38544 34742 38596
rect 41774 38544 41826 38596
rect 42326 38544 42378 38596
rect 47570 38544 47622 38596
rect 48030 38544 48082 38596
rect 51342 38544 51394 38596
rect 53918 38544 53970 38596
rect 34874 38476 34926 38528
rect 43522 38476 43574 38528
rect 18590 38204 18642 38256
rect 29722 38340 29774 38392
rect 24662 38315 24714 38324
rect 24662 38281 24671 38315
rect 24671 38281 24705 38315
rect 24705 38281 24714 38315
rect 24662 38272 24714 38281
rect 29630 38204 29682 38256
rect 39474 38451 39526 38460
rect 39474 38417 39483 38451
rect 39483 38417 39517 38451
rect 39517 38417 39526 38451
rect 39474 38408 39526 38417
rect 40026 38451 40078 38460
rect 40026 38417 40035 38451
rect 40035 38417 40069 38451
rect 40069 38417 40078 38451
rect 40026 38408 40078 38417
rect 33586 38383 33638 38392
rect 33586 38349 33595 38383
rect 33595 38349 33629 38383
rect 33629 38349 33638 38383
rect 33586 38340 33638 38349
rect 40302 38383 40354 38392
rect 40302 38349 40311 38383
rect 40311 38349 40345 38383
rect 40345 38349 40354 38383
rect 40302 38340 40354 38349
rect 39934 38272 39986 38324
rect 33954 38204 34006 38256
rect 34874 38247 34926 38256
rect 34874 38213 34883 38247
rect 34883 38213 34917 38247
rect 34917 38213 34926 38247
rect 34874 38204 34926 38213
rect 40854 38204 40906 38256
rect 44718 38451 44770 38460
rect 44718 38417 44727 38451
rect 44727 38417 44761 38451
rect 44761 38417 44770 38451
rect 44718 38408 44770 38417
rect 48122 38408 48174 38460
rect 41314 38204 41366 38256
rect 45454 38204 45506 38256
rect 46006 38247 46058 38256
rect 46006 38213 46015 38247
rect 46015 38213 46049 38247
rect 46049 38213 46058 38247
rect 46006 38204 46058 38213
rect 46098 38204 46150 38256
rect 48122 38247 48174 38256
rect 48122 38213 48131 38247
rect 48131 38213 48165 38247
rect 48165 38213 48174 38247
rect 48122 38204 48174 38213
rect 51986 38451 52038 38460
rect 51986 38417 51995 38451
rect 51995 38417 52029 38451
rect 52029 38417 52038 38451
rect 51986 38408 52038 38417
rect 54194 38476 54246 38528
rect 54654 38519 54706 38528
rect 54654 38485 54663 38519
rect 54663 38485 54697 38519
rect 54697 38485 54706 38519
rect 54654 38476 54706 38485
rect 55206 38408 55258 38460
rect 55390 38476 55442 38528
rect 59070 38408 59122 38460
rect 61646 38544 61698 38596
rect 63670 38587 63722 38596
rect 63670 38553 63679 38587
rect 63679 38553 63713 38587
rect 63713 38553 63722 38587
rect 63670 38544 63722 38553
rect 68638 38544 68690 38596
rect 72410 38544 72462 38596
rect 61370 38476 61422 38528
rect 74250 38544 74302 38596
rect 76458 38544 76510 38596
rect 77102 38544 77154 38596
rect 88418 38544 88470 38596
rect 73422 38519 73474 38528
rect 60634 38383 60686 38392
rect 52446 38315 52498 38324
rect 52446 38281 52455 38315
rect 52455 38281 52489 38315
rect 52489 38281 52498 38315
rect 52446 38272 52498 38281
rect 53918 38204 53970 38256
rect 60634 38349 60643 38383
rect 60643 38349 60677 38383
rect 60677 38349 60686 38383
rect 60634 38340 60686 38349
rect 57966 38204 58018 38256
rect 61738 38247 61790 38256
rect 61738 38213 61747 38247
rect 61747 38213 61781 38247
rect 61781 38213 61790 38247
rect 61738 38204 61790 38213
rect 63210 38204 63262 38256
rect 64130 38408 64182 38460
rect 73422 38485 73431 38519
rect 73431 38485 73465 38519
rect 73465 38485 73474 38519
rect 73422 38476 73474 38485
rect 73790 38476 73842 38528
rect 67810 38451 67862 38460
rect 67810 38417 67819 38451
rect 67819 38417 67853 38451
rect 67853 38417 67862 38451
rect 68362 38451 68414 38460
rect 67810 38408 67862 38417
rect 68362 38417 68371 38451
rect 68371 38417 68405 38451
rect 68405 38417 68414 38451
rect 68362 38408 68414 38417
rect 69098 38451 69150 38460
rect 69098 38417 69107 38451
rect 69107 38417 69141 38451
rect 69141 38417 69150 38451
rect 69098 38408 69150 38417
rect 72594 38408 72646 38460
rect 73698 38408 73750 38460
rect 74986 38408 75038 38460
rect 75446 38408 75498 38460
rect 80414 38408 80466 38460
rect 82806 38408 82858 38460
rect 83266 38451 83318 38460
rect 83266 38417 83275 38451
rect 83275 38417 83309 38451
rect 83309 38417 83318 38451
rect 83266 38408 83318 38417
rect 74710 38340 74762 38392
rect 86394 38408 86446 38460
rect 90718 38544 90770 38596
rect 89890 38451 89942 38460
rect 85106 38340 85158 38392
rect 88694 38340 88746 38392
rect 89890 38417 89899 38451
rect 89899 38417 89933 38451
rect 89933 38417 89942 38451
rect 89890 38408 89942 38417
rect 91454 38451 91506 38460
rect 91454 38417 91463 38451
rect 91463 38417 91497 38451
rect 91497 38417 91506 38451
rect 91454 38408 91506 38417
rect 68270 38204 68322 38256
rect 68546 38204 68598 38256
rect 69650 38204 69702 38256
rect 72226 38247 72278 38256
rect 72226 38213 72235 38247
rect 72235 38213 72269 38247
rect 72269 38213 72278 38247
rect 72226 38204 72278 38213
rect 77470 38204 77522 38256
rect 79218 38204 79270 38256
rect 85290 38204 85342 38256
rect 3680 38102 3732 38154
rect 3744 38102 3796 38154
rect 3808 38102 3860 38154
rect 3872 38102 3924 38154
rect 9008 38102 9060 38154
rect 9072 38102 9124 38154
rect 9136 38102 9188 38154
rect 9200 38102 9252 38154
rect 14336 38102 14388 38154
rect 14400 38102 14452 38154
rect 14464 38102 14516 38154
rect 14528 38102 14580 38154
rect 19664 38102 19716 38154
rect 19728 38102 19780 38154
rect 19792 38102 19844 38154
rect 19856 38102 19908 38154
rect 24992 38102 25044 38154
rect 25056 38102 25108 38154
rect 25120 38102 25172 38154
rect 25184 38102 25236 38154
rect 30320 38102 30372 38154
rect 30384 38102 30436 38154
rect 30448 38102 30500 38154
rect 30512 38102 30564 38154
rect 35648 38102 35700 38154
rect 35712 38102 35764 38154
rect 35776 38102 35828 38154
rect 35840 38102 35892 38154
rect 40976 38102 41028 38154
rect 41040 38102 41092 38154
rect 41104 38102 41156 38154
rect 41168 38102 41220 38154
rect 46304 38102 46356 38154
rect 46368 38102 46420 38154
rect 46432 38102 46484 38154
rect 46496 38102 46548 38154
rect 51632 38102 51684 38154
rect 51696 38102 51748 38154
rect 51760 38102 51812 38154
rect 51824 38102 51876 38154
rect 56960 38102 57012 38154
rect 57024 38102 57076 38154
rect 57088 38102 57140 38154
rect 57152 38102 57204 38154
rect 62288 38102 62340 38154
rect 62352 38102 62404 38154
rect 62416 38102 62468 38154
rect 62480 38102 62532 38154
rect 67616 38102 67668 38154
rect 67680 38102 67732 38154
rect 67744 38102 67796 38154
rect 67808 38102 67860 38154
rect 72944 38102 72996 38154
rect 73008 38102 73060 38154
rect 73072 38102 73124 38154
rect 73136 38102 73188 38154
rect 78272 38102 78324 38154
rect 78336 38102 78388 38154
rect 78400 38102 78452 38154
rect 78464 38102 78516 38154
rect 83600 38102 83652 38154
rect 83664 38102 83716 38154
rect 83728 38102 83780 38154
rect 83792 38102 83844 38154
rect 88928 38102 88980 38154
rect 88992 38102 89044 38154
rect 89056 38102 89108 38154
rect 89120 38102 89172 38154
rect 9298 38043 9350 38052
rect 9298 38009 9307 38043
rect 9307 38009 9341 38043
rect 9341 38009 9350 38043
rect 9298 38000 9350 38009
rect 9758 38000 9810 38052
rect 10402 38000 10454 38052
rect 17578 38000 17630 38052
rect 20246 38000 20298 38052
rect 27422 38000 27474 38052
rect 33586 38000 33638 38052
rect 40026 38000 40078 38052
rect 8654 37932 8706 37984
rect 9114 37932 9166 37984
rect 8102 37864 8154 37916
rect 11966 37864 12018 37916
rect 17762 37932 17814 37984
rect 29630 37932 29682 37984
rect 2214 37796 2266 37848
rect 2398 37839 2450 37848
rect 2398 37805 2407 37839
rect 2407 37805 2441 37839
rect 2441 37805 2450 37839
rect 2398 37796 2450 37805
rect 7458 37839 7510 37848
rect 7458 37805 7467 37839
rect 7467 37805 7501 37839
rect 7501 37805 7510 37839
rect 7458 37796 7510 37805
rect 12794 37839 12846 37848
rect 4422 37728 4474 37780
rect 3962 37703 4014 37712
rect 3962 37669 3971 37703
rect 3971 37669 4005 37703
rect 4005 37669 4014 37703
rect 3962 37660 4014 37669
rect 12794 37805 12803 37839
rect 12803 37805 12837 37839
rect 12837 37805 12846 37839
rect 12794 37796 12846 37805
rect 17946 37864 17998 37916
rect 20614 37864 20666 37916
rect 21074 37864 21126 37916
rect 24662 37864 24714 37916
rect 25674 37907 25726 37916
rect 25674 37873 25683 37907
rect 25683 37873 25717 37907
rect 25717 37873 25726 37907
rect 25674 37864 25726 37873
rect 27974 37864 28026 37916
rect 20430 37839 20482 37848
rect 14174 37771 14226 37780
rect 14174 37737 14183 37771
rect 14183 37737 14217 37771
rect 14217 37737 14226 37771
rect 14174 37728 14226 37737
rect 15830 37728 15882 37780
rect 16014 37771 16066 37780
rect 16014 37737 16023 37771
rect 16023 37737 16057 37771
rect 16057 37737 16066 37771
rect 16014 37728 16066 37737
rect 17670 37771 17722 37780
rect 17670 37737 17679 37771
rect 17679 37737 17713 37771
rect 17713 37737 17722 37771
rect 17670 37728 17722 37737
rect 20430 37805 20439 37839
rect 20439 37805 20473 37839
rect 20473 37805 20482 37839
rect 20430 37796 20482 37805
rect 25582 37839 25634 37848
rect 25582 37805 25591 37839
rect 25591 37805 25625 37839
rect 25625 37805 25634 37839
rect 25582 37796 25634 37805
rect 27330 37796 27382 37848
rect 17946 37728 17998 37780
rect 20338 37771 20390 37780
rect 20338 37737 20347 37771
rect 20347 37737 20381 37771
rect 20381 37737 20390 37771
rect 20338 37728 20390 37737
rect 27054 37728 27106 37780
rect 29722 37796 29774 37848
rect 34874 37932 34926 37984
rect 42326 38000 42378 38052
rect 69098 38000 69150 38052
rect 72226 38000 72278 38052
rect 82070 38000 82122 38052
rect 86394 38043 86446 38052
rect 86394 38009 86403 38043
rect 86403 38009 86437 38043
rect 86437 38009 86446 38043
rect 86394 38000 86446 38009
rect 90166 38043 90218 38052
rect 90166 38009 90175 38043
rect 90175 38009 90209 38043
rect 90209 38009 90218 38043
rect 90166 38000 90218 38009
rect 45362 37932 45414 37984
rect 47386 37932 47438 37984
rect 31930 37864 31982 37916
rect 34046 37864 34098 37916
rect 34966 37864 35018 37916
rect 36622 37907 36674 37916
rect 36622 37873 36631 37907
rect 36631 37873 36665 37907
rect 36665 37873 36674 37907
rect 36622 37864 36674 37873
rect 37818 37864 37870 37916
rect 32298 37728 32350 37780
rect 33402 37796 33454 37848
rect 33586 37796 33638 37848
rect 35150 37796 35202 37848
rect 14082 37660 14134 37712
rect 27330 37703 27382 37712
rect 27330 37669 27339 37703
rect 27339 37669 27373 37703
rect 27373 37669 27382 37703
rect 27330 37660 27382 37669
rect 28894 37703 28946 37712
rect 28894 37669 28903 37703
rect 28903 37669 28937 37703
rect 28937 37669 28946 37703
rect 28894 37660 28946 37669
rect 29722 37703 29774 37712
rect 29722 37669 29731 37703
rect 29731 37669 29765 37703
rect 29765 37669 29774 37703
rect 29722 37660 29774 37669
rect 33586 37703 33638 37712
rect 33586 37669 33595 37703
rect 33595 37669 33629 37703
rect 33629 37669 33638 37703
rect 33586 37660 33638 37669
rect 34966 37703 35018 37712
rect 34966 37669 34975 37703
rect 34975 37669 35009 37703
rect 35009 37669 35018 37703
rect 34966 37660 35018 37669
rect 35058 37660 35110 37712
rect 40394 37796 40446 37848
rect 40578 37864 40630 37916
rect 47478 37907 47530 37916
rect 37634 37728 37686 37780
rect 37818 37771 37870 37780
rect 37818 37737 37827 37771
rect 37827 37737 37861 37771
rect 37861 37737 37870 37771
rect 37818 37728 37870 37737
rect 40578 37771 40630 37780
rect 39566 37660 39618 37712
rect 39842 37660 39894 37712
rect 40578 37737 40587 37771
rect 40587 37737 40621 37771
rect 40621 37737 40630 37771
rect 40578 37728 40630 37737
rect 41222 37796 41274 37848
rect 41774 37796 41826 37848
rect 43522 37796 43574 37848
rect 45454 37796 45506 37848
rect 46834 37796 46886 37848
rect 47478 37873 47487 37907
rect 47487 37873 47521 37907
rect 47521 37873 47530 37907
rect 47478 37864 47530 37873
rect 51250 37907 51302 37916
rect 51250 37873 51259 37907
rect 51259 37873 51293 37907
rect 51293 37873 51302 37907
rect 51250 37864 51302 37873
rect 53918 37932 53970 37984
rect 60542 37932 60594 37984
rect 69006 37932 69058 37984
rect 73054 37932 73106 37984
rect 73790 37932 73842 37984
rect 48490 37839 48542 37848
rect 40486 37660 40538 37712
rect 41038 37660 41090 37712
rect 41222 37703 41274 37712
rect 41222 37669 41231 37703
rect 41231 37669 41265 37703
rect 41265 37669 41274 37703
rect 41222 37660 41274 37669
rect 41774 37703 41826 37712
rect 41774 37669 41783 37703
rect 41783 37669 41817 37703
rect 41817 37669 41826 37703
rect 41774 37660 41826 37669
rect 45546 37660 45598 37712
rect 47386 37728 47438 37780
rect 48490 37805 48499 37839
rect 48499 37805 48533 37839
rect 48533 37805 48542 37839
rect 48490 37796 48542 37805
rect 51894 37839 51946 37848
rect 51894 37805 51903 37839
rect 51903 37805 51937 37839
rect 51937 37805 51946 37839
rect 51894 37796 51946 37805
rect 52262 37796 52314 37848
rect 54746 37796 54798 37848
rect 55206 37796 55258 37848
rect 56862 37796 56914 37848
rect 55298 37728 55350 37780
rect 52354 37703 52406 37712
rect 52354 37669 52363 37703
rect 52363 37669 52397 37703
rect 52397 37669 52406 37703
rect 52354 37660 52406 37669
rect 55022 37660 55074 37712
rect 56126 37703 56178 37712
rect 56126 37669 56135 37703
rect 56135 37669 56169 37703
rect 56169 37669 56178 37703
rect 56126 37660 56178 37669
rect 57138 37864 57190 37916
rect 57690 37864 57742 37916
rect 60634 37864 60686 37916
rect 67994 37907 68046 37916
rect 58058 37796 58110 37848
rect 58150 37796 58202 37848
rect 58886 37796 58938 37848
rect 59070 37796 59122 37848
rect 59438 37796 59490 37848
rect 61738 37796 61790 37848
rect 62106 37796 62158 37848
rect 62474 37796 62526 37848
rect 67994 37873 68003 37907
rect 68003 37873 68037 37907
rect 68037 37873 68046 37907
rect 67994 37864 68046 37873
rect 68270 37907 68322 37916
rect 68270 37873 68279 37907
rect 68279 37873 68313 37907
rect 68313 37873 68322 37907
rect 68270 37864 68322 37873
rect 69926 37864 69978 37916
rect 73974 37839 74026 37848
rect 58058 37703 58110 37712
rect 58058 37669 58067 37703
rect 58067 37669 58101 37703
rect 58101 37669 58110 37703
rect 58058 37660 58110 37669
rect 59070 37660 59122 37712
rect 61370 37703 61422 37712
rect 61370 37669 61379 37703
rect 61379 37669 61413 37703
rect 61413 37669 61422 37703
rect 61370 37660 61422 37669
rect 62106 37703 62158 37712
rect 62106 37669 62115 37703
rect 62115 37669 62149 37703
rect 62149 37669 62158 37703
rect 62106 37660 62158 37669
rect 63762 37703 63814 37712
rect 63762 37669 63771 37703
rect 63771 37669 63805 37703
rect 63805 37669 63814 37703
rect 63762 37660 63814 37669
rect 72226 37660 72278 37712
rect 73974 37805 73983 37839
rect 73983 37805 74017 37839
rect 74017 37805 74026 37839
rect 73974 37796 74026 37805
rect 72778 37728 72830 37780
rect 73882 37728 73934 37780
rect 74158 37796 74210 37848
rect 74710 37839 74762 37848
rect 74710 37805 74719 37839
rect 74719 37805 74753 37839
rect 74753 37805 74762 37839
rect 74710 37796 74762 37805
rect 74066 37660 74118 37712
rect 74158 37660 74210 37712
rect 74986 37796 75038 37848
rect 76642 37864 76694 37916
rect 76826 37864 76878 37916
rect 77930 37864 77982 37916
rect 82806 37932 82858 37984
rect 85106 37907 85158 37916
rect 85106 37873 85115 37907
rect 85115 37873 85149 37907
rect 85149 37873 85158 37907
rect 85106 37864 85158 37873
rect 88602 37907 88654 37916
rect 88602 37873 88611 37907
rect 88611 37873 88645 37907
rect 88645 37873 88654 37907
rect 88602 37864 88654 37873
rect 89522 37864 89574 37916
rect 76458 37839 76510 37848
rect 76458 37805 76467 37839
rect 76467 37805 76501 37839
rect 76501 37805 76510 37839
rect 76458 37796 76510 37805
rect 79218 37839 79270 37848
rect 79218 37805 79227 37839
rect 79227 37805 79261 37839
rect 79261 37805 79270 37839
rect 79218 37796 79270 37805
rect 82162 37796 82214 37848
rect 75354 37771 75406 37780
rect 75354 37737 75363 37771
rect 75363 37737 75397 37771
rect 75397 37737 75406 37771
rect 75354 37728 75406 37737
rect 76366 37660 76418 37712
rect 76734 37660 76786 37712
rect 84922 37796 84974 37848
rect 88510 37796 88562 37848
rect 84278 37728 84330 37780
rect 86578 37728 86630 37780
rect 89246 37728 89298 37780
rect 89890 37796 89942 37848
rect 90350 37796 90402 37848
rect 90718 37839 90770 37848
rect 90718 37805 90727 37839
rect 90727 37805 90761 37839
rect 90761 37805 90770 37839
rect 90718 37796 90770 37805
rect 84002 37703 84054 37712
rect 84002 37669 84011 37703
rect 84011 37669 84045 37703
rect 84045 37669 84054 37703
rect 84002 37660 84054 37669
rect 91362 37660 91414 37712
rect 6344 37558 6396 37610
rect 6408 37558 6460 37610
rect 6472 37558 6524 37610
rect 6536 37558 6588 37610
rect 11672 37558 11724 37610
rect 11736 37558 11788 37610
rect 11800 37558 11852 37610
rect 11864 37558 11916 37610
rect 17000 37558 17052 37610
rect 17064 37558 17116 37610
rect 17128 37558 17180 37610
rect 17192 37558 17244 37610
rect 22328 37558 22380 37610
rect 22392 37558 22444 37610
rect 22456 37558 22508 37610
rect 22520 37558 22572 37610
rect 27656 37558 27708 37610
rect 27720 37558 27772 37610
rect 27784 37558 27836 37610
rect 27848 37558 27900 37610
rect 32984 37558 33036 37610
rect 33048 37558 33100 37610
rect 33112 37558 33164 37610
rect 33176 37558 33228 37610
rect 38312 37558 38364 37610
rect 38376 37558 38428 37610
rect 38440 37558 38492 37610
rect 38504 37558 38556 37610
rect 43640 37558 43692 37610
rect 43704 37558 43756 37610
rect 43768 37558 43820 37610
rect 43832 37558 43884 37610
rect 48968 37558 49020 37610
rect 49032 37558 49084 37610
rect 49096 37558 49148 37610
rect 49160 37558 49212 37610
rect 54296 37558 54348 37610
rect 54360 37558 54412 37610
rect 54424 37558 54476 37610
rect 54488 37558 54540 37610
rect 59624 37558 59676 37610
rect 59688 37558 59740 37610
rect 59752 37558 59804 37610
rect 59816 37558 59868 37610
rect 64952 37558 65004 37610
rect 65016 37558 65068 37610
rect 65080 37558 65132 37610
rect 65144 37558 65196 37610
rect 70280 37558 70332 37610
rect 70344 37558 70396 37610
rect 70408 37558 70460 37610
rect 70472 37558 70524 37610
rect 75608 37558 75660 37610
rect 75672 37558 75724 37610
rect 75736 37558 75788 37610
rect 75800 37558 75852 37610
rect 80936 37558 80988 37610
rect 81000 37558 81052 37610
rect 81064 37558 81116 37610
rect 81128 37558 81180 37610
rect 86264 37558 86316 37610
rect 86328 37558 86380 37610
rect 86392 37558 86444 37610
rect 86456 37558 86508 37610
rect 91592 37558 91644 37610
rect 91656 37558 91708 37610
rect 91720 37558 91772 37610
rect 91784 37558 91836 37610
rect 3134 37456 3186 37508
rect 3962 37456 4014 37508
rect 5894 37456 5946 37508
rect 7458 37456 7510 37508
rect 10310 37456 10362 37508
rect 10494 37456 10546 37508
rect 7642 37388 7694 37440
rect 12794 37456 12846 37508
rect 19418 37456 19470 37508
rect 27054 37456 27106 37508
rect 27238 37499 27290 37508
rect 27238 37465 27247 37499
rect 27247 37465 27281 37499
rect 27281 37465 27290 37499
rect 27238 37456 27290 37465
rect 28894 37456 28946 37508
rect 32114 37499 32166 37508
rect 32114 37465 32123 37499
rect 32123 37465 32157 37499
rect 32157 37465 32166 37499
rect 32114 37456 32166 37465
rect 4422 37363 4474 37372
rect 4422 37329 4431 37363
rect 4431 37329 4465 37363
rect 4465 37329 4474 37363
rect 4422 37320 4474 37329
rect 10770 37363 10822 37372
rect 10770 37329 10779 37363
rect 10779 37329 10813 37363
rect 10813 37329 10822 37363
rect 10770 37320 10822 37329
rect 12058 37388 12110 37440
rect 11506 37320 11558 37372
rect 14174 37388 14226 37440
rect 16014 37388 16066 37440
rect 17670 37388 17722 37440
rect 27514 37388 27566 37440
rect 15830 37363 15882 37372
rect 15830 37329 15839 37363
rect 15839 37329 15873 37363
rect 15873 37329 15882 37363
rect 15830 37320 15882 37329
rect 17210 37363 17262 37372
rect 17210 37329 17219 37363
rect 17219 37329 17253 37363
rect 17253 37329 17262 37363
rect 17210 37320 17262 37329
rect 16474 37252 16526 37304
rect 20890 37320 20942 37372
rect 27422 37320 27474 37372
rect 32758 37388 32810 37440
rect 28802 37320 28854 37372
rect 21350 37252 21402 37304
rect 27698 37295 27750 37304
rect 27698 37261 27707 37295
rect 27707 37261 27741 37295
rect 27741 37261 27750 37295
rect 27698 37252 27750 37261
rect 31930 37320 31982 37372
rect 32666 37363 32718 37372
rect 32666 37329 32675 37363
rect 32675 37329 32709 37363
rect 32709 37329 32718 37363
rect 32666 37320 32718 37329
rect 29814 37252 29866 37304
rect 35058 37456 35110 37508
rect 35150 37456 35202 37508
rect 37726 37456 37778 37508
rect 36622 37388 36674 37440
rect 17578 37184 17630 37236
rect 32666 37184 32718 37236
rect 34966 37320 35018 37372
rect 40486 37456 40538 37508
rect 38002 37388 38054 37440
rect 37910 37363 37962 37372
rect 37910 37329 37919 37363
rect 37919 37329 37953 37363
rect 37953 37329 37962 37363
rect 40302 37388 40354 37440
rect 37910 37320 37962 37329
rect 39290 37320 39342 37372
rect 39750 37320 39802 37372
rect 47386 37456 47438 37508
rect 48490 37456 48542 37508
rect 40486 37295 40538 37304
rect 40486 37261 40495 37295
rect 40495 37261 40529 37295
rect 40529 37261 40538 37295
rect 42142 37320 42194 37372
rect 43614 37320 43666 37372
rect 45086 37320 45138 37372
rect 45362 37363 45414 37372
rect 45362 37329 45371 37363
rect 45371 37329 45405 37363
rect 45405 37329 45414 37363
rect 45362 37320 45414 37329
rect 40486 37252 40538 37261
rect 42878 37295 42930 37304
rect 38002 37184 38054 37236
rect 38094 37184 38146 37236
rect 39474 37184 39526 37236
rect 42878 37261 42887 37295
rect 42887 37261 42921 37295
rect 42921 37261 42930 37295
rect 42878 37252 42930 37261
rect 43062 37184 43114 37236
rect 17394 37116 17446 37168
rect 21534 37116 21586 37168
rect 29630 37159 29682 37168
rect 29630 37125 29639 37159
rect 29639 37125 29673 37159
rect 29673 37125 29682 37159
rect 29630 37116 29682 37125
rect 29814 37116 29866 37168
rect 39106 37116 39158 37168
rect 39290 37159 39342 37168
rect 39290 37125 39299 37159
rect 39299 37125 39333 37159
rect 39333 37125 39342 37159
rect 39290 37116 39342 37125
rect 39842 37116 39894 37168
rect 40394 37116 40446 37168
rect 42142 37116 42194 37168
rect 44166 37116 44218 37168
rect 45454 37116 45506 37168
rect 46558 37320 46610 37372
rect 46742 37363 46794 37372
rect 46742 37329 46751 37363
rect 46751 37329 46785 37363
rect 46785 37329 46794 37363
rect 46742 37320 46794 37329
rect 46926 37388 46978 37440
rect 48214 37252 48266 37304
rect 50606 37295 50658 37304
rect 50606 37261 50615 37295
rect 50615 37261 50649 37295
rect 50649 37261 50658 37295
rect 50606 37252 50658 37261
rect 51894 37388 51946 37440
rect 54930 37388 54982 37440
rect 52354 37320 52406 37372
rect 55022 37363 55074 37372
rect 55022 37329 55031 37363
rect 55031 37329 55065 37363
rect 55065 37329 55074 37363
rect 55022 37320 55074 37329
rect 55298 37456 55350 37508
rect 60358 37456 60410 37508
rect 61370 37456 61422 37508
rect 55206 37388 55258 37440
rect 58242 37388 58294 37440
rect 55482 37363 55534 37372
rect 55482 37329 55491 37363
rect 55491 37329 55525 37363
rect 55525 37329 55534 37363
rect 55482 37320 55534 37329
rect 55574 37363 55626 37372
rect 55574 37329 55583 37363
rect 55583 37329 55617 37363
rect 55617 37329 55626 37363
rect 55574 37320 55626 37329
rect 57966 37363 58018 37372
rect 57966 37329 57975 37363
rect 57975 37329 58009 37363
rect 58009 37329 58018 37363
rect 58610 37363 58662 37372
rect 57966 37320 58018 37329
rect 58610 37329 58619 37363
rect 58619 37329 58653 37363
rect 58653 37329 58662 37363
rect 58610 37320 58662 37329
rect 58886 37320 58938 37372
rect 54746 37252 54798 37304
rect 54838 37252 54890 37304
rect 48122 37184 48174 37236
rect 50422 37184 50474 37236
rect 56770 37252 56822 37304
rect 57138 37295 57190 37304
rect 57138 37261 57147 37295
rect 57147 37261 57181 37295
rect 57181 37261 57190 37295
rect 57138 37252 57190 37261
rect 59622 37295 59674 37304
rect 59622 37261 59631 37295
rect 59631 37261 59665 37295
rect 59665 37261 59674 37295
rect 59622 37252 59674 37261
rect 57966 37184 58018 37236
rect 47478 37116 47530 37168
rect 52170 37159 52222 37168
rect 52170 37125 52179 37159
rect 52179 37125 52213 37159
rect 52213 37125 52222 37159
rect 52170 37116 52222 37125
rect 52354 37159 52406 37168
rect 52354 37125 52363 37159
rect 52363 37125 52397 37159
rect 52397 37125 52406 37159
rect 52354 37116 52406 37125
rect 52538 37116 52590 37168
rect 59438 37184 59490 37236
rect 60174 37320 60226 37372
rect 60358 37363 60410 37372
rect 60358 37329 60367 37363
rect 60367 37329 60401 37363
rect 60401 37329 60410 37363
rect 60358 37320 60410 37329
rect 60542 37363 60594 37372
rect 60542 37329 60551 37363
rect 60551 37329 60585 37363
rect 60585 37329 60594 37363
rect 60542 37320 60594 37329
rect 62474 37388 62526 37440
rect 67074 37363 67126 37372
rect 67074 37329 67083 37363
rect 67083 37329 67117 37363
rect 67117 37329 67126 37363
rect 67074 37320 67126 37329
rect 69006 37388 69058 37440
rect 71582 37388 71634 37440
rect 72502 37388 72554 37440
rect 74434 37388 74486 37440
rect 75446 37456 75498 37508
rect 83266 37456 83318 37508
rect 88418 37456 88470 37508
rect 75906 37388 75958 37440
rect 68362 37320 68414 37372
rect 69190 37363 69242 37372
rect 69190 37329 69199 37363
rect 69199 37329 69233 37363
rect 69233 37329 69242 37363
rect 69190 37320 69242 37329
rect 69282 37320 69334 37372
rect 69650 37320 69702 37372
rect 72594 37320 72646 37372
rect 73054 37363 73106 37372
rect 73054 37329 73063 37363
rect 73063 37329 73097 37363
rect 73097 37329 73106 37363
rect 73054 37320 73106 37329
rect 73698 37320 73750 37372
rect 73882 37320 73934 37372
rect 74250 37363 74302 37372
rect 74250 37329 74259 37363
rect 74259 37329 74293 37363
rect 74293 37329 74302 37363
rect 74250 37320 74302 37329
rect 62106 37252 62158 37304
rect 68178 37252 68230 37304
rect 68270 37252 68322 37304
rect 68546 37295 68598 37304
rect 68546 37261 68555 37295
rect 68555 37261 68589 37295
rect 68589 37261 68598 37295
rect 68546 37252 68598 37261
rect 73606 37252 73658 37304
rect 73974 37252 74026 37304
rect 74986 37363 75038 37372
rect 74986 37329 74995 37363
rect 74995 37329 75029 37363
rect 75029 37329 75038 37363
rect 74986 37320 75038 37329
rect 75354 37320 75406 37372
rect 77470 37252 77522 37304
rect 60358 37184 60410 37236
rect 58242 37116 58294 37168
rect 60542 37116 60594 37168
rect 61186 37159 61238 37168
rect 61186 37125 61195 37159
rect 61195 37125 61229 37159
rect 61229 37125 61238 37159
rect 61186 37116 61238 37125
rect 62106 37116 62158 37168
rect 68454 37184 68506 37236
rect 69282 37184 69334 37236
rect 74250 37184 74302 37236
rect 63210 37116 63262 37168
rect 64038 37159 64090 37168
rect 64038 37125 64047 37159
rect 64047 37125 64081 37159
rect 64081 37125 64090 37159
rect 64038 37116 64090 37125
rect 67074 37116 67126 37168
rect 68638 37116 68690 37168
rect 70018 37116 70070 37168
rect 76642 37116 76694 37168
rect 76734 37116 76786 37168
rect 77470 37159 77522 37168
rect 77470 37125 77479 37159
rect 77479 37125 77513 37159
rect 77513 37125 77522 37159
rect 77470 37116 77522 37125
rect 82070 37363 82122 37372
rect 82070 37329 82079 37363
rect 82079 37329 82113 37363
rect 82113 37329 82122 37363
rect 82070 37320 82122 37329
rect 84278 37363 84330 37372
rect 84278 37329 84287 37363
rect 84287 37329 84321 37363
rect 84321 37329 84330 37363
rect 84278 37320 84330 37329
rect 90718 37456 90770 37508
rect 88326 37252 88378 37304
rect 89522 37363 89574 37372
rect 89522 37329 89531 37363
rect 89531 37329 89565 37363
rect 89565 37329 89574 37363
rect 89522 37320 89574 37329
rect 91362 37320 91414 37372
rect 89522 37184 89574 37236
rect 90258 37184 90310 37236
rect 78114 37116 78166 37168
rect 79218 37159 79270 37168
rect 79218 37125 79227 37159
rect 79227 37125 79261 37159
rect 79261 37125 79270 37159
rect 79218 37116 79270 37125
rect 80322 37159 80374 37168
rect 80322 37125 80331 37159
rect 80331 37125 80365 37159
rect 80365 37125 80374 37159
rect 80322 37116 80374 37125
rect 82714 37116 82766 37168
rect 83910 37159 83962 37168
rect 83910 37125 83919 37159
rect 83919 37125 83953 37159
rect 83953 37125 83962 37159
rect 83910 37116 83962 37125
rect 86578 37159 86630 37168
rect 86578 37125 86587 37159
rect 86587 37125 86621 37159
rect 86621 37125 86630 37159
rect 86578 37116 86630 37125
rect 3680 37014 3732 37066
rect 3744 37014 3796 37066
rect 3808 37014 3860 37066
rect 3872 37014 3924 37066
rect 9008 37014 9060 37066
rect 9072 37014 9124 37066
rect 9136 37014 9188 37066
rect 9200 37014 9252 37066
rect 14336 37014 14388 37066
rect 14400 37014 14452 37066
rect 14464 37014 14516 37066
rect 14528 37014 14580 37066
rect 19664 37014 19716 37066
rect 19728 37014 19780 37066
rect 19792 37014 19844 37066
rect 19856 37014 19908 37066
rect 24992 37014 25044 37066
rect 25056 37014 25108 37066
rect 25120 37014 25172 37066
rect 25184 37014 25236 37066
rect 30320 37014 30372 37066
rect 30384 37014 30436 37066
rect 30448 37014 30500 37066
rect 30512 37014 30564 37066
rect 35648 37014 35700 37066
rect 35712 37014 35764 37066
rect 35776 37014 35828 37066
rect 35840 37014 35892 37066
rect 40976 37014 41028 37066
rect 41040 37014 41092 37066
rect 41104 37014 41156 37066
rect 41168 37014 41220 37066
rect 46304 37014 46356 37066
rect 46368 37014 46420 37066
rect 46432 37014 46484 37066
rect 46496 37014 46548 37066
rect 51632 37014 51684 37066
rect 51696 37014 51748 37066
rect 51760 37014 51812 37066
rect 51824 37014 51876 37066
rect 56960 37014 57012 37066
rect 57024 37014 57076 37066
rect 57088 37014 57140 37066
rect 57152 37014 57204 37066
rect 62288 37014 62340 37066
rect 62352 37014 62404 37066
rect 62416 37014 62468 37066
rect 62480 37014 62532 37066
rect 67616 37014 67668 37066
rect 67680 37014 67732 37066
rect 67744 37014 67796 37066
rect 67808 37014 67860 37066
rect 72944 37014 72996 37066
rect 73008 37014 73060 37066
rect 73072 37014 73124 37066
rect 73136 37014 73188 37066
rect 78272 37014 78324 37066
rect 78336 37014 78388 37066
rect 78400 37014 78452 37066
rect 78464 37014 78516 37066
rect 83600 37014 83652 37066
rect 83664 37014 83716 37066
rect 83728 37014 83780 37066
rect 83792 37014 83844 37066
rect 88928 37014 88980 37066
rect 88992 37014 89044 37066
rect 89056 37014 89108 37066
rect 89120 37014 89172 37066
rect 2398 36912 2450 36964
rect 16014 36912 16066 36964
rect 17210 36912 17262 36964
rect 21350 36955 21402 36964
rect 21350 36921 21359 36955
rect 21359 36921 21393 36955
rect 21393 36921 21402 36955
rect 21350 36912 21402 36921
rect 27698 36912 27750 36964
rect 28250 36912 28302 36964
rect 29722 36912 29774 36964
rect 51434 36912 51486 36964
rect 51986 36912 52038 36964
rect 52170 36912 52222 36964
rect 52354 36912 52406 36964
rect 22822 36844 22874 36896
rect 27330 36844 27382 36896
rect 39290 36844 39342 36896
rect 40486 36887 40538 36896
rect 40486 36853 40495 36887
rect 40495 36853 40529 36887
rect 40529 36853 40538 36887
rect 40486 36844 40538 36853
rect 43062 36844 43114 36896
rect 43982 36887 44034 36896
rect 43982 36853 43991 36887
rect 43991 36853 44025 36887
rect 44025 36853 44034 36887
rect 43982 36844 44034 36853
rect 45546 36887 45598 36896
rect 45546 36853 45555 36887
rect 45555 36853 45589 36887
rect 45589 36853 45598 36887
rect 45546 36844 45598 36853
rect 51342 36844 51394 36896
rect 3134 36819 3186 36828
rect 3134 36785 3143 36819
rect 3143 36785 3177 36819
rect 3177 36785 3186 36819
rect 3134 36776 3186 36785
rect 15830 36776 15882 36828
rect 2490 36708 2542 36760
rect 3410 36751 3462 36760
rect 3410 36717 3419 36751
rect 3419 36717 3453 36751
rect 3453 36717 3462 36751
rect 3410 36708 3462 36717
rect 20338 36819 20390 36828
rect 5802 36640 5854 36692
rect 17670 36751 17722 36760
rect 17670 36717 17679 36751
rect 17679 36717 17713 36751
rect 17713 36717 17722 36751
rect 17670 36708 17722 36717
rect 20338 36785 20347 36819
rect 20347 36785 20381 36819
rect 20381 36785 20390 36819
rect 20338 36776 20390 36785
rect 31378 36819 31430 36828
rect 31378 36785 31387 36819
rect 31387 36785 31421 36819
rect 31421 36785 31430 36819
rect 31378 36776 31430 36785
rect 32114 36819 32166 36828
rect 32114 36785 32123 36819
rect 32123 36785 32157 36819
rect 32157 36785 32166 36819
rect 32114 36776 32166 36785
rect 32298 36776 32350 36828
rect 21258 36751 21310 36760
rect 21258 36717 21267 36751
rect 21267 36717 21301 36751
rect 21301 36717 21310 36751
rect 21258 36708 21310 36717
rect 28986 36708 29038 36760
rect 31930 36708 31982 36760
rect 32482 36708 32534 36760
rect 33494 36708 33546 36760
rect 33586 36708 33638 36760
rect 37542 36708 37594 36760
rect 43706 36776 43758 36828
rect 21534 36640 21586 36692
rect 32206 36640 32258 36692
rect 37450 36640 37502 36692
rect 4974 36615 5026 36624
rect 4974 36581 4983 36615
rect 4983 36581 5017 36615
rect 5017 36581 5026 36615
rect 4974 36572 5026 36581
rect 9482 36615 9534 36624
rect 9482 36581 9491 36615
rect 9491 36581 9525 36615
rect 9525 36581 9534 36615
rect 9482 36572 9534 36581
rect 10494 36572 10546 36624
rect 16198 36572 16250 36624
rect 28802 36615 28854 36624
rect 28802 36581 28811 36615
rect 28811 36581 28845 36615
rect 28845 36581 28854 36615
rect 28802 36572 28854 36581
rect 32022 36572 32074 36624
rect 32114 36572 32166 36624
rect 32758 36572 32810 36624
rect 34782 36572 34834 36624
rect 40854 36708 40906 36760
rect 42694 36751 42746 36760
rect 42694 36717 42703 36751
rect 42703 36717 42737 36751
rect 42737 36717 42746 36751
rect 42694 36708 42746 36717
rect 42878 36708 42930 36760
rect 43062 36708 43114 36760
rect 43246 36751 43298 36760
rect 43246 36717 43255 36751
rect 43255 36717 43289 36751
rect 43289 36717 43298 36751
rect 43246 36708 43298 36717
rect 45546 36708 45598 36760
rect 46558 36708 46610 36760
rect 46742 36751 46794 36760
rect 46742 36717 46751 36751
rect 46751 36717 46785 36751
rect 46785 36717 46794 36751
rect 46742 36708 46794 36717
rect 46834 36751 46886 36760
rect 46834 36717 46843 36751
rect 46843 36717 46877 36751
rect 46877 36717 46886 36751
rect 46834 36708 46886 36717
rect 47662 36708 47714 36760
rect 44074 36640 44126 36692
rect 50422 36640 50474 36692
rect 37726 36572 37778 36624
rect 37910 36572 37962 36624
rect 42694 36572 42746 36624
rect 43246 36572 43298 36624
rect 47662 36572 47714 36624
rect 50606 36640 50658 36692
rect 51802 36708 51854 36760
rect 52446 36776 52498 36828
rect 54930 36912 54982 36964
rect 57966 36912 58018 36964
rect 58058 36912 58110 36964
rect 62014 36912 62066 36964
rect 72502 36912 72554 36964
rect 72594 36912 72646 36964
rect 80322 36912 80374 36964
rect 82162 36912 82214 36964
rect 88326 36912 88378 36964
rect 88786 36912 88838 36964
rect 55482 36844 55534 36896
rect 61186 36844 61238 36896
rect 56126 36776 56178 36828
rect 65602 36776 65654 36828
rect 68086 36844 68138 36896
rect 68178 36844 68230 36896
rect 68730 36844 68782 36896
rect 57138 36708 57190 36760
rect 57782 36708 57834 36760
rect 58058 36751 58110 36760
rect 58058 36717 58067 36751
rect 58067 36717 58101 36751
rect 58101 36717 58110 36751
rect 58058 36708 58110 36717
rect 62934 36708 62986 36760
rect 63762 36708 63814 36760
rect 64038 36751 64090 36760
rect 64038 36717 64047 36751
rect 64047 36717 64081 36751
rect 64081 36717 64090 36751
rect 64038 36708 64090 36717
rect 69190 36819 69242 36828
rect 69190 36785 69199 36819
rect 69199 36785 69233 36819
rect 69233 36785 69242 36819
rect 69190 36776 69242 36785
rect 68362 36708 68414 36760
rect 68730 36751 68782 36760
rect 68730 36717 68739 36751
rect 68739 36717 68773 36751
rect 68773 36717 68782 36751
rect 73974 36844 74026 36896
rect 74066 36844 74118 36896
rect 72226 36776 72278 36828
rect 74710 36776 74762 36828
rect 79310 36819 79362 36828
rect 79310 36785 79319 36819
rect 79319 36785 79353 36819
rect 79353 36785 79362 36819
rect 79310 36776 79362 36785
rect 68730 36708 68782 36717
rect 52722 36640 52774 36692
rect 57690 36640 57742 36692
rect 58426 36640 58478 36692
rect 68914 36640 68966 36692
rect 51802 36572 51854 36624
rect 53366 36572 53418 36624
rect 53458 36572 53510 36624
rect 57782 36572 57834 36624
rect 58610 36572 58662 36624
rect 62474 36572 62526 36624
rect 65970 36572 66022 36624
rect 76458 36708 76510 36760
rect 79218 36751 79270 36760
rect 79218 36717 79227 36751
rect 79227 36717 79261 36751
rect 79261 36717 79270 36751
rect 79218 36708 79270 36717
rect 84002 36844 84054 36896
rect 84462 36776 84514 36828
rect 85474 36844 85526 36896
rect 88510 36844 88562 36896
rect 86578 36776 86630 36828
rect 82714 36708 82766 36760
rect 85474 36751 85526 36760
rect 85474 36717 85483 36751
rect 85483 36717 85517 36751
rect 85517 36717 85526 36751
rect 85474 36708 85526 36717
rect 85934 36751 85986 36760
rect 85934 36717 85943 36751
rect 85943 36717 85977 36751
rect 85977 36717 85986 36751
rect 88786 36751 88838 36760
rect 85934 36708 85986 36717
rect 88786 36717 88795 36751
rect 88795 36717 88829 36751
rect 88829 36717 88838 36751
rect 88786 36708 88838 36717
rect 89246 36708 89298 36760
rect 89522 36751 89574 36760
rect 89522 36717 89531 36751
rect 89531 36717 89565 36751
rect 89565 36717 89574 36751
rect 89522 36708 89574 36717
rect 86026 36640 86078 36692
rect 86394 36640 86446 36692
rect 76734 36572 76786 36624
rect 83082 36572 83134 36624
rect 85290 36572 85342 36624
rect 85934 36572 85986 36624
rect 6344 36470 6396 36522
rect 6408 36470 6460 36522
rect 6472 36470 6524 36522
rect 6536 36470 6588 36522
rect 11672 36470 11724 36522
rect 11736 36470 11788 36522
rect 11800 36470 11852 36522
rect 11864 36470 11916 36522
rect 17000 36470 17052 36522
rect 17064 36470 17116 36522
rect 17128 36470 17180 36522
rect 17192 36470 17244 36522
rect 22328 36470 22380 36522
rect 22392 36470 22444 36522
rect 22456 36470 22508 36522
rect 22520 36470 22572 36522
rect 27656 36470 27708 36522
rect 27720 36470 27772 36522
rect 27784 36470 27836 36522
rect 27848 36470 27900 36522
rect 32984 36470 33036 36522
rect 33048 36470 33100 36522
rect 33112 36470 33164 36522
rect 33176 36470 33228 36522
rect 38312 36470 38364 36522
rect 38376 36470 38428 36522
rect 38440 36470 38492 36522
rect 38504 36470 38556 36522
rect 43640 36470 43692 36522
rect 43704 36470 43756 36522
rect 43768 36470 43820 36522
rect 43832 36470 43884 36522
rect 48968 36470 49020 36522
rect 49032 36470 49084 36522
rect 49096 36470 49148 36522
rect 49160 36470 49212 36522
rect 54296 36470 54348 36522
rect 54360 36470 54412 36522
rect 54424 36470 54476 36522
rect 54488 36470 54540 36522
rect 59624 36470 59676 36522
rect 59688 36470 59740 36522
rect 59752 36470 59804 36522
rect 59816 36470 59868 36522
rect 64952 36470 65004 36522
rect 65016 36470 65068 36522
rect 65080 36470 65132 36522
rect 65144 36470 65196 36522
rect 70280 36470 70332 36522
rect 70344 36470 70396 36522
rect 70408 36470 70460 36522
rect 70472 36470 70524 36522
rect 75608 36470 75660 36522
rect 75672 36470 75724 36522
rect 75736 36470 75788 36522
rect 75800 36470 75852 36522
rect 80936 36470 80988 36522
rect 81000 36470 81052 36522
rect 81064 36470 81116 36522
rect 81128 36470 81180 36522
rect 86264 36470 86316 36522
rect 86328 36470 86380 36522
rect 86392 36470 86444 36522
rect 86456 36470 86508 36522
rect 91592 36470 91644 36522
rect 91656 36470 91708 36522
rect 91720 36470 91772 36522
rect 91784 36470 91836 36522
rect 2490 36411 2542 36420
rect 2490 36377 2499 36411
rect 2499 36377 2533 36411
rect 2533 36377 2542 36411
rect 2490 36368 2542 36377
rect 3410 36368 3462 36420
rect 4974 36368 5026 36420
rect 7458 36368 7510 36420
rect 9758 36411 9810 36420
rect 9758 36377 9767 36411
rect 9767 36377 9801 36411
rect 9801 36377 9810 36411
rect 9758 36368 9810 36377
rect 14910 36368 14962 36420
rect 17670 36368 17722 36420
rect 5802 36275 5854 36284
rect 5802 36241 5811 36275
rect 5811 36241 5845 36275
rect 5845 36241 5854 36275
rect 5802 36232 5854 36241
rect 10218 36232 10270 36284
rect 10494 36232 10546 36284
rect 11506 36232 11558 36284
rect 2674 36164 2726 36216
rect 16106 36232 16158 36284
rect 21534 36232 21586 36284
rect 24018 36275 24070 36284
rect 24018 36241 24027 36275
rect 24027 36241 24061 36275
rect 24061 36241 24070 36275
rect 24018 36232 24070 36241
rect 25674 36232 25726 36284
rect 12058 36207 12110 36216
rect 12058 36173 12067 36207
rect 12067 36173 12101 36207
rect 12101 36173 12110 36207
rect 12058 36164 12110 36173
rect 12610 36096 12662 36148
rect 12150 36028 12202 36080
rect 15554 36028 15606 36080
rect 16750 36207 16802 36216
rect 16750 36173 16759 36207
rect 16759 36173 16793 36207
rect 16793 36173 16802 36207
rect 16750 36164 16802 36173
rect 29354 36368 29406 36420
rect 29906 36368 29958 36420
rect 29078 36300 29130 36352
rect 39198 36343 39250 36352
rect 32114 36232 32166 36284
rect 28066 36164 28118 36216
rect 28342 36164 28394 36216
rect 32850 36207 32902 36216
rect 32850 36173 32859 36207
rect 32859 36173 32893 36207
rect 32893 36173 32902 36207
rect 32850 36164 32902 36173
rect 27054 36096 27106 36148
rect 20154 36028 20206 36080
rect 21534 36028 21586 36080
rect 23374 36028 23426 36080
rect 24570 36028 24622 36080
rect 29906 36096 29958 36148
rect 33586 36232 33638 36284
rect 39198 36309 39207 36343
rect 39207 36309 39241 36343
rect 39241 36309 39250 36343
rect 39198 36300 39250 36309
rect 40486 36343 40538 36352
rect 35058 36164 35110 36216
rect 38186 36164 38238 36216
rect 28986 36071 29038 36080
rect 28986 36037 28995 36071
rect 28995 36037 29029 36071
rect 29029 36037 29038 36071
rect 28986 36028 29038 36037
rect 29262 36028 29314 36080
rect 34506 36096 34558 36148
rect 37634 36096 37686 36148
rect 39842 36275 39894 36284
rect 39842 36241 39851 36275
rect 39851 36241 39885 36275
rect 39885 36241 39894 36275
rect 39842 36232 39894 36241
rect 40486 36309 40495 36343
rect 40495 36309 40529 36343
rect 40529 36309 40538 36343
rect 40486 36300 40538 36309
rect 40578 36300 40630 36352
rect 49318 36300 49370 36352
rect 51342 36300 51394 36352
rect 52262 36300 52314 36352
rect 61462 36300 61514 36352
rect 45362 36275 45414 36284
rect 45362 36241 45371 36275
rect 45371 36241 45405 36275
rect 45405 36241 45414 36275
rect 45362 36232 45414 36241
rect 45638 36275 45690 36284
rect 45638 36241 45647 36275
rect 45647 36241 45681 36275
rect 45681 36241 45690 36275
rect 45638 36232 45690 36241
rect 39658 36207 39710 36216
rect 39658 36173 39667 36207
rect 39667 36173 39701 36207
rect 39701 36173 39710 36207
rect 39658 36164 39710 36173
rect 40118 36207 40170 36216
rect 40118 36173 40127 36207
rect 40127 36173 40161 36207
rect 40161 36173 40170 36207
rect 40118 36164 40170 36173
rect 45086 36164 45138 36216
rect 48858 36164 48910 36216
rect 51342 36164 51394 36216
rect 51618 36275 51670 36284
rect 51618 36241 51627 36275
rect 51627 36241 51661 36275
rect 51661 36241 51670 36275
rect 51618 36232 51670 36241
rect 52722 36232 52774 36284
rect 53366 36232 53418 36284
rect 56770 36275 56822 36284
rect 56770 36241 56779 36275
rect 56779 36241 56813 36275
rect 56813 36241 56822 36275
rect 56770 36232 56822 36241
rect 61830 36275 61882 36284
rect 61830 36241 61839 36275
rect 61839 36241 61873 36275
rect 61873 36241 61882 36275
rect 61830 36232 61882 36241
rect 51894 36207 51946 36216
rect 51526 36096 51578 36148
rect 51618 36096 51670 36148
rect 51894 36173 51903 36207
rect 51903 36173 51937 36207
rect 51937 36173 51946 36207
rect 51894 36164 51946 36173
rect 52078 36164 52130 36216
rect 56126 36164 56178 36216
rect 57138 36164 57190 36216
rect 61554 36207 61606 36216
rect 33954 36028 34006 36080
rect 34138 36028 34190 36080
rect 39842 36028 39894 36080
rect 42878 36028 42930 36080
rect 48398 36028 48450 36080
rect 52354 36071 52406 36080
rect 52354 36037 52363 36071
rect 52363 36037 52397 36071
rect 52397 36037 52406 36071
rect 52354 36028 52406 36037
rect 52722 36028 52774 36080
rect 61554 36173 61563 36207
rect 61563 36173 61597 36207
rect 61597 36173 61606 36207
rect 61554 36164 61606 36173
rect 58058 36139 58110 36148
rect 58058 36105 58067 36139
rect 58067 36105 58101 36139
rect 58101 36105 58110 36139
rect 58058 36096 58110 36105
rect 61462 36096 61514 36148
rect 61738 36164 61790 36216
rect 63302 36232 63354 36284
rect 59070 36028 59122 36080
rect 62566 36096 62618 36148
rect 65602 36368 65654 36420
rect 68178 36368 68230 36420
rect 82162 36368 82214 36420
rect 82530 36368 82582 36420
rect 88234 36368 88286 36420
rect 69190 36232 69242 36284
rect 73330 36275 73382 36284
rect 73330 36241 73339 36275
rect 73339 36241 73373 36275
rect 73373 36241 73382 36275
rect 73330 36232 73382 36241
rect 73606 36232 73658 36284
rect 74158 36232 74210 36284
rect 75262 36232 75314 36284
rect 66522 36096 66574 36148
rect 63026 36028 63078 36080
rect 63210 36071 63262 36080
rect 63210 36037 63219 36071
rect 63219 36037 63253 36071
rect 63253 36037 63262 36071
rect 63210 36028 63262 36037
rect 64130 36028 64182 36080
rect 69650 36164 69702 36216
rect 69374 36096 69426 36148
rect 70110 36096 70162 36148
rect 82714 36275 82766 36284
rect 82714 36241 82723 36275
rect 82723 36241 82757 36275
rect 82757 36241 82766 36275
rect 82714 36232 82766 36241
rect 83082 36275 83134 36284
rect 83082 36241 83091 36275
rect 83091 36241 83125 36275
rect 83125 36241 83134 36275
rect 83082 36232 83134 36241
rect 86026 36232 86078 36284
rect 88694 36232 88746 36284
rect 82530 36207 82582 36216
rect 82530 36173 82539 36207
rect 82539 36173 82573 36207
rect 82573 36173 82582 36207
rect 82530 36164 82582 36173
rect 89522 36275 89574 36284
rect 89522 36241 89531 36275
rect 89531 36241 89565 36275
rect 89565 36241 89574 36275
rect 91362 36275 91414 36284
rect 89522 36232 89574 36241
rect 82714 36096 82766 36148
rect 69006 36071 69058 36080
rect 69006 36037 69015 36071
rect 69015 36037 69049 36071
rect 69049 36037 69058 36071
rect 69006 36028 69058 36037
rect 74526 36071 74578 36080
rect 74526 36037 74535 36071
rect 74535 36037 74569 36071
rect 74569 36037 74578 36071
rect 74526 36028 74578 36037
rect 85658 36028 85710 36080
rect 91362 36241 91371 36275
rect 91371 36241 91405 36275
rect 91405 36241 91414 36275
rect 91362 36232 91414 36241
rect 90442 36096 90494 36148
rect 90718 36028 90770 36080
rect 3680 35926 3732 35978
rect 3744 35926 3796 35978
rect 3808 35926 3860 35978
rect 3872 35926 3924 35978
rect 9008 35926 9060 35978
rect 9072 35926 9124 35978
rect 9136 35926 9188 35978
rect 9200 35926 9252 35978
rect 14336 35926 14388 35978
rect 14400 35926 14452 35978
rect 14464 35926 14516 35978
rect 14528 35926 14580 35978
rect 19664 35926 19716 35978
rect 19728 35926 19780 35978
rect 19792 35926 19844 35978
rect 19856 35926 19908 35978
rect 24992 35926 25044 35978
rect 25056 35926 25108 35978
rect 25120 35926 25172 35978
rect 25184 35926 25236 35978
rect 30320 35926 30372 35978
rect 30384 35926 30436 35978
rect 30448 35926 30500 35978
rect 30512 35926 30564 35978
rect 35648 35926 35700 35978
rect 35712 35926 35764 35978
rect 35776 35926 35828 35978
rect 35840 35926 35892 35978
rect 40976 35926 41028 35978
rect 41040 35926 41092 35978
rect 41104 35926 41156 35978
rect 41168 35926 41220 35978
rect 46304 35926 46356 35978
rect 46368 35926 46420 35978
rect 46432 35926 46484 35978
rect 46496 35926 46548 35978
rect 51632 35926 51684 35978
rect 51696 35926 51748 35978
rect 51760 35926 51812 35978
rect 51824 35926 51876 35978
rect 56960 35926 57012 35978
rect 57024 35926 57076 35978
rect 57088 35926 57140 35978
rect 57152 35926 57204 35978
rect 62288 35926 62340 35978
rect 62352 35926 62404 35978
rect 62416 35926 62468 35978
rect 62480 35926 62532 35978
rect 67616 35926 67668 35978
rect 67680 35926 67732 35978
rect 67744 35926 67796 35978
rect 67808 35926 67860 35978
rect 72944 35926 72996 35978
rect 73008 35926 73060 35978
rect 73072 35926 73124 35978
rect 73136 35926 73188 35978
rect 78272 35926 78324 35978
rect 78336 35926 78388 35978
rect 78400 35926 78452 35978
rect 78464 35926 78516 35978
rect 83600 35926 83652 35978
rect 83664 35926 83716 35978
rect 83728 35926 83780 35978
rect 83792 35926 83844 35978
rect 88928 35926 88980 35978
rect 88992 35926 89044 35978
rect 89056 35926 89108 35978
rect 89120 35926 89172 35978
rect 16750 35824 16802 35876
rect 10218 35756 10270 35808
rect 2674 35731 2726 35740
rect 2674 35697 2683 35731
rect 2683 35697 2717 35731
rect 2717 35697 2726 35731
rect 2674 35688 2726 35697
rect 10494 35688 10546 35740
rect 10586 35620 10638 35672
rect 18498 35756 18550 35808
rect 12150 35731 12202 35740
rect 12150 35697 12159 35731
rect 12159 35697 12193 35731
rect 12193 35697 12202 35731
rect 12150 35688 12202 35697
rect 11322 35620 11374 35672
rect 11414 35552 11466 35604
rect 3962 35527 4014 35536
rect 3962 35493 3971 35527
rect 3971 35493 4005 35527
rect 4005 35493 4014 35527
rect 3962 35484 4014 35493
rect 4238 35527 4290 35536
rect 4238 35493 4247 35527
rect 4247 35493 4281 35527
rect 4281 35493 4290 35527
rect 4238 35484 4290 35493
rect 10126 35484 10178 35536
rect 12610 35484 12662 35536
rect 16106 35620 16158 35672
rect 21626 35824 21678 35876
rect 22822 35824 22874 35876
rect 40578 35824 40630 35876
rect 48398 35867 48450 35876
rect 27054 35756 27106 35808
rect 30458 35756 30510 35808
rect 23374 35731 23426 35740
rect 17578 35663 17630 35672
rect 17578 35629 17587 35663
rect 17587 35629 17621 35663
rect 17621 35629 17630 35663
rect 17578 35620 17630 35629
rect 23374 35697 23383 35731
rect 23383 35697 23417 35731
rect 23417 35697 23426 35731
rect 23374 35688 23426 35697
rect 32850 35756 32902 35808
rect 34046 35756 34098 35808
rect 34506 35799 34558 35808
rect 34506 35765 34515 35799
rect 34515 35765 34549 35799
rect 34549 35765 34558 35799
rect 34506 35756 34558 35765
rect 34782 35799 34834 35808
rect 34782 35765 34791 35799
rect 34791 35765 34825 35799
rect 34825 35765 34834 35799
rect 34782 35756 34834 35765
rect 39566 35756 39618 35808
rect 48398 35833 48407 35867
rect 48407 35833 48441 35867
rect 48441 35833 48450 35867
rect 48398 35824 48450 35833
rect 21074 35663 21126 35672
rect 14082 35484 14134 35536
rect 15554 35484 15606 35536
rect 16842 35484 16894 35536
rect 20522 35552 20574 35604
rect 21074 35629 21083 35663
rect 21083 35629 21117 35663
rect 21117 35629 21126 35663
rect 21074 35620 21126 35629
rect 38094 35688 38146 35740
rect 21534 35552 21586 35604
rect 22822 35552 22874 35604
rect 25674 35663 25726 35672
rect 25674 35629 25683 35663
rect 25683 35629 25717 35663
rect 25717 35629 25726 35663
rect 25674 35620 25726 35629
rect 28250 35620 28302 35672
rect 29354 35663 29406 35672
rect 29354 35629 29363 35663
rect 29363 35629 29397 35663
rect 29397 35629 29406 35663
rect 29354 35620 29406 35629
rect 30274 35620 30326 35672
rect 32114 35663 32166 35672
rect 32114 35629 32123 35663
rect 32123 35629 32157 35663
rect 32157 35629 32166 35663
rect 32114 35620 32166 35629
rect 32022 35552 32074 35604
rect 32758 35620 32810 35672
rect 33310 35552 33362 35604
rect 18498 35527 18550 35536
rect 18498 35493 18507 35527
rect 18507 35493 18541 35527
rect 18541 35493 18550 35527
rect 18498 35484 18550 35493
rect 23834 35484 23886 35536
rect 29078 35484 29130 35536
rect 29354 35484 29406 35536
rect 30090 35527 30142 35536
rect 30090 35493 30099 35527
rect 30099 35493 30133 35527
rect 30133 35493 30142 35527
rect 30090 35484 30142 35493
rect 34782 35620 34834 35672
rect 37174 35620 37226 35672
rect 42878 35688 42930 35740
rect 44074 35688 44126 35740
rect 47662 35688 47714 35740
rect 35518 35552 35570 35604
rect 40026 35620 40078 35672
rect 39842 35552 39894 35604
rect 36070 35484 36122 35536
rect 37174 35527 37226 35536
rect 37174 35493 37183 35527
rect 37183 35493 37217 35527
rect 37217 35493 37226 35527
rect 37174 35484 37226 35493
rect 40762 35484 40814 35536
rect 44626 35595 44678 35604
rect 44626 35561 44635 35595
rect 44635 35561 44669 35595
rect 44669 35561 44678 35595
rect 46742 35620 46794 35672
rect 48398 35620 48450 35672
rect 48858 35663 48910 35672
rect 48858 35629 48867 35663
rect 48867 35629 48901 35663
rect 48901 35629 48910 35663
rect 48858 35620 48910 35629
rect 54194 35824 54246 35876
rect 53182 35620 53234 35672
rect 53458 35620 53510 35672
rect 80690 35824 80742 35876
rect 85842 35824 85894 35876
rect 91362 35824 91414 35876
rect 55574 35756 55626 35808
rect 56678 35620 56730 35672
rect 57874 35688 57926 35740
rect 58334 35663 58386 35672
rect 58334 35629 58343 35663
rect 58343 35629 58377 35663
rect 58377 35629 58386 35663
rect 58334 35620 58386 35629
rect 58886 35663 58938 35672
rect 44626 35552 44678 35561
rect 43062 35484 43114 35536
rect 43982 35484 44034 35536
rect 49410 35552 49462 35604
rect 51986 35552 52038 35604
rect 54654 35552 54706 35604
rect 58886 35629 58895 35663
rect 58895 35629 58929 35663
rect 58929 35629 58938 35663
rect 58886 35620 58938 35629
rect 59070 35663 59122 35672
rect 59070 35629 59079 35663
rect 59079 35629 59113 35663
rect 59113 35629 59122 35663
rect 59070 35620 59122 35629
rect 59990 35688 60042 35740
rect 61830 35688 61882 35740
rect 60174 35620 60226 35672
rect 62382 35663 62434 35672
rect 62382 35629 62391 35663
rect 62391 35629 62425 35663
rect 62425 35629 62434 35663
rect 62382 35620 62434 35629
rect 62566 35663 62618 35672
rect 62566 35629 62575 35663
rect 62575 35629 62609 35663
rect 62609 35629 62618 35663
rect 62566 35620 62618 35629
rect 46650 35484 46702 35536
rect 47110 35484 47162 35536
rect 51894 35484 51946 35536
rect 52354 35484 52406 35536
rect 52630 35484 52682 35536
rect 53274 35484 53326 35536
rect 54010 35484 54062 35536
rect 54194 35484 54246 35536
rect 60266 35552 60318 35604
rect 63302 35620 63354 35672
rect 67442 35756 67494 35808
rect 68362 35756 68414 35808
rect 75262 35756 75314 35808
rect 63946 35731 63998 35740
rect 63946 35697 63955 35731
rect 63955 35697 63989 35731
rect 63989 35697 63998 35731
rect 63946 35688 63998 35697
rect 67902 35688 67954 35740
rect 69282 35731 69334 35740
rect 69282 35697 69291 35731
rect 69291 35697 69325 35731
rect 69325 35697 69334 35731
rect 69282 35688 69334 35697
rect 66890 35552 66942 35604
rect 61922 35484 61974 35536
rect 62106 35527 62158 35536
rect 62106 35493 62115 35527
rect 62115 35493 62149 35527
rect 62149 35493 62158 35527
rect 62106 35484 62158 35493
rect 62566 35484 62618 35536
rect 63210 35484 63262 35536
rect 63578 35527 63630 35536
rect 63578 35493 63587 35527
rect 63587 35493 63621 35527
rect 63621 35493 63630 35527
rect 63578 35484 63630 35493
rect 64130 35527 64182 35536
rect 64130 35493 64139 35527
rect 64139 35493 64173 35527
rect 64173 35493 64182 35527
rect 64130 35484 64182 35493
rect 68914 35620 68966 35672
rect 73238 35688 73290 35740
rect 73330 35688 73382 35740
rect 73698 35688 73750 35740
rect 69558 35620 69610 35672
rect 73790 35663 73842 35672
rect 70662 35595 70714 35604
rect 70662 35561 70671 35595
rect 70671 35561 70705 35595
rect 70705 35561 70714 35595
rect 70662 35552 70714 35561
rect 70110 35484 70162 35536
rect 73790 35629 73799 35663
rect 73799 35629 73833 35663
rect 73833 35629 73842 35663
rect 73790 35620 73842 35629
rect 85474 35688 85526 35740
rect 74342 35663 74394 35672
rect 74342 35629 74351 35663
rect 74351 35629 74385 35663
rect 74385 35629 74394 35663
rect 74342 35620 74394 35629
rect 74066 35484 74118 35536
rect 74158 35484 74210 35536
rect 75446 35484 75498 35536
rect 81794 35620 81846 35672
rect 82070 35663 82122 35672
rect 82070 35629 82079 35663
rect 82079 35629 82113 35663
rect 82113 35629 82122 35663
rect 82070 35620 82122 35629
rect 82714 35663 82766 35672
rect 82714 35629 82723 35663
rect 82723 35629 82757 35663
rect 82757 35629 82766 35663
rect 82714 35620 82766 35629
rect 85658 35620 85710 35672
rect 86578 35688 86630 35740
rect 88234 35731 88286 35740
rect 88234 35697 88243 35731
rect 88243 35697 88277 35731
rect 88277 35697 88286 35731
rect 88234 35688 88286 35697
rect 90718 35731 90770 35740
rect 90718 35697 90727 35731
rect 90727 35697 90761 35731
rect 90761 35697 90770 35731
rect 90718 35688 90770 35697
rect 80230 35484 80282 35536
rect 81702 35527 81754 35536
rect 81702 35493 81711 35527
rect 81711 35493 81745 35527
rect 81745 35493 81754 35527
rect 81702 35484 81754 35493
rect 83542 35552 83594 35604
rect 86026 35620 86078 35672
rect 88326 35663 88378 35672
rect 86578 35552 86630 35604
rect 88326 35629 88335 35663
rect 88335 35629 88369 35663
rect 88369 35629 88378 35663
rect 88326 35620 88378 35629
rect 88786 35663 88838 35672
rect 88786 35629 88795 35663
rect 88795 35629 88829 35663
rect 88829 35629 88838 35663
rect 88786 35620 88838 35629
rect 87774 35552 87826 35604
rect 89982 35552 90034 35604
rect 86670 35527 86722 35536
rect 86670 35493 86679 35527
rect 86679 35493 86713 35527
rect 86713 35493 86722 35527
rect 86670 35484 86722 35493
rect 89522 35484 89574 35536
rect 6344 35382 6396 35434
rect 6408 35382 6460 35434
rect 6472 35382 6524 35434
rect 6536 35382 6588 35434
rect 11672 35382 11724 35434
rect 11736 35382 11788 35434
rect 11800 35382 11852 35434
rect 11864 35382 11916 35434
rect 17000 35382 17052 35434
rect 17064 35382 17116 35434
rect 17128 35382 17180 35434
rect 17192 35382 17244 35434
rect 22328 35382 22380 35434
rect 22392 35382 22444 35434
rect 22456 35382 22508 35434
rect 22520 35382 22572 35434
rect 27656 35382 27708 35434
rect 27720 35382 27772 35434
rect 27784 35382 27836 35434
rect 27848 35382 27900 35434
rect 32984 35382 33036 35434
rect 33048 35382 33100 35434
rect 33112 35382 33164 35434
rect 33176 35382 33228 35434
rect 38312 35382 38364 35434
rect 38376 35382 38428 35434
rect 38440 35382 38492 35434
rect 38504 35382 38556 35434
rect 43640 35382 43692 35434
rect 43704 35382 43756 35434
rect 43768 35382 43820 35434
rect 43832 35382 43884 35434
rect 48968 35382 49020 35434
rect 49032 35382 49084 35434
rect 49096 35382 49148 35434
rect 49160 35382 49212 35434
rect 54296 35382 54348 35434
rect 54360 35382 54412 35434
rect 54424 35382 54476 35434
rect 54488 35382 54540 35434
rect 59624 35382 59676 35434
rect 59688 35382 59740 35434
rect 59752 35382 59804 35434
rect 59816 35382 59868 35434
rect 64952 35382 65004 35434
rect 65016 35382 65068 35434
rect 65080 35382 65132 35434
rect 65144 35382 65196 35434
rect 70280 35382 70332 35434
rect 70344 35382 70396 35434
rect 70408 35382 70460 35434
rect 70472 35382 70524 35434
rect 75608 35382 75660 35434
rect 75672 35382 75724 35434
rect 75736 35382 75788 35434
rect 75800 35382 75852 35434
rect 80936 35382 80988 35434
rect 81000 35382 81052 35434
rect 81064 35382 81116 35434
rect 81128 35382 81180 35434
rect 86264 35382 86316 35434
rect 86328 35382 86380 35434
rect 86392 35382 86444 35434
rect 86456 35382 86508 35434
rect 91592 35382 91644 35434
rect 91656 35382 91708 35434
rect 91720 35382 91772 35434
rect 91784 35382 91836 35434
rect 2674 35280 2726 35332
rect 10586 35280 10638 35332
rect 11966 35280 12018 35332
rect 12794 35280 12846 35332
rect 15554 35323 15606 35332
rect 15554 35289 15563 35323
rect 15563 35289 15597 35323
rect 15597 35289 15606 35323
rect 15554 35280 15606 35289
rect 18958 35280 19010 35332
rect 19418 35323 19470 35332
rect 19418 35289 19427 35323
rect 19427 35289 19461 35323
rect 19461 35289 19470 35323
rect 19418 35280 19470 35289
rect 21166 35280 21218 35332
rect 23834 35280 23886 35332
rect 24018 35323 24070 35332
rect 24018 35289 24027 35323
rect 24027 35289 24061 35323
rect 24061 35289 24070 35323
rect 24018 35280 24070 35289
rect 28066 35280 28118 35332
rect 15094 35255 15146 35264
rect 2582 35144 2634 35196
rect 3962 35144 4014 35196
rect 10126 35187 10178 35196
rect 10126 35153 10135 35187
rect 10135 35153 10169 35187
rect 10169 35153 10178 35187
rect 10126 35144 10178 35153
rect 11414 35144 11466 35196
rect 15094 35221 15103 35255
rect 15103 35221 15137 35255
rect 15137 35221 15146 35255
rect 15094 35212 15146 35221
rect 17578 35212 17630 35264
rect 14726 35187 14778 35196
rect 4238 35076 4290 35128
rect 11322 35076 11374 35128
rect 14726 35153 14735 35187
rect 14735 35153 14769 35187
rect 14769 35153 14778 35187
rect 14726 35144 14778 35153
rect 20154 35212 20206 35264
rect 15554 35076 15606 35128
rect 16014 35119 16066 35128
rect 16014 35085 16023 35119
rect 16023 35085 16057 35119
rect 16057 35085 16066 35119
rect 16014 35076 16066 35085
rect 18958 35144 19010 35196
rect 21074 35144 21126 35196
rect 21718 35144 21770 35196
rect 24570 35212 24622 35264
rect 29262 35280 29314 35332
rect 35518 35280 35570 35332
rect 23282 35144 23334 35196
rect 23834 35187 23886 35196
rect 23834 35153 23843 35187
rect 23843 35153 23877 35187
rect 23877 35153 23886 35187
rect 23834 35144 23886 35153
rect 27054 35187 27106 35196
rect 27054 35153 27063 35187
rect 27063 35153 27097 35187
rect 27097 35153 27106 35187
rect 27054 35144 27106 35153
rect 28986 35212 29038 35264
rect 28802 35144 28854 35196
rect 30274 35187 30326 35196
rect 30274 35153 30283 35187
rect 30283 35153 30317 35187
rect 30317 35153 30326 35187
rect 30274 35144 30326 35153
rect 30458 35212 30510 35264
rect 32022 35144 32074 35196
rect 33126 35187 33178 35196
rect 33126 35153 33135 35187
rect 33135 35153 33169 35187
rect 33169 35153 33178 35187
rect 33126 35144 33178 35153
rect 30090 35076 30142 35128
rect 30734 35076 30786 35128
rect 33402 35187 33454 35196
rect 33402 35153 33411 35187
rect 33411 35153 33445 35187
rect 33445 35153 33454 35187
rect 33402 35144 33454 35153
rect 34230 35144 34282 35196
rect 40026 35280 40078 35332
rect 43062 35323 43114 35332
rect 43062 35289 43071 35323
rect 43071 35289 43105 35323
rect 43105 35289 43114 35323
rect 43062 35280 43114 35289
rect 46098 35280 46150 35332
rect 48214 35280 48266 35332
rect 49318 35323 49370 35332
rect 49318 35289 49327 35323
rect 49327 35289 49361 35323
rect 49361 35289 49370 35323
rect 49318 35280 49370 35289
rect 49410 35280 49462 35332
rect 62106 35280 62158 35332
rect 64038 35280 64090 35332
rect 64130 35280 64182 35332
rect 69558 35280 69610 35332
rect 69650 35280 69702 35332
rect 75446 35280 75498 35332
rect 80690 35280 80742 35332
rect 40578 35212 40630 35264
rect 36070 35144 36122 35196
rect 37818 35187 37870 35196
rect 37818 35153 37827 35187
rect 37827 35153 37861 35187
rect 37861 35153 37870 35187
rect 37818 35144 37870 35153
rect 39842 35144 39894 35196
rect 47478 35212 47530 35264
rect 44166 35144 44218 35196
rect 45178 35144 45230 35196
rect 47570 35144 47622 35196
rect 49318 35144 49370 35196
rect 51894 35187 51946 35196
rect 51894 35153 51903 35187
rect 51903 35153 51937 35187
rect 51937 35153 51946 35187
rect 51894 35144 51946 35153
rect 22730 35051 22782 35060
rect 7090 34983 7142 34992
rect 7090 34949 7099 34983
rect 7099 34949 7133 34983
rect 7133 34949 7142 34983
rect 7090 34940 7142 34949
rect 8378 34940 8430 34992
rect 11322 34940 11374 34992
rect 13530 34983 13582 34992
rect 13530 34949 13539 34983
rect 13539 34949 13573 34983
rect 13573 34949 13582 34983
rect 13530 34940 13582 34949
rect 17302 34983 17354 34992
rect 17302 34949 17311 34983
rect 17311 34949 17345 34983
rect 17345 34949 17354 34983
rect 17302 34940 17354 34949
rect 22730 35017 22739 35051
rect 22739 35017 22773 35051
rect 22773 35017 22782 35051
rect 22730 35008 22782 35017
rect 34598 35008 34650 35060
rect 37174 35008 37226 35060
rect 40118 35076 40170 35128
rect 43430 35076 43482 35128
rect 46098 35076 46150 35128
rect 52078 35144 52130 35196
rect 24294 34940 24346 34992
rect 30642 34940 30694 34992
rect 39474 34940 39526 34992
rect 41314 34940 41366 34992
rect 53366 35144 53418 35196
rect 52722 35076 52774 35128
rect 54102 35212 54154 35264
rect 60818 35212 60870 35264
rect 63302 35212 63354 35264
rect 80874 35212 80926 35264
rect 82070 35212 82122 35264
rect 62566 35144 62618 35196
rect 63118 35187 63170 35196
rect 63118 35153 63127 35187
rect 63127 35153 63161 35187
rect 63161 35153 63170 35187
rect 63118 35144 63170 35153
rect 63210 35187 63262 35196
rect 63210 35153 63219 35187
rect 63219 35153 63253 35187
rect 63253 35153 63262 35187
rect 65878 35187 65930 35196
rect 63210 35144 63262 35153
rect 54654 35119 54706 35128
rect 54654 35085 54663 35119
rect 54663 35085 54697 35119
rect 54697 35085 54706 35119
rect 54654 35076 54706 35085
rect 55850 35076 55902 35128
rect 62106 35076 62158 35128
rect 65878 35153 65887 35187
rect 65887 35153 65921 35187
rect 65921 35153 65930 35187
rect 65878 35144 65930 35153
rect 68362 35144 68414 35196
rect 70662 35144 70714 35196
rect 73238 35144 73290 35196
rect 73974 35144 74026 35196
rect 74158 35187 74210 35196
rect 74158 35153 74167 35187
rect 74167 35153 74201 35187
rect 74201 35153 74210 35187
rect 74158 35144 74210 35153
rect 67902 35076 67954 35128
rect 68178 35076 68230 35128
rect 69282 35119 69334 35128
rect 63394 35008 63446 35060
rect 69282 35085 69291 35119
rect 69291 35085 69325 35119
rect 69325 35085 69334 35119
rect 69282 35076 69334 35085
rect 69926 35119 69978 35128
rect 69926 35085 69935 35119
rect 69935 35085 69969 35119
rect 69969 35085 69978 35119
rect 69926 35076 69978 35085
rect 76734 35076 76786 35128
rect 81150 35144 81202 35196
rect 83910 35280 83962 35332
rect 89522 35323 89574 35332
rect 89522 35289 89531 35323
rect 89531 35289 89565 35323
rect 89565 35289 89574 35323
rect 89522 35280 89574 35289
rect 83542 35187 83594 35196
rect 83542 35153 83551 35187
rect 83551 35153 83585 35187
rect 83585 35153 83594 35187
rect 83542 35144 83594 35153
rect 89982 35187 90034 35196
rect 89982 35153 89991 35187
rect 89991 35153 90025 35187
rect 90025 35153 90034 35187
rect 89982 35144 90034 35153
rect 46926 34940 46978 34992
rect 52630 34983 52682 34992
rect 52630 34949 52639 34983
rect 52639 34949 52673 34983
rect 52673 34949 52682 34983
rect 52630 34940 52682 34949
rect 52722 34983 52774 34992
rect 52722 34949 52731 34983
rect 52731 34949 52765 34983
rect 52765 34949 52774 34983
rect 52722 34940 52774 34949
rect 54102 34940 54154 34992
rect 54286 34983 54338 34992
rect 54286 34949 54295 34983
rect 54295 34949 54329 34983
rect 54329 34949 54338 34983
rect 54286 34940 54338 34949
rect 55298 34940 55350 34992
rect 63854 34940 63906 34992
rect 65970 34983 66022 34992
rect 65970 34949 65979 34983
rect 65979 34949 66013 34983
rect 66013 34949 66022 34983
rect 65970 34940 66022 34949
rect 68362 34983 68414 34992
rect 68362 34949 68371 34983
rect 68371 34949 68405 34983
rect 68405 34949 68414 34983
rect 68362 34940 68414 34949
rect 69742 35008 69794 35060
rect 75446 34940 75498 34992
rect 84278 35008 84330 35060
rect 82898 34940 82950 34992
rect 84646 34983 84698 34992
rect 84646 34949 84655 34983
rect 84655 34949 84689 34983
rect 84689 34949 84698 34983
rect 84646 34940 84698 34949
rect 90626 34940 90678 34992
rect 91086 34983 91138 34992
rect 91086 34949 91095 34983
rect 91095 34949 91129 34983
rect 91129 34949 91138 34983
rect 91086 34940 91138 34949
rect 3680 34838 3732 34890
rect 3744 34838 3796 34890
rect 3808 34838 3860 34890
rect 3872 34838 3924 34890
rect 9008 34838 9060 34890
rect 9072 34838 9124 34890
rect 9136 34838 9188 34890
rect 9200 34838 9252 34890
rect 14336 34838 14388 34890
rect 14400 34838 14452 34890
rect 14464 34838 14516 34890
rect 14528 34838 14580 34890
rect 19664 34838 19716 34890
rect 19728 34838 19780 34890
rect 19792 34838 19844 34890
rect 19856 34838 19908 34890
rect 24992 34838 25044 34890
rect 25056 34838 25108 34890
rect 25120 34838 25172 34890
rect 25184 34838 25236 34890
rect 30320 34838 30372 34890
rect 30384 34838 30436 34890
rect 30448 34838 30500 34890
rect 30512 34838 30564 34890
rect 35648 34838 35700 34890
rect 35712 34838 35764 34890
rect 35776 34838 35828 34890
rect 35840 34838 35892 34890
rect 40976 34838 41028 34890
rect 41040 34838 41092 34890
rect 41104 34838 41156 34890
rect 41168 34838 41220 34890
rect 46304 34838 46356 34890
rect 46368 34838 46420 34890
rect 46432 34838 46484 34890
rect 46496 34838 46548 34890
rect 51632 34838 51684 34890
rect 51696 34838 51748 34890
rect 51760 34838 51812 34890
rect 51824 34838 51876 34890
rect 56960 34838 57012 34890
rect 57024 34838 57076 34890
rect 57088 34838 57140 34890
rect 57152 34838 57204 34890
rect 62288 34838 62340 34890
rect 62352 34838 62404 34890
rect 62416 34838 62468 34890
rect 62480 34838 62532 34890
rect 67616 34838 67668 34890
rect 67680 34838 67732 34890
rect 67744 34838 67796 34890
rect 67808 34838 67860 34890
rect 72944 34838 72996 34890
rect 73008 34838 73060 34890
rect 73072 34838 73124 34890
rect 73136 34838 73188 34890
rect 78272 34838 78324 34890
rect 78336 34838 78388 34890
rect 78400 34838 78452 34890
rect 78464 34838 78516 34890
rect 83600 34838 83652 34890
rect 83664 34838 83716 34890
rect 83728 34838 83780 34890
rect 83792 34838 83844 34890
rect 88928 34838 88980 34890
rect 88992 34838 89044 34890
rect 89056 34838 89108 34890
rect 89120 34838 89172 34890
rect 4238 34736 4290 34788
rect 12794 34779 12846 34788
rect 12794 34745 12803 34779
rect 12803 34745 12837 34779
rect 12837 34745 12846 34779
rect 12794 34736 12846 34745
rect 16106 34736 16158 34788
rect 16842 34600 16894 34652
rect 2582 34575 2634 34584
rect 2582 34541 2591 34575
rect 2591 34541 2625 34575
rect 2625 34541 2634 34575
rect 2582 34532 2634 34541
rect 3226 34532 3278 34584
rect 9114 34532 9166 34584
rect 9482 34532 9534 34584
rect 12794 34532 12846 34584
rect 6630 34464 6682 34516
rect 3870 34439 3922 34448
rect 3870 34405 3879 34439
rect 3879 34405 3913 34439
rect 3913 34405 3922 34439
rect 3870 34396 3922 34405
rect 13070 34439 13122 34448
rect 13070 34405 13079 34439
rect 13079 34405 13113 34439
rect 13113 34405 13122 34439
rect 13070 34396 13122 34405
rect 16842 34396 16894 34448
rect 21166 34736 21218 34788
rect 22822 34736 22874 34788
rect 30642 34736 30694 34788
rect 33126 34736 33178 34788
rect 33402 34736 33454 34788
rect 34598 34779 34650 34788
rect 34598 34745 34607 34779
rect 34607 34745 34641 34779
rect 34641 34745 34650 34779
rect 34598 34736 34650 34745
rect 35518 34736 35570 34788
rect 40118 34736 40170 34788
rect 40210 34736 40262 34788
rect 55298 34736 55350 34788
rect 55390 34736 55442 34788
rect 61002 34736 61054 34788
rect 63394 34736 63446 34788
rect 21258 34643 21310 34652
rect 21258 34609 21267 34643
rect 21267 34609 21301 34643
rect 21301 34609 21310 34643
rect 21258 34600 21310 34609
rect 20522 34575 20574 34584
rect 20522 34541 20531 34575
rect 20531 34541 20565 34575
rect 20565 34541 20574 34575
rect 20522 34532 20574 34541
rect 20614 34575 20666 34584
rect 20614 34541 20623 34575
rect 20623 34541 20657 34575
rect 20657 34541 20666 34575
rect 20614 34532 20666 34541
rect 23282 34532 23334 34584
rect 24938 34464 24990 34516
rect 17670 34396 17722 34448
rect 18406 34439 18458 34448
rect 18406 34405 18415 34439
rect 18415 34405 18449 34439
rect 18449 34405 18458 34439
rect 18406 34396 18458 34405
rect 20614 34396 20666 34448
rect 23006 34396 23058 34448
rect 25858 34600 25910 34652
rect 26226 34643 26278 34652
rect 26226 34609 26235 34643
rect 26235 34609 26269 34643
rect 26269 34609 26278 34643
rect 29814 34668 29866 34720
rect 29906 34711 29958 34720
rect 29906 34677 29915 34711
rect 29915 34677 29949 34711
rect 29949 34677 29958 34711
rect 29906 34668 29958 34677
rect 26226 34600 26278 34609
rect 25490 34575 25542 34584
rect 25490 34541 25499 34575
rect 25499 34541 25533 34575
rect 25533 34541 25542 34575
rect 25490 34532 25542 34541
rect 26870 34600 26922 34652
rect 39382 34668 39434 34720
rect 48214 34668 48266 34720
rect 40026 34643 40078 34652
rect 40026 34609 40035 34643
rect 40035 34609 40069 34643
rect 40069 34609 40078 34643
rect 40026 34600 40078 34609
rect 41314 34600 41366 34652
rect 47662 34643 47714 34652
rect 29814 34532 29866 34584
rect 34138 34575 34190 34584
rect 34138 34541 34147 34575
rect 34147 34541 34181 34575
rect 34181 34541 34190 34575
rect 34138 34532 34190 34541
rect 34598 34532 34650 34584
rect 35058 34575 35110 34584
rect 35058 34541 35067 34575
rect 35067 34541 35101 34575
rect 35101 34541 35110 34575
rect 35058 34532 35110 34541
rect 40118 34575 40170 34584
rect 40118 34541 40127 34575
rect 40127 34541 40161 34575
rect 40161 34541 40170 34575
rect 40118 34532 40170 34541
rect 40578 34575 40630 34584
rect 40578 34541 40587 34575
rect 40587 34541 40621 34575
rect 40621 34541 40630 34575
rect 40578 34532 40630 34541
rect 40670 34575 40722 34584
rect 40670 34541 40679 34575
rect 40679 34541 40713 34575
rect 40713 34541 40722 34575
rect 40670 34532 40722 34541
rect 46098 34532 46150 34584
rect 46834 34532 46886 34584
rect 40302 34464 40354 34516
rect 44442 34464 44494 34516
rect 25766 34439 25818 34448
rect 25766 34405 25775 34439
rect 25775 34405 25809 34439
rect 25809 34405 25818 34439
rect 25766 34396 25818 34405
rect 25858 34396 25910 34448
rect 26778 34396 26830 34448
rect 27054 34439 27106 34448
rect 27054 34405 27063 34439
rect 27063 34405 27097 34439
rect 27097 34405 27106 34439
rect 27054 34396 27106 34405
rect 31838 34396 31890 34448
rect 32482 34396 32534 34448
rect 38186 34396 38238 34448
rect 40210 34396 40262 34448
rect 43522 34396 43574 34448
rect 46926 34396 46978 34448
rect 47662 34609 47671 34643
rect 47671 34609 47705 34643
rect 47705 34609 47714 34643
rect 47662 34600 47714 34609
rect 51894 34668 51946 34720
rect 52814 34668 52866 34720
rect 53182 34668 53234 34720
rect 47570 34464 47622 34516
rect 53274 34600 53326 34652
rect 54010 34668 54062 34720
rect 64774 34668 64826 34720
rect 67994 34711 68046 34720
rect 67994 34677 68003 34711
rect 68003 34677 68037 34711
rect 68037 34677 68046 34711
rect 67994 34668 68046 34677
rect 69282 34711 69334 34720
rect 69282 34677 69291 34711
rect 69291 34677 69325 34711
rect 69325 34677 69334 34711
rect 69282 34668 69334 34677
rect 69466 34736 69518 34788
rect 84278 34736 84330 34788
rect 88786 34736 88838 34788
rect 90718 34736 90770 34788
rect 74158 34668 74210 34720
rect 57782 34600 57834 34652
rect 59438 34643 59490 34652
rect 59438 34609 59447 34643
rect 59447 34609 59481 34643
rect 59481 34609 59490 34643
rect 59438 34600 59490 34609
rect 59990 34600 60042 34652
rect 62106 34600 62158 34652
rect 54010 34575 54062 34584
rect 54010 34541 54019 34575
rect 54019 34541 54053 34575
rect 54053 34541 54062 34575
rect 54010 34532 54062 34541
rect 51526 34439 51578 34448
rect 51526 34405 51535 34439
rect 51535 34405 51569 34439
rect 51569 34405 51578 34439
rect 51526 34396 51578 34405
rect 54286 34464 54338 34516
rect 54194 34396 54246 34448
rect 54654 34396 54706 34448
rect 57414 34532 57466 34584
rect 58334 34575 58386 34584
rect 58334 34541 58343 34575
rect 58343 34541 58377 34575
rect 58377 34541 58386 34575
rect 58334 34532 58386 34541
rect 58426 34575 58478 34584
rect 58426 34541 58435 34575
rect 58435 34541 58469 34575
rect 58469 34541 58478 34575
rect 58886 34575 58938 34584
rect 58426 34532 58478 34541
rect 58886 34541 58895 34575
rect 58895 34541 58929 34575
rect 58929 34541 58938 34575
rect 58886 34532 58938 34541
rect 60174 34532 60226 34584
rect 62566 34575 62618 34584
rect 62566 34541 62575 34575
rect 62575 34541 62609 34575
rect 62609 34541 62618 34575
rect 62566 34532 62618 34541
rect 63210 34575 63262 34584
rect 63210 34541 63215 34575
rect 63215 34541 63249 34575
rect 63249 34541 63262 34575
rect 63210 34532 63262 34541
rect 67810 34575 67862 34584
rect 67810 34541 67819 34575
rect 67819 34541 67853 34575
rect 67853 34541 67862 34575
rect 67810 34532 67862 34541
rect 68178 34575 68230 34584
rect 68178 34541 68187 34575
rect 68187 34541 68221 34575
rect 68221 34541 68230 34575
rect 68178 34532 68230 34541
rect 68270 34532 68322 34584
rect 73974 34600 74026 34652
rect 74526 34643 74578 34652
rect 68914 34575 68966 34584
rect 68914 34541 68923 34575
rect 68923 34541 68957 34575
rect 68957 34541 68966 34575
rect 68914 34532 68966 34541
rect 69650 34532 69702 34584
rect 74526 34609 74535 34643
rect 74535 34609 74569 34643
rect 74569 34609 74578 34643
rect 74526 34600 74578 34609
rect 80874 34668 80926 34720
rect 81150 34711 81202 34720
rect 81150 34677 81159 34711
rect 81159 34677 81193 34711
rect 81193 34677 81202 34711
rect 81150 34668 81202 34677
rect 81334 34600 81386 34652
rect 80230 34575 80282 34584
rect 80230 34541 80239 34575
rect 80239 34541 80273 34575
rect 80273 34541 80282 34575
rect 80782 34575 80834 34584
rect 80230 34532 80282 34541
rect 80782 34541 80791 34575
rect 80791 34541 80825 34575
rect 80825 34541 80834 34575
rect 80782 34532 80834 34541
rect 81242 34532 81294 34584
rect 82530 34532 82582 34584
rect 62566 34396 62618 34448
rect 63210 34396 63262 34448
rect 63486 34396 63538 34448
rect 63670 34396 63722 34448
rect 69466 34396 69518 34448
rect 69650 34439 69702 34448
rect 69650 34405 69659 34439
rect 69659 34405 69693 34439
rect 69693 34405 69702 34439
rect 69650 34396 69702 34405
rect 74342 34464 74394 34516
rect 84646 34532 84698 34584
rect 86578 34575 86630 34584
rect 75354 34396 75406 34448
rect 80782 34396 80834 34448
rect 81334 34396 81386 34448
rect 82346 34396 82398 34448
rect 82714 34396 82766 34448
rect 86578 34541 86587 34575
rect 86587 34541 86621 34575
rect 86621 34541 86630 34575
rect 86578 34532 86630 34541
rect 87774 34532 87826 34584
rect 91086 34575 91138 34584
rect 91086 34541 91095 34575
rect 91095 34541 91129 34575
rect 91129 34541 91138 34575
rect 91086 34532 91138 34541
rect 87958 34464 88010 34516
rect 86026 34396 86078 34448
rect 86578 34396 86630 34448
rect 6344 34294 6396 34346
rect 6408 34294 6460 34346
rect 6472 34294 6524 34346
rect 6536 34294 6588 34346
rect 11672 34294 11724 34346
rect 11736 34294 11788 34346
rect 11800 34294 11852 34346
rect 11864 34294 11916 34346
rect 17000 34294 17052 34346
rect 17064 34294 17116 34346
rect 17128 34294 17180 34346
rect 17192 34294 17244 34346
rect 22328 34294 22380 34346
rect 22392 34294 22444 34346
rect 22456 34294 22508 34346
rect 22520 34294 22572 34346
rect 27656 34294 27708 34346
rect 27720 34294 27772 34346
rect 27784 34294 27836 34346
rect 27848 34294 27900 34346
rect 32984 34294 33036 34346
rect 33048 34294 33100 34346
rect 33112 34294 33164 34346
rect 33176 34294 33228 34346
rect 38312 34294 38364 34346
rect 38376 34294 38428 34346
rect 38440 34294 38492 34346
rect 38504 34294 38556 34346
rect 43640 34294 43692 34346
rect 43704 34294 43756 34346
rect 43768 34294 43820 34346
rect 43832 34294 43884 34346
rect 48968 34294 49020 34346
rect 49032 34294 49084 34346
rect 49096 34294 49148 34346
rect 49160 34294 49212 34346
rect 54296 34294 54348 34346
rect 54360 34294 54412 34346
rect 54424 34294 54476 34346
rect 54488 34294 54540 34346
rect 59624 34294 59676 34346
rect 59688 34294 59740 34346
rect 59752 34294 59804 34346
rect 59816 34294 59868 34346
rect 64952 34294 65004 34346
rect 65016 34294 65068 34346
rect 65080 34294 65132 34346
rect 65144 34294 65196 34346
rect 70280 34294 70332 34346
rect 70344 34294 70396 34346
rect 70408 34294 70460 34346
rect 70472 34294 70524 34346
rect 75608 34294 75660 34346
rect 75672 34294 75724 34346
rect 75736 34294 75788 34346
rect 75800 34294 75852 34346
rect 80936 34294 80988 34346
rect 81000 34294 81052 34346
rect 81064 34294 81116 34346
rect 81128 34294 81180 34346
rect 86264 34294 86316 34346
rect 86328 34294 86380 34346
rect 86392 34294 86444 34346
rect 86456 34294 86508 34346
rect 91592 34294 91644 34346
rect 91656 34294 91708 34346
rect 91720 34294 91772 34346
rect 91784 34294 91836 34346
rect 10218 34192 10270 34244
rect 15738 34192 15790 34244
rect 6630 34124 6682 34176
rect 3870 34056 3922 34108
rect 9114 34056 9166 34108
rect 16014 34192 16066 34244
rect 17578 34192 17630 34244
rect 26870 34192 26922 34244
rect 27054 34192 27106 34244
rect 51526 34192 51578 34244
rect 52814 34235 52866 34244
rect 52814 34201 52823 34235
rect 52823 34201 52857 34235
rect 52857 34201 52866 34235
rect 52814 34192 52866 34201
rect 54194 34192 54246 34244
rect 60450 34192 60502 34244
rect 61002 34192 61054 34244
rect 63762 34192 63814 34244
rect 64774 34192 64826 34244
rect 4698 33988 4750 34040
rect 7090 33920 7142 33972
rect 16014 34056 16066 34108
rect 17762 34124 17814 34176
rect 18406 34124 18458 34176
rect 23006 34124 23058 34176
rect 10402 33920 10454 33972
rect 17578 34056 17630 34108
rect 20154 34056 20206 34108
rect 17486 33988 17538 34040
rect 22730 34056 22782 34108
rect 23374 34056 23426 34108
rect 25490 34056 25542 34108
rect 25950 34099 26002 34108
rect 25950 34065 25959 34099
rect 25959 34065 25993 34099
rect 25993 34065 26002 34099
rect 25950 34056 26002 34065
rect 28894 34099 28946 34108
rect 28894 34065 28903 34099
rect 28903 34065 28937 34099
rect 28937 34065 28946 34099
rect 28894 34056 28946 34065
rect 29814 34056 29866 34108
rect 32482 34056 32534 34108
rect 34046 34099 34098 34108
rect 21718 33920 21770 33972
rect 24938 33920 24990 33972
rect 26870 33963 26922 33972
rect 9390 33895 9442 33904
rect 9390 33861 9399 33895
rect 9399 33861 9433 33895
rect 9433 33861 9442 33895
rect 9390 33852 9442 33861
rect 17670 33852 17722 33904
rect 25398 33852 25450 33904
rect 26870 33929 26879 33963
rect 26879 33929 26913 33963
rect 26913 33929 26922 33963
rect 26870 33920 26922 33929
rect 29078 33963 29130 33972
rect 29078 33929 29087 33963
rect 29087 33929 29121 33963
rect 29121 33929 29130 33963
rect 29078 33920 29130 33929
rect 26226 33895 26278 33904
rect 26226 33861 26235 33895
rect 26235 33861 26269 33895
rect 26269 33861 26278 33895
rect 26226 33852 26278 33861
rect 31470 33852 31522 33904
rect 34046 34065 34055 34099
rect 34055 34065 34089 34099
rect 34089 34065 34098 34099
rect 34046 34056 34098 34065
rect 35518 34056 35570 34108
rect 40118 34124 40170 34176
rect 40670 34124 40722 34176
rect 45086 34167 45138 34176
rect 45086 34133 45095 34167
rect 45095 34133 45129 34167
rect 45129 34133 45138 34167
rect 45086 34124 45138 34133
rect 46650 34124 46702 34176
rect 39934 34099 39986 34108
rect 39934 34065 39943 34099
rect 39943 34065 39977 34099
rect 39977 34065 39986 34099
rect 39934 34056 39986 34065
rect 40302 34099 40354 34108
rect 40302 34065 40311 34099
rect 40311 34065 40345 34099
rect 40345 34065 40354 34099
rect 40302 34056 40354 34065
rect 40394 34099 40446 34108
rect 40394 34065 40403 34099
rect 40403 34065 40437 34099
rect 40437 34065 40446 34099
rect 40394 34056 40446 34065
rect 33954 33920 34006 33972
rect 34414 33963 34466 33972
rect 34414 33929 34423 33963
rect 34423 33929 34457 33963
rect 34457 33929 34466 33963
rect 34414 33920 34466 33929
rect 45178 34056 45230 34108
rect 46558 34056 46610 34108
rect 47662 34124 47714 34176
rect 47018 34056 47070 34108
rect 52446 34056 52498 34108
rect 63578 34167 63630 34176
rect 63578 34133 63587 34167
rect 63587 34133 63621 34167
rect 63621 34133 63630 34167
rect 63578 34124 63630 34133
rect 64130 34124 64182 34176
rect 52814 34056 52866 34108
rect 54654 33988 54706 34040
rect 55390 34056 55442 34108
rect 63670 34056 63722 34108
rect 63854 34056 63906 34108
rect 59806 33988 59858 34040
rect 35058 33895 35110 33904
rect 35058 33861 35067 33895
rect 35067 33861 35101 33895
rect 35101 33861 35110 33895
rect 35058 33852 35110 33861
rect 43338 33852 43390 33904
rect 43522 33852 43574 33904
rect 47202 33852 47254 33904
rect 59438 33920 59490 33972
rect 60082 33920 60134 33972
rect 65602 33988 65654 34040
rect 67626 34056 67678 34108
rect 68270 34124 68322 34176
rect 69650 34124 69702 34176
rect 73698 34124 73750 34176
rect 68638 34099 68690 34108
rect 68638 34065 68647 34099
rect 68647 34065 68681 34099
rect 68681 34065 68690 34099
rect 68638 34056 68690 34065
rect 73882 34056 73934 34108
rect 75446 34056 75498 34108
rect 76090 34056 76142 34108
rect 77930 34099 77982 34108
rect 77930 34065 77939 34099
rect 77939 34065 77973 34099
rect 77973 34065 77982 34099
rect 77930 34056 77982 34065
rect 78574 34056 78626 34108
rect 79954 34124 80006 34176
rect 80414 34056 80466 34108
rect 73698 33988 73750 34040
rect 74066 34031 74118 34040
rect 74066 33997 74075 34031
rect 74075 33997 74109 34031
rect 74109 33997 74118 34031
rect 74066 33988 74118 33997
rect 80690 34192 80742 34244
rect 81242 34124 81294 34176
rect 90258 34124 90310 34176
rect 89798 34056 89850 34108
rect 88418 33988 88470 34040
rect 90258 34031 90310 34040
rect 90258 33997 90267 34031
rect 90267 33997 90301 34031
rect 90301 33997 90310 34031
rect 90258 33988 90310 33997
rect 64130 33920 64182 33972
rect 66062 33920 66114 33972
rect 67902 33920 67954 33972
rect 68638 33920 68690 33972
rect 68730 33920 68782 33972
rect 52814 33852 52866 33904
rect 52906 33852 52958 33904
rect 53458 33852 53510 33904
rect 54654 33895 54706 33904
rect 54654 33861 54663 33895
rect 54663 33861 54697 33895
rect 54697 33861 54706 33895
rect 54654 33852 54706 33861
rect 59530 33852 59582 33904
rect 59990 33852 60042 33904
rect 91362 33963 91414 33972
rect 91362 33929 91371 33963
rect 91371 33929 91405 33963
rect 91405 33929 91414 33963
rect 91362 33920 91414 33929
rect 73882 33852 73934 33904
rect 74342 33852 74394 33904
rect 78942 33852 78994 33904
rect 3680 33750 3732 33802
rect 3744 33750 3796 33802
rect 3808 33750 3860 33802
rect 3872 33750 3924 33802
rect 9008 33750 9060 33802
rect 9072 33750 9124 33802
rect 9136 33750 9188 33802
rect 9200 33750 9252 33802
rect 14336 33750 14388 33802
rect 14400 33750 14452 33802
rect 14464 33750 14516 33802
rect 14528 33750 14580 33802
rect 19664 33750 19716 33802
rect 19728 33750 19780 33802
rect 19792 33750 19844 33802
rect 19856 33750 19908 33802
rect 24992 33750 25044 33802
rect 25056 33750 25108 33802
rect 25120 33750 25172 33802
rect 25184 33750 25236 33802
rect 30320 33750 30372 33802
rect 30384 33750 30436 33802
rect 30448 33750 30500 33802
rect 30512 33750 30564 33802
rect 35648 33750 35700 33802
rect 35712 33750 35764 33802
rect 35776 33750 35828 33802
rect 35840 33750 35892 33802
rect 40976 33750 41028 33802
rect 41040 33750 41092 33802
rect 41104 33750 41156 33802
rect 41168 33750 41220 33802
rect 46304 33750 46356 33802
rect 46368 33750 46420 33802
rect 46432 33750 46484 33802
rect 46496 33750 46548 33802
rect 51632 33750 51684 33802
rect 51696 33750 51748 33802
rect 51760 33750 51812 33802
rect 51824 33750 51876 33802
rect 56960 33750 57012 33802
rect 57024 33750 57076 33802
rect 57088 33750 57140 33802
rect 57152 33750 57204 33802
rect 62288 33750 62340 33802
rect 62352 33750 62404 33802
rect 62416 33750 62468 33802
rect 62480 33750 62532 33802
rect 67616 33750 67668 33802
rect 67680 33750 67732 33802
rect 67744 33750 67796 33802
rect 67808 33750 67860 33802
rect 72944 33750 72996 33802
rect 73008 33750 73060 33802
rect 73072 33750 73124 33802
rect 73136 33750 73188 33802
rect 78272 33750 78324 33802
rect 78336 33750 78388 33802
rect 78400 33750 78452 33802
rect 78464 33750 78516 33802
rect 83600 33750 83652 33802
rect 83664 33750 83716 33802
rect 83728 33750 83780 33802
rect 83792 33750 83844 33802
rect 88928 33750 88980 33802
rect 88992 33750 89044 33802
rect 89056 33750 89108 33802
rect 89120 33750 89172 33802
rect 2582 33648 2634 33700
rect 17578 33691 17630 33700
rect 17578 33657 17587 33691
rect 17587 33657 17621 33691
rect 17621 33657 17630 33691
rect 17578 33648 17630 33657
rect 23282 33691 23334 33700
rect 23282 33657 23291 33691
rect 23291 33657 23325 33691
rect 23325 33657 23334 33691
rect 23282 33648 23334 33657
rect 25398 33648 25450 33700
rect 28342 33648 28394 33700
rect 29722 33648 29774 33700
rect 30182 33648 30234 33700
rect 39290 33648 39342 33700
rect 39658 33648 39710 33700
rect 40670 33648 40722 33700
rect 46006 33648 46058 33700
rect 49318 33648 49370 33700
rect 9390 33512 9442 33564
rect 13070 33580 13122 33632
rect 3502 33444 3554 33496
rect 5158 33487 5210 33496
rect 3226 33376 3278 33428
rect 5158 33453 5167 33487
rect 5167 33453 5201 33487
rect 5201 33453 5210 33487
rect 5158 33444 5210 33453
rect 6630 33444 6682 33496
rect 7090 33444 7142 33496
rect 10034 33444 10086 33496
rect 12518 33487 12570 33496
rect 12518 33453 12527 33487
rect 12527 33453 12561 33487
rect 12561 33453 12570 33487
rect 12518 33444 12570 33453
rect 6170 33376 6222 33428
rect 10402 33419 10454 33428
rect 10402 33385 10411 33419
rect 10411 33385 10445 33419
rect 10445 33385 10454 33419
rect 10402 33376 10454 33385
rect 12426 33376 12478 33428
rect 4974 33308 5026 33360
rect 11506 33308 11558 33360
rect 24294 33555 24346 33564
rect 24294 33521 24303 33555
rect 24303 33521 24337 33555
rect 24337 33521 24346 33555
rect 24294 33512 24346 33521
rect 13898 33487 13950 33496
rect 13898 33453 13907 33487
rect 13907 33453 13941 33487
rect 13941 33453 13950 33487
rect 13898 33444 13950 33453
rect 17302 33444 17354 33496
rect 18774 33487 18826 33496
rect 18774 33453 18783 33487
rect 18783 33453 18817 33487
rect 18817 33453 18826 33487
rect 18774 33444 18826 33453
rect 20798 33444 20850 33496
rect 23374 33444 23426 33496
rect 24018 33444 24070 33496
rect 26134 33444 26186 33496
rect 30366 33555 30418 33564
rect 30366 33521 30375 33555
rect 30375 33521 30409 33555
rect 30409 33521 30418 33555
rect 30366 33512 30418 33521
rect 33954 33512 34006 33564
rect 35058 33512 35110 33564
rect 35242 33512 35294 33564
rect 44442 33580 44494 33632
rect 53642 33580 53694 33632
rect 28894 33444 28946 33496
rect 30182 33444 30234 33496
rect 31470 33487 31522 33496
rect 31470 33453 31479 33487
rect 31479 33453 31513 33487
rect 31513 33453 31522 33487
rect 31470 33444 31522 33453
rect 31838 33444 31890 33496
rect 32114 33444 32166 33496
rect 32574 33444 32626 33496
rect 35426 33487 35478 33496
rect 35426 33453 35435 33487
rect 35435 33453 35469 33487
rect 35469 33453 35478 33487
rect 35426 33444 35478 33453
rect 35518 33487 35570 33496
rect 35518 33453 35527 33487
rect 35527 33453 35561 33487
rect 35561 33453 35570 33487
rect 52538 33512 52590 33564
rect 54654 33648 54706 33700
rect 58886 33648 58938 33700
rect 59990 33648 60042 33700
rect 60082 33648 60134 33700
rect 60266 33691 60318 33700
rect 60266 33657 60275 33691
rect 60275 33657 60309 33691
rect 60309 33657 60318 33691
rect 60450 33691 60502 33700
rect 60266 33648 60318 33657
rect 60450 33657 60459 33691
rect 60459 33657 60493 33691
rect 60493 33657 60502 33691
rect 60450 33648 60502 33657
rect 63486 33691 63538 33700
rect 63486 33657 63495 33691
rect 63495 33657 63529 33691
rect 63529 33657 63538 33691
rect 63486 33648 63538 33657
rect 64130 33691 64182 33700
rect 54010 33580 54062 33632
rect 62658 33580 62710 33632
rect 64130 33657 64139 33691
rect 64139 33657 64173 33691
rect 64173 33657 64182 33691
rect 64130 33648 64182 33657
rect 63762 33580 63814 33632
rect 65970 33648 66022 33700
rect 66062 33580 66114 33632
rect 73606 33648 73658 33700
rect 81518 33648 81570 33700
rect 85290 33648 85342 33700
rect 85658 33691 85710 33700
rect 85658 33657 85667 33691
rect 85667 33657 85701 33691
rect 85701 33657 85710 33691
rect 85658 33648 85710 33657
rect 35518 33444 35570 33453
rect 18682 33376 18734 33428
rect 20798 33351 20850 33360
rect 20798 33317 20807 33351
rect 20807 33317 20841 33351
rect 20841 33317 20850 33351
rect 20798 33308 20850 33317
rect 21626 33308 21678 33360
rect 25490 33308 25542 33360
rect 31838 33308 31890 33360
rect 32574 33308 32626 33360
rect 39658 33376 39710 33428
rect 39934 33419 39986 33428
rect 39934 33385 39943 33419
rect 39943 33385 39977 33419
rect 39977 33385 39986 33419
rect 39934 33376 39986 33385
rect 40578 33487 40630 33496
rect 40578 33453 40587 33487
rect 40587 33453 40621 33487
rect 40621 33453 40630 33487
rect 40578 33444 40630 33453
rect 40670 33444 40722 33496
rect 43522 33444 43574 33496
rect 43982 33444 44034 33496
rect 46926 33419 46978 33428
rect 46926 33385 46935 33419
rect 46935 33385 46969 33419
rect 46969 33385 46978 33419
rect 46926 33376 46978 33385
rect 47110 33487 47162 33496
rect 47110 33453 47119 33487
rect 47119 33453 47153 33487
rect 47153 33453 47162 33487
rect 47110 33444 47162 33453
rect 48858 33444 48910 33496
rect 52262 33444 52314 33496
rect 47478 33419 47530 33428
rect 39566 33308 39618 33360
rect 43982 33351 44034 33360
rect 43982 33317 43991 33351
rect 43991 33317 44025 33351
rect 44025 33317 44034 33351
rect 43982 33308 44034 33317
rect 44718 33308 44770 33360
rect 46650 33308 46702 33360
rect 47018 33308 47070 33360
rect 47478 33385 47487 33419
rect 47487 33385 47521 33419
rect 47521 33385 47530 33419
rect 47478 33376 47530 33385
rect 49686 33376 49738 33428
rect 52906 33487 52958 33496
rect 52906 33453 52915 33487
rect 52915 33453 52949 33487
rect 52949 33453 52958 33487
rect 52906 33444 52958 33453
rect 53458 33487 53510 33496
rect 53458 33453 53467 33487
rect 53467 33453 53501 33487
rect 53501 33453 53510 33487
rect 53458 33444 53510 33453
rect 57874 33444 57926 33496
rect 58426 33487 58478 33496
rect 58426 33453 58435 33487
rect 58435 33453 58469 33487
rect 58469 33453 58478 33487
rect 58426 33444 58478 33453
rect 58518 33487 58570 33496
rect 58518 33453 58527 33487
rect 58527 33453 58561 33487
rect 58561 33453 58570 33487
rect 58518 33444 58570 33453
rect 62842 33512 62894 33564
rect 65970 33555 66022 33564
rect 59346 33444 59398 33496
rect 60910 33487 60962 33496
rect 59162 33376 59214 33428
rect 57598 33351 57650 33360
rect 57598 33317 57607 33351
rect 57607 33317 57641 33351
rect 57641 33317 57650 33351
rect 57598 33308 57650 33317
rect 57966 33308 58018 33360
rect 59438 33351 59490 33360
rect 59438 33317 59447 33351
rect 59447 33317 59481 33351
rect 59481 33317 59490 33351
rect 59438 33308 59490 33317
rect 60910 33453 60919 33487
rect 60919 33453 60953 33487
rect 60953 33453 60962 33487
rect 60910 33444 60962 33453
rect 63026 33444 63078 33496
rect 65970 33521 65979 33555
rect 65979 33521 66013 33555
rect 66013 33521 66022 33555
rect 65970 33512 66022 33521
rect 68730 33555 68782 33564
rect 68730 33521 68739 33555
rect 68739 33521 68773 33555
rect 68773 33521 68782 33555
rect 68730 33512 68782 33521
rect 63946 33487 63998 33496
rect 63946 33453 63955 33487
rect 63955 33453 63989 33487
rect 63989 33453 63998 33487
rect 63946 33444 63998 33453
rect 65510 33376 65562 33428
rect 68638 33487 68690 33496
rect 68638 33453 68647 33487
rect 68647 33453 68681 33487
rect 68681 33453 68690 33487
rect 68638 33444 68690 33453
rect 69006 33487 69058 33496
rect 69006 33453 69015 33487
rect 69015 33453 69049 33487
rect 69049 33453 69058 33487
rect 69006 33444 69058 33453
rect 69098 33376 69150 33428
rect 61922 33308 61974 33360
rect 65970 33308 66022 33360
rect 67534 33308 67586 33360
rect 68638 33308 68690 33360
rect 81702 33580 81754 33632
rect 73606 33555 73658 33564
rect 73606 33521 73615 33555
rect 73615 33521 73649 33555
rect 73649 33521 73658 33555
rect 73606 33512 73658 33521
rect 74158 33555 74210 33564
rect 74158 33521 74167 33555
rect 74167 33521 74201 33555
rect 74201 33521 74210 33555
rect 74158 33512 74210 33521
rect 78574 33512 78626 33564
rect 73882 33444 73934 33496
rect 74434 33444 74486 33496
rect 75354 33444 75406 33496
rect 79310 33444 79362 33496
rect 80414 33512 80466 33564
rect 79862 33487 79914 33496
rect 79862 33453 79871 33487
rect 79871 33453 79905 33487
rect 79905 33453 79914 33487
rect 79862 33444 79914 33453
rect 79954 33487 80006 33496
rect 79954 33453 79963 33487
rect 79963 33453 79997 33487
rect 79997 33453 80006 33487
rect 79954 33444 80006 33453
rect 80598 33444 80650 33496
rect 82346 33487 82398 33496
rect 82346 33453 82355 33487
rect 82355 33453 82389 33487
rect 82389 33453 82398 33487
rect 82346 33444 82398 33453
rect 86026 33487 86078 33496
rect 86026 33453 86035 33487
rect 86035 33453 86069 33487
rect 86069 33453 86078 33487
rect 86026 33444 86078 33453
rect 90626 33580 90678 33632
rect 90350 33512 90402 33564
rect 82254 33376 82306 33428
rect 82714 33419 82766 33428
rect 82714 33385 82723 33419
rect 82723 33385 82757 33419
rect 82757 33385 82766 33419
rect 82714 33376 82766 33385
rect 86670 33376 86722 33428
rect 89798 33444 89850 33496
rect 69926 33308 69978 33360
rect 72134 33308 72186 33360
rect 73882 33308 73934 33360
rect 84186 33308 84238 33360
rect 87590 33308 87642 33360
rect 6344 33206 6396 33258
rect 6408 33206 6460 33258
rect 6472 33206 6524 33258
rect 6536 33206 6588 33258
rect 11672 33206 11724 33258
rect 11736 33206 11788 33258
rect 11800 33206 11852 33258
rect 11864 33206 11916 33258
rect 17000 33206 17052 33258
rect 17064 33206 17116 33258
rect 17128 33206 17180 33258
rect 17192 33206 17244 33258
rect 22328 33206 22380 33258
rect 22392 33206 22444 33258
rect 22456 33206 22508 33258
rect 22520 33206 22572 33258
rect 27656 33206 27708 33258
rect 27720 33206 27772 33258
rect 27784 33206 27836 33258
rect 27848 33206 27900 33258
rect 32984 33206 33036 33258
rect 33048 33206 33100 33258
rect 33112 33206 33164 33258
rect 33176 33206 33228 33258
rect 38312 33206 38364 33258
rect 38376 33206 38428 33258
rect 38440 33206 38492 33258
rect 38504 33206 38556 33258
rect 43640 33206 43692 33258
rect 43704 33206 43756 33258
rect 43768 33206 43820 33258
rect 43832 33206 43884 33258
rect 48968 33206 49020 33258
rect 49032 33206 49084 33258
rect 49096 33206 49148 33258
rect 49160 33206 49212 33258
rect 54296 33206 54348 33258
rect 54360 33206 54412 33258
rect 54424 33206 54476 33258
rect 54488 33206 54540 33258
rect 59624 33206 59676 33258
rect 59688 33206 59740 33258
rect 59752 33206 59804 33258
rect 59816 33206 59868 33258
rect 64952 33206 65004 33258
rect 65016 33206 65068 33258
rect 65080 33206 65132 33258
rect 65144 33206 65196 33258
rect 70280 33206 70332 33258
rect 70344 33206 70396 33258
rect 70408 33206 70460 33258
rect 70472 33206 70524 33258
rect 75608 33206 75660 33258
rect 75672 33206 75724 33258
rect 75736 33206 75788 33258
rect 75800 33206 75852 33258
rect 80936 33206 80988 33258
rect 81000 33206 81052 33258
rect 81064 33206 81116 33258
rect 81128 33206 81180 33258
rect 86264 33206 86316 33258
rect 86328 33206 86380 33258
rect 86392 33206 86444 33258
rect 86456 33206 86508 33258
rect 91592 33206 91644 33258
rect 91656 33206 91708 33258
rect 91720 33206 91772 33258
rect 91784 33206 91836 33258
rect 7090 33104 7142 33156
rect 4698 33011 4750 33020
rect 4698 32977 4707 33011
rect 4707 32977 4741 33011
rect 4741 32977 4750 33011
rect 4698 32968 4750 32977
rect 4974 33011 5026 33020
rect 4974 32977 4983 33011
rect 4983 32977 5017 33011
rect 5017 32977 5026 33011
rect 4974 32968 5026 32977
rect 10034 33011 10086 33020
rect 10034 32977 10043 33011
rect 10043 32977 10077 33011
rect 10077 32977 10086 33011
rect 10034 32968 10086 32977
rect 11322 32968 11374 33020
rect 12426 32968 12478 33020
rect 13162 32968 13214 33020
rect 15094 33104 15146 33156
rect 15830 33104 15882 33156
rect 18682 33104 18734 33156
rect 21626 33104 21678 33156
rect 18958 33036 19010 33088
rect 19326 33036 19378 33088
rect 17302 32943 17354 32952
rect 17302 32909 17311 32943
rect 17311 32909 17345 32943
rect 17345 32909 17354 32943
rect 17302 32900 17354 32909
rect 6262 32807 6314 32816
rect 6262 32773 6271 32807
rect 6271 32773 6305 32807
rect 6305 32773 6314 32807
rect 6262 32764 6314 32773
rect 10402 32764 10454 32816
rect 14174 32832 14226 32884
rect 18682 32968 18734 33020
rect 18866 32832 18918 32884
rect 24294 33104 24346 33156
rect 28802 33104 28854 33156
rect 28894 33104 28946 33156
rect 33402 33147 33454 33156
rect 25950 33079 26002 33088
rect 25950 33045 25959 33079
rect 25959 33045 25993 33079
rect 25993 33045 26002 33079
rect 25950 33036 26002 33045
rect 23374 32900 23426 32952
rect 25398 32832 25450 32884
rect 11230 32764 11282 32816
rect 13622 32807 13674 32816
rect 13622 32773 13631 32807
rect 13631 32773 13665 32807
rect 13665 32773 13674 32807
rect 13622 32764 13674 32773
rect 16106 32764 16158 32816
rect 21074 32807 21126 32816
rect 21074 32773 21083 32807
rect 21083 32773 21117 32807
rect 21117 32773 21126 32807
rect 21074 32764 21126 32773
rect 25766 32968 25818 33020
rect 26134 32900 26186 32952
rect 26778 32968 26830 33020
rect 26870 32943 26922 32952
rect 26870 32909 26879 32943
rect 26879 32909 26913 32943
rect 26913 32909 26922 32943
rect 26870 32900 26922 32909
rect 29170 32968 29222 33020
rect 33402 33113 33411 33147
rect 33411 33113 33445 33147
rect 33445 33113 33454 33147
rect 33402 33104 33454 33113
rect 35426 33147 35478 33156
rect 31838 33011 31890 33020
rect 31838 32977 31847 33011
rect 31847 32977 31881 33011
rect 31881 32977 31890 33011
rect 31838 32968 31890 32977
rect 35426 33113 35435 33147
rect 35435 33113 35469 33147
rect 35469 33113 35478 33147
rect 35426 33104 35478 33113
rect 39290 33147 39342 33156
rect 39290 33113 39299 33147
rect 39299 33113 39333 33147
rect 39333 33113 39342 33147
rect 39290 33104 39342 33113
rect 43982 33104 44034 33156
rect 34414 32968 34466 33020
rect 37818 32968 37870 33020
rect 39750 32900 39802 32952
rect 40026 32968 40078 33020
rect 41130 33011 41182 33020
rect 41130 32977 41139 33011
rect 41139 32977 41173 33011
rect 41173 32977 41182 33011
rect 44074 33036 44126 33088
rect 47478 33036 47530 33088
rect 49318 33104 49370 33156
rect 57598 33104 57650 33156
rect 58426 33104 58478 33156
rect 59346 33104 59398 33156
rect 60082 33104 60134 33156
rect 60910 33104 60962 33156
rect 65418 33104 65470 33156
rect 65510 33104 65562 33156
rect 65970 33104 66022 33156
rect 82898 33147 82950 33156
rect 82898 33113 82907 33147
rect 82907 33113 82941 33147
rect 82941 33113 82950 33147
rect 82898 33104 82950 33113
rect 41130 32968 41182 32977
rect 40670 32900 40722 32952
rect 40762 32900 40814 32952
rect 44442 32968 44494 33020
rect 44718 32968 44770 33020
rect 47202 32968 47254 33020
rect 61094 33036 61146 33088
rect 61278 33036 61330 33088
rect 77838 33036 77890 33088
rect 49686 33011 49738 33020
rect 44994 32943 45046 32952
rect 37818 32875 37870 32884
rect 37818 32841 37827 32875
rect 37827 32841 37861 32875
rect 37861 32841 37870 32875
rect 37818 32832 37870 32841
rect 25766 32764 25818 32816
rect 26778 32764 26830 32816
rect 27514 32807 27566 32816
rect 27514 32773 27523 32807
rect 27523 32773 27557 32807
rect 27557 32773 27566 32807
rect 27514 32764 27566 32773
rect 33034 32764 33086 32816
rect 37726 32764 37778 32816
rect 40854 32764 40906 32816
rect 41130 32832 41182 32884
rect 41774 32875 41826 32884
rect 41774 32841 41783 32875
rect 41783 32841 41817 32875
rect 41817 32841 41826 32875
rect 41774 32832 41826 32841
rect 44994 32909 45003 32943
rect 45003 32909 45037 32943
rect 45037 32909 45046 32943
rect 44994 32900 45046 32909
rect 47294 32900 47346 32952
rect 49686 32977 49695 33011
rect 49695 32977 49729 33011
rect 49729 32977 49738 33011
rect 49686 32968 49738 32977
rect 51434 32900 51486 32952
rect 42326 32832 42378 32884
rect 44902 32875 44954 32884
rect 44902 32841 44911 32875
rect 44911 32841 44945 32875
rect 44945 32841 44954 32875
rect 44902 32832 44954 32841
rect 44166 32764 44218 32816
rect 44442 32807 44494 32816
rect 44442 32773 44451 32807
rect 44451 32773 44485 32807
rect 44485 32773 44494 32807
rect 44442 32764 44494 32773
rect 44810 32764 44862 32816
rect 46742 32807 46794 32816
rect 46742 32773 46751 32807
rect 46751 32773 46785 32807
rect 46785 32773 46794 32807
rect 46742 32764 46794 32773
rect 46834 32764 46886 32816
rect 47570 32807 47622 32816
rect 47570 32773 47579 32807
rect 47579 32773 47613 32807
rect 47613 32773 47622 32807
rect 47570 32764 47622 32773
rect 47662 32764 47714 32816
rect 48582 32764 48634 32816
rect 50606 32832 50658 32884
rect 52906 32764 52958 32816
rect 54194 32832 54246 32884
rect 57414 32968 57466 33020
rect 57966 32968 58018 33020
rect 58058 33011 58110 33020
rect 58058 32977 58067 33011
rect 58067 32977 58101 33011
rect 58101 32977 58110 33011
rect 58242 33011 58294 33020
rect 58058 32968 58110 32977
rect 58242 32977 58251 33011
rect 58251 32977 58285 33011
rect 58285 32977 58294 33011
rect 58242 32968 58294 32977
rect 56586 32900 56638 32952
rect 57322 32943 57374 32952
rect 57322 32909 57331 32943
rect 57331 32909 57365 32943
rect 57365 32909 57374 32943
rect 57322 32900 57374 32909
rect 59438 32968 59490 33020
rect 60174 32968 60226 33020
rect 60358 33011 60410 33020
rect 60358 32977 60367 33011
rect 60367 32977 60401 33011
rect 60401 32977 60410 33011
rect 60358 32968 60410 32977
rect 60910 32968 60962 33020
rect 62750 32968 62802 33020
rect 62934 33011 62986 33020
rect 62934 32977 62943 33011
rect 62943 32977 62977 33011
rect 62977 32977 62986 33011
rect 62934 32968 62986 32977
rect 63210 32968 63262 33020
rect 59806 32832 59858 32884
rect 58242 32764 58294 32816
rect 58334 32764 58386 32816
rect 58794 32807 58846 32816
rect 58794 32773 58803 32807
rect 58803 32773 58837 32807
rect 58837 32773 58846 32807
rect 58794 32764 58846 32773
rect 59346 32764 59398 32816
rect 60358 32764 60410 32816
rect 61370 32807 61422 32816
rect 61370 32773 61379 32807
rect 61379 32773 61413 32807
rect 61413 32773 61422 32807
rect 61370 32764 61422 32773
rect 63854 32832 63906 32884
rect 65050 32968 65102 33020
rect 65786 32968 65838 33020
rect 66522 33011 66574 33020
rect 66522 32977 66531 33011
rect 66531 32977 66565 33011
rect 66565 32977 66574 33011
rect 66522 32968 66574 32977
rect 67074 33011 67126 33020
rect 67074 32977 67083 33011
rect 67083 32977 67117 33011
rect 67117 32977 67126 33011
rect 67074 32968 67126 32977
rect 65602 32943 65654 32952
rect 65602 32909 65611 32943
rect 65611 32909 65645 32943
rect 65645 32909 65654 32943
rect 66890 32943 66942 32952
rect 65602 32900 65654 32909
rect 66890 32909 66899 32943
rect 66899 32909 66933 32943
rect 66933 32909 66942 32943
rect 66890 32900 66942 32909
rect 64130 32832 64182 32884
rect 64682 32875 64734 32884
rect 64682 32841 64691 32875
rect 64691 32841 64725 32875
rect 64725 32841 64734 32875
rect 64682 32832 64734 32841
rect 65050 32875 65102 32884
rect 65050 32841 65059 32875
rect 65059 32841 65093 32875
rect 65093 32841 65102 32875
rect 65050 32832 65102 32841
rect 67442 32968 67494 33020
rect 68546 32968 68598 33020
rect 69098 33011 69150 33020
rect 69098 32977 69107 33011
rect 69107 32977 69141 33011
rect 69141 32977 69150 33011
rect 69098 32968 69150 32977
rect 74434 33011 74486 33020
rect 74434 32977 74443 33011
rect 74443 32977 74477 33011
rect 74477 32977 74486 33011
rect 74434 32968 74486 32977
rect 74710 32968 74762 33020
rect 76826 32968 76878 33020
rect 77930 33011 77982 33020
rect 77930 32977 77939 33011
rect 77939 32977 77973 33011
rect 77973 32977 77982 33011
rect 77930 32968 77982 32977
rect 78574 33036 78626 33088
rect 78206 32968 78258 33020
rect 82806 32968 82858 33020
rect 83266 33011 83318 33020
rect 83266 32977 83275 33011
rect 83275 32977 83309 33011
rect 83309 32977 83318 33011
rect 83266 32968 83318 32977
rect 83634 32968 83686 33020
rect 83910 32968 83962 33020
rect 75354 32943 75406 32952
rect 65234 32764 65286 32816
rect 65970 32764 66022 32816
rect 66706 32807 66758 32816
rect 66706 32773 66715 32807
rect 66715 32773 66749 32807
rect 66749 32773 66758 32807
rect 66706 32764 66758 32773
rect 68086 32807 68138 32816
rect 68086 32773 68095 32807
rect 68095 32773 68129 32807
rect 68129 32773 68138 32807
rect 68086 32764 68138 32773
rect 68546 32832 68598 32884
rect 69282 32832 69334 32884
rect 69374 32832 69426 32884
rect 71214 32832 71266 32884
rect 74342 32832 74394 32884
rect 68730 32764 68782 32816
rect 69742 32764 69794 32816
rect 75354 32909 75363 32943
rect 75363 32909 75397 32943
rect 75397 32909 75406 32943
rect 75354 32900 75406 32909
rect 74526 32832 74578 32884
rect 81518 32832 81570 32884
rect 83450 32832 83502 32884
rect 83634 32832 83686 32884
rect 87498 32968 87550 33020
rect 87958 33011 88010 33020
rect 87958 32977 87967 33011
rect 87967 32977 88001 33011
rect 88001 32977 88010 33011
rect 87958 32968 88010 32977
rect 87406 32900 87458 32952
rect 86118 32832 86170 32884
rect 75630 32807 75682 32816
rect 75630 32773 75639 32807
rect 75639 32773 75673 32807
rect 75673 32773 75682 32807
rect 75630 32764 75682 32773
rect 75906 32764 75958 32816
rect 76642 32764 76694 32816
rect 81426 32764 81478 32816
rect 83082 32764 83134 32816
rect 84094 32764 84146 32816
rect 84278 32807 84330 32816
rect 84278 32773 84287 32807
rect 84287 32773 84321 32807
rect 84321 32773 84330 32807
rect 84278 32764 84330 32773
rect 86670 32807 86722 32816
rect 86670 32773 86679 32807
rect 86679 32773 86713 32807
rect 86713 32773 86722 32807
rect 86670 32764 86722 32773
rect 87406 32807 87458 32816
rect 87406 32773 87415 32807
rect 87415 32773 87449 32807
rect 87449 32773 87458 32807
rect 87406 32764 87458 32773
rect 3680 32662 3732 32714
rect 3744 32662 3796 32714
rect 3808 32662 3860 32714
rect 3872 32662 3924 32714
rect 9008 32662 9060 32714
rect 9072 32662 9124 32714
rect 9136 32662 9188 32714
rect 9200 32662 9252 32714
rect 14336 32662 14388 32714
rect 14400 32662 14452 32714
rect 14464 32662 14516 32714
rect 14528 32662 14580 32714
rect 19664 32662 19716 32714
rect 19728 32662 19780 32714
rect 19792 32662 19844 32714
rect 19856 32662 19908 32714
rect 24992 32662 25044 32714
rect 25056 32662 25108 32714
rect 25120 32662 25172 32714
rect 25184 32662 25236 32714
rect 30320 32662 30372 32714
rect 30384 32662 30436 32714
rect 30448 32662 30500 32714
rect 30512 32662 30564 32714
rect 35648 32662 35700 32714
rect 35712 32662 35764 32714
rect 35776 32662 35828 32714
rect 35840 32662 35892 32714
rect 40976 32662 41028 32714
rect 41040 32662 41092 32714
rect 41104 32662 41156 32714
rect 41168 32662 41220 32714
rect 46304 32662 46356 32714
rect 46368 32662 46420 32714
rect 46432 32662 46484 32714
rect 46496 32662 46548 32714
rect 51632 32662 51684 32714
rect 51696 32662 51748 32714
rect 51760 32662 51812 32714
rect 51824 32662 51876 32714
rect 56960 32662 57012 32714
rect 57024 32662 57076 32714
rect 57088 32662 57140 32714
rect 57152 32662 57204 32714
rect 62288 32662 62340 32714
rect 62352 32662 62404 32714
rect 62416 32662 62468 32714
rect 62480 32662 62532 32714
rect 67616 32662 67668 32714
rect 67680 32662 67732 32714
rect 67744 32662 67796 32714
rect 67808 32662 67860 32714
rect 72944 32662 72996 32714
rect 73008 32662 73060 32714
rect 73072 32662 73124 32714
rect 73136 32662 73188 32714
rect 78272 32662 78324 32714
rect 78336 32662 78388 32714
rect 78400 32662 78452 32714
rect 78464 32662 78516 32714
rect 83600 32662 83652 32714
rect 83664 32662 83716 32714
rect 83728 32662 83780 32714
rect 83792 32662 83844 32714
rect 88928 32662 88980 32714
rect 88992 32662 89044 32714
rect 89056 32662 89108 32714
rect 89120 32662 89172 32714
rect 5158 32560 5210 32612
rect 6262 32560 6314 32612
rect 16106 32603 16158 32612
rect 4698 32492 4750 32544
rect 5066 32535 5118 32544
rect 5066 32501 5075 32535
rect 5075 32501 5109 32535
rect 5109 32501 5118 32535
rect 5066 32492 5118 32501
rect 7918 32492 7970 32544
rect 1662 32288 1714 32340
rect 2766 32399 2818 32408
rect 2766 32365 2775 32399
rect 2775 32365 2809 32399
rect 2809 32365 2818 32399
rect 2766 32356 2818 32365
rect 6630 32356 6682 32408
rect 6998 32399 7050 32408
rect 6998 32365 7007 32399
rect 7007 32365 7041 32399
rect 7041 32365 7050 32399
rect 6998 32356 7050 32365
rect 12886 32399 12938 32408
rect 12886 32365 12895 32399
rect 12895 32365 12929 32399
rect 12929 32365 12938 32399
rect 16106 32569 16115 32603
rect 16115 32569 16149 32603
rect 16149 32569 16158 32603
rect 16106 32560 16158 32569
rect 16474 32603 16526 32612
rect 16474 32569 16483 32603
rect 16483 32569 16517 32603
rect 16517 32569 16526 32603
rect 16474 32560 16526 32569
rect 18774 32560 18826 32612
rect 20430 32560 20482 32612
rect 26870 32560 26922 32612
rect 32574 32560 32626 32612
rect 35150 32560 35202 32612
rect 39934 32560 39986 32612
rect 40578 32560 40630 32612
rect 15554 32492 15606 32544
rect 12886 32356 12938 32365
rect 13346 32399 13398 32408
rect 13346 32365 13355 32399
rect 13355 32365 13389 32399
rect 13389 32365 13398 32399
rect 13346 32356 13398 32365
rect 14174 32399 14226 32408
rect 14174 32365 14183 32399
rect 14183 32365 14217 32399
rect 14217 32365 14226 32399
rect 14174 32356 14226 32365
rect 14266 32399 14318 32408
rect 14266 32365 14275 32399
rect 14275 32365 14309 32399
rect 14309 32365 14318 32399
rect 14266 32356 14318 32365
rect 16290 32356 16342 32408
rect 22086 32492 22138 32544
rect 28802 32492 28854 32544
rect 34874 32492 34926 32544
rect 35058 32492 35110 32544
rect 38094 32492 38146 32544
rect 40670 32492 40722 32544
rect 44166 32560 44218 32612
rect 60082 32560 60134 32612
rect 65786 32603 65838 32612
rect 65786 32569 65795 32603
rect 65795 32569 65829 32603
rect 65829 32569 65838 32603
rect 65786 32560 65838 32569
rect 21074 32467 21126 32476
rect 21074 32433 21083 32467
rect 21083 32433 21117 32467
rect 21117 32433 21126 32467
rect 21074 32424 21126 32433
rect 25490 32467 25542 32476
rect 25490 32433 25499 32467
rect 25499 32433 25533 32467
rect 25533 32433 25542 32467
rect 25490 32424 25542 32433
rect 17486 32399 17538 32408
rect 17486 32365 17495 32399
rect 17495 32365 17529 32399
rect 17529 32365 17538 32399
rect 17486 32356 17538 32365
rect 18222 32356 18274 32408
rect 21350 32356 21402 32408
rect 13622 32288 13674 32340
rect 16198 32288 16250 32340
rect 19142 32220 19194 32272
rect 23834 32288 23886 32340
rect 24846 32220 24898 32272
rect 33034 32399 33086 32408
rect 33034 32365 33043 32399
rect 33043 32365 33077 32399
rect 33077 32365 33086 32399
rect 33034 32356 33086 32365
rect 34690 32399 34742 32408
rect 34690 32365 34699 32399
rect 34699 32365 34733 32399
rect 34733 32365 34742 32399
rect 34690 32356 34742 32365
rect 35150 32356 35202 32408
rect 39290 32424 39342 32476
rect 39474 32356 39526 32408
rect 26962 32288 27014 32340
rect 27514 32288 27566 32340
rect 26318 32220 26370 32272
rect 34322 32220 34374 32272
rect 40026 32424 40078 32476
rect 44442 32492 44494 32544
rect 40394 32356 40446 32408
rect 40670 32356 40722 32408
rect 42326 32424 42378 32476
rect 48398 32492 48450 32544
rect 48582 32492 48634 32544
rect 50606 32492 50658 32544
rect 52262 32492 52314 32544
rect 53182 32492 53234 32544
rect 58426 32535 58478 32544
rect 58426 32501 58435 32535
rect 58435 32501 58469 32535
rect 58469 32501 58478 32535
rect 58426 32492 58478 32501
rect 41682 32399 41734 32408
rect 41682 32365 41691 32399
rect 41691 32365 41725 32399
rect 41725 32365 41734 32399
rect 41682 32356 41734 32365
rect 48030 32424 48082 32476
rect 48858 32467 48910 32476
rect 48858 32433 48867 32467
rect 48867 32433 48901 32467
rect 48901 32433 48910 32467
rect 48858 32424 48910 32433
rect 44074 32356 44126 32408
rect 46742 32356 46794 32408
rect 47018 32356 47070 32408
rect 47202 32399 47254 32408
rect 47202 32365 47211 32399
rect 47211 32365 47245 32399
rect 47245 32365 47254 32399
rect 47478 32399 47530 32408
rect 47202 32356 47254 32365
rect 47478 32365 47487 32399
rect 47487 32365 47521 32399
rect 47521 32365 47530 32399
rect 47478 32356 47530 32365
rect 43982 32288 44034 32340
rect 46466 32331 46518 32340
rect 46466 32297 46475 32331
rect 46475 32297 46509 32331
rect 46509 32297 46518 32331
rect 46466 32288 46518 32297
rect 47570 32220 47622 32272
rect 48398 32288 48450 32340
rect 47754 32263 47806 32272
rect 47754 32229 47763 32263
rect 47763 32229 47797 32263
rect 47797 32229 47806 32263
rect 47938 32263 47990 32272
rect 47754 32220 47806 32229
rect 47938 32229 47947 32263
rect 47947 32229 47981 32263
rect 47981 32229 47990 32263
rect 47938 32220 47990 32229
rect 48030 32220 48082 32272
rect 49686 32424 49738 32476
rect 57322 32424 57374 32476
rect 58334 32424 58386 32476
rect 59530 32492 59582 32544
rect 62750 32492 62802 32544
rect 51066 32356 51118 32408
rect 51526 32399 51578 32408
rect 51526 32365 51535 32399
rect 51535 32365 51569 32399
rect 51569 32365 51578 32399
rect 51526 32356 51578 32365
rect 51986 32356 52038 32408
rect 58058 32356 58110 32408
rect 58518 32356 58570 32408
rect 59346 32399 59398 32408
rect 59346 32365 59355 32399
rect 59355 32365 59389 32399
rect 59389 32365 59398 32399
rect 59346 32356 59398 32365
rect 60358 32399 60410 32408
rect 60358 32365 60367 32399
rect 60367 32365 60401 32399
rect 60401 32365 60410 32399
rect 60358 32356 60410 32365
rect 61370 32356 61422 32408
rect 63302 32399 63354 32408
rect 63302 32365 63311 32399
rect 63311 32365 63345 32399
rect 63345 32365 63354 32399
rect 63302 32356 63354 32365
rect 63394 32399 63446 32408
rect 63394 32365 63403 32399
rect 63403 32365 63437 32399
rect 63437 32365 63446 32399
rect 63854 32399 63906 32408
rect 63394 32356 63446 32365
rect 63854 32365 63863 32399
rect 63863 32365 63897 32399
rect 63897 32365 63906 32399
rect 63854 32356 63906 32365
rect 64498 32492 64550 32544
rect 74526 32560 74578 32612
rect 76274 32560 76326 32612
rect 83082 32560 83134 32612
rect 84278 32560 84330 32612
rect 64682 32467 64734 32476
rect 64682 32433 64691 32467
rect 64691 32433 64725 32467
rect 64725 32433 64734 32467
rect 65970 32492 66022 32544
rect 68546 32492 68598 32544
rect 71214 32535 71266 32544
rect 64682 32424 64734 32433
rect 71214 32501 71223 32535
rect 71223 32501 71257 32535
rect 71257 32501 71266 32535
rect 71214 32492 71266 32501
rect 81426 32492 81478 32544
rect 83542 32535 83594 32544
rect 83542 32501 83551 32535
rect 83551 32501 83585 32535
rect 83585 32501 83594 32535
rect 83542 32492 83594 32501
rect 86578 32492 86630 32544
rect 65234 32356 65286 32408
rect 65970 32356 66022 32408
rect 52630 32220 52682 32272
rect 58426 32220 58478 32272
rect 64590 32288 64642 32340
rect 65142 32288 65194 32340
rect 65418 32288 65470 32340
rect 68822 32356 68874 32408
rect 69374 32356 69426 32408
rect 69742 32399 69794 32408
rect 69742 32365 69751 32399
rect 69751 32365 69785 32399
rect 69785 32365 69794 32399
rect 69742 32356 69794 32365
rect 69834 32356 69886 32408
rect 74618 32424 74670 32476
rect 75906 32467 75958 32476
rect 75906 32433 75915 32467
rect 75915 32433 75949 32467
rect 75949 32433 75958 32467
rect 75906 32424 75958 32433
rect 76090 32467 76142 32476
rect 76090 32433 76099 32467
rect 76099 32433 76133 32467
rect 76133 32433 76142 32467
rect 76090 32424 76142 32433
rect 79862 32424 79914 32476
rect 82622 32424 82674 32476
rect 89062 32424 89114 32476
rect 71214 32356 71266 32408
rect 73698 32356 73750 32408
rect 73974 32356 74026 32408
rect 74158 32356 74210 32408
rect 75354 32356 75406 32408
rect 75630 32356 75682 32408
rect 76274 32399 76326 32408
rect 76274 32365 76283 32399
rect 76283 32365 76317 32399
rect 76317 32365 76326 32399
rect 76274 32356 76326 32365
rect 76642 32356 76694 32408
rect 76826 32399 76878 32408
rect 76826 32365 76835 32399
rect 76835 32365 76869 32399
rect 76869 32365 76878 32399
rect 76826 32356 76878 32365
rect 80414 32356 80466 32408
rect 66890 32288 66942 32340
rect 69190 32288 69242 32340
rect 62106 32220 62158 32272
rect 64682 32220 64734 32272
rect 65510 32220 65562 32272
rect 81334 32288 81386 32340
rect 82530 32356 82582 32408
rect 82714 32356 82766 32408
rect 83634 32356 83686 32408
rect 86118 32399 86170 32408
rect 86118 32365 86127 32399
rect 86127 32365 86161 32399
rect 86161 32365 86170 32399
rect 86118 32356 86170 32365
rect 82254 32288 82306 32340
rect 82990 32288 83042 32340
rect 83450 32288 83502 32340
rect 87406 32356 87458 32408
rect 87590 32356 87642 32408
rect 74986 32263 75038 32272
rect 74986 32229 74995 32263
rect 74995 32229 75029 32263
rect 75029 32229 75038 32263
rect 74986 32220 75038 32229
rect 76918 32220 76970 32272
rect 87498 32220 87550 32272
rect 6344 32118 6396 32170
rect 6408 32118 6460 32170
rect 6472 32118 6524 32170
rect 6536 32118 6588 32170
rect 11672 32118 11724 32170
rect 11736 32118 11788 32170
rect 11800 32118 11852 32170
rect 11864 32118 11916 32170
rect 17000 32118 17052 32170
rect 17064 32118 17116 32170
rect 17128 32118 17180 32170
rect 17192 32118 17244 32170
rect 22328 32118 22380 32170
rect 22392 32118 22444 32170
rect 22456 32118 22508 32170
rect 22520 32118 22572 32170
rect 27656 32118 27708 32170
rect 27720 32118 27772 32170
rect 27784 32118 27836 32170
rect 27848 32118 27900 32170
rect 32984 32118 33036 32170
rect 33048 32118 33100 32170
rect 33112 32118 33164 32170
rect 33176 32118 33228 32170
rect 38312 32118 38364 32170
rect 38376 32118 38428 32170
rect 38440 32118 38492 32170
rect 38504 32118 38556 32170
rect 43640 32118 43692 32170
rect 43704 32118 43756 32170
rect 43768 32118 43820 32170
rect 43832 32118 43884 32170
rect 48968 32118 49020 32170
rect 49032 32118 49084 32170
rect 49096 32118 49148 32170
rect 49160 32118 49212 32170
rect 54296 32118 54348 32170
rect 54360 32118 54412 32170
rect 54424 32118 54476 32170
rect 54488 32118 54540 32170
rect 59624 32118 59676 32170
rect 59688 32118 59740 32170
rect 59752 32118 59804 32170
rect 59816 32118 59868 32170
rect 64952 32118 65004 32170
rect 65016 32118 65068 32170
rect 65080 32118 65132 32170
rect 65144 32118 65196 32170
rect 70280 32118 70332 32170
rect 70344 32118 70396 32170
rect 70408 32118 70460 32170
rect 70472 32118 70524 32170
rect 75608 32118 75660 32170
rect 75672 32118 75724 32170
rect 75736 32118 75788 32170
rect 75800 32118 75852 32170
rect 80936 32118 80988 32170
rect 81000 32118 81052 32170
rect 81064 32118 81116 32170
rect 81128 32118 81180 32170
rect 86264 32118 86316 32170
rect 86328 32118 86380 32170
rect 86392 32118 86444 32170
rect 86456 32118 86508 32170
rect 91592 32118 91644 32170
rect 91656 32118 91708 32170
rect 91720 32118 91772 32170
rect 91784 32118 91836 32170
rect 5342 32016 5394 32068
rect 4974 31880 5026 31932
rect 6078 32016 6130 32068
rect 12886 32059 12938 32068
rect 6170 31948 6222 32000
rect 12518 31948 12570 32000
rect 12886 32025 12895 32059
rect 12895 32025 12929 32059
rect 12929 32025 12938 32059
rect 12886 32016 12938 32025
rect 26318 32016 26370 32068
rect 28618 32016 28670 32068
rect 28894 32016 28946 32068
rect 36070 32016 36122 32068
rect 40762 32016 40814 32068
rect 41682 32016 41734 32068
rect 46926 32016 46978 32068
rect 16014 31948 16066 32000
rect 18222 31991 18274 32000
rect 8470 31880 8522 31932
rect 11046 31880 11098 31932
rect 11230 31923 11282 31932
rect 11230 31889 11239 31923
rect 11239 31889 11273 31923
rect 11273 31889 11282 31923
rect 11230 31880 11282 31889
rect 11506 31880 11558 31932
rect 13070 31880 13122 31932
rect 14266 31880 14318 31932
rect 17854 31923 17906 31932
rect 17854 31889 17863 31923
rect 17863 31889 17897 31923
rect 17897 31889 17906 31923
rect 17854 31880 17906 31889
rect 18222 31957 18231 31991
rect 18231 31957 18265 31991
rect 18265 31957 18274 31991
rect 18222 31948 18274 31957
rect 18682 31948 18734 32000
rect 18958 31880 19010 31932
rect 19142 31923 19194 31932
rect 19142 31889 19151 31923
rect 19151 31889 19185 31923
rect 19185 31889 19194 31923
rect 19142 31880 19194 31889
rect 6998 31812 7050 31864
rect 3502 31744 3554 31796
rect 6078 31744 6130 31796
rect 6630 31744 6682 31796
rect 13530 31812 13582 31864
rect 17302 31812 17354 31864
rect 18130 31812 18182 31864
rect 21810 31923 21862 31932
rect 21810 31889 21819 31923
rect 21819 31889 21853 31923
rect 21853 31889 21862 31923
rect 21810 31880 21862 31889
rect 19418 31812 19470 31864
rect 21534 31812 21586 31864
rect 6170 31719 6222 31728
rect 6170 31685 6179 31719
rect 6179 31685 6213 31719
rect 6213 31685 6222 31719
rect 6170 31676 6222 31685
rect 8194 31676 8246 31728
rect 16106 31676 16158 31728
rect 17854 31744 17906 31796
rect 18682 31744 18734 31796
rect 20798 31744 20850 31796
rect 24570 31948 24622 32000
rect 35334 31948 35386 32000
rect 39474 31991 39526 32000
rect 39474 31957 39483 31991
rect 39483 31957 39517 31991
rect 39517 31957 39526 31991
rect 39474 31948 39526 31957
rect 23742 31880 23794 31932
rect 26870 31880 26922 31932
rect 28158 31880 28210 31932
rect 28710 31880 28762 31932
rect 28894 31923 28946 31932
rect 28894 31889 28903 31923
rect 28903 31889 28937 31923
rect 28937 31889 28946 31923
rect 28894 31880 28946 31889
rect 30090 31880 30142 31932
rect 39566 31923 39618 31932
rect 39566 31889 39575 31923
rect 39575 31889 39609 31923
rect 39609 31889 39618 31923
rect 39566 31880 39618 31889
rect 44810 31948 44862 32000
rect 47478 31991 47530 32000
rect 24478 31812 24530 31864
rect 25858 31812 25910 31864
rect 27146 31812 27198 31864
rect 28526 31812 28578 31864
rect 29170 31812 29222 31864
rect 40854 31880 40906 31932
rect 43522 31880 43574 31932
rect 44718 31923 44770 31932
rect 44718 31889 44727 31923
rect 44727 31889 44761 31923
rect 44761 31889 44770 31923
rect 44718 31880 44770 31889
rect 40762 31812 40814 31864
rect 47478 31957 47487 31991
rect 47487 31957 47521 31991
rect 47521 31957 47530 31991
rect 47478 31948 47530 31957
rect 45178 31923 45230 31932
rect 45178 31889 45187 31923
rect 45187 31889 45221 31923
rect 45221 31889 45230 31923
rect 45178 31880 45230 31889
rect 46098 31880 46150 31932
rect 46742 31923 46794 31932
rect 46742 31889 46751 31923
rect 46751 31889 46785 31923
rect 46785 31889 46794 31923
rect 46742 31880 46794 31889
rect 48398 31923 48450 31932
rect 48398 31889 48407 31923
rect 48407 31889 48441 31923
rect 48441 31889 48450 31923
rect 48398 31880 48450 31889
rect 50790 31880 50842 31932
rect 47662 31812 47714 31864
rect 32482 31744 32534 31796
rect 32574 31744 32626 31796
rect 19326 31719 19378 31728
rect 19326 31685 19335 31719
rect 19335 31685 19369 31719
rect 19369 31685 19378 31719
rect 19326 31676 19378 31685
rect 21534 31719 21586 31728
rect 21534 31685 21543 31719
rect 21543 31685 21577 31719
rect 21577 31685 21586 31719
rect 21534 31676 21586 31685
rect 21810 31676 21862 31728
rect 23742 31719 23794 31728
rect 23742 31685 23751 31719
rect 23751 31685 23785 31719
rect 23785 31685 23794 31719
rect 23742 31676 23794 31685
rect 24018 31719 24070 31728
rect 24018 31685 24027 31719
rect 24027 31685 24061 31719
rect 24061 31685 24070 31719
rect 24018 31676 24070 31685
rect 26134 31676 26186 31728
rect 27698 31719 27750 31728
rect 27698 31685 27707 31719
rect 27707 31685 27741 31719
rect 27741 31685 27750 31719
rect 27698 31676 27750 31685
rect 28158 31676 28210 31728
rect 37542 31676 37594 31728
rect 39750 31719 39802 31728
rect 39750 31685 39759 31719
rect 39759 31685 39793 31719
rect 39793 31685 39802 31719
rect 39750 31676 39802 31685
rect 46098 31719 46150 31728
rect 46098 31685 46107 31719
rect 46107 31685 46141 31719
rect 46141 31685 46150 31719
rect 46098 31676 46150 31685
rect 58610 31948 58662 32000
rect 58702 31948 58754 32000
rect 53642 31880 53694 31932
rect 54102 31880 54154 31932
rect 57598 31880 57650 31932
rect 51066 31812 51118 31864
rect 57690 31812 57742 31864
rect 60174 31880 60226 31932
rect 68362 31880 68414 31932
rect 53918 31744 53970 31796
rect 58150 31744 58202 31796
rect 58334 31812 58386 31864
rect 58518 31812 58570 31864
rect 63946 31855 63998 31864
rect 63946 31821 63955 31855
rect 63955 31821 63989 31855
rect 63989 31821 63998 31855
rect 63946 31812 63998 31821
rect 64130 31855 64182 31864
rect 64130 31821 64139 31855
rect 64139 31821 64173 31855
rect 64173 31821 64182 31855
rect 64130 31812 64182 31821
rect 64682 31812 64734 31864
rect 69006 31880 69058 31932
rect 69190 31923 69242 31932
rect 69190 31889 69199 31923
rect 69199 31889 69233 31923
rect 69233 31889 69242 31923
rect 69190 31880 69242 31889
rect 69374 31923 69426 31932
rect 69374 31889 69383 31923
rect 69383 31889 69417 31923
rect 69417 31889 69426 31923
rect 69374 31880 69426 31889
rect 69650 31948 69702 32000
rect 69834 31880 69886 31932
rect 70018 31923 70070 31932
rect 70018 31889 70027 31923
rect 70027 31889 70061 31923
rect 70061 31889 70070 31923
rect 70018 31880 70070 31889
rect 68822 31812 68874 31864
rect 50974 31676 51026 31728
rect 51986 31676 52038 31728
rect 52722 31676 52774 31728
rect 53826 31676 53878 31728
rect 54010 31676 54062 31728
rect 54194 31676 54246 31728
rect 58610 31676 58662 31728
rect 58794 31719 58846 31728
rect 58794 31685 58803 31719
rect 58803 31685 58837 31719
rect 58837 31685 58846 31719
rect 58794 31676 58846 31685
rect 58886 31676 58938 31728
rect 63210 31676 63262 31728
rect 63394 31719 63446 31728
rect 63394 31685 63403 31719
rect 63403 31685 63437 31719
rect 63437 31685 63446 31719
rect 63394 31676 63446 31685
rect 66890 31676 66942 31728
rect 68638 31744 68690 31796
rect 74710 31948 74762 32000
rect 71766 31923 71818 31932
rect 71766 31889 71775 31923
rect 71775 31889 71809 31923
rect 71809 31889 71818 31923
rect 71766 31880 71818 31889
rect 72134 31880 72186 31932
rect 74250 31923 74302 31932
rect 74250 31889 74259 31923
rect 74259 31889 74293 31923
rect 74293 31889 74302 31923
rect 74250 31880 74302 31889
rect 74986 31880 75038 31932
rect 76826 31948 76878 32000
rect 77470 31948 77522 32000
rect 77378 31923 77430 31932
rect 75446 31812 75498 31864
rect 77378 31889 77387 31923
rect 77387 31889 77421 31923
rect 77421 31889 77430 31923
rect 77378 31880 77430 31889
rect 78574 31948 78626 32000
rect 82806 31991 82858 32000
rect 82806 31957 82815 31991
rect 82815 31957 82849 31991
rect 82849 31957 82858 31991
rect 82806 31948 82858 31957
rect 83266 32016 83318 32068
rect 84830 32016 84882 32068
rect 87406 32016 87458 32068
rect 79310 31880 79362 31932
rect 79678 31880 79730 31932
rect 80414 31923 80466 31932
rect 80414 31889 80423 31923
rect 80423 31889 80457 31923
rect 80457 31889 80466 31923
rect 80414 31880 80466 31889
rect 83266 31923 83318 31932
rect 83266 31889 83275 31923
rect 83275 31889 83309 31923
rect 83309 31889 83318 31923
rect 83266 31880 83318 31889
rect 83634 31880 83686 31932
rect 83910 31880 83962 31932
rect 89062 32016 89114 32068
rect 90442 31880 90494 31932
rect 91362 31880 91414 31932
rect 91546 31923 91598 31932
rect 91546 31889 91555 31923
rect 91555 31889 91589 31923
rect 91589 31889 91598 31923
rect 91546 31880 91598 31889
rect 78850 31812 78902 31864
rect 83450 31812 83502 31864
rect 89706 31812 89758 31864
rect 68822 31676 68874 31728
rect 68914 31676 68966 31728
rect 84370 31744 84422 31796
rect 69834 31676 69886 31728
rect 73882 31676 73934 31728
rect 75354 31676 75406 31728
rect 77102 31676 77154 31728
rect 78666 31719 78718 31728
rect 78666 31685 78675 31719
rect 78675 31685 78709 31719
rect 78709 31685 78718 31719
rect 78666 31676 78718 31685
rect 80598 31719 80650 31728
rect 80598 31685 80607 31719
rect 80607 31685 80641 31719
rect 80641 31685 80650 31719
rect 80598 31676 80650 31685
rect 84278 31719 84330 31728
rect 84278 31685 84287 31719
rect 84287 31685 84321 31719
rect 84321 31685 84330 31719
rect 84278 31676 84330 31685
rect 88326 31676 88378 31728
rect 3680 31574 3732 31626
rect 3744 31574 3796 31626
rect 3808 31574 3860 31626
rect 3872 31574 3924 31626
rect 9008 31574 9060 31626
rect 9072 31574 9124 31626
rect 9136 31574 9188 31626
rect 9200 31574 9252 31626
rect 14336 31574 14388 31626
rect 14400 31574 14452 31626
rect 14464 31574 14516 31626
rect 14528 31574 14580 31626
rect 19664 31574 19716 31626
rect 19728 31574 19780 31626
rect 19792 31574 19844 31626
rect 19856 31574 19908 31626
rect 24992 31574 25044 31626
rect 25056 31574 25108 31626
rect 25120 31574 25172 31626
rect 25184 31574 25236 31626
rect 30320 31574 30372 31626
rect 30384 31574 30436 31626
rect 30448 31574 30500 31626
rect 30512 31574 30564 31626
rect 35648 31574 35700 31626
rect 35712 31574 35764 31626
rect 35776 31574 35828 31626
rect 35840 31574 35892 31626
rect 40976 31574 41028 31626
rect 41040 31574 41092 31626
rect 41104 31574 41156 31626
rect 41168 31574 41220 31626
rect 46304 31574 46356 31626
rect 46368 31574 46420 31626
rect 46432 31574 46484 31626
rect 46496 31574 46548 31626
rect 51632 31574 51684 31626
rect 51696 31574 51748 31626
rect 51760 31574 51812 31626
rect 51824 31574 51876 31626
rect 56960 31574 57012 31626
rect 57024 31574 57076 31626
rect 57088 31574 57140 31626
rect 57152 31574 57204 31626
rect 62288 31574 62340 31626
rect 62352 31574 62404 31626
rect 62416 31574 62468 31626
rect 62480 31574 62532 31626
rect 67616 31574 67668 31626
rect 67680 31574 67732 31626
rect 67744 31574 67796 31626
rect 67808 31574 67860 31626
rect 72944 31574 72996 31626
rect 73008 31574 73060 31626
rect 73072 31574 73124 31626
rect 73136 31574 73188 31626
rect 78272 31574 78324 31626
rect 78336 31574 78388 31626
rect 78400 31574 78452 31626
rect 78464 31574 78516 31626
rect 83600 31574 83652 31626
rect 83664 31574 83716 31626
rect 83728 31574 83780 31626
rect 83792 31574 83844 31626
rect 88928 31574 88980 31626
rect 88992 31574 89044 31626
rect 89056 31574 89108 31626
rect 89120 31574 89172 31626
rect 834 31472 886 31524
rect 2766 31472 2818 31524
rect 3502 31515 3554 31524
rect 3502 31481 3511 31515
rect 3511 31481 3545 31515
rect 3545 31481 3554 31515
rect 3502 31472 3554 31481
rect 5158 31472 5210 31524
rect 6446 31472 6498 31524
rect 11046 31472 11098 31524
rect 19142 31472 19194 31524
rect 22086 31515 22138 31524
rect 22086 31481 22095 31515
rect 22095 31481 22129 31515
rect 22129 31481 22138 31515
rect 22086 31472 22138 31481
rect 24570 31515 24622 31524
rect 24570 31481 24579 31515
rect 24579 31481 24613 31515
rect 24613 31481 24622 31515
rect 24570 31472 24622 31481
rect 1662 31379 1714 31388
rect 1662 31345 1671 31379
rect 1671 31345 1705 31379
rect 1705 31345 1714 31379
rect 1662 31336 1714 31345
rect 3502 31336 3554 31388
rect 6170 31404 6222 31456
rect 25858 31404 25910 31456
rect 6998 31336 7050 31388
rect 12334 31336 12386 31388
rect 4882 31200 4934 31252
rect 6446 31311 6498 31320
rect 6446 31277 6455 31311
rect 6455 31277 6489 31311
rect 6489 31277 6498 31311
rect 6446 31268 6498 31277
rect 6722 31268 6774 31320
rect 9298 31268 9350 31320
rect 12426 31311 12478 31320
rect 12426 31277 12435 31311
rect 12435 31277 12469 31311
rect 12469 31277 12478 31311
rect 12426 31268 12478 31277
rect 13346 31336 13398 31388
rect 6814 31200 6866 31252
rect 16658 31336 16710 31388
rect 18866 31336 18918 31388
rect 13070 31200 13122 31252
rect 17762 31268 17814 31320
rect 18958 31268 19010 31320
rect 26134 31336 26186 31388
rect 23282 31268 23334 31320
rect 23834 31311 23886 31320
rect 23834 31277 23843 31311
rect 23843 31277 23877 31311
rect 23877 31277 23886 31311
rect 23834 31268 23886 31277
rect 24110 31268 24162 31320
rect 24570 31268 24622 31320
rect 8102 31175 8154 31184
rect 8102 31141 8111 31175
rect 8111 31141 8145 31175
rect 8145 31141 8154 31175
rect 8102 31132 8154 31141
rect 12150 31132 12202 31184
rect 20706 31200 20758 31252
rect 32298 31472 32350 31524
rect 32482 31472 32534 31524
rect 39842 31472 39894 31524
rect 40026 31515 40078 31524
rect 40026 31481 40035 31515
rect 40035 31481 40069 31515
rect 40069 31481 40078 31515
rect 40026 31472 40078 31481
rect 47018 31515 47070 31524
rect 47018 31481 47027 31515
rect 47027 31481 47061 31515
rect 47061 31481 47070 31515
rect 47018 31472 47070 31481
rect 51526 31472 51578 31524
rect 26962 31404 27014 31456
rect 27698 31404 27750 31456
rect 28158 31404 28210 31456
rect 28434 31404 28486 31456
rect 30090 31447 30142 31456
rect 30090 31413 30099 31447
rect 30099 31413 30133 31447
rect 30133 31413 30142 31447
rect 30090 31404 30142 31413
rect 44442 31404 44494 31456
rect 44718 31404 44770 31456
rect 50882 31404 50934 31456
rect 54102 31472 54154 31524
rect 26778 31200 26830 31252
rect 28526 31336 28578 31388
rect 28986 31379 29038 31388
rect 28986 31345 28995 31379
rect 28995 31345 29029 31379
rect 29029 31345 29038 31379
rect 28986 31336 29038 31345
rect 18130 31132 18182 31184
rect 18682 31175 18734 31184
rect 18682 31141 18691 31175
rect 18691 31141 18725 31175
rect 18725 31141 18734 31175
rect 18682 31132 18734 31141
rect 18958 31175 19010 31184
rect 18958 31141 18967 31175
rect 18967 31141 19001 31175
rect 19001 31141 19010 31175
rect 18958 31132 19010 31141
rect 19878 31175 19930 31184
rect 19878 31141 19887 31175
rect 19887 31141 19921 31175
rect 19921 31141 19930 31175
rect 19878 31132 19930 31141
rect 22914 31175 22966 31184
rect 22914 31141 22923 31175
rect 22923 31141 22957 31175
rect 22957 31141 22966 31175
rect 22914 31132 22966 31141
rect 24110 31132 24162 31184
rect 31470 31268 31522 31320
rect 32206 31311 32258 31320
rect 32206 31277 32215 31311
rect 32215 31277 32249 31311
rect 32249 31277 32258 31311
rect 32206 31268 32258 31277
rect 32298 31311 32350 31320
rect 32298 31277 32307 31311
rect 32307 31277 32341 31311
rect 32341 31277 32350 31311
rect 32298 31268 32350 31277
rect 32666 31268 32718 31320
rect 33126 31200 33178 31252
rect 33310 31243 33362 31252
rect 33310 31209 33319 31243
rect 33319 31209 33353 31243
rect 33353 31209 33362 31243
rect 33310 31200 33362 31209
rect 28802 31132 28854 31184
rect 29262 31132 29314 31184
rect 32206 31132 32258 31184
rect 32666 31132 32718 31184
rect 33494 31132 33546 31184
rect 34414 31132 34466 31184
rect 35426 31132 35478 31184
rect 37358 31268 37410 31320
rect 39934 31311 39986 31320
rect 39934 31277 39943 31311
rect 39943 31277 39977 31311
rect 39977 31277 39986 31311
rect 39934 31268 39986 31277
rect 40854 31268 40906 31320
rect 46466 31336 46518 31388
rect 48858 31336 48910 31388
rect 63394 31472 63446 31524
rect 68638 31515 68690 31524
rect 68638 31481 68647 31515
rect 68647 31481 68681 31515
rect 68681 31481 68690 31515
rect 68638 31472 68690 31481
rect 54286 31404 54338 31456
rect 54654 31404 54706 31456
rect 62014 31404 62066 31456
rect 46926 31311 46978 31320
rect 46926 31277 46935 31311
rect 46935 31277 46969 31311
rect 46969 31277 46978 31311
rect 46926 31268 46978 31277
rect 51434 31311 51486 31320
rect 51434 31277 51443 31311
rect 51443 31277 51477 31311
rect 51477 31277 51486 31311
rect 51434 31268 51486 31277
rect 53642 31268 53694 31320
rect 54010 31268 54062 31320
rect 54746 31336 54798 31388
rect 36990 31243 37042 31252
rect 36990 31209 36999 31243
rect 36999 31209 37033 31243
rect 37033 31209 37042 31243
rect 36990 31200 37042 31209
rect 51066 31200 51118 31252
rect 57506 31268 57558 31320
rect 57874 31311 57926 31320
rect 54654 31200 54706 31252
rect 47386 31132 47438 31184
rect 49778 31132 49830 31184
rect 50882 31132 50934 31184
rect 54102 31132 54154 31184
rect 54838 31175 54890 31184
rect 54838 31141 54847 31175
rect 54847 31141 54881 31175
rect 54881 31141 54890 31175
rect 54838 31132 54890 31141
rect 57874 31277 57883 31311
rect 57883 31277 57917 31311
rect 57917 31277 57926 31311
rect 57874 31268 57926 31277
rect 58610 31336 58662 31388
rect 67902 31404 67954 31456
rect 68362 31404 68414 31456
rect 69190 31472 69242 31524
rect 71674 31472 71726 31524
rect 73974 31472 74026 31524
rect 78666 31472 78718 31524
rect 82990 31472 83042 31524
rect 88326 31472 88378 31524
rect 88418 31515 88470 31524
rect 88418 31481 88427 31515
rect 88427 31481 88461 31515
rect 88461 31481 88470 31515
rect 88418 31472 88470 31481
rect 68822 31404 68874 31456
rect 63210 31336 63262 31388
rect 60174 31311 60226 31320
rect 60174 31277 60183 31311
rect 60183 31277 60217 31311
rect 60217 31277 60226 31311
rect 60174 31268 60226 31277
rect 62750 31268 62802 31320
rect 61830 31200 61882 31252
rect 68086 31268 68138 31320
rect 73790 31336 73842 31388
rect 71766 31268 71818 31320
rect 60358 31132 60410 31184
rect 65878 31175 65930 31184
rect 65878 31141 65887 31175
rect 65887 31141 65921 31175
rect 65921 31141 65930 31175
rect 65878 31132 65930 31141
rect 66062 31175 66114 31184
rect 66062 31141 66071 31175
rect 66071 31141 66105 31175
rect 66105 31141 66114 31175
rect 66062 31132 66114 31141
rect 68178 31175 68230 31184
rect 68178 31141 68187 31175
rect 68187 31141 68221 31175
rect 68221 31141 68230 31175
rect 68178 31132 68230 31141
rect 73238 31132 73290 31184
rect 74158 31268 74210 31320
rect 75354 31311 75406 31320
rect 75354 31277 75363 31311
rect 75363 31277 75397 31311
rect 75397 31277 75406 31311
rect 75354 31268 75406 31277
rect 76550 31268 76602 31320
rect 74342 31200 74394 31252
rect 81518 31311 81570 31320
rect 80598 31200 80650 31252
rect 81518 31277 81527 31311
rect 81527 31277 81561 31311
rect 81561 31277 81570 31311
rect 81518 31268 81570 31277
rect 82622 31311 82674 31320
rect 82622 31277 82631 31311
rect 82631 31277 82665 31311
rect 82665 31277 82674 31311
rect 82622 31268 82674 31277
rect 84278 31404 84330 31456
rect 84370 31404 84422 31456
rect 89338 31404 89390 31456
rect 90718 31379 90770 31388
rect 88326 31311 88378 31320
rect 88326 31277 88335 31311
rect 88335 31277 88369 31311
rect 88369 31277 88378 31311
rect 88326 31268 88378 31277
rect 90718 31345 90727 31379
rect 90727 31345 90761 31379
rect 90761 31345 90770 31379
rect 90718 31336 90770 31345
rect 90902 31311 90954 31320
rect 90902 31277 90911 31311
rect 90911 31277 90945 31311
rect 90945 31277 90954 31311
rect 90902 31268 90954 31277
rect 91454 31311 91506 31320
rect 91454 31277 91463 31311
rect 91463 31277 91497 31311
rect 91497 31277 91506 31311
rect 91454 31268 91506 31277
rect 80322 31132 80374 31184
rect 80506 31175 80558 31184
rect 80506 31141 80515 31175
rect 80515 31141 80549 31175
rect 80549 31141 80558 31175
rect 80506 31132 80558 31141
rect 80782 31175 80834 31184
rect 80782 31141 80791 31175
rect 80791 31141 80825 31175
rect 80825 31141 80834 31175
rect 80782 31132 80834 31141
rect 6344 31030 6396 31082
rect 6408 31030 6460 31082
rect 6472 31030 6524 31082
rect 6536 31030 6588 31082
rect 11672 31030 11724 31082
rect 11736 31030 11788 31082
rect 11800 31030 11852 31082
rect 11864 31030 11916 31082
rect 17000 31030 17052 31082
rect 17064 31030 17116 31082
rect 17128 31030 17180 31082
rect 17192 31030 17244 31082
rect 22328 31030 22380 31082
rect 22392 31030 22444 31082
rect 22456 31030 22508 31082
rect 22520 31030 22572 31082
rect 27656 31030 27708 31082
rect 27720 31030 27772 31082
rect 27784 31030 27836 31082
rect 27848 31030 27900 31082
rect 32984 31030 33036 31082
rect 33048 31030 33100 31082
rect 33112 31030 33164 31082
rect 33176 31030 33228 31082
rect 38312 31030 38364 31082
rect 38376 31030 38428 31082
rect 38440 31030 38492 31082
rect 38504 31030 38556 31082
rect 43640 31030 43692 31082
rect 43704 31030 43756 31082
rect 43768 31030 43820 31082
rect 43832 31030 43884 31082
rect 48968 31030 49020 31082
rect 49032 31030 49084 31082
rect 49096 31030 49148 31082
rect 49160 31030 49212 31082
rect 54296 31030 54348 31082
rect 54360 31030 54412 31082
rect 54424 31030 54476 31082
rect 54488 31030 54540 31082
rect 59624 31030 59676 31082
rect 59688 31030 59740 31082
rect 59752 31030 59804 31082
rect 59816 31030 59868 31082
rect 64952 31030 65004 31082
rect 65016 31030 65068 31082
rect 65080 31030 65132 31082
rect 65144 31030 65196 31082
rect 70280 31030 70332 31082
rect 70344 31030 70396 31082
rect 70408 31030 70460 31082
rect 70472 31030 70524 31082
rect 75608 31030 75660 31082
rect 75672 31030 75724 31082
rect 75736 31030 75788 31082
rect 75800 31030 75852 31082
rect 80936 31030 80988 31082
rect 81000 31030 81052 31082
rect 81064 31030 81116 31082
rect 81128 31030 81180 31082
rect 86264 31030 86316 31082
rect 86328 31030 86380 31082
rect 86392 31030 86444 31082
rect 86456 31030 86508 31082
rect 91592 31030 91644 31082
rect 91656 31030 91708 31082
rect 91720 31030 91772 31082
rect 91784 31030 91836 31082
rect 4974 30928 5026 30980
rect 5066 30928 5118 30980
rect 14726 30928 14778 30980
rect 15922 30971 15974 30980
rect 15922 30937 15931 30971
rect 15931 30937 15965 30971
rect 15965 30937 15974 30971
rect 15922 30928 15974 30937
rect 17670 30928 17722 30980
rect 11506 30860 11558 30912
rect 6262 30724 6314 30776
rect 6630 30835 6682 30844
rect 6630 30801 6639 30835
rect 6639 30801 6673 30835
rect 6673 30801 6682 30835
rect 6630 30792 6682 30801
rect 6906 30792 6958 30844
rect 10310 30835 10362 30844
rect 10310 30801 10319 30835
rect 10319 30801 10353 30835
rect 10353 30801 10362 30835
rect 10310 30792 10362 30801
rect 10402 30835 10454 30844
rect 10402 30801 10411 30835
rect 10411 30801 10445 30835
rect 10445 30801 10454 30835
rect 10402 30792 10454 30801
rect 11414 30792 11466 30844
rect 12334 30835 12386 30844
rect 12334 30801 12343 30835
rect 12343 30801 12377 30835
rect 12377 30801 12386 30835
rect 12334 30792 12386 30801
rect 12426 30792 12478 30844
rect 12794 30792 12846 30844
rect 19878 30860 19930 30912
rect 14818 30792 14870 30844
rect 15922 30792 15974 30844
rect 16750 30835 16802 30844
rect 16750 30801 16759 30835
rect 16759 30801 16793 30835
rect 16793 30801 16802 30835
rect 16750 30792 16802 30801
rect 17578 30792 17630 30844
rect 18866 30792 18918 30844
rect 5066 30656 5118 30708
rect 9482 30724 9534 30776
rect 10126 30767 10178 30776
rect 10126 30733 10135 30767
rect 10135 30733 10169 30767
rect 10169 30733 10178 30767
rect 10126 30724 10178 30733
rect 11506 30724 11558 30776
rect 8194 30656 8246 30708
rect 6906 30588 6958 30640
rect 7090 30588 7142 30640
rect 13162 30588 13214 30640
rect 18038 30724 18090 30776
rect 29262 30928 29314 30980
rect 29354 30928 29406 30980
rect 30918 30860 30970 30912
rect 38646 30928 38698 30980
rect 68178 30928 68230 30980
rect 52170 30860 52222 30912
rect 23926 30792 23978 30844
rect 24846 30792 24898 30844
rect 28802 30792 28854 30844
rect 23098 30724 23150 30776
rect 27514 30724 27566 30776
rect 27698 30724 27750 30776
rect 33310 30792 33362 30844
rect 16382 30656 16434 30708
rect 19510 30656 19562 30708
rect 23742 30656 23794 30708
rect 27330 30656 27382 30708
rect 17578 30631 17630 30640
rect 17578 30597 17587 30631
rect 17587 30597 17621 30631
rect 17621 30597 17630 30631
rect 17578 30588 17630 30597
rect 18866 30588 18918 30640
rect 23650 30631 23702 30640
rect 23650 30597 23659 30631
rect 23659 30597 23693 30631
rect 23693 30597 23702 30631
rect 23650 30588 23702 30597
rect 28710 30631 28762 30640
rect 28710 30597 28719 30631
rect 28719 30597 28753 30631
rect 28753 30597 28762 30631
rect 28710 30588 28762 30597
rect 34506 30724 34558 30776
rect 34046 30631 34098 30640
rect 34046 30597 34055 30631
rect 34055 30597 34089 30631
rect 34089 30597 34098 30631
rect 34046 30588 34098 30597
rect 34230 30656 34282 30708
rect 34690 30656 34742 30708
rect 36990 30792 37042 30844
rect 43614 30792 43666 30844
rect 44442 30835 44494 30844
rect 44442 30801 44451 30835
rect 44451 30801 44485 30835
rect 44485 30801 44494 30835
rect 44442 30792 44494 30801
rect 44626 30792 44678 30844
rect 53826 30860 53878 30912
rect 35058 30656 35110 30708
rect 37818 30724 37870 30776
rect 42878 30724 42930 30776
rect 43430 30724 43482 30776
rect 47662 30724 47714 30776
rect 48858 30767 48910 30776
rect 48858 30733 48867 30767
rect 48867 30733 48901 30767
rect 48901 30733 48910 30767
rect 48858 30724 48910 30733
rect 50698 30724 50750 30776
rect 54102 30792 54154 30844
rect 57874 30860 57926 30912
rect 62106 30860 62158 30912
rect 54838 30792 54890 30844
rect 58150 30835 58202 30844
rect 52814 30767 52866 30776
rect 52814 30733 52823 30767
rect 52823 30733 52857 30767
rect 52857 30733 52866 30767
rect 52814 30724 52866 30733
rect 52906 30724 52958 30776
rect 58150 30801 58159 30835
rect 58159 30801 58193 30835
rect 58193 30801 58202 30835
rect 58150 30792 58202 30801
rect 58334 30792 58386 30844
rect 58518 30792 58570 30844
rect 62014 30792 62066 30844
rect 63394 30860 63446 30912
rect 62658 30792 62710 30844
rect 63026 30792 63078 30844
rect 69926 30792 69978 30844
rect 71214 30792 71266 30844
rect 74158 30835 74210 30844
rect 46098 30656 46150 30708
rect 36990 30588 37042 30640
rect 45454 30631 45506 30640
rect 45454 30597 45463 30631
rect 45463 30597 45497 30631
rect 45497 30597 45506 30631
rect 45454 30588 45506 30597
rect 48306 30588 48358 30640
rect 48674 30631 48726 30640
rect 48674 30597 48683 30631
rect 48683 30597 48717 30631
rect 48717 30597 48726 30631
rect 54010 30656 54062 30708
rect 48674 30588 48726 30597
rect 49410 30588 49462 30640
rect 59622 30588 59674 30640
rect 66522 30767 66574 30776
rect 66522 30733 66531 30767
rect 66531 30733 66565 30767
rect 66565 30733 66574 30767
rect 66522 30724 66574 30733
rect 66798 30767 66850 30776
rect 66798 30733 66807 30767
rect 66807 30733 66841 30767
rect 66841 30733 66850 30767
rect 66798 30724 66850 30733
rect 66982 30724 67034 30776
rect 71398 30767 71450 30776
rect 71398 30733 71407 30767
rect 71407 30733 71441 30767
rect 71441 30733 71450 30767
rect 71398 30724 71450 30733
rect 71766 30724 71818 30776
rect 72318 30724 72370 30776
rect 74158 30801 74167 30835
rect 74167 30801 74201 30835
rect 74201 30801 74210 30835
rect 74158 30792 74210 30801
rect 75262 30860 75314 30912
rect 79678 30928 79730 30980
rect 84830 30971 84882 30980
rect 84830 30937 84839 30971
rect 84839 30937 84873 30971
rect 84873 30937 84882 30971
rect 84830 30928 84882 30937
rect 75078 30792 75130 30844
rect 75538 30792 75590 30844
rect 77470 30792 77522 30844
rect 77102 30767 77154 30776
rect 77102 30733 77111 30767
rect 77111 30733 77145 30767
rect 77145 30733 77154 30767
rect 77102 30724 77154 30733
rect 78114 30724 78166 30776
rect 80782 30792 80834 30844
rect 80966 30835 81018 30844
rect 80966 30801 80975 30835
rect 80975 30801 81009 30835
rect 81009 30801 81018 30835
rect 80966 30792 81018 30801
rect 81518 30792 81570 30844
rect 82070 30835 82122 30844
rect 82070 30801 82079 30835
rect 82079 30801 82113 30835
rect 82113 30801 82122 30835
rect 82070 30792 82122 30801
rect 87682 30928 87734 30980
rect 89706 30971 89758 30980
rect 89706 30937 89715 30971
rect 89715 30937 89749 30971
rect 89749 30937 89758 30971
rect 89706 30928 89758 30937
rect 89246 30860 89298 30912
rect 88418 30835 88470 30844
rect 81058 30724 81110 30776
rect 88418 30801 88427 30835
rect 88427 30801 88461 30835
rect 88461 30801 88470 30835
rect 88418 30792 88470 30801
rect 88786 30792 88838 30844
rect 89614 30835 89666 30844
rect 89614 30801 89623 30835
rect 89623 30801 89657 30835
rect 89657 30801 89666 30835
rect 89614 30792 89666 30801
rect 90902 30792 90954 30844
rect 91362 30835 91414 30844
rect 91362 30801 91371 30835
rect 91371 30801 91405 30835
rect 91405 30801 91414 30835
rect 91362 30792 91414 30801
rect 61278 30656 61330 30708
rect 66062 30656 66114 30708
rect 74342 30656 74394 30708
rect 74434 30656 74486 30708
rect 67258 30588 67310 30640
rect 69190 30631 69242 30640
rect 69190 30597 69199 30631
rect 69199 30597 69233 30631
rect 69233 30597 69242 30631
rect 69190 30588 69242 30597
rect 75446 30656 75498 30708
rect 77010 30656 77062 30708
rect 80598 30656 80650 30708
rect 86762 30724 86814 30776
rect 77746 30588 77798 30640
rect 78022 30588 78074 30640
rect 78850 30631 78902 30640
rect 78850 30597 78859 30631
rect 78859 30597 78893 30631
rect 78893 30597 78902 30631
rect 78850 30588 78902 30597
rect 86118 30588 86170 30640
rect 91454 30588 91506 30640
rect 3680 30486 3732 30538
rect 3744 30486 3796 30538
rect 3808 30486 3860 30538
rect 3872 30486 3924 30538
rect 9008 30486 9060 30538
rect 9072 30486 9124 30538
rect 9136 30486 9188 30538
rect 9200 30486 9252 30538
rect 14336 30486 14388 30538
rect 14400 30486 14452 30538
rect 14464 30486 14516 30538
rect 14528 30486 14580 30538
rect 19664 30486 19716 30538
rect 19728 30486 19780 30538
rect 19792 30486 19844 30538
rect 19856 30486 19908 30538
rect 24992 30486 25044 30538
rect 25056 30486 25108 30538
rect 25120 30486 25172 30538
rect 25184 30486 25236 30538
rect 30320 30486 30372 30538
rect 30384 30486 30436 30538
rect 30448 30486 30500 30538
rect 30512 30486 30564 30538
rect 35648 30486 35700 30538
rect 35712 30486 35764 30538
rect 35776 30486 35828 30538
rect 35840 30486 35892 30538
rect 40976 30486 41028 30538
rect 41040 30486 41092 30538
rect 41104 30486 41156 30538
rect 41168 30486 41220 30538
rect 46304 30486 46356 30538
rect 46368 30486 46420 30538
rect 46432 30486 46484 30538
rect 46496 30486 46548 30538
rect 51632 30486 51684 30538
rect 51696 30486 51748 30538
rect 51760 30486 51812 30538
rect 51824 30486 51876 30538
rect 56960 30486 57012 30538
rect 57024 30486 57076 30538
rect 57088 30486 57140 30538
rect 57152 30486 57204 30538
rect 62288 30486 62340 30538
rect 62352 30486 62404 30538
rect 62416 30486 62468 30538
rect 62480 30486 62532 30538
rect 67616 30486 67668 30538
rect 67680 30486 67732 30538
rect 67744 30486 67796 30538
rect 67808 30486 67860 30538
rect 72944 30486 72996 30538
rect 73008 30486 73060 30538
rect 73072 30486 73124 30538
rect 73136 30486 73188 30538
rect 78272 30486 78324 30538
rect 78336 30486 78388 30538
rect 78400 30486 78452 30538
rect 78464 30486 78516 30538
rect 83600 30486 83652 30538
rect 83664 30486 83716 30538
rect 83728 30486 83780 30538
rect 83792 30486 83844 30538
rect 88928 30486 88980 30538
rect 88992 30486 89044 30538
rect 89056 30486 89108 30538
rect 89120 30486 89172 30538
rect 3226 30427 3278 30436
rect 3226 30393 3235 30427
rect 3235 30393 3269 30427
rect 3269 30393 3278 30427
rect 3226 30384 3278 30393
rect 5710 30384 5762 30436
rect 8102 30316 8154 30368
rect 8286 30316 8338 30368
rect 2398 30248 2450 30300
rect 3042 30180 3094 30232
rect 6906 30248 6958 30300
rect 7090 30291 7142 30300
rect 7090 30257 7099 30291
rect 7099 30257 7133 30291
rect 7133 30257 7142 30291
rect 7090 30248 7142 30257
rect 9298 30248 9350 30300
rect 12610 30316 12662 30368
rect 12334 30248 12386 30300
rect 5066 30223 5118 30232
rect 5066 30189 5075 30223
rect 5075 30189 5109 30223
rect 5109 30189 5118 30223
rect 5066 30180 5118 30189
rect 6262 30180 6314 30232
rect 6814 30180 6866 30232
rect 7734 30180 7786 30232
rect 7918 30223 7970 30232
rect 7918 30189 7927 30223
rect 7927 30189 7961 30223
rect 7961 30189 7970 30223
rect 7918 30180 7970 30189
rect 8194 30223 8246 30232
rect 8194 30189 8203 30223
rect 8203 30189 8237 30223
rect 8237 30189 8246 30223
rect 8194 30180 8246 30189
rect 9482 30223 9534 30232
rect 9482 30189 9491 30223
rect 9491 30189 9525 30223
rect 9525 30189 9534 30223
rect 9482 30180 9534 30189
rect 12518 30223 12570 30232
rect 12518 30189 12527 30223
rect 12527 30189 12561 30223
rect 12561 30189 12570 30223
rect 12518 30180 12570 30189
rect 12794 30223 12846 30232
rect 12794 30189 12803 30223
rect 12803 30189 12837 30223
rect 12837 30189 12846 30223
rect 12794 30180 12846 30189
rect 2950 30044 3002 30096
rect 6722 30044 6774 30096
rect 11414 30112 11466 30164
rect 11966 30155 12018 30164
rect 11966 30121 11975 30155
rect 11975 30121 12009 30155
rect 12009 30121 12018 30155
rect 11966 30112 12018 30121
rect 18866 30384 18918 30436
rect 23834 30384 23886 30436
rect 27146 30384 27198 30436
rect 27974 30384 28026 30436
rect 36806 30384 36858 30436
rect 38646 30384 38698 30436
rect 42786 30384 42838 30436
rect 23650 30316 23702 30368
rect 24018 30316 24070 30368
rect 18682 30248 18734 30300
rect 19602 30291 19654 30300
rect 19602 30257 19611 30291
rect 19611 30257 19645 30291
rect 19645 30257 19654 30291
rect 19602 30248 19654 30257
rect 23098 30291 23150 30300
rect 23098 30257 23107 30291
rect 23107 30257 23141 30291
rect 23141 30257 23150 30291
rect 23098 30248 23150 30257
rect 27698 30316 27750 30368
rect 28342 30316 28394 30368
rect 29354 30316 29406 30368
rect 30090 30316 30142 30368
rect 34046 30248 34098 30300
rect 40946 30316 40998 30368
rect 43706 30316 43758 30368
rect 43982 30359 44034 30368
rect 43982 30325 43991 30359
rect 43991 30325 44025 30359
rect 44025 30325 44034 30359
rect 43982 30316 44034 30325
rect 17486 30180 17538 30232
rect 18038 30180 18090 30232
rect 14726 30112 14778 30164
rect 17762 30155 17814 30164
rect 17762 30121 17771 30155
rect 17771 30121 17805 30155
rect 17805 30121 17814 30155
rect 17762 30112 17814 30121
rect 13162 30044 13214 30096
rect 15922 30044 15974 30096
rect 17394 30044 17446 30096
rect 23650 30180 23702 30232
rect 22822 30155 22874 30164
rect 22822 30121 22831 30155
rect 22831 30121 22865 30155
rect 22865 30121 22874 30155
rect 23834 30180 23886 30232
rect 24294 30180 24346 30232
rect 24478 30223 24530 30232
rect 24478 30189 24487 30223
rect 24487 30189 24521 30223
rect 24521 30189 24530 30223
rect 24478 30180 24530 30189
rect 27054 30180 27106 30232
rect 27330 30180 27382 30232
rect 34230 30180 34282 30232
rect 22822 30112 22874 30121
rect 23006 30044 23058 30096
rect 27422 30112 27474 30164
rect 36898 30223 36950 30232
rect 36898 30189 36907 30223
rect 36907 30189 36941 30223
rect 36941 30189 36950 30223
rect 36898 30180 36950 30189
rect 28894 30044 28946 30096
rect 34414 30087 34466 30096
rect 34414 30053 34423 30087
rect 34423 30053 34457 30087
rect 34457 30053 34466 30087
rect 34414 30044 34466 30053
rect 48674 30384 48726 30436
rect 62106 30384 62158 30436
rect 67350 30384 67402 30436
rect 53642 30359 53694 30368
rect 53642 30325 53651 30359
rect 53651 30325 53685 30359
rect 53685 30325 53694 30359
rect 53642 30316 53694 30325
rect 60174 30359 60226 30368
rect 43706 30223 43758 30232
rect 38186 30044 38238 30096
rect 38646 30087 38698 30096
rect 38646 30053 38655 30087
rect 38655 30053 38689 30087
rect 38689 30053 38698 30087
rect 38646 30044 38698 30053
rect 39750 30044 39802 30096
rect 43062 30087 43114 30096
rect 43062 30053 43071 30087
rect 43071 30053 43105 30087
rect 43105 30053 43114 30087
rect 43062 30044 43114 30053
rect 43706 30189 43715 30223
rect 43715 30189 43749 30223
rect 43749 30189 43758 30223
rect 43706 30180 43758 30189
rect 44074 30112 44126 30164
rect 44166 30044 44218 30096
rect 45362 30044 45414 30096
rect 53918 30248 53970 30300
rect 59622 30291 59674 30300
rect 47846 30223 47898 30232
rect 47846 30189 47855 30223
rect 47855 30189 47889 30223
rect 47889 30189 47898 30223
rect 47846 30180 47898 30189
rect 51066 30180 51118 30232
rect 51986 30180 52038 30232
rect 48858 30112 48910 30164
rect 52630 30180 52682 30232
rect 54010 30180 54062 30232
rect 54194 30112 54246 30164
rect 59622 30257 59631 30291
rect 59631 30257 59665 30291
rect 59665 30257 59674 30291
rect 59622 30248 59674 30257
rect 60174 30325 60183 30359
rect 60183 30325 60217 30359
rect 60217 30325 60226 30359
rect 60174 30316 60226 30325
rect 63026 30316 63078 30368
rect 66062 30316 66114 30368
rect 70754 30384 70806 30436
rect 71030 30384 71082 30436
rect 74434 30384 74486 30436
rect 74526 30384 74578 30436
rect 76918 30384 76970 30436
rect 77102 30384 77154 30436
rect 78022 30384 78074 30436
rect 82070 30384 82122 30436
rect 86762 30427 86814 30436
rect 86762 30393 86771 30427
rect 86771 30393 86805 30427
rect 86805 30393 86814 30427
rect 86762 30384 86814 30393
rect 89614 30384 89666 30436
rect 91362 30384 91414 30436
rect 62290 30248 62342 30300
rect 66522 30248 66574 30300
rect 66614 30248 66666 30300
rect 69834 30248 69886 30300
rect 70846 30248 70898 30300
rect 58610 30223 58662 30232
rect 58610 30189 58619 30223
rect 58619 30189 58653 30223
rect 58653 30189 58662 30223
rect 58610 30180 58662 30189
rect 59162 30223 59214 30232
rect 59162 30189 59171 30223
rect 59171 30189 59205 30223
rect 59205 30189 59214 30223
rect 59990 30223 60042 30232
rect 59162 30180 59214 30189
rect 59990 30189 59999 30223
rect 59999 30189 60033 30223
rect 60033 30189 60042 30223
rect 59990 30180 60042 30189
rect 62658 30223 62710 30232
rect 54010 30087 54062 30096
rect 54010 30053 54019 30087
rect 54019 30053 54053 30087
rect 54053 30053 54062 30087
rect 54010 30044 54062 30053
rect 54102 30044 54154 30096
rect 55022 30087 55074 30096
rect 55022 30053 55031 30087
rect 55031 30053 55065 30087
rect 55065 30053 55074 30087
rect 55022 30044 55074 30053
rect 59530 30112 59582 30164
rect 62658 30189 62667 30223
rect 62667 30189 62701 30223
rect 62701 30189 62710 30223
rect 62658 30180 62710 30189
rect 65786 30180 65838 30232
rect 66890 30223 66942 30232
rect 66890 30189 66899 30223
rect 66899 30189 66933 30223
rect 66933 30189 66942 30223
rect 66890 30180 66942 30189
rect 69926 30223 69978 30232
rect 62566 30155 62618 30164
rect 62566 30121 62575 30155
rect 62575 30121 62609 30155
rect 62609 30121 62618 30155
rect 62566 30112 62618 30121
rect 63118 30155 63170 30164
rect 63118 30121 63127 30155
rect 63127 30121 63161 30155
rect 63161 30121 63170 30155
rect 63118 30112 63170 30121
rect 63946 30112 63998 30164
rect 65418 30112 65470 30164
rect 67166 30112 67218 30164
rect 67258 30112 67310 30164
rect 68638 30112 68690 30164
rect 69926 30189 69935 30223
rect 69935 30189 69969 30223
rect 69969 30189 69978 30223
rect 69926 30180 69978 30189
rect 71030 30223 71082 30232
rect 71030 30189 71039 30223
rect 71039 30189 71073 30223
rect 71073 30189 71082 30223
rect 71030 30180 71082 30189
rect 75538 30248 75590 30300
rect 72318 30223 72370 30232
rect 72318 30189 72327 30223
rect 72327 30189 72361 30223
rect 72361 30189 72370 30223
rect 72318 30180 72370 30189
rect 72778 30180 72830 30232
rect 73882 30223 73934 30232
rect 73882 30189 73891 30223
rect 73891 30189 73925 30223
rect 73925 30189 73934 30223
rect 73882 30180 73934 30189
rect 75998 30180 76050 30232
rect 76182 30223 76234 30232
rect 76182 30189 76191 30223
rect 76191 30189 76225 30223
rect 76225 30189 76234 30223
rect 76918 30248 76970 30300
rect 77746 30248 77798 30300
rect 93294 30248 93346 30300
rect 76182 30180 76234 30189
rect 76642 30223 76694 30232
rect 76642 30189 76651 30223
rect 76651 30189 76685 30223
rect 76685 30189 76694 30223
rect 76642 30180 76694 30189
rect 77470 30223 77522 30232
rect 77470 30189 77479 30223
rect 77479 30189 77513 30223
rect 77513 30189 77522 30223
rect 77470 30180 77522 30189
rect 81058 30223 81110 30232
rect 75078 30112 75130 30164
rect 78022 30112 78074 30164
rect 63394 30044 63446 30096
rect 67718 30044 67770 30096
rect 70018 30044 70070 30096
rect 70754 30044 70806 30096
rect 74158 30044 74210 30096
rect 74342 30087 74394 30096
rect 74342 30053 74351 30087
rect 74351 30053 74385 30087
rect 74385 30053 74394 30087
rect 74342 30044 74394 30053
rect 74710 30044 74762 30096
rect 75354 30087 75406 30096
rect 75354 30053 75363 30087
rect 75363 30053 75397 30087
rect 75397 30053 75406 30087
rect 75354 30044 75406 30053
rect 75906 30044 75958 30096
rect 79770 30112 79822 30164
rect 79494 30044 79546 30096
rect 81058 30189 81067 30223
rect 81067 30189 81101 30223
rect 81101 30189 81110 30223
rect 81058 30180 81110 30189
rect 86026 30180 86078 30232
rect 88510 30223 88562 30232
rect 88510 30189 88519 30223
rect 88519 30189 88553 30223
rect 88553 30189 88562 30223
rect 88510 30180 88562 30189
rect 85198 30087 85250 30096
rect 85198 30053 85207 30087
rect 85207 30053 85241 30087
rect 85241 30053 85250 30087
rect 85198 30044 85250 30053
rect 87590 30044 87642 30096
rect 88786 30180 88838 30232
rect 89246 30180 89298 30232
rect 90442 30180 90494 30232
rect 90994 30223 91046 30232
rect 90994 30189 91003 30223
rect 91003 30189 91037 30223
rect 91037 30189 91046 30223
rect 90994 30180 91046 30189
rect 6344 29942 6396 29994
rect 6408 29942 6460 29994
rect 6472 29942 6524 29994
rect 6536 29942 6588 29994
rect 11672 29942 11724 29994
rect 11736 29942 11788 29994
rect 11800 29942 11852 29994
rect 11864 29942 11916 29994
rect 17000 29942 17052 29994
rect 17064 29942 17116 29994
rect 17128 29942 17180 29994
rect 17192 29942 17244 29994
rect 22328 29942 22380 29994
rect 22392 29942 22444 29994
rect 22456 29942 22508 29994
rect 22520 29942 22572 29994
rect 27656 29942 27708 29994
rect 27720 29942 27772 29994
rect 27784 29942 27836 29994
rect 27848 29942 27900 29994
rect 32984 29942 33036 29994
rect 33048 29942 33100 29994
rect 33112 29942 33164 29994
rect 33176 29942 33228 29994
rect 38312 29942 38364 29994
rect 38376 29942 38428 29994
rect 38440 29942 38492 29994
rect 38504 29942 38556 29994
rect 43640 29942 43692 29994
rect 43704 29942 43756 29994
rect 43768 29942 43820 29994
rect 43832 29942 43884 29994
rect 48968 29942 49020 29994
rect 49032 29942 49084 29994
rect 49096 29942 49148 29994
rect 49160 29942 49212 29994
rect 54296 29942 54348 29994
rect 54360 29942 54412 29994
rect 54424 29942 54476 29994
rect 54488 29942 54540 29994
rect 59624 29942 59676 29994
rect 59688 29942 59740 29994
rect 59752 29942 59804 29994
rect 59816 29942 59868 29994
rect 64952 29942 65004 29994
rect 65016 29942 65068 29994
rect 65080 29942 65132 29994
rect 65144 29942 65196 29994
rect 70280 29942 70332 29994
rect 70344 29942 70396 29994
rect 70408 29942 70460 29994
rect 70472 29942 70524 29994
rect 75608 29942 75660 29994
rect 75672 29942 75724 29994
rect 75736 29942 75788 29994
rect 75800 29942 75852 29994
rect 80936 29942 80988 29994
rect 81000 29942 81052 29994
rect 81064 29942 81116 29994
rect 81128 29942 81180 29994
rect 86264 29942 86316 29994
rect 86328 29942 86380 29994
rect 86392 29942 86444 29994
rect 86456 29942 86508 29994
rect 91592 29942 91644 29994
rect 91656 29942 91708 29994
rect 91720 29942 91772 29994
rect 91784 29942 91836 29994
rect 11414 29840 11466 29892
rect 5710 29815 5762 29824
rect 5710 29781 5719 29815
rect 5719 29781 5753 29815
rect 5753 29781 5762 29815
rect 5710 29772 5762 29781
rect 8102 29772 8154 29824
rect 9482 29815 9534 29824
rect 9482 29781 9491 29815
rect 9491 29781 9525 29815
rect 9525 29781 9534 29815
rect 9482 29772 9534 29781
rect 10310 29772 10362 29824
rect 6170 29747 6222 29756
rect 6170 29713 6179 29747
rect 6179 29713 6213 29747
rect 6213 29713 6222 29747
rect 6170 29704 6222 29713
rect 6354 29747 6406 29756
rect 6354 29713 6363 29747
rect 6363 29713 6397 29747
rect 6397 29713 6406 29747
rect 6354 29704 6406 29713
rect 6446 29704 6498 29756
rect 6722 29704 6774 29756
rect 8010 29704 8062 29756
rect 8194 29704 8246 29756
rect 9390 29747 9442 29756
rect 9390 29713 9399 29747
rect 9399 29713 9433 29747
rect 9433 29713 9442 29747
rect 9390 29704 9442 29713
rect 17486 29883 17538 29892
rect 17486 29849 17495 29883
rect 17495 29849 17529 29883
rect 17529 29849 17538 29883
rect 17486 29840 17538 29849
rect 18958 29840 19010 29892
rect 22730 29840 22782 29892
rect 12794 29704 12846 29756
rect 9850 29679 9902 29688
rect 9850 29645 9859 29679
rect 9859 29645 9893 29679
rect 9893 29645 9902 29679
rect 9850 29636 9902 29645
rect 9298 29568 9350 29620
rect 10126 29568 10178 29620
rect 13162 29704 13214 29756
rect 15922 29704 15974 29756
rect 4330 29500 4382 29552
rect 8470 29500 8522 29552
rect 9482 29500 9534 29552
rect 12886 29500 12938 29552
rect 15830 29500 15882 29552
rect 22822 29772 22874 29824
rect 16382 29747 16434 29756
rect 16382 29713 16391 29747
rect 16391 29713 16425 29747
rect 16425 29713 16434 29747
rect 16382 29704 16434 29713
rect 19602 29704 19654 29756
rect 23742 29747 23794 29756
rect 17670 29636 17722 29688
rect 21810 29636 21862 29688
rect 23742 29713 23751 29747
rect 23751 29713 23785 29747
rect 23785 29713 23794 29747
rect 23742 29704 23794 29713
rect 24294 29772 24346 29824
rect 27514 29815 27566 29824
rect 27514 29781 27523 29815
rect 27523 29781 27557 29815
rect 27557 29781 27566 29815
rect 27514 29772 27566 29781
rect 27606 29772 27658 29824
rect 28894 29840 28946 29892
rect 24478 29704 24530 29756
rect 24110 29636 24162 29688
rect 27054 29636 27106 29688
rect 27606 29636 27658 29688
rect 27974 29747 28026 29756
rect 27974 29713 27983 29747
rect 27983 29713 28017 29747
rect 28017 29713 28026 29747
rect 28158 29747 28210 29756
rect 27974 29704 28026 29713
rect 28158 29713 28167 29747
rect 28167 29713 28201 29747
rect 28201 29713 28210 29747
rect 28158 29704 28210 29713
rect 28618 29772 28670 29824
rect 28710 29747 28762 29756
rect 28710 29713 28719 29747
rect 28719 29713 28753 29747
rect 28753 29713 28762 29747
rect 28710 29704 28762 29713
rect 29078 29704 29130 29756
rect 29170 29636 29222 29688
rect 30090 29772 30142 29824
rect 34230 29840 34282 29892
rect 30826 29772 30878 29824
rect 34966 29840 35018 29892
rect 37358 29883 37410 29892
rect 37358 29849 37367 29883
rect 37367 29849 37401 29883
rect 37401 29849 37410 29883
rect 37358 29840 37410 29849
rect 40946 29840 40998 29892
rect 43062 29840 43114 29892
rect 43982 29883 44034 29892
rect 34414 29772 34466 29824
rect 30090 29636 30142 29688
rect 36898 29704 36950 29756
rect 37358 29704 37410 29756
rect 38830 29704 38882 29756
rect 34506 29636 34558 29688
rect 17302 29568 17354 29620
rect 22822 29568 22874 29620
rect 23190 29568 23242 29620
rect 24662 29568 24714 29620
rect 25858 29568 25910 29620
rect 27974 29568 28026 29620
rect 28158 29568 28210 29620
rect 36346 29568 36398 29620
rect 18314 29500 18366 29552
rect 28986 29500 29038 29552
rect 29078 29500 29130 29552
rect 37818 29500 37870 29552
rect 39198 29747 39250 29756
rect 39198 29713 39207 29747
rect 39207 29713 39241 29747
rect 39241 29713 39250 29747
rect 39198 29704 39250 29713
rect 39474 29704 39526 29756
rect 42786 29747 42838 29756
rect 42786 29713 42795 29747
rect 42795 29713 42829 29747
rect 42829 29713 42838 29747
rect 42786 29704 42838 29713
rect 43062 29704 43114 29756
rect 43430 29747 43482 29756
rect 43430 29713 43439 29747
rect 43439 29713 43473 29747
rect 43473 29713 43482 29747
rect 43430 29704 43482 29713
rect 43522 29747 43574 29756
rect 43522 29713 43531 29747
rect 43531 29713 43565 29747
rect 43565 29713 43574 29747
rect 43982 29849 43991 29883
rect 43991 29849 44025 29883
rect 44025 29849 44034 29883
rect 43982 29840 44034 29849
rect 44166 29840 44218 29892
rect 49410 29840 49462 29892
rect 54102 29840 54154 29892
rect 54194 29840 54246 29892
rect 54654 29840 54706 29892
rect 50790 29772 50842 29824
rect 52446 29772 52498 29824
rect 43522 29704 43574 29713
rect 50698 29704 50750 29756
rect 50882 29704 50934 29756
rect 55022 29772 55074 29824
rect 58610 29840 58662 29892
rect 60174 29840 60226 29892
rect 60358 29883 60410 29892
rect 60358 29849 60367 29883
rect 60367 29849 60401 29883
rect 60401 29849 60410 29883
rect 60358 29840 60410 29849
rect 61186 29840 61238 29892
rect 66798 29883 66850 29892
rect 66798 29849 66807 29883
rect 66807 29849 66841 29883
rect 66841 29849 66850 29883
rect 66798 29840 66850 29849
rect 65786 29815 65838 29824
rect 52814 29704 52866 29756
rect 53826 29704 53878 29756
rect 39750 29568 39802 29620
rect 52262 29568 52314 29620
rect 53918 29568 53970 29620
rect 54102 29704 54154 29756
rect 56402 29704 56454 29756
rect 65786 29781 65795 29815
rect 65795 29781 65829 29815
rect 65829 29781 65838 29815
rect 65786 29772 65838 29781
rect 61278 29636 61330 29688
rect 63118 29704 63170 29756
rect 65326 29747 65378 29756
rect 65326 29713 65335 29747
rect 65335 29713 65369 29747
rect 65369 29713 65378 29747
rect 65326 29704 65378 29713
rect 54378 29568 54430 29620
rect 54470 29568 54522 29620
rect 60450 29568 60502 29620
rect 61186 29568 61238 29620
rect 62290 29568 62342 29620
rect 62750 29636 62802 29688
rect 68638 29772 68690 29824
rect 67442 29704 67494 29756
rect 67718 29747 67770 29756
rect 67718 29713 67727 29747
rect 67727 29713 67761 29747
rect 67761 29713 67770 29747
rect 67718 29704 67770 29713
rect 69006 29704 69058 29756
rect 69098 29747 69150 29756
rect 69098 29713 69107 29747
rect 69107 29713 69141 29747
rect 69141 29713 69150 29747
rect 71398 29772 71450 29824
rect 74158 29772 74210 29824
rect 77378 29840 77430 29892
rect 77746 29840 77798 29892
rect 78114 29883 78166 29892
rect 78114 29849 78123 29883
rect 78123 29849 78157 29883
rect 78157 29849 78166 29883
rect 78114 29840 78166 29849
rect 79126 29840 79178 29892
rect 69098 29704 69150 29713
rect 68638 29636 68690 29688
rect 70846 29747 70898 29756
rect 70846 29713 70855 29747
rect 70855 29713 70889 29747
rect 70889 29713 70898 29747
rect 70846 29704 70898 29713
rect 69650 29679 69702 29688
rect 69650 29645 69659 29679
rect 69659 29645 69693 29679
rect 69693 29645 69702 29679
rect 69650 29636 69702 29645
rect 70018 29636 70070 29688
rect 72778 29747 72830 29756
rect 72778 29713 72787 29747
rect 72787 29713 72821 29747
rect 72821 29713 72830 29747
rect 72778 29704 72830 29713
rect 74342 29704 74394 29756
rect 75906 29772 75958 29824
rect 75998 29772 76050 29824
rect 76274 29772 76326 29824
rect 79678 29772 79730 29824
rect 74986 29747 75038 29756
rect 74986 29713 74995 29747
rect 74995 29713 75029 29747
rect 75029 29713 75038 29747
rect 74986 29704 75038 29713
rect 75170 29747 75222 29756
rect 75170 29713 75180 29747
rect 75180 29713 75214 29747
rect 75214 29713 75222 29747
rect 78022 29747 78074 29756
rect 75170 29704 75222 29713
rect 78022 29713 78031 29747
rect 78031 29713 78065 29747
rect 78065 29713 78074 29747
rect 78022 29704 78074 29713
rect 78942 29704 78994 29756
rect 84094 29840 84146 29892
rect 84554 29840 84606 29892
rect 87774 29883 87826 29892
rect 87774 29849 87783 29883
rect 87783 29849 87817 29883
rect 87817 29849 87826 29883
rect 87774 29840 87826 29849
rect 88510 29840 88562 29892
rect 80322 29772 80374 29824
rect 86670 29772 86722 29824
rect 84186 29747 84238 29756
rect 84186 29713 84195 29747
rect 84195 29713 84229 29747
rect 84229 29713 84238 29747
rect 84186 29704 84238 29713
rect 86118 29747 86170 29756
rect 86118 29713 86127 29747
rect 86127 29713 86161 29747
rect 86161 29713 86170 29747
rect 87682 29747 87734 29756
rect 86118 29704 86170 29713
rect 87682 29713 87691 29747
rect 87691 29713 87725 29747
rect 87725 29713 87734 29747
rect 87682 29704 87734 29713
rect 90534 29747 90586 29756
rect 90534 29713 90543 29747
rect 90543 29713 90577 29747
rect 90577 29713 90586 29747
rect 90534 29704 90586 29713
rect 90626 29704 90678 29756
rect 39198 29500 39250 29552
rect 46834 29500 46886 29552
rect 47846 29500 47898 29552
rect 48398 29500 48450 29552
rect 52446 29500 52498 29552
rect 52630 29500 52682 29552
rect 54010 29500 54062 29552
rect 62842 29500 62894 29552
rect 63946 29500 63998 29552
rect 67166 29500 67218 29552
rect 67350 29500 67402 29552
rect 68086 29568 68138 29620
rect 68178 29568 68230 29620
rect 74710 29636 74762 29688
rect 75078 29636 75130 29688
rect 75538 29636 75590 29688
rect 75998 29636 76050 29688
rect 69558 29500 69610 29552
rect 69742 29500 69794 29552
rect 71030 29543 71082 29552
rect 71030 29509 71039 29543
rect 71039 29509 71073 29543
rect 71073 29509 71082 29543
rect 71030 29500 71082 29509
rect 75170 29568 75222 29620
rect 76918 29636 76970 29688
rect 77010 29636 77062 29688
rect 79126 29679 79178 29688
rect 79126 29645 79135 29679
rect 79135 29645 79169 29679
rect 79169 29645 79178 29679
rect 79126 29636 79178 29645
rect 80598 29679 80650 29688
rect 80598 29645 80607 29679
rect 80607 29645 80641 29679
rect 80641 29645 80650 29679
rect 80598 29636 80650 29645
rect 76550 29568 76602 29620
rect 83174 29568 83226 29620
rect 85842 29679 85894 29688
rect 85842 29645 85851 29679
rect 85851 29645 85885 29679
rect 85885 29645 85894 29679
rect 85842 29636 85894 29645
rect 86026 29636 86078 29688
rect 73238 29500 73290 29552
rect 76274 29500 76326 29552
rect 76918 29543 76970 29552
rect 76918 29509 76927 29543
rect 76927 29509 76961 29543
rect 76961 29509 76970 29543
rect 76918 29500 76970 29509
rect 90810 29543 90862 29552
rect 90810 29509 90819 29543
rect 90819 29509 90853 29543
rect 90853 29509 90862 29543
rect 90810 29500 90862 29509
rect 3680 29398 3732 29450
rect 3744 29398 3796 29450
rect 3808 29398 3860 29450
rect 3872 29398 3924 29450
rect 9008 29398 9060 29450
rect 9072 29398 9124 29450
rect 9136 29398 9188 29450
rect 9200 29398 9252 29450
rect 14336 29398 14388 29450
rect 14400 29398 14452 29450
rect 14464 29398 14516 29450
rect 14528 29398 14580 29450
rect 19664 29398 19716 29450
rect 19728 29398 19780 29450
rect 19792 29398 19844 29450
rect 19856 29398 19908 29450
rect 24992 29398 25044 29450
rect 25056 29398 25108 29450
rect 25120 29398 25172 29450
rect 25184 29398 25236 29450
rect 30320 29398 30372 29450
rect 30384 29398 30436 29450
rect 30448 29398 30500 29450
rect 30512 29398 30564 29450
rect 35648 29398 35700 29450
rect 35712 29398 35764 29450
rect 35776 29398 35828 29450
rect 35840 29398 35892 29450
rect 40976 29398 41028 29450
rect 41040 29398 41092 29450
rect 41104 29398 41156 29450
rect 41168 29398 41220 29450
rect 46304 29398 46356 29450
rect 46368 29398 46420 29450
rect 46432 29398 46484 29450
rect 46496 29398 46548 29450
rect 51632 29398 51684 29450
rect 51696 29398 51748 29450
rect 51760 29398 51812 29450
rect 51824 29398 51876 29450
rect 56960 29398 57012 29450
rect 57024 29398 57076 29450
rect 57088 29398 57140 29450
rect 57152 29398 57204 29450
rect 62288 29398 62340 29450
rect 62352 29398 62404 29450
rect 62416 29398 62468 29450
rect 62480 29398 62532 29450
rect 67616 29398 67668 29450
rect 67680 29398 67732 29450
rect 67744 29398 67796 29450
rect 67808 29398 67860 29450
rect 72944 29398 72996 29450
rect 73008 29398 73060 29450
rect 73072 29398 73124 29450
rect 73136 29398 73188 29450
rect 78272 29398 78324 29450
rect 78336 29398 78388 29450
rect 78400 29398 78452 29450
rect 78464 29398 78516 29450
rect 83600 29398 83652 29450
rect 83664 29398 83716 29450
rect 83728 29398 83780 29450
rect 83792 29398 83844 29450
rect 88928 29398 88980 29450
rect 88992 29398 89044 29450
rect 89056 29398 89108 29450
rect 89120 29398 89172 29450
rect 3042 29339 3094 29348
rect 3042 29305 3051 29339
rect 3051 29305 3085 29339
rect 3085 29305 3094 29339
rect 3042 29296 3094 29305
rect 8010 29296 8062 29348
rect 8286 29339 8338 29348
rect 8286 29305 8295 29339
rect 8295 29305 8329 29339
rect 8329 29305 8338 29339
rect 8286 29296 8338 29305
rect 9390 29296 9442 29348
rect 10402 29296 10454 29348
rect 12886 29296 12938 29348
rect 4698 29228 4750 29280
rect 6446 29203 6498 29212
rect 6446 29169 6455 29203
rect 6455 29169 6489 29203
rect 6489 29169 6498 29203
rect 6446 29160 6498 29169
rect 7734 29160 7786 29212
rect 8194 29160 8246 29212
rect 10126 29160 10178 29212
rect 3042 29092 3094 29144
rect 6354 29092 6406 29144
rect 6906 29092 6958 29144
rect 8102 29135 8154 29144
rect 8102 29101 8111 29135
rect 8111 29101 8145 29135
rect 8145 29101 8154 29135
rect 8102 29092 8154 29101
rect 9482 29024 9534 29076
rect 10954 29067 11006 29076
rect 10954 29033 10963 29067
rect 10963 29033 10997 29067
rect 10997 29033 11006 29067
rect 10954 29024 11006 29033
rect 13530 29296 13582 29348
rect 19326 29296 19378 29348
rect 19970 29296 20022 29348
rect 23006 29296 23058 29348
rect 23466 29339 23518 29348
rect 23466 29305 23475 29339
rect 23475 29305 23509 29339
rect 23509 29305 23518 29339
rect 23466 29296 23518 29305
rect 23742 29296 23794 29348
rect 24846 29296 24898 29348
rect 36346 29339 36398 29348
rect 18774 29228 18826 29280
rect 18958 29271 19010 29280
rect 18958 29237 18967 29271
rect 18967 29237 19001 29271
rect 19001 29237 19010 29271
rect 18958 29228 19010 29237
rect 28158 29228 28210 29280
rect 28894 29271 28946 29280
rect 28894 29237 28903 29271
rect 28903 29237 28937 29271
rect 28937 29237 28946 29271
rect 28894 29228 28946 29237
rect 28986 29228 29038 29280
rect 32298 29228 32350 29280
rect 34138 29228 34190 29280
rect 36346 29305 36355 29339
rect 36355 29305 36389 29339
rect 36389 29305 36398 29339
rect 36346 29296 36398 29305
rect 37726 29339 37778 29348
rect 37726 29305 37735 29339
rect 37735 29305 37769 29339
rect 37769 29305 37778 29339
rect 37726 29296 37778 29305
rect 37818 29296 37870 29348
rect 42234 29296 42286 29348
rect 44074 29296 44126 29348
rect 47294 29296 47346 29348
rect 48122 29296 48174 29348
rect 48306 29339 48358 29348
rect 48306 29305 48315 29339
rect 48315 29305 48349 29339
rect 48349 29305 48358 29339
rect 48306 29296 48358 29305
rect 48398 29296 48450 29348
rect 48582 29296 48634 29348
rect 50882 29296 50934 29348
rect 50974 29296 51026 29348
rect 54102 29296 54154 29348
rect 54286 29296 54338 29348
rect 60358 29296 60410 29348
rect 60726 29296 60778 29348
rect 62934 29296 62986 29348
rect 67258 29296 67310 29348
rect 68086 29296 68138 29348
rect 36254 29228 36306 29280
rect 16106 29160 16158 29212
rect 22730 29160 22782 29212
rect 17486 29135 17538 29144
rect 17486 29101 17495 29135
rect 17495 29101 17529 29135
rect 17529 29101 17538 29135
rect 17486 29092 17538 29101
rect 18774 29092 18826 29144
rect 23006 29092 23058 29144
rect 23190 29135 23242 29144
rect 23190 29101 23199 29135
rect 23199 29101 23233 29135
rect 23233 29101 23242 29135
rect 23190 29092 23242 29101
rect 23374 29160 23426 29212
rect 24018 29160 24070 29212
rect 24202 29160 24254 29212
rect 28710 29160 28762 29212
rect 23742 29092 23794 29144
rect 24662 29092 24714 29144
rect 28526 29092 28578 29144
rect 29078 29135 29130 29144
rect 29078 29101 29087 29135
rect 29087 29101 29121 29135
rect 29121 29101 29130 29135
rect 29078 29092 29130 29101
rect 29538 29160 29590 29212
rect 30182 29160 30234 29212
rect 32022 29203 32074 29212
rect 29998 29092 30050 29144
rect 30458 29135 30510 29144
rect 30458 29101 30467 29135
rect 30467 29101 30501 29135
rect 30501 29101 30510 29135
rect 30458 29092 30510 29101
rect 30826 29135 30878 29144
rect 30826 29101 30835 29135
rect 30835 29101 30869 29135
rect 30869 29101 30878 29135
rect 30826 29092 30878 29101
rect 32022 29169 32031 29203
rect 32031 29169 32065 29203
rect 32065 29169 32074 29203
rect 32022 29160 32074 29169
rect 37266 29228 37318 29280
rect 38646 29228 38698 29280
rect 31286 29092 31338 29144
rect 33954 29092 34006 29144
rect 35886 29092 35938 29144
rect 36162 29092 36214 29144
rect 36714 29135 36766 29144
rect 36714 29101 36723 29135
rect 36723 29101 36757 29135
rect 36757 29101 36766 29135
rect 36714 29092 36766 29101
rect 37818 29160 37870 29212
rect 37266 29135 37318 29144
rect 37266 29101 37275 29135
rect 37275 29101 37309 29135
rect 37309 29101 37318 29135
rect 37266 29092 37318 29101
rect 38830 29092 38882 29144
rect 41774 29135 41826 29144
rect 41774 29101 41783 29135
rect 41783 29101 41817 29135
rect 41817 29101 41826 29135
rect 41774 29092 41826 29101
rect 42234 29135 42286 29144
rect 42234 29101 42243 29135
rect 42243 29101 42277 29135
rect 42277 29101 42286 29135
rect 42234 29092 42286 29101
rect 42326 29135 42378 29144
rect 42326 29101 42335 29135
rect 42335 29101 42369 29135
rect 42369 29101 42378 29135
rect 42326 29092 42378 29101
rect 42970 29092 43022 29144
rect 44994 29228 45046 29280
rect 45822 29271 45874 29280
rect 45822 29237 45831 29271
rect 45831 29237 45865 29271
rect 45865 29237 45874 29271
rect 45822 29228 45874 29237
rect 46006 29228 46058 29280
rect 45454 29160 45506 29212
rect 46834 29203 46886 29212
rect 46834 29169 46843 29203
rect 46843 29169 46877 29203
rect 46877 29169 46886 29203
rect 46834 29160 46886 29169
rect 47294 29135 47346 29144
rect 47294 29101 47303 29135
rect 47303 29101 47337 29135
rect 47337 29101 47346 29135
rect 48306 29160 48358 29212
rect 48490 29160 48542 29212
rect 47294 29092 47346 29101
rect 48674 29092 48726 29144
rect 52354 29160 52406 29212
rect 51158 29135 51210 29144
rect 51158 29101 51167 29135
rect 51167 29101 51201 29135
rect 51201 29101 51210 29135
rect 51158 29092 51210 29101
rect 51802 29092 51854 29144
rect 54286 29203 54338 29212
rect 54286 29169 54295 29203
rect 54295 29169 54329 29203
rect 54329 29169 54338 29203
rect 54286 29160 54338 29169
rect 54930 29228 54982 29280
rect 60174 29228 60226 29280
rect 86394 29296 86446 29348
rect 86670 29339 86722 29348
rect 86670 29305 86679 29339
rect 86679 29305 86713 29339
rect 86713 29305 86722 29339
rect 86670 29296 86722 29305
rect 86762 29296 86814 29348
rect 90994 29339 91046 29348
rect 90994 29305 91003 29339
rect 91003 29305 91037 29339
rect 91037 29305 91046 29339
rect 90994 29296 91046 29305
rect 52538 29092 52590 29144
rect 53642 29135 53694 29144
rect 53642 29101 53651 29135
rect 53651 29101 53685 29135
rect 53685 29101 53694 29135
rect 53642 29092 53694 29101
rect 54102 29092 54154 29144
rect 54378 29092 54430 29144
rect 2306 28956 2358 29008
rect 2950 28956 3002 29008
rect 6722 28999 6774 29008
rect 6722 28965 6731 28999
rect 6731 28965 6765 28999
rect 6765 28965 6774 28999
rect 6722 28956 6774 28965
rect 11322 28956 11374 29008
rect 17578 28999 17630 29008
rect 17578 28965 17587 28999
rect 17587 28965 17621 28999
rect 17621 28965 17630 28999
rect 33218 29024 33270 29076
rect 37726 29024 37778 29076
rect 38278 29024 38330 29076
rect 45362 29024 45414 29076
rect 45546 29067 45598 29076
rect 45546 29033 45555 29067
rect 45555 29033 45589 29067
rect 45589 29033 45598 29067
rect 45546 29024 45598 29033
rect 52630 29024 52682 29076
rect 55298 29092 55350 29144
rect 17578 28956 17630 28965
rect 19326 28956 19378 29008
rect 24662 28956 24714 29008
rect 24754 28999 24806 29008
rect 24754 28965 24763 28999
rect 24763 28965 24797 28999
rect 24797 28965 24806 28999
rect 30274 28999 30326 29008
rect 24754 28956 24806 28965
rect 30274 28965 30283 28999
rect 30283 28965 30317 28999
rect 30317 28965 30326 28999
rect 30274 28956 30326 28965
rect 30366 28956 30418 29008
rect 34046 28956 34098 29008
rect 35426 28956 35478 29008
rect 36714 28956 36766 29008
rect 38186 28956 38238 29008
rect 39014 28956 39066 29008
rect 42326 28956 42378 29008
rect 43430 28956 43482 29008
rect 48674 28999 48726 29008
rect 48674 28965 48683 28999
rect 48683 28965 48717 28999
rect 48717 28965 48726 28999
rect 48674 28956 48726 28965
rect 49686 28956 49738 29008
rect 49962 28956 50014 29008
rect 53826 28956 53878 29008
rect 57506 29024 57558 29076
rect 58610 29160 58662 29212
rect 59438 29160 59490 29212
rect 61830 29160 61882 29212
rect 58886 29135 58938 29144
rect 58886 29101 58895 29135
rect 58895 29101 58929 29135
rect 58929 29101 58938 29135
rect 58886 29092 58938 29101
rect 59162 29092 59214 29144
rect 60450 29135 60502 29144
rect 59438 29024 59490 29076
rect 60450 29101 60459 29135
rect 60459 29101 60493 29135
rect 60493 29101 60502 29135
rect 60450 29092 60502 29101
rect 60726 29024 60778 29076
rect 58886 28956 58938 29008
rect 62842 29092 62894 29144
rect 67442 29160 67494 29212
rect 69098 29203 69150 29212
rect 69098 29169 69107 29203
rect 69107 29169 69141 29203
rect 69141 29169 69150 29203
rect 69098 29160 69150 29169
rect 69466 29228 69518 29280
rect 65326 29092 65378 29144
rect 67902 29092 67954 29144
rect 68178 29092 68230 29144
rect 68638 29135 68690 29144
rect 68638 29101 68647 29135
rect 68647 29101 68681 29135
rect 68681 29101 68690 29135
rect 68638 29092 68690 29101
rect 69006 29135 69058 29144
rect 62106 29024 62158 29076
rect 64498 29024 64550 29076
rect 69006 29101 69015 29135
rect 69015 29101 69049 29135
rect 69049 29101 69058 29135
rect 69006 29092 69058 29101
rect 69558 29092 69610 29144
rect 62658 28956 62710 29008
rect 63210 28999 63262 29008
rect 63210 28965 63219 28999
rect 63219 28965 63253 28999
rect 63253 28965 63262 28999
rect 63210 28956 63262 28965
rect 64406 28999 64458 29008
rect 64406 28965 64415 28999
rect 64415 28965 64449 28999
rect 64449 28965 64458 28999
rect 64406 28956 64458 28965
rect 69190 28956 69242 29008
rect 69466 29024 69518 29076
rect 71122 29135 71174 29144
rect 71122 29101 71131 29135
rect 71131 29101 71165 29135
rect 71165 29101 71174 29135
rect 74986 29160 75038 29212
rect 76918 29228 76970 29280
rect 84922 29271 84974 29280
rect 78942 29160 78994 29212
rect 84922 29237 84931 29271
rect 84931 29237 84965 29271
rect 84965 29237 84974 29271
rect 84922 29228 84974 29237
rect 85842 29228 85894 29280
rect 91086 29160 91138 29212
rect 71122 29092 71174 29101
rect 74250 29092 74302 29144
rect 77746 29135 77798 29144
rect 74618 29067 74670 29076
rect 74618 29033 74627 29067
rect 74627 29033 74661 29067
rect 74661 29033 74670 29067
rect 77746 29101 77755 29135
rect 77755 29101 77789 29135
rect 77789 29101 77798 29135
rect 77746 29092 77798 29101
rect 79862 29135 79914 29144
rect 79862 29101 79871 29135
rect 79871 29101 79905 29135
rect 79905 29101 79914 29135
rect 79862 29092 79914 29101
rect 81242 29135 81294 29144
rect 81242 29101 81251 29135
rect 81251 29101 81285 29135
rect 81285 29101 81294 29135
rect 81242 29092 81294 29101
rect 84830 29092 84882 29144
rect 74618 29024 74670 29033
rect 80138 29024 80190 29076
rect 80322 29024 80374 29076
rect 81426 29024 81478 29076
rect 84094 29024 84146 29076
rect 84554 29067 84606 29076
rect 84554 29033 84563 29067
rect 84563 29033 84597 29067
rect 84597 29033 84606 29067
rect 86762 29092 86814 29144
rect 90810 29135 90862 29144
rect 90810 29101 90819 29135
rect 90819 29101 90853 29135
rect 90853 29101 90862 29135
rect 90810 29092 90862 29101
rect 91454 29092 91506 29144
rect 91914 29092 91966 29144
rect 84554 29024 84606 29033
rect 87774 29024 87826 29076
rect 90718 29067 90770 29076
rect 90718 29033 90727 29067
rect 90727 29033 90761 29067
rect 90761 29033 90770 29067
rect 90718 29024 90770 29033
rect 73698 28999 73750 29008
rect 73698 28965 73707 28999
rect 73707 28965 73741 28999
rect 73741 28965 73750 28999
rect 77562 28999 77614 29008
rect 73698 28956 73750 28965
rect 77562 28965 77571 28999
rect 77571 28965 77605 28999
rect 77605 28965 77614 28999
rect 77562 28956 77614 28965
rect 79494 28956 79546 29008
rect 81334 28999 81386 29008
rect 81334 28965 81343 28999
rect 81343 28965 81377 28999
rect 81377 28965 81386 28999
rect 81334 28956 81386 28965
rect 90626 28956 90678 29008
rect 6344 28854 6396 28906
rect 6408 28854 6460 28906
rect 6472 28854 6524 28906
rect 6536 28854 6588 28906
rect 11672 28854 11724 28906
rect 11736 28854 11788 28906
rect 11800 28854 11852 28906
rect 11864 28854 11916 28906
rect 17000 28854 17052 28906
rect 17064 28854 17116 28906
rect 17128 28854 17180 28906
rect 17192 28854 17244 28906
rect 22328 28854 22380 28906
rect 22392 28854 22444 28906
rect 22456 28854 22508 28906
rect 22520 28854 22572 28906
rect 27656 28854 27708 28906
rect 27720 28854 27772 28906
rect 27784 28854 27836 28906
rect 27848 28854 27900 28906
rect 32984 28854 33036 28906
rect 33048 28854 33100 28906
rect 33112 28854 33164 28906
rect 33176 28854 33228 28906
rect 38312 28854 38364 28906
rect 38376 28854 38428 28906
rect 38440 28854 38492 28906
rect 38504 28854 38556 28906
rect 43640 28854 43692 28906
rect 43704 28854 43756 28906
rect 43768 28854 43820 28906
rect 43832 28854 43884 28906
rect 48968 28854 49020 28906
rect 49032 28854 49084 28906
rect 49096 28854 49148 28906
rect 49160 28854 49212 28906
rect 54296 28854 54348 28906
rect 54360 28854 54412 28906
rect 54424 28854 54476 28906
rect 54488 28854 54540 28906
rect 59624 28854 59676 28906
rect 59688 28854 59740 28906
rect 59752 28854 59804 28906
rect 59816 28854 59868 28906
rect 64952 28854 65004 28906
rect 65016 28854 65068 28906
rect 65080 28854 65132 28906
rect 65144 28854 65196 28906
rect 70280 28854 70332 28906
rect 70344 28854 70396 28906
rect 70408 28854 70460 28906
rect 70472 28854 70524 28906
rect 75608 28854 75660 28906
rect 75672 28854 75724 28906
rect 75736 28854 75788 28906
rect 75800 28854 75852 28906
rect 80936 28854 80988 28906
rect 81000 28854 81052 28906
rect 81064 28854 81116 28906
rect 81128 28854 81180 28906
rect 86264 28854 86316 28906
rect 86328 28854 86380 28906
rect 86392 28854 86444 28906
rect 86456 28854 86508 28906
rect 91592 28854 91644 28906
rect 91656 28854 91708 28906
rect 91720 28854 91772 28906
rect 91784 28854 91836 28906
rect 6722 28795 6774 28804
rect 6722 28761 6731 28795
rect 6731 28761 6765 28795
rect 6765 28761 6774 28795
rect 6722 28752 6774 28761
rect 6170 28616 6222 28668
rect 9298 28752 9350 28804
rect 9482 28727 9534 28736
rect 9482 28693 9491 28727
rect 9491 28693 9525 28727
rect 9525 28693 9534 28727
rect 9482 28684 9534 28693
rect 10954 28684 11006 28736
rect 12978 28727 13030 28736
rect 8102 28616 8154 28668
rect 9390 28659 9442 28668
rect 9390 28625 9399 28659
rect 9399 28625 9433 28659
rect 9433 28625 9442 28659
rect 11506 28659 11558 28668
rect 9390 28616 9442 28625
rect 11506 28625 11515 28659
rect 11515 28625 11549 28659
rect 11549 28625 11558 28659
rect 11506 28616 11558 28625
rect 12978 28693 12987 28727
rect 12987 28693 13021 28727
rect 13021 28693 13030 28727
rect 12978 28684 13030 28693
rect 12058 28659 12110 28668
rect 12058 28625 12067 28659
rect 12067 28625 12101 28659
rect 12101 28625 12110 28659
rect 12058 28616 12110 28625
rect 13530 28752 13582 28804
rect 17302 28752 17354 28804
rect 17854 28752 17906 28804
rect 24662 28752 24714 28804
rect 16658 28684 16710 28736
rect 14726 28659 14778 28668
rect 10954 28548 11006 28600
rect 5986 28480 6038 28532
rect 11322 28480 11374 28532
rect 11506 28480 11558 28532
rect 14726 28625 14735 28659
rect 14735 28625 14769 28659
rect 14769 28625 14778 28659
rect 14726 28616 14778 28625
rect 15922 28616 15974 28668
rect 16750 28548 16802 28600
rect 18590 28684 18642 28736
rect 25490 28684 25542 28736
rect 25766 28727 25818 28736
rect 17302 28616 17354 28668
rect 17670 28548 17722 28600
rect 15094 28412 15146 28464
rect 16106 28412 16158 28464
rect 16290 28455 16342 28464
rect 16290 28421 16299 28455
rect 16299 28421 16333 28455
rect 16333 28421 16342 28455
rect 16290 28412 16342 28421
rect 18958 28659 19010 28668
rect 18958 28625 18967 28659
rect 18967 28625 19001 28659
rect 19001 28625 19010 28659
rect 18958 28616 19010 28625
rect 22730 28659 22782 28668
rect 22730 28625 22739 28659
rect 22739 28625 22773 28659
rect 22773 28625 22782 28659
rect 23466 28659 23518 28668
rect 22730 28616 22782 28625
rect 23098 28591 23150 28600
rect 23098 28557 23107 28591
rect 23107 28557 23141 28591
rect 23141 28557 23150 28591
rect 23098 28548 23150 28557
rect 23466 28625 23475 28659
rect 23475 28625 23509 28659
rect 23509 28625 23518 28659
rect 23466 28616 23518 28625
rect 23834 28659 23886 28668
rect 23834 28625 23843 28659
rect 23843 28625 23877 28659
rect 23877 28625 23886 28659
rect 23834 28616 23886 28625
rect 23742 28548 23794 28600
rect 18222 28480 18274 28532
rect 20982 28480 21034 28532
rect 24846 28616 24898 28668
rect 25766 28693 25775 28727
rect 25775 28693 25809 28727
rect 25809 28693 25818 28727
rect 25766 28684 25818 28693
rect 26502 28684 26554 28736
rect 27146 28616 27198 28668
rect 27422 28684 27474 28736
rect 28342 28684 28394 28736
rect 28526 28752 28578 28804
rect 30366 28752 30418 28804
rect 30458 28752 30510 28804
rect 34046 28752 34098 28804
rect 34506 28752 34558 28804
rect 37726 28752 37778 28804
rect 42878 28795 42930 28804
rect 42878 28761 42887 28795
rect 42887 28761 42921 28795
rect 42921 28761 42930 28795
rect 42878 28752 42930 28761
rect 36162 28727 36214 28736
rect 36162 28693 36171 28727
rect 36171 28693 36205 28727
rect 36205 28693 36214 28727
rect 36162 28684 36214 28693
rect 36254 28684 36306 28736
rect 39566 28684 39618 28736
rect 43062 28684 43114 28736
rect 22638 28412 22690 28464
rect 23742 28412 23794 28464
rect 26502 28480 26554 28532
rect 27698 28548 27750 28600
rect 28710 28616 28762 28668
rect 29814 28659 29866 28668
rect 29814 28625 29823 28659
rect 29823 28625 29857 28659
rect 29857 28625 29866 28659
rect 29814 28616 29866 28625
rect 30090 28616 30142 28668
rect 31562 28659 31614 28668
rect 27882 28548 27934 28600
rect 29538 28548 29590 28600
rect 29722 28548 29774 28600
rect 30274 28591 30326 28600
rect 30274 28557 30283 28591
rect 30283 28557 30317 28591
rect 30317 28557 30326 28591
rect 30274 28548 30326 28557
rect 31562 28625 31571 28659
rect 31571 28625 31605 28659
rect 31605 28625 31614 28659
rect 31562 28616 31614 28625
rect 32022 28616 32074 28668
rect 33954 28548 34006 28600
rect 34414 28591 34466 28600
rect 34414 28557 34423 28591
rect 34423 28557 34457 28591
rect 34457 28557 34466 28591
rect 34414 28548 34466 28557
rect 35426 28548 35478 28600
rect 35518 28548 35570 28600
rect 37450 28548 37502 28600
rect 38554 28591 38606 28600
rect 38554 28557 38563 28591
rect 38563 28557 38597 28591
rect 38597 28557 38606 28591
rect 38554 28548 38606 28557
rect 38830 28616 38882 28668
rect 39198 28659 39250 28668
rect 39198 28625 39207 28659
rect 39207 28625 39241 28659
rect 39241 28625 39250 28659
rect 39198 28616 39250 28625
rect 39474 28616 39526 28668
rect 40670 28616 40722 28668
rect 43798 28684 43850 28736
rect 27974 28480 28026 28532
rect 31102 28480 31154 28532
rect 35886 28480 35938 28532
rect 36898 28480 36950 28532
rect 39842 28480 39894 28532
rect 43522 28616 43574 28668
rect 45546 28752 45598 28804
rect 54930 28752 54982 28804
rect 56402 28795 56454 28804
rect 49318 28659 49370 28668
rect 49318 28625 49327 28659
rect 49327 28625 49361 28659
rect 49361 28625 49370 28659
rect 49318 28616 49370 28625
rect 47938 28548 47990 28600
rect 49686 28659 49738 28668
rect 49686 28625 49695 28659
rect 49695 28625 49729 28659
rect 49729 28625 49738 28659
rect 49686 28616 49738 28625
rect 50054 28616 50106 28668
rect 50330 28684 50382 28736
rect 56402 28761 56411 28795
rect 56411 28761 56445 28795
rect 56445 28761 56454 28795
rect 56402 28752 56454 28761
rect 56586 28684 56638 28736
rect 62750 28684 62802 28736
rect 64406 28684 64458 28736
rect 67902 28752 67954 28804
rect 67994 28752 68046 28804
rect 69006 28752 69058 28804
rect 69466 28684 69518 28736
rect 51894 28616 51946 28668
rect 52078 28659 52130 28668
rect 52078 28625 52087 28659
rect 52087 28625 52121 28659
rect 52121 28625 52130 28659
rect 52078 28616 52130 28625
rect 52814 28659 52866 28668
rect 51802 28548 51854 28600
rect 50422 28480 50474 28532
rect 50882 28523 50934 28532
rect 50882 28489 50891 28523
rect 50891 28489 50925 28523
rect 50925 28489 50934 28523
rect 50882 28480 50934 28489
rect 25398 28455 25450 28464
rect 25398 28421 25407 28455
rect 25407 28421 25441 28455
rect 25441 28421 25450 28455
rect 25398 28412 25450 28421
rect 25490 28412 25542 28464
rect 28342 28455 28394 28464
rect 28342 28421 28351 28455
rect 28351 28421 28385 28455
rect 28385 28421 28394 28455
rect 28342 28412 28394 28421
rect 28526 28412 28578 28464
rect 29722 28412 29774 28464
rect 30826 28412 30878 28464
rect 31010 28412 31062 28464
rect 38370 28455 38422 28464
rect 38370 28421 38379 28455
rect 38379 28421 38413 28455
rect 38413 28421 38422 28455
rect 38370 28412 38422 28421
rect 39198 28412 39250 28464
rect 39750 28455 39802 28464
rect 39750 28421 39759 28455
rect 39759 28421 39793 28455
rect 39793 28421 39802 28455
rect 39750 28412 39802 28421
rect 42878 28412 42930 28464
rect 45270 28412 45322 28464
rect 47754 28412 47806 28464
rect 48858 28412 48910 28464
rect 52354 28548 52406 28600
rect 52814 28625 52823 28659
rect 52823 28625 52857 28659
rect 52857 28625 52866 28659
rect 52814 28616 52866 28625
rect 53826 28616 53878 28668
rect 54194 28616 54246 28668
rect 55298 28659 55350 28668
rect 55298 28625 55307 28659
rect 55307 28625 55341 28659
rect 55341 28625 55350 28659
rect 55298 28616 55350 28625
rect 57506 28659 57558 28668
rect 57506 28625 57515 28659
rect 57515 28625 57549 28659
rect 57549 28625 57558 28659
rect 57506 28616 57558 28625
rect 59530 28616 59582 28668
rect 52998 28591 53050 28600
rect 52998 28557 53007 28591
rect 53007 28557 53041 28591
rect 53041 28557 53050 28591
rect 52998 28548 53050 28557
rect 53826 28480 53878 28532
rect 53642 28412 53694 28464
rect 54286 28548 54338 28600
rect 56494 28548 56546 28600
rect 63210 28616 63262 28668
rect 63302 28616 63354 28668
rect 67166 28659 67218 28668
rect 67166 28625 67175 28659
rect 67175 28625 67209 28659
rect 67209 28625 67218 28659
rect 67166 28616 67218 28625
rect 69374 28659 69426 28668
rect 69374 28625 69383 28659
rect 69383 28625 69417 28659
rect 69417 28625 69426 28659
rect 69374 28616 69426 28625
rect 61186 28548 61238 28600
rect 64222 28548 64274 28600
rect 74618 28752 74670 28804
rect 81242 28752 81294 28804
rect 84186 28752 84238 28804
rect 89246 28752 89298 28804
rect 90718 28752 90770 28804
rect 73238 28727 73290 28736
rect 73238 28693 73247 28727
rect 73247 28693 73281 28727
rect 73281 28693 73290 28727
rect 73238 28684 73290 28693
rect 71674 28616 71726 28668
rect 73882 28684 73934 28736
rect 73606 28659 73658 28668
rect 73606 28625 73615 28659
rect 73615 28625 73649 28659
rect 73649 28625 73658 28659
rect 73606 28616 73658 28625
rect 79218 28616 79270 28668
rect 79494 28659 79546 28668
rect 79494 28625 79503 28659
rect 79503 28625 79537 28659
rect 79537 28625 79546 28659
rect 79494 28616 79546 28625
rect 90074 28659 90126 28668
rect 90074 28625 90083 28659
rect 90083 28625 90117 28659
rect 90117 28625 90126 28659
rect 90074 28616 90126 28625
rect 90350 28659 90402 28668
rect 90350 28625 90359 28659
rect 90359 28625 90393 28659
rect 90393 28625 90402 28659
rect 90350 28616 90402 28625
rect 91086 28616 91138 28668
rect 91822 28659 91874 28668
rect 91822 28625 91831 28659
rect 91831 28625 91865 28659
rect 91865 28625 91874 28659
rect 91822 28616 91874 28625
rect 74066 28591 74118 28600
rect 74066 28557 74075 28591
rect 74075 28557 74109 28591
rect 74109 28557 74118 28591
rect 74066 28548 74118 28557
rect 80414 28548 80466 28600
rect 84554 28591 84606 28600
rect 62658 28523 62710 28532
rect 62658 28489 62667 28523
rect 62667 28489 62701 28523
rect 62701 28489 62710 28523
rect 62658 28480 62710 28489
rect 57598 28412 57650 28464
rect 59806 28455 59858 28464
rect 59806 28421 59815 28455
rect 59815 28421 59849 28455
rect 59849 28421 59858 28455
rect 59806 28412 59858 28421
rect 64774 28480 64826 28532
rect 69742 28480 69794 28532
rect 64130 28412 64182 28464
rect 72686 28412 72738 28464
rect 84554 28557 84563 28591
rect 84563 28557 84597 28591
rect 84597 28557 84606 28591
rect 84554 28548 84606 28557
rect 90626 28480 90678 28532
rect 85198 28412 85250 28464
rect 85566 28412 85618 28464
rect 3680 28310 3732 28362
rect 3744 28310 3796 28362
rect 3808 28310 3860 28362
rect 3872 28310 3924 28362
rect 9008 28310 9060 28362
rect 9072 28310 9124 28362
rect 9136 28310 9188 28362
rect 9200 28310 9252 28362
rect 14336 28310 14388 28362
rect 14400 28310 14452 28362
rect 14464 28310 14516 28362
rect 14528 28310 14580 28362
rect 19664 28310 19716 28362
rect 19728 28310 19780 28362
rect 19792 28310 19844 28362
rect 19856 28310 19908 28362
rect 24992 28310 25044 28362
rect 25056 28310 25108 28362
rect 25120 28310 25172 28362
rect 25184 28310 25236 28362
rect 30320 28310 30372 28362
rect 30384 28310 30436 28362
rect 30448 28310 30500 28362
rect 30512 28310 30564 28362
rect 35648 28310 35700 28362
rect 35712 28310 35764 28362
rect 35776 28310 35828 28362
rect 35840 28310 35892 28362
rect 40976 28310 41028 28362
rect 41040 28310 41092 28362
rect 41104 28310 41156 28362
rect 41168 28310 41220 28362
rect 46304 28310 46356 28362
rect 46368 28310 46420 28362
rect 46432 28310 46484 28362
rect 46496 28310 46548 28362
rect 51632 28310 51684 28362
rect 51696 28310 51748 28362
rect 51760 28310 51812 28362
rect 51824 28310 51876 28362
rect 56960 28310 57012 28362
rect 57024 28310 57076 28362
rect 57088 28310 57140 28362
rect 57152 28310 57204 28362
rect 62288 28310 62340 28362
rect 62352 28310 62404 28362
rect 62416 28310 62468 28362
rect 62480 28310 62532 28362
rect 67616 28310 67668 28362
rect 67680 28310 67732 28362
rect 67744 28310 67796 28362
rect 67808 28310 67860 28362
rect 72944 28310 72996 28362
rect 73008 28310 73060 28362
rect 73072 28310 73124 28362
rect 73136 28310 73188 28362
rect 78272 28310 78324 28362
rect 78336 28310 78388 28362
rect 78400 28310 78452 28362
rect 78464 28310 78516 28362
rect 83600 28310 83652 28362
rect 83664 28310 83716 28362
rect 83728 28310 83780 28362
rect 83792 28310 83844 28362
rect 88928 28310 88980 28362
rect 88992 28310 89044 28362
rect 89056 28310 89108 28362
rect 89120 28310 89172 28362
rect 3042 28251 3094 28260
rect 3042 28217 3051 28251
rect 3051 28217 3085 28251
rect 3085 28217 3094 28251
rect 3042 28208 3094 28217
rect 12886 28208 12938 28260
rect 13530 28251 13582 28260
rect 13530 28217 13539 28251
rect 13539 28217 13573 28251
rect 13573 28217 13582 28251
rect 13530 28208 13582 28217
rect 15094 28251 15146 28260
rect 15094 28217 15103 28251
rect 15103 28217 15137 28251
rect 15137 28217 15146 28251
rect 15094 28208 15146 28217
rect 15922 28208 15974 28260
rect 20982 28208 21034 28260
rect 8102 28140 8154 28192
rect 13254 28183 13306 28192
rect 926 28072 978 28124
rect 2306 28072 2358 28124
rect 6170 28072 6222 28124
rect 8562 28072 8614 28124
rect 11966 28072 12018 28124
rect 1938 28047 1990 28056
rect 1938 28013 1947 28047
rect 1947 28013 1981 28047
rect 1981 28013 1990 28047
rect 1938 28004 1990 28013
rect 7734 28004 7786 28056
rect 9482 28004 9534 28056
rect 10954 28004 11006 28056
rect 12242 28004 12294 28056
rect 12702 28047 12754 28056
rect 12702 28013 12711 28047
rect 12711 28013 12745 28047
rect 12745 28013 12754 28047
rect 12702 28004 12754 28013
rect 12886 28047 12938 28056
rect 12886 28013 12895 28047
rect 12895 28013 12929 28047
rect 12929 28013 12938 28047
rect 12886 28004 12938 28013
rect 4054 27868 4106 27920
rect 13254 28149 13263 28183
rect 13263 28149 13297 28183
rect 13297 28149 13306 28183
rect 13254 28140 13306 28149
rect 15186 28140 15238 28192
rect 15738 28004 15790 28056
rect 17394 28140 17446 28192
rect 16198 28072 16250 28124
rect 16658 28072 16710 28124
rect 17762 28115 17814 28124
rect 17762 28081 17771 28115
rect 17771 28081 17805 28115
rect 17805 28081 17814 28115
rect 17762 28072 17814 28081
rect 18222 28115 18274 28124
rect 18222 28081 18231 28115
rect 18231 28081 18265 28115
rect 18265 28081 18274 28115
rect 18222 28072 18274 28081
rect 19326 28115 19378 28124
rect 19326 28081 19335 28115
rect 19335 28081 19369 28115
rect 19369 28081 19378 28115
rect 19326 28072 19378 28081
rect 23926 28140 23978 28192
rect 27698 28183 27750 28192
rect 27698 28149 27707 28183
rect 27707 28149 27741 28183
rect 27741 28149 27750 28183
rect 27698 28140 27750 28149
rect 28342 28208 28394 28260
rect 35150 28208 35202 28260
rect 30734 28140 30786 28192
rect 24386 28072 24438 28124
rect 30642 28072 30694 28124
rect 35426 28183 35478 28192
rect 35426 28149 35435 28183
rect 35435 28149 35469 28183
rect 35469 28149 35478 28183
rect 35426 28140 35478 28149
rect 36898 28208 36950 28260
rect 40578 28208 40630 28260
rect 46098 28208 46150 28260
rect 38186 28140 38238 28192
rect 39198 28140 39250 28192
rect 16106 28004 16158 28056
rect 18866 28004 18918 28056
rect 20982 28047 21034 28056
rect 20982 28013 20991 28047
rect 20991 28013 21025 28047
rect 21025 28013 21034 28047
rect 20982 28004 21034 28013
rect 21350 28004 21402 28056
rect 23558 28004 23610 28056
rect 24018 28004 24070 28056
rect 24754 28004 24806 28056
rect 25858 28047 25910 28056
rect 25858 28013 25867 28047
rect 25867 28013 25901 28047
rect 25901 28013 25910 28047
rect 25858 28004 25910 28013
rect 29446 28004 29498 28056
rect 29538 28047 29590 28056
rect 29538 28013 29547 28047
rect 29547 28013 29581 28047
rect 29581 28013 29590 28047
rect 29722 28047 29774 28056
rect 29538 28004 29590 28013
rect 29722 28013 29731 28047
rect 29731 28013 29765 28047
rect 29765 28013 29774 28047
rect 29722 28004 29774 28013
rect 29906 28047 29958 28056
rect 29906 28013 29915 28047
rect 29915 28013 29949 28047
rect 29949 28013 29958 28047
rect 29906 28004 29958 28013
rect 29998 28004 30050 28056
rect 30182 28004 30234 28056
rect 30826 28047 30878 28056
rect 30826 28013 30835 28047
rect 30835 28013 30869 28047
rect 30869 28013 30878 28047
rect 30826 28004 30878 28013
rect 19050 27936 19102 27988
rect 8562 27868 8614 27920
rect 9298 27868 9350 27920
rect 14818 27868 14870 27920
rect 15370 27868 15422 27920
rect 17302 27868 17354 27920
rect 17394 27868 17446 27920
rect 20890 27868 20942 27920
rect 23282 27911 23334 27920
rect 23282 27877 23291 27911
rect 23291 27877 23325 27911
rect 23325 27877 23334 27911
rect 23282 27868 23334 27877
rect 23466 27936 23518 27988
rect 24110 27936 24162 27988
rect 31102 28004 31154 28056
rect 34046 28072 34098 28124
rect 34598 28072 34650 28124
rect 44994 28140 45046 28192
rect 49318 28208 49370 28260
rect 49962 28208 50014 28260
rect 50330 28208 50382 28260
rect 50422 28208 50474 28260
rect 52078 28208 52130 28260
rect 53826 28251 53878 28260
rect 53826 28217 53835 28251
rect 53835 28217 53869 28251
rect 53869 28217 53878 28251
rect 53826 28208 53878 28217
rect 53918 28208 53970 28260
rect 59806 28208 59858 28260
rect 63946 28251 63998 28260
rect 63946 28217 63955 28251
rect 63955 28217 63989 28251
rect 63989 28217 63998 28251
rect 63946 28208 63998 28217
rect 64222 28208 64274 28260
rect 74250 28208 74302 28260
rect 80414 28251 80466 28260
rect 80414 28217 80423 28251
rect 80423 28217 80457 28251
rect 80457 28217 80466 28251
rect 80414 28208 80466 28217
rect 90350 28208 90402 28260
rect 31378 28004 31430 28056
rect 33954 28047 34006 28056
rect 33954 28013 33963 28047
rect 33963 28013 33997 28047
rect 33997 28013 34006 28047
rect 33954 28004 34006 28013
rect 34230 28004 34282 28056
rect 35242 28047 35294 28056
rect 35242 28013 35251 28047
rect 35251 28013 35285 28047
rect 35285 28013 35294 28047
rect 35242 28004 35294 28013
rect 31194 27936 31246 27988
rect 35794 27936 35846 27988
rect 36162 28004 36214 28056
rect 38554 28004 38606 28056
rect 40670 28004 40722 28056
rect 36714 27936 36766 27988
rect 38370 27936 38422 27988
rect 38646 27936 38698 27988
rect 41774 28004 41826 28056
rect 42970 28072 43022 28124
rect 45822 28072 45874 28124
rect 43062 28047 43114 28056
rect 43062 28013 43071 28047
rect 43071 28013 43105 28047
rect 43105 28013 43114 28047
rect 43062 28004 43114 28013
rect 43430 28004 43482 28056
rect 42510 27936 42562 27988
rect 43798 28047 43850 28056
rect 43798 28013 43807 28047
rect 43807 28013 43841 28047
rect 43841 28013 43850 28047
rect 43798 28004 43850 28013
rect 44442 28004 44494 28056
rect 47846 28004 47898 28056
rect 48306 28072 48358 28124
rect 51526 28140 51578 28192
rect 57506 28140 57558 28192
rect 46282 27979 46334 27988
rect 46282 27945 46291 27979
rect 46291 27945 46325 27979
rect 46325 27945 46334 27979
rect 46282 27936 46334 27945
rect 25858 27868 25910 27920
rect 31286 27868 31338 27920
rect 31378 27868 31430 27920
rect 38738 27868 38790 27920
rect 42878 27911 42930 27920
rect 42878 27877 42887 27911
rect 42887 27877 42921 27911
rect 42921 27877 42930 27911
rect 42878 27868 42930 27877
rect 43246 27868 43298 27920
rect 48214 27868 48266 27920
rect 48398 27868 48450 27920
rect 50054 28047 50106 28056
rect 50054 28013 50063 28047
rect 50063 28013 50097 28047
rect 50097 28013 50106 28047
rect 50054 28004 50106 28013
rect 50790 28004 50842 28056
rect 52538 28072 52590 28124
rect 52906 28072 52958 28124
rect 57598 28072 57650 28124
rect 58426 28072 58478 28124
rect 52078 28004 52130 28056
rect 52354 28004 52406 28056
rect 53458 28004 53510 28056
rect 57414 28047 57466 28056
rect 57414 28013 57423 28047
rect 57423 28013 57457 28047
rect 57457 28013 57466 28047
rect 57414 28004 57466 28013
rect 50422 27979 50474 27988
rect 50422 27945 50431 27979
rect 50431 27945 50465 27979
rect 50465 27945 50474 27979
rect 50422 27936 50474 27945
rect 56862 27979 56914 27988
rect 51066 27868 51118 27920
rect 51250 27868 51302 27920
rect 53366 27911 53418 27920
rect 53366 27877 53375 27911
rect 53375 27877 53409 27911
rect 53409 27877 53418 27911
rect 56862 27945 56871 27979
rect 56871 27945 56905 27979
rect 56905 27945 56914 27979
rect 56862 27936 56914 27945
rect 56954 27936 57006 27988
rect 58334 28004 58386 28056
rect 65878 28140 65930 28192
rect 62658 28047 62710 28056
rect 62658 28013 62667 28047
rect 62667 28013 62701 28047
rect 62701 28013 62710 28047
rect 62658 28004 62710 28013
rect 62934 28047 62986 28056
rect 62934 28013 62943 28047
rect 62943 28013 62977 28047
rect 62977 28013 62986 28047
rect 62934 28004 62986 28013
rect 64130 27979 64182 27988
rect 53366 27868 53418 27877
rect 64130 27945 64139 27979
rect 64139 27945 64173 27979
rect 64173 27945 64182 27979
rect 64130 27936 64182 27945
rect 58794 27868 58846 27920
rect 71030 28140 71082 28192
rect 73330 28140 73382 28192
rect 79126 28140 79178 28192
rect 81242 28140 81294 28192
rect 67994 28072 68046 28124
rect 73606 28072 73658 28124
rect 74066 28072 74118 28124
rect 79770 28072 79822 28124
rect 83174 28183 83226 28192
rect 83174 28149 83183 28183
rect 83183 28149 83217 28183
rect 83217 28149 83226 28183
rect 83174 28140 83226 28149
rect 69558 28047 69610 28056
rect 69558 28013 69567 28047
rect 69567 28013 69601 28047
rect 69601 28013 69610 28047
rect 69558 28004 69610 28013
rect 69742 28047 69794 28056
rect 69742 28013 69751 28047
rect 69751 28013 69785 28047
rect 69785 28013 69794 28047
rect 69742 28004 69794 28013
rect 72686 28047 72738 28056
rect 68638 27936 68690 27988
rect 70110 27979 70162 27988
rect 70110 27945 70119 27979
rect 70119 27945 70153 27979
rect 70153 27945 70162 27979
rect 72686 28013 72695 28047
rect 72695 28013 72729 28047
rect 72729 28013 72738 28047
rect 72686 28004 72738 28013
rect 73698 28004 73750 28056
rect 73790 28004 73842 28056
rect 77562 28004 77614 28056
rect 81334 28004 81386 28056
rect 84554 28072 84606 28124
rect 90074 28140 90126 28192
rect 87590 28072 87642 28124
rect 70110 27936 70162 27945
rect 73054 27936 73106 27988
rect 80138 27979 80190 27988
rect 80138 27945 80147 27979
rect 80147 27945 80181 27979
rect 80181 27945 80190 27979
rect 80138 27936 80190 27945
rect 81242 27936 81294 27988
rect 68270 27911 68322 27920
rect 68270 27877 68279 27911
rect 68279 27877 68313 27911
rect 68313 27877 68322 27911
rect 68270 27868 68322 27877
rect 79862 27868 79914 27920
rect 84922 28004 84974 28056
rect 85014 28004 85066 28056
rect 85750 28004 85802 28056
rect 86118 28047 86170 28056
rect 86118 28013 86127 28047
rect 86127 28013 86161 28047
rect 86161 28013 86170 28047
rect 86118 28004 86170 28013
rect 89338 28047 89390 28056
rect 89338 28013 89347 28047
rect 89347 28013 89381 28047
rect 89381 28013 89390 28047
rect 89614 28047 89666 28056
rect 89338 28004 89390 28013
rect 89614 28013 89623 28047
rect 89623 28013 89657 28047
rect 89657 28013 89666 28047
rect 89614 28004 89666 28013
rect 90350 28072 90402 28124
rect 91086 28047 91138 28056
rect 83266 27936 83318 27988
rect 86578 27936 86630 27988
rect 89246 27936 89298 27988
rect 91086 28013 91095 28047
rect 91095 28013 91129 28047
rect 91129 28013 91138 28047
rect 91086 28004 91138 28013
rect 6344 27766 6396 27818
rect 6408 27766 6460 27818
rect 6472 27766 6524 27818
rect 6536 27766 6588 27818
rect 11672 27766 11724 27818
rect 11736 27766 11788 27818
rect 11800 27766 11852 27818
rect 11864 27766 11916 27818
rect 17000 27766 17052 27818
rect 17064 27766 17116 27818
rect 17128 27766 17180 27818
rect 17192 27766 17244 27818
rect 22328 27766 22380 27818
rect 22392 27766 22444 27818
rect 22456 27766 22508 27818
rect 22520 27766 22572 27818
rect 27656 27766 27708 27818
rect 27720 27766 27772 27818
rect 27784 27766 27836 27818
rect 27848 27766 27900 27818
rect 32984 27766 33036 27818
rect 33048 27766 33100 27818
rect 33112 27766 33164 27818
rect 33176 27766 33228 27818
rect 38312 27766 38364 27818
rect 38376 27766 38428 27818
rect 38440 27766 38492 27818
rect 38504 27766 38556 27818
rect 43640 27766 43692 27818
rect 43704 27766 43756 27818
rect 43768 27766 43820 27818
rect 43832 27766 43884 27818
rect 48968 27766 49020 27818
rect 49032 27766 49084 27818
rect 49096 27766 49148 27818
rect 49160 27766 49212 27818
rect 54296 27766 54348 27818
rect 54360 27766 54412 27818
rect 54424 27766 54476 27818
rect 54488 27766 54540 27818
rect 59624 27766 59676 27818
rect 59688 27766 59740 27818
rect 59752 27766 59804 27818
rect 59816 27766 59868 27818
rect 64952 27766 65004 27818
rect 65016 27766 65068 27818
rect 65080 27766 65132 27818
rect 65144 27766 65196 27818
rect 70280 27766 70332 27818
rect 70344 27766 70396 27818
rect 70408 27766 70460 27818
rect 70472 27766 70524 27818
rect 75608 27766 75660 27818
rect 75672 27766 75724 27818
rect 75736 27766 75788 27818
rect 75800 27766 75852 27818
rect 80936 27766 80988 27818
rect 81000 27766 81052 27818
rect 81064 27766 81116 27818
rect 81128 27766 81180 27818
rect 86264 27766 86316 27818
rect 86328 27766 86380 27818
rect 86392 27766 86444 27818
rect 86456 27766 86508 27818
rect 91592 27766 91644 27818
rect 91656 27766 91708 27818
rect 91720 27766 91772 27818
rect 91784 27766 91836 27818
rect 1938 27664 1990 27716
rect 7734 27707 7786 27716
rect 7734 27673 7743 27707
rect 7743 27673 7777 27707
rect 7777 27673 7786 27707
rect 7734 27664 7786 27673
rect 8102 27707 8154 27716
rect 8102 27673 8111 27707
rect 8111 27673 8145 27707
rect 8145 27673 8154 27707
rect 8102 27664 8154 27673
rect 15370 27664 15422 27716
rect 926 27571 978 27580
rect 926 27537 935 27571
rect 935 27537 969 27571
rect 969 27537 978 27571
rect 926 27528 978 27537
rect 8562 27596 8614 27648
rect 15830 27664 15882 27716
rect 16658 27664 16710 27716
rect 17670 27664 17722 27716
rect 23098 27664 23150 27716
rect 23650 27664 23702 27716
rect 15738 27596 15790 27648
rect 17578 27596 17630 27648
rect 8102 27528 8154 27580
rect 4790 27392 4842 27444
rect 10310 27460 10362 27512
rect 11874 27571 11926 27580
rect 11874 27537 11883 27571
rect 11883 27537 11917 27571
rect 11917 27537 11926 27571
rect 11874 27528 11926 27537
rect 12242 27528 12294 27580
rect 12610 27528 12662 27580
rect 15646 27571 15698 27580
rect 15646 27537 15655 27571
rect 15655 27537 15689 27571
rect 15689 27537 15698 27571
rect 15646 27528 15698 27537
rect 2950 27367 3002 27376
rect 2950 27333 2959 27367
rect 2959 27333 2993 27367
rect 2993 27333 3002 27367
rect 2950 27324 3002 27333
rect 4238 27324 4290 27376
rect 9298 27392 9350 27444
rect 12426 27392 12478 27444
rect 13162 27392 13214 27444
rect 15186 27392 15238 27444
rect 16106 27571 16158 27580
rect 16106 27537 16115 27571
rect 16115 27537 16149 27571
rect 16149 27537 16158 27571
rect 16474 27571 16526 27580
rect 16106 27528 16158 27537
rect 16474 27537 16483 27571
rect 16483 27537 16517 27571
rect 16517 27537 16526 27571
rect 16474 27528 16526 27537
rect 16566 27571 16618 27580
rect 16566 27537 16575 27571
rect 16575 27537 16609 27571
rect 16609 27537 16618 27571
rect 16566 27528 16618 27537
rect 18590 27528 18642 27580
rect 18774 27571 18826 27580
rect 18774 27537 18783 27571
rect 18783 27537 18817 27571
rect 18817 27537 18826 27571
rect 23926 27596 23978 27648
rect 18774 27528 18826 27537
rect 22546 27571 22598 27580
rect 22546 27537 22555 27571
rect 22555 27537 22589 27571
rect 22589 27537 22598 27571
rect 22546 27528 22598 27537
rect 22638 27528 22690 27580
rect 24570 27664 24622 27716
rect 24754 27707 24806 27716
rect 24754 27673 24763 27707
rect 24763 27673 24797 27707
rect 24797 27673 24806 27707
rect 24754 27664 24806 27673
rect 24110 27528 24162 27580
rect 25214 27596 25266 27648
rect 27146 27596 27198 27648
rect 29814 27664 29866 27716
rect 30642 27664 30694 27716
rect 38646 27664 38698 27716
rect 38830 27664 38882 27716
rect 42510 27707 42562 27716
rect 42510 27673 42519 27707
rect 42519 27673 42553 27707
rect 42553 27673 42562 27707
rect 42510 27664 42562 27673
rect 42786 27664 42838 27716
rect 43522 27664 43574 27716
rect 44350 27664 44402 27716
rect 48214 27664 48266 27716
rect 30366 27596 30418 27648
rect 31562 27596 31614 27648
rect 33770 27596 33822 27648
rect 36990 27596 37042 27648
rect 17670 27460 17722 27512
rect 20890 27460 20942 27512
rect 23374 27460 23426 27512
rect 23650 27503 23702 27512
rect 23650 27469 23659 27503
rect 23659 27469 23693 27503
rect 23693 27469 23702 27503
rect 23650 27460 23702 27469
rect 23834 27460 23886 27512
rect 19142 27392 19194 27444
rect 27422 27528 27474 27580
rect 28802 27528 28854 27580
rect 29722 27528 29774 27580
rect 31838 27528 31890 27580
rect 24754 27460 24806 27512
rect 27054 27503 27106 27512
rect 27054 27469 27063 27503
rect 27063 27469 27097 27503
rect 27097 27469 27106 27503
rect 27054 27460 27106 27469
rect 27238 27460 27290 27512
rect 31010 27460 31062 27512
rect 31286 27460 31338 27512
rect 33126 27528 33178 27580
rect 35242 27528 35294 27580
rect 36162 27528 36214 27580
rect 39750 27596 39802 27648
rect 46282 27596 46334 27648
rect 48490 27639 48542 27648
rect 48490 27605 48499 27639
rect 48499 27605 48533 27639
rect 48533 27605 48542 27639
rect 48490 27596 48542 27605
rect 50146 27639 50198 27648
rect 50146 27605 50155 27639
rect 50155 27605 50189 27639
rect 50189 27605 50198 27639
rect 52170 27664 52222 27716
rect 56954 27664 57006 27716
rect 57414 27664 57466 27716
rect 67902 27707 67954 27716
rect 67902 27673 67911 27707
rect 67911 27673 67945 27707
rect 67945 27673 67954 27707
rect 67902 27664 67954 27673
rect 69742 27664 69794 27716
rect 76182 27664 76234 27716
rect 50146 27596 50198 27605
rect 38830 27528 38882 27580
rect 42786 27571 42838 27580
rect 42786 27537 42795 27571
rect 42795 27537 42829 27571
rect 42829 27537 42838 27571
rect 42786 27528 42838 27537
rect 42970 27571 43022 27580
rect 42970 27537 42979 27571
rect 42979 27537 43013 27571
rect 43013 27537 43022 27571
rect 42970 27528 43022 27537
rect 43062 27528 43114 27580
rect 43522 27571 43574 27580
rect 43522 27537 43531 27571
rect 43531 27537 43565 27571
rect 43565 27537 43574 27571
rect 43522 27528 43574 27537
rect 43706 27528 43758 27580
rect 45546 27528 45598 27580
rect 47754 27528 47806 27580
rect 48398 27571 48450 27580
rect 48398 27537 48407 27571
rect 48407 27537 48441 27571
rect 48441 27537 48450 27571
rect 48398 27528 48450 27537
rect 49778 27528 49830 27580
rect 50238 27571 50290 27580
rect 50238 27537 50247 27571
rect 50247 27537 50281 27571
rect 50281 27537 50290 27571
rect 50238 27528 50290 27537
rect 24846 27392 24898 27444
rect 26962 27392 27014 27444
rect 28618 27435 28670 27444
rect 28618 27401 28627 27435
rect 28627 27401 28661 27435
rect 28661 27401 28670 27435
rect 28618 27392 28670 27401
rect 31378 27392 31430 27444
rect 7550 27324 7602 27376
rect 10586 27324 10638 27376
rect 11874 27324 11926 27376
rect 12150 27324 12202 27376
rect 15278 27324 15330 27376
rect 16014 27324 16066 27376
rect 17026 27367 17078 27376
rect 17026 27333 17035 27367
rect 17035 27333 17069 27367
rect 17069 27333 17078 27367
rect 17026 27324 17078 27333
rect 17118 27324 17170 27376
rect 22914 27324 22966 27376
rect 23374 27324 23426 27376
rect 35242 27392 35294 27444
rect 35794 27435 35846 27444
rect 35794 27401 35803 27435
rect 35803 27401 35837 27435
rect 35837 27401 35846 27435
rect 35794 27392 35846 27401
rect 31746 27367 31798 27376
rect 31746 27333 31755 27367
rect 31755 27333 31789 27367
rect 31789 27333 31798 27367
rect 31746 27324 31798 27333
rect 33126 27324 33178 27376
rect 34414 27324 34466 27376
rect 42234 27460 42286 27512
rect 45362 27503 45414 27512
rect 45362 27469 45371 27503
rect 45371 27469 45405 27503
rect 45405 27469 45414 27503
rect 45362 27460 45414 27469
rect 51250 27528 51302 27580
rect 53734 27596 53786 27648
rect 53826 27596 53878 27648
rect 51618 27528 51670 27580
rect 53366 27528 53418 27580
rect 54010 27571 54062 27580
rect 54010 27537 54019 27571
rect 54019 27537 54053 27571
rect 54053 27537 54062 27571
rect 54010 27528 54062 27537
rect 58794 27596 58846 27648
rect 62106 27596 62158 27648
rect 57690 27528 57742 27580
rect 44350 27435 44402 27444
rect 36162 27367 36214 27376
rect 36162 27333 36171 27367
rect 36171 27333 36205 27367
rect 36205 27333 36214 27367
rect 36162 27324 36214 27333
rect 42970 27324 43022 27376
rect 43706 27324 43758 27376
rect 44350 27401 44359 27435
rect 44359 27401 44393 27435
rect 44393 27401 44402 27435
rect 44350 27392 44402 27401
rect 45270 27435 45322 27444
rect 45270 27401 45279 27435
rect 45279 27401 45313 27435
rect 45313 27401 45322 27435
rect 45270 27392 45322 27401
rect 51434 27460 51486 27512
rect 52354 27460 52406 27512
rect 55298 27460 55350 27512
rect 63302 27528 63354 27580
rect 58426 27503 58478 27512
rect 45546 27324 45598 27376
rect 48674 27324 48726 27376
rect 49778 27324 49830 27376
rect 50790 27367 50842 27376
rect 50790 27333 50799 27367
rect 50799 27333 50833 27367
rect 50833 27333 50842 27367
rect 50790 27324 50842 27333
rect 51158 27324 51210 27376
rect 51526 27324 51578 27376
rect 56954 27392 57006 27444
rect 58426 27469 58435 27503
rect 58435 27469 58469 27503
rect 58469 27469 58478 27503
rect 58426 27460 58478 27469
rect 62658 27460 62710 27512
rect 63394 27503 63446 27512
rect 63394 27469 63403 27503
rect 63403 27469 63437 27503
rect 63437 27469 63446 27503
rect 63394 27460 63446 27469
rect 64130 27528 64182 27580
rect 70110 27596 70162 27648
rect 73054 27596 73106 27648
rect 68270 27571 68322 27580
rect 68270 27537 68279 27571
rect 68279 27537 68313 27571
rect 68313 27537 68322 27571
rect 68270 27528 68322 27537
rect 71674 27528 71726 27580
rect 65418 27460 65470 27512
rect 67074 27460 67126 27512
rect 67994 27460 68046 27512
rect 72318 27503 72370 27512
rect 66154 27392 66206 27444
rect 70018 27392 70070 27444
rect 68270 27324 68322 27376
rect 68730 27324 68782 27376
rect 71950 27324 72002 27376
rect 72318 27469 72327 27503
rect 72327 27469 72361 27503
rect 72361 27469 72370 27503
rect 72318 27460 72370 27469
rect 73698 27528 73750 27580
rect 78666 27528 78718 27580
rect 75630 27460 75682 27512
rect 80138 27664 80190 27716
rect 80598 27664 80650 27716
rect 81426 27596 81478 27648
rect 90074 27664 90126 27716
rect 90534 27707 90586 27716
rect 84830 27596 84882 27648
rect 89798 27596 89850 27648
rect 90534 27673 90543 27707
rect 90543 27673 90577 27707
rect 90577 27673 90586 27707
rect 90534 27664 90586 27673
rect 91086 27664 91138 27716
rect 79954 27528 80006 27580
rect 80322 27528 80374 27580
rect 75538 27392 75590 27444
rect 79770 27392 79822 27444
rect 73790 27367 73842 27376
rect 73790 27333 73799 27367
rect 73799 27333 73833 27367
rect 73833 27333 73842 27367
rect 73790 27324 73842 27333
rect 73882 27324 73934 27376
rect 79034 27324 79086 27376
rect 80230 27503 80282 27512
rect 80230 27469 80239 27503
rect 80239 27469 80273 27503
rect 80273 27469 80282 27503
rect 83266 27528 83318 27580
rect 80230 27460 80282 27469
rect 80506 27392 80558 27444
rect 84094 27503 84146 27512
rect 84094 27469 84103 27503
rect 84103 27469 84137 27503
rect 84137 27469 84146 27503
rect 84094 27460 84146 27469
rect 86118 27528 86170 27580
rect 87682 27571 87734 27580
rect 87682 27537 87691 27571
rect 87691 27537 87725 27571
rect 87725 27537 87734 27571
rect 87682 27528 87734 27537
rect 89246 27571 89298 27580
rect 89246 27537 89255 27571
rect 89255 27537 89289 27571
rect 89289 27537 89298 27571
rect 89246 27528 89298 27537
rect 90350 27528 90402 27580
rect 85750 27503 85802 27512
rect 85750 27469 85759 27503
rect 85759 27469 85793 27503
rect 85793 27469 85802 27503
rect 85750 27460 85802 27469
rect 85014 27435 85066 27444
rect 85014 27401 85023 27435
rect 85023 27401 85057 27435
rect 85057 27401 85066 27435
rect 85014 27392 85066 27401
rect 87590 27324 87642 27376
rect 89338 27367 89390 27376
rect 89338 27333 89347 27367
rect 89347 27333 89381 27367
rect 89381 27333 89390 27367
rect 89338 27324 89390 27333
rect 3680 27222 3732 27274
rect 3744 27222 3796 27274
rect 3808 27222 3860 27274
rect 3872 27222 3924 27274
rect 9008 27222 9060 27274
rect 9072 27222 9124 27274
rect 9136 27222 9188 27274
rect 9200 27222 9252 27274
rect 14336 27222 14388 27274
rect 14400 27222 14452 27274
rect 14464 27222 14516 27274
rect 14528 27222 14580 27274
rect 19664 27222 19716 27274
rect 19728 27222 19780 27274
rect 19792 27222 19844 27274
rect 19856 27222 19908 27274
rect 24992 27222 25044 27274
rect 25056 27222 25108 27274
rect 25120 27222 25172 27274
rect 25184 27222 25236 27274
rect 30320 27222 30372 27274
rect 30384 27222 30436 27274
rect 30448 27222 30500 27274
rect 30512 27222 30564 27274
rect 35648 27222 35700 27274
rect 35712 27222 35764 27274
rect 35776 27222 35828 27274
rect 35840 27222 35892 27274
rect 40976 27222 41028 27274
rect 41040 27222 41092 27274
rect 41104 27222 41156 27274
rect 41168 27222 41220 27274
rect 46304 27222 46356 27274
rect 46368 27222 46420 27274
rect 46432 27222 46484 27274
rect 46496 27222 46548 27274
rect 51632 27222 51684 27274
rect 51696 27222 51748 27274
rect 51760 27222 51812 27274
rect 51824 27222 51876 27274
rect 56960 27222 57012 27274
rect 57024 27222 57076 27274
rect 57088 27222 57140 27274
rect 57152 27222 57204 27274
rect 62288 27222 62340 27274
rect 62352 27222 62404 27274
rect 62416 27222 62468 27274
rect 62480 27222 62532 27274
rect 67616 27222 67668 27274
rect 67680 27222 67732 27274
rect 67744 27222 67796 27274
rect 67808 27222 67860 27274
rect 72944 27222 72996 27274
rect 73008 27222 73060 27274
rect 73072 27222 73124 27274
rect 73136 27222 73188 27274
rect 78272 27222 78324 27274
rect 78336 27222 78388 27274
rect 78400 27222 78452 27274
rect 78464 27222 78516 27274
rect 83600 27222 83652 27274
rect 83664 27222 83716 27274
rect 83728 27222 83780 27274
rect 83792 27222 83844 27274
rect 88928 27222 88980 27274
rect 88992 27222 89044 27274
rect 89056 27222 89108 27274
rect 89120 27222 89172 27274
rect 4054 27120 4106 27172
rect 9298 27163 9350 27172
rect 9298 27129 9307 27163
rect 9307 27129 9341 27163
rect 9341 27129 9350 27163
rect 9298 27120 9350 27129
rect 12150 27120 12202 27172
rect 12702 27120 12754 27172
rect 13162 27163 13214 27172
rect 13162 27129 13171 27163
rect 13171 27129 13205 27163
rect 13205 27129 13214 27163
rect 13162 27120 13214 27129
rect 16474 27163 16526 27172
rect 4606 27052 4658 27104
rect 2950 26984 3002 27036
rect 10586 27052 10638 27104
rect 4054 26916 4106 26968
rect 4422 26916 4474 26968
rect 4698 26916 4750 26968
rect 9298 26916 9350 26968
rect 10126 26959 10178 26968
rect 10126 26925 10135 26959
rect 10135 26925 10169 26959
rect 10169 26925 10178 26959
rect 10126 26916 10178 26925
rect 10310 26959 10362 26968
rect 10310 26925 10319 26959
rect 10319 26925 10353 26959
rect 10353 26925 10362 26959
rect 10310 26916 10362 26925
rect 5526 26848 5578 26900
rect 9022 26848 9074 26900
rect 10678 26891 10730 26900
rect 4790 26780 4842 26832
rect 10678 26857 10687 26891
rect 10687 26857 10721 26891
rect 10721 26857 10730 26891
rect 10678 26848 10730 26857
rect 12058 26984 12110 27036
rect 12426 26959 12478 26968
rect 12426 26925 12435 26959
rect 12435 26925 12469 26959
rect 12469 26925 12478 26959
rect 12426 26916 12478 26925
rect 12702 26959 12754 26968
rect 12702 26925 12711 26959
rect 12711 26925 12745 26959
rect 12745 26925 12754 26959
rect 12702 26916 12754 26925
rect 16474 27129 16483 27163
rect 16483 27129 16517 27163
rect 16517 27129 16526 27163
rect 16474 27120 16526 27129
rect 16566 27120 16618 27172
rect 15646 26984 15698 27036
rect 17578 27052 17630 27104
rect 17762 27052 17814 27104
rect 16566 26916 16618 26968
rect 17026 26984 17078 27036
rect 17670 26916 17722 26968
rect 17762 26916 17814 26968
rect 19142 26916 19194 26968
rect 23742 27052 23794 27104
rect 22546 26984 22598 27036
rect 24478 27052 24530 27104
rect 24662 27120 24714 27172
rect 24110 27027 24162 27036
rect 24110 26993 24119 27027
rect 24119 26993 24153 27027
rect 24153 26993 24162 27027
rect 24110 26984 24162 26993
rect 25858 27052 25910 27104
rect 26962 27052 27014 27104
rect 22914 26959 22966 26968
rect 22914 26925 22923 26959
rect 22923 26925 22957 26959
rect 22957 26925 22966 26959
rect 22914 26916 22966 26925
rect 23650 26848 23702 26900
rect 18774 26780 18826 26832
rect 24018 26916 24070 26968
rect 24662 26916 24714 26968
rect 25858 26916 25910 26968
rect 27606 26959 27658 26968
rect 27606 26925 27615 26959
rect 27615 26925 27649 26959
rect 27649 26925 27658 26959
rect 27606 26916 27658 26925
rect 23926 26848 23978 26900
rect 27974 27095 28026 27104
rect 27974 27061 27983 27095
rect 27983 27061 28017 27095
rect 28017 27061 28026 27095
rect 27974 27052 28026 27061
rect 28618 27052 28670 27104
rect 30734 27120 30786 27172
rect 33770 27120 33822 27172
rect 33954 27163 34006 27172
rect 33954 27129 33963 27163
rect 33963 27129 33997 27163
rect 33997 27129 34006 27163
rect 33954 27120 34006 27129
rect 34138 27120 34190 27172
rect 35242 27120 35294 27172
rect 29446 27027 29498 27036
rect 29446 26993 29455 27027
rect 29455 26993 29489 27027
rect 29489 26993 29498 27027
rect 29446 26984 29498 26993
rect 30826 27052 30878 27104
rect 31470 27052 31522 27104
rect 31654 27052 31706 27104
rect 33126 27052 33178 27104
rect 35610 27052 35662 27104
rect 29814 26916 29866 26968
rect 29354 26848 29406 26900
rect 30274 26916 30326 26968
rect 30734 26959 30786 26968
rect 30734 26925 30743 26959
rect 30743 26925 30777 26959
rect 30777 26925 30786 26959
rect 30734 26916 30786 26925
rect 31286 26984 31338 27036
rect 31194 26916 31246 26968
rect 36162 27052 36214 27104
rect 43246 27120 43298 27172
rect 45362 27120 45414 27172
rect 48674 27120 48726 27172
rect 55298 27120 55350 27172
rect 56494 27163 56546 27172
rect 56494 27129 56503 27163
rect 56503 27129 56537 27163
rect 56537 27129 56546 27163
rect 56494 27120 56546 27129
rect 58334 27163 58386 27172
rect 39014 26984 39066 27036
rect 51158 27052 51210 27104
rect 52906 27095 52958 27104
rect 52906 27061 52915 27095
rect 52915 27061 52949 27095
rect 52949 27061 52958 27095
rect 52906 27052 52958 27061
rect 53734 27052 53786 27104
rect 58334 27129 58343 27163
rect 58343 27129 58377 27163
rect 58377 27129 58386 27163
rect 58334 27120 58386 27129
rect 91178 27120 91230 27172
rect 63394 27052 63446 27104
rect 66154 27095 66206 27104
rect 66154 27061 66163 27095
rect 66163 27061 66197 27095
rect 66197 27061 66206 27095
rect 66154 27052 66206 27061
rect 69374 27095 69426 27104
rect 69374 27061 69383 27095
rect 69383 27061 69417 27095
rect 69417 27061 69426 27095
rect 69374 27052 69426 27061
rect 71122 27052 71174 27104
rect 35150 26916 35202 26968
rect 36346 26959 36398 26968
rect 36346 26925 36355 26959
rect 36355 26925 36389 26959
rect 36389 26925 36398 26959
rect 36346 26916 36398 26925
rect 36530 26959 36582 26968
rect 36530 26925 36539 26959
rect 36539 26925 36573 26959
rect 36573 26925 36582 26959
rect 36530 26916 36582 26925
rect 36714 26916 36766 26968
rect 39290 26916 39342 26968
rect 34966 26848 35018 26900
rect 35610 26891 35662 26900
rect 35610 26857 35619 26891
rect 35619 26857 35653 26891
rect 35653 26857 35662 26891
rect 42510 26959 42562 26968
rect 42510 26925 42519 26959
rect 42519 26925 42553 26959
rect 42553 26925 42562 26959
rect 42510 26916 42562 26925
rect 44166 26984 44218 27036
rect 44350 26984 44402 27036
rect 48398 26984 48450 27036
rect 50146 27027 50198 27036
rect 48582 26916 48634 26968
rect 50146 26993 50155 27027
rect 50155 26993 50189 27027
rect 50189 26993 50198 27027
rect 50146 26984 50198 26993
rect 51434 27027 51486 27036
rect 35610 26848 35662 26857
rect 49318 26848 49370 26900
rect 50238 26916 50290 26968
rect 50422 26916 50474 26968
rect 51066 26916 51118 26968
rect 51434 26993 51443 27027
rect 51443 26993 51477 27027
rect 51477 26993 51486 27027
rect 51434 26984 51486 26993
rect 52170 26984 52222 27036
rect 56494 26984 56546 27036
rect 61186 26984 61238 27036
rect 62658 27027 62710 27036
rect 62658 26993 62667 27027
rect 62667 26993 62701 27027
rect 62701 26993 62710 27027
rect 62658 26984 62710 26993
rect 63302 26984 63354 27036
rect 64130 26984 64182 27036
rect 34414 26780 34466 26832
rect 56862 26916 56914 26968
rect 65418 26959 65470 26968
rect 53458 26848 53510 26900
rect 65418 26925 65427 26959
rect 65427 26925 65461 26959
rect 65461 26925 65470 26959
rect 65418 26916 65470 26925
rect 67994 27027 68046 27036
rect 67994 26993 68003 27027
rect 68003 26993 68037 27027
rect 68037 26993 68046 27027
rect 67994 26984 68046 26993
rect 68270 27027 68322 27036
rect 68270 26993 68279 27027
rect 68279 26993 68313 27027
rect 68313 26993 68322 27027
rect 68270 26984 68322 26993
rect 68454 26984 68506 27036
rect 70110 27027 70162 27036
rect 70110 26993 70119 27027
rect 70119 26993 70153 27027
rect 70153 26993 70162 27027
rect 70110 26984 70162 26993
rect 72318 26984 72370 27036
rect 68362 26916 68414 26968
rect 75630 27095 75682 27104
rect 73606 26984 73658 27036
rect 73330 26959 73382 26968
rect 70018 26848 70070 26900
rect 70846 26848 70898 26900
rect 70938 26891 70990 26900
rect 70938 26857 70947 26891
rect 70947 26857 70981 26891
rect 70981 26857 70990 26891
rect 71214 26891 71266 26900
rect 70938 26848 70990 26857
rect 71214 26857 71223 26891
rect 71223 26857 71257 26891
rect 71257 26857 71266 26891
rect 71214 26848 71266 26857
rect 71306 26891 71358 26900
rect 71306 26857 71315 26891
rect 71315 26857 71349 26891
rect 71349 26857 71358 26891
rect 71490 26891 71542 26900
rect 71306 26848 71358 26857
rect 71490 26857 71499 26891
rect 71499 26857 71533 26891
rect 71533 26857 71542 26891
rect 71490 26848 71542 26857
rect 71950 26848 72002 26900
rect 73330 26925 73339 26959
rect 73339 26925 73373 26959
rect 73373 26925 73382 26959
rect 73330 26916 73382 26925
rect 73882 26916 73934 26968
rect 75630 27061 75639 27095
rect 75639 27061 75673 27095
rect 75673 27061 75682 27095
rect 75630 27052 75682 27061
rect 79218 27052 79270 27104
rect 87682 27095 87734 27104
rect 87682 27061 87691 27095
rect 87691 27061 87725 27095
rect 87725 27061 87734 27095
rect 87682 27052 87734 27061
rect 75538 26959 75590 26968
rect 75538 26925 75547 26959
rect 75547 26925 75581 26959
rect 75581 26925 75590 26959
rect 75538 26916 75590 26925
rect 79034 26916 79086 26968
rect 79218 26959 79270 26968
rect 79218 26925 79227 26959
rect 79227 26925 79261 26959
rect 79261 26925 79270 26959
rect 79218 26916 79270 26925
rect 85750 26984 85802 27036
rect 86578 27027 86630 27036
rect 86578 26993 86587 27027
rect 86587 26993 86621 27027
rect 86621 26993 86630 27027
rect 86578 26984 86630 26993
rect 89338 26984 89390 27036
rect 50330 26780 50382 26832
rect 50422 26780 50474 26832
rect 69926 26823 69978 26832
rect 69926 26789 69935 26823
rect 69935 26789 69969 26823
rect 69969 26789 69978 26823
rect 69926 26780 69978 26789
rect 78666 26848 78718 26900
rect 84094 26916 84146 26968
rect 85566 26916 85618 26968
rect 90442 26959 90494 26968
rect 90442 26925 90451 26959
rect 90451 26925 90485 26959
rect 90485 26925 90494 26959
rect 90442 26916 90494 26925
rect 80506 26848 80558 26900
rect 84830 26891 84882 26900
rect 84830 26857 84839 26891
rect 84839 26857 84873 26891
rect 84873 26857 84882 26891
rect 84830 26848 84882 26857
rect 89614 26848 89666 26900
rect 6344 26678 6396 26730
rect 6408 26678 6460 26730
rect 6472 26678 6524 26730
rect 6536 26678 6588 26730
rect 11672 26678 11724 26730
rect 11736 26678 11788 26730
rect 11800 26678 11852 26730
rect 11864 26678 11916 26730
rect 17000 26678 17052 26730
rect 17064 26678 17116 26730
rect 17128 26678 17180 26730
rect 17192 26678 17244 26730
rect 22328 26678 22380 26730
rect 22392 26678 22444 26730
rect 22456 26678 22508 26730
rect 22520 26678 22572 26730
rect 27656 26678 27708 26730
rect 27720 26678 27772 26730
rect 27784 26678 27836 26730
rect 27848 26678 27900 26730
rect 32984 26678 33036 26730
rect 33048 26678 33100 26730
rect 33112 26678 33164 26730
rect 33176 26678 33228 26730
rect 38312 26678 38364 26730
rect 38376 26678 38428 26730
rect 38440 26678 38492 26730
rect 38504 26678 38556 26730
rect 43640 26678 43692 26730
rect 43704 26678 43756 26730
rect 43768 26678 43820 26730
rect 43832 26678 43884 26730
rect 48968 26678 49020 26730
rect 49032 26678 49084 26730
rect 49096 26678 49148 26730
rect 49160 26678 49212 26730
rect 54296 26678 54348 26730
rect 54360 26678 54412 26730
rect 54424 26678 54476 26730
rect 54488 26678 54540 26730
rect 59624 26678 59676 26730
rect 59688 26678 59740 26730
rect 59752 26678 59804 26730
rect 59816 26678 59868 26730
rect 64952 26678 65004 26730
rect 65016 26678 65068 26730
rect 65080 26678 65132 26730
rect 65144 26678 65196 26730
rect 70280 26678 70332 26730
rect 70344 26678 70396 26730
rect 70408 26678 70460 26730
rect 70472 26678 70524 26730
rect 75608 26678 75660 26730
rect 75672 26678 75724 26730
rect 75736 26678 75788 26730
rect 75800 26678 75852 26730
rect 80936 26678 80988 26730
rect 81000 26678 81052 26730
rect 81064 26678 81116 26730
rect 81128 26678 81180 26730
rect 86264 26678 86316 26730
rect 86328 26678 86380 26730
rect 86392 26678 86444 26730
rect 86456 26678 86508 26730
rect 91592 26678 91644 26730
rect 91656 26678 91708 26730
rect 91720 26678 91772 26730
rect 91784 26678 91836 26730
rect 3962 26619 4014 26628
rect 3962 26585 3971 26619
rect 3971 26585 4005 26619
rect 4005 26585 4014 26619
rect 3962 26576 4014 26585
rect 5526 26576 5578 26628
rect 6170 26576 6222 26628
rect 23650 26576 23702 26628
rect 25398 26576 25450 26628
rect 38094 26619 38146 26628
rect 38094 26585 38103 26619
rect 38103 26585 38137 26619
rect 38137 26585 38146 26619
rect 38094 26576 38146 26585
rect 39382 26576 39434 26628
rect 31378 26508 31430 26560
rect 34138 26440 34190 26492
rect 42878 26508 42930 26560
rect 5802 26415 5854 26424
rect 5802 26381 5811 26415
rect 5811 26381 5845 26415
rect 5845 26381 5854 26415
rect 5802 26372 5854 26381
rect 33954 26372 34006 26424
rect 35978 26440 36030 26492
rect 38094 26440 38146 26492
rect 39290 26483 39342 26492
rect 39290 26449 39299 26483
rect 39299 26449 39333 26483
rect 39333 26449 39342 26483
rect 39290 26440 39342 26449
rect 39382 26483 39434 26492
rect 39382 26449 39391 26483
rect 39391 26449 39425 26483
rect 39425 26449 39434 26483
rect 39382 26440 39434 26449
rect 38554 26415 38606 26424
rect 38554 26381 38563 26415
rect 38563 26381 38597 26415
rect 38597 26381 38606 26415
rect 38554 26372 38606 26381
rect 6630 26304 6682 26356
rect 11506 26304 11558 26356
rect 3502 26236 3554 26288
rect 34690 26236 34742 26288
rect 36806 26236 36858 26288
rect 37726 26236 37778 26288
rect 38554 26236 38606 26288
rect 40854 26236 40906 26288
rect 67074 26236 67126 26288
rect 69926 26236 69978 26288
rect 3680 26134 3732 26186
rect 3744 26134 3796 26186
rect 3808 26134 3860 26186
rect 3872 26134 3924 26186
rect 35648 26134 35700 26186
rect 35712 26134 35764 26186
rect 35776 26134 35828 26186
rect 35840 26134 35892 26186
rect 40976 26134 41028 26186
rect 41040 26134 41092 26186
rect 41104 26134 41156 26186
rect 41168 26134 41220 26186
rect 4054 26032 4106 26084
rect 6630 26075 6682 26084
rect 6630 26041 6639 26075
rect 6639 26041 6673 26075
rect 6673 26041 6682 26075
rect 6630 26032 6682 26041
rect 35978 26075 36030 26084
rect 35978 26041 35987 26075
rect 35987 26041 36021 26075
rect 36021 26041 36030 26075
rect 35978 26032 36030 26041
rect 36530 26032 36582 26084
rect 4238 25964 4290 26016
rect 4514 25964 4566 26016
rect 2766 25828 2818 25880
rect 3502 25828 3554 25880
rect 39290 26032 39342 26084
rect 31838 25896 31890 25948
rect 34690 25939 34742 25948
rect 34414 25871 34466 25880
rect 34414 25837 34423 25871
rect 34423 25837 34457 25871
rect 34457 25837 34466 25871
rect 34414 25828 34466 25837
rect 34690 25905 34699 25939
rect 34699 25905 34733 25939
rect 34733 25905 34742 25939
rect 34690 25896 34742 25905
rect 36714 25896 36766 25948
rect 42510 25896 42562 25948
rect 6630 25760 6682 25812
rect 37174 25760 37226 25812
rect 42234 25828 42286 25880
rect 38830 25692 38882 25744
rect 6344 25590 6396 25642
rect 6408 25590 6460 25642
rect 6472 25590 6524 25642
rect 6536 25590 6588 25642
rect 38312 25590 38364 25642
rect 38376 25590 38428 25642
rect 38440 25590 38492 25642
rect 38504 25590 38556 25642
rect 16750 25488 16802 25540
rect 70202 25488 70254 25540
rect 2766 25420 2818 25472
rect 4238 25420 4290 25472
rect 5802 25463 5854 25472
rect 5802 25429 5811 25463
rect 5811 25429 5845 25463
rect 5845 25429 5854 25463
rect 5802 25420 5854 25429
rect 34414 25463 34466 25472
rect 34414 25429 34423 25463
rect 34423 25429 34457 25463
rect 34457 25429 34466 25463
rect 34414 25420 34466 25429
rect 36806 25420 36858 25472
rect 6630 25352 6682 25404
rect 38094 25395 38146 25404
rect 38094 25361 38103 25395
rect 38103 25361 38137 25395
rect 38137 25361 38146 25395
rect 38094 25352 38146 25361
rect 38830 25395 38882 25404
rect 38830 25361 38839 25395
rect 38839 25361 38873 25395
rect 38873 25361 38882 25395
rect 38830 25352 38882 25361
rect 42510 25420 42562 25472
rect 4606 25327 4658 25336
rect 4606 25293 4615 25327
rect 4615 25293 4649 25327
rect 4649 25293 4658 25327
rect 4606 25284 4658 25293
rect 37542 25284 37594 25336
rect 4146 25216 4198 25268
rect 4054 25148 4106 25200
rect 23834 25148 23886 25200
rect 39290 25148 39342 25200
rect 3680 25046 3732 25098
rect 3744 25046 3796 25098
rect 3808 25046 3860 25098
rect 3872 25046 3924 25098
rect 35648 25046 35700 25098
rect 35712 25046 35764 25098
rect 35776 25046 35828 25098
rect 35840 25046 35892 25098
rect 40976 25046 41028 25098
rect 41040 25046 41092 25098
rect 41104 25046 41156 25098
rect 41168 25046 41220 25098
rect 2766 24944 2818 24996
rect 7090 24944 7142 24996
rect 35150 24987 35202 24996
rect 35150 24953 35159 24987
rect 35159 24953 35193 24987
rect 35193 24953 35202 24987
rect 35150 24944 35202 24953
rect 42234 24987 42286 24996
rect 42234 24953 42243 24987
rect 42243 24953 42277 24987
rect 42277 24953 42286 24987
rect 42234 24944 42286 24953
rect 3410 24808 3462 24860
rect 5066 24808 5118 24860
rect 34874 24876 34926 24928
rect 4698 24740 4750 24792
rect 7090 24783 7142 24792
rect 7090 24749 7099 24783
rect 7099 24749 7133 24783
rect 7133 24749 7142 24783
rect 7090 24740 7142 24749
rect 4054 24672 4106 24724
rect 16750 24672 16802 24724
rect 34414 24740 34466 24792
rect 38186 24808 38238 24860
rect 38830 24808 38882 24860
rect 40854 24808 40906 24860
rect 36898 24783 36950 24792
rect 25398 24672 25450 24724
rect 36898 24749 36907 24783
rect 36907 24749 36941 24783
rect 36941 24749 36950 24783
rect 36898 24740 36950 24749
rect 37082 24783 37134 24792
rect 37082 24749 37091 24783
rect 37091 24749 37125 24783
rect 37125 24749 37134 24783
rect 37082 24740 37134 24749
rect 38186 24672 38238 24724
rect 3686 24604 3738 24656
rect 6722 24604 6774 24656
rect 9850 24604 9902 24656
rect 36714 24604 36766 24656
rect 6344 24502 6396 24554
rect 6408 24502 6460 24554
rect 6472 24502 6524 24554
rect 6536 24502 6588 24554
rect 38312 24502 38364 24554
rect 38376 24502 38428 24554
rect 38440 24502 38492 24554
rect 38504 24502 38556 24554
rect 4698 24443 4750 24452
rect 4698 24409 4707 24443
rect 4707 24409 4741 24443
rect 4741 24409 4750 24443
rect 4698 24400 4750 24409
rect 2490 24332 2542 24384
rect 5066 24375 5118 24384
rect 3686 24307 3738 24316
rect 3686 24273 3695 24307
rect 3695 24273 3729 24307
rect 3729 24273 3738 24307
rect 3686 24264 3738 24273
rect 5066 24341 5075 24375
rect 5075 24341 5109 24375
rect 5109 24341 5118 24375
rect 5066 24332 5118 24341
rect 7550 24375 7602 24384
rect 7550 24341 7559 24375
rect 7559 24341 7593 24375
rect 7593 24341 7602 24375
rect 7550 24332 7602 24341
rect 37082 24400 37134 24452
rect 15278 24332 15330 24384
rect 4146 24307 4198 24316
rect 4146 24273 4155 24307
rect 4155 24273 4189 24307
rect 4189 24273 4198 24307
rect 4146 24264 4198 24273
rect 4238 24307 4290 24316
rect 4238 24273 4247 24307
rect 4247 24273 4281 24307
rect 4281 24273 4290 24307
rect 4238 24264 4290 24273
rect 10678 24264 10730 24316
rect 35150 24264 35202 24316
rect 36990 24264 37042 24316
rect 39474 24264 39526 24316
rect 6722 24196 6774 24248
rect 7550 24196 7602 24248
rect 36714 24128 36766 24180
rect 39474 24128 39526 24180
rect 70018 24128 70070 24180
rect 7274 24103 7326 24112
rect 7274 24069 7283 24103
rect 7283 24069 7317 24103
rect 7317 24069 7326 24103
rect 7274 24060 7326 24069
rect 3680 23958 3732 24010
rect 3744 23958 3796 24010
rect 3808 23958 3860 24010
rect 3872 23958 3924 24010
rect 7274 23856 7326 23908
rect 30274 24060 30326 24112
rect 35648 23958 35700 24010
rect 35712 23958 35764 24010
rect 35776 23958 35828 24010
rect 35840 23958 35892 24010
rect 40976 23958 41028 24010
rect 41040 23958 41092 24010
rect 41104 23958 41156 24010
rect 41168 23958 41220 24010
rect 6906 23788 6958 23840
rect 33954 23856 34006 23908
rect 34046 23856 34098 23908
rect 34874 23899 34926 23908
rect 6630 23720 6682 23772
rect 31378 23720 31430 23772
rect 2490 23652 2542 23704
rect 2674 23652 2726 23704
rect 3594 23652 3646 23704
rect 7274 23652 7326 23704
rect 34598 23652 34650 23704
rect 34874 23865 34883 23899
rect 34883 23865 34917 23899
rect 34917 23865 34926 23899
rect 34874 23856 34926 23865
rect 36806 23856 36858 23908
rect 35610 23652 35662 23704
rect 42326 23720 42378 23772
rect 68270 23720 68322 23772
rect 70938 23720 70990 23772
rect 36806 23652 36858 23704
rect 36530 23627 36582 23636
rect 36530 23593 36539 23627
rect 36539 23593 36573 23627
rect 36573 23593 36582 23627
rect 36530 23584 36582 23593
rect 3318 23559 3370 23568
rect 3318 23525 3327 23559
rect 3327 23525 3361 23559
rect 3361 23525 3370 23559
rect 3318 23516 3370 23525
rect 9022 23516 9074 23568
rect 38646 23516 38698 23568
rect 43522 23516 43574 23568
rect 6344 23414 6396 23466
rect 6408 23414 6460 23466
rect 6472 23414 6524 23466
rect 6536 23414 6588 23466
rect 38312 23414 38364 23466
rect 38376 23414 38428 23466
rect 38440 23414 38492 23466
rect 38504 23414 38556 23466
rect 3594 23355 3646 23364
rect 3594 23321 3603 23355
rect 3603 23321 3637 23355
rect 3637 23321 3646 23355
rect 3594 23312 3646 23321
rect 3410 23244 3462 23296
rect 6722 23312 6774 23364
rect 39474 23355 39526 23364
rect 39474 23321 39483 23355
rect 39483 23321 39517 23355
rect 39517 23321 39526 23355
rect 39474 23312 39526 23321
rect 3502 23219 3554 23228
rect 3502 23185 3511 23219
rect 3511 23185 3545 23219
rect 3545 23185 3554 23219
rect 3502 23176 3554 23185
rect 6630 23244 6682 23296
rect 39566 23244 39618 23296
rect 34414 23219 34466 23228
rect 34414 23185 34423 23219
rect 34423 23185 34457 23219
rect 34457 23185 34466 23219
rect 34414 23176 34466 23185
rect 38186 23219 38238 23228
rect 38186 23185 38195 23219
rect 38195 23185 38229 23219
rect 38229 23185 38238 23219
rect 38186 23176 38238 23185
rect 7182 23108 7234 23160
rect 3502 22972 3554 23024
rect 35334 22972 35386 23024
rect 36714 22972 36766 23024
rect 42326 23108 42378 23160
rect 40670 22972 40722 23024
rect 3680 22870 3732 22922
rect 3744 22870 3796 22922
rect 3808 22870 3860 22922
rect 3872 22870 3924 22922
rect 35648 22870 35700 22922
rect 35712 22870 35764 22922
rect 35776 22870 35828 22922
rect 35840 22870 35892 22922
rect 40976 22870 41028 22922
rect 41040 22870 41092 22922
rect 41104 22870 41156 22922
rect 41168 22870 41220 22922
rect 6630 22811 6682 22820
rect 6630 22777 6639 22811
rect 6639 22777 6673 22811
rect 6673 22777 6682 22811
rect 6630 22768 6682 22777
rect 34598 22811 34650 22820
rect 34598 22777 34607 22811
rect 34607 22777 34641 22811
rect 34641 22777 34650 22811
rect 34598 22768 34650 22777
rect 3502 22700 3554 22752
rect 3318 22632 3370 22684
rect 3410 22675 3462 22684
rect 3410 22641 3419 22675
rect 3419 22641 3453 22675
rect 3453 22641 3462 22675
rect 3410 22632 3462 22641
rect 3594 22564 3646 22616
rect 4422 22564 4474 22616
rect 30366 22632 30418 22684
rect 42326 22675 42378 22684
rect 30918 22564 30970 22616
rect 36898 22564 36950 22616
rect 38646 22607 38698 22616
rect 38646 22573 38655 22607
rect 38655 22573 38689 22607
rect 38689 22573 38698 22607
rect 38646 22564 38698 22573
rect 6630 22496 6682 22548
rect 36530 22496 36582 22548
rect 4422 22471 4474 22480
rect 4422 22437 4431 22471
rect 4431 22437 4465 22471
rect 4465 22437 4474 22471
rect 4422 22428 4474 22437
rect 34782 22471 34834 22480
rect 34782 22437 34791 22471
rect 34791 22437 34825 22471
rect 34825 22437 34834 22471
rect 34782 22428 34834 22437
rect 38094 22428 38146 22480
rect 39658 22428 39710 22480
rect 42326 22641 42335 22675
rect 42335 22641 42369 22675
rect 42369 22641 42378 22675
rect 42326 22632 42378 22641
rect 40946 22607 40998 22616
rect 40946 22573 40955 22607
rect 40955 22573 40989 22607
rect 40989 22573 40998 22607
rect 40946 22564 40998 22573
rect 43062 22471 43114 22480
rect 43062 22437 43071 22471
rect 43071 22437 43105 22471
rect 43105 22437 43114 22471
rect 43062 22428 43114 22437
rect 6344 22326 6396 22378
rect 6408 22326 6460 22378
rect 6472 22326 6524 22378
rect 6536 22326 6588 22378
rect 38312 22326 38364 22378
rect 38376 22326 38428 22378
rect 38440 22326 38492 22378
rect 38504 22326 38556 22378
rect 3870 22224 3922 22276
rect 4606 22224 4658 22276
rect 7182 22267 7234 22276
rect 7182 22233 7191 22267
rect 7191 22233 7225 22267
rect 7225 22233 7234 22267
rect 7182 22224 7234 22233
rect 39290 22224 39342 22276
rect 40946 22267 40998 22276
rect 40946 22233 40955 22267
rect 40955 22233 40989 22267
rect 40989 22233 40998 22267
rect 40946 22224 40998 22233
rect 2674 22156 2726 22208
rect 4422 22156 4474 22208
rect 2766 22088 2818 22140
rect 6078 22088 6130 22140
rect 6630 22131 6682 22140
rect 3594 22020 3646 22072
rect 3870 22063 3922 22072
rect 3870 22029 3879 22063
rect 3879 22029 3913 22063
rect 3913 22029 3922 22063
rect 3870 22020 3922 22029
rect 6630 22097 6639 22131
rect 6639 22097 6673 22131
rect 6673 22097 6682 22131
rect 6630 22088 6682 22097
rect 35426 22088 35478 22140
rect 36530 22088 36582 22140
rect 36622 22088 36674 22140
rect 40670 22131 40722 22140
rect 40670 22097 40679 22131
rect 40679 22097 40713 22131
rect 40713 22097 40722 22131
rect 40670 22088 40722 22097
rect 39290 22020 39342 22072
rect 8378 21952 8430 22004
rect 2766 21884 2818 21936
rect 4974 21927 5026 21936
rect 4974 21893 4983 21927
rect 4983 21893 5017 21927
rect 5017 21893 5026 21927
rect 4974 21884 5026 21893
rect 35426 21927 35478 21936
rect 35426 21893 35435 21927
rect 35435 21893 35469 21927
rect 35469 21893 35478 21927
rect 35426 21884 35478 21893
rect 3680 21782 3732 21834
rect 3744 21782 3796 21834
rect 3808 21782 3860 21834
rect 3872 21782 3924 21834
rect 35648 21782 35700 21834
rect 35712 21782 35764 21834
rect 35776 21782 35828 21834
rect 35840 21782 35892 21834
rect 40976 21782 41028 21834
rect 41040 21782 41092 21834
rect 41104 21782 41156 21834
rect 41168 21782 41220 21834
rect 67074 21748 67126 21800
rect 71214 21748 71266 21800
rect 4514 21680 4566 21732
rect 2674 21519 2726 21528
rect 2674 21485 2683 21519
rect 2683 21485 2717 21519
rect 2717 21485 2726 21519
rect 2674 21476 2726 21485
rect 2766 21476 2818 21528
rect 6170 21476 6222 21528
rect 36714 21680 36766 21732
rect 39658 21680 39710 21732
rect 38738 21612 38790 21664
rect 43062 21612 43114 21664
rect 36530 21544 36582 21596
rect 36990 21587 37042 21596
rect 36990 21553 36999 21587
rect 36999 21553 37033 21587
rect 37033 21553 37042 21587
rect 36990 21544 37042 21553
rect 35886 21519 35938 21528
rect 35886 21485 35895 21519
rect 35895 21485 35929 21519
rect 35929 21485 35938 21519
rect 35886 21476 35938 21485
rect 39842 21519 39894 21528
rect 39842 21485 39851 21519
rect 39851 21485 39885 21519
rect 39885 21485 39894 21519
rect 39842 21476 39894 21485
rect 41498 21476 41550 21528
rect 5066 21451 5118 21460
rect 5066 21417 5075 21451
rect 5075 21417 5109 21451
rect 5109 21417 5118 21451
rect 5066 21408 5118 21417
rect 3318 21340 3370 21392
rect 34598 21383 34650 21392
rect 34598 21349 34607 21383
rect 34607 21349 34641 21383
rect 34641 21349 34650 21383
rect 34598 21340 34650 21349
rect 34782 21383 34834 21392
rect 34782 21349 34791 21383
rect 34791 21349 34825 21383
rect 34825 21349 34834 21383
rect 34782 21340 34834 21349
rect 39474 21340 39526 21392
rect 43062 21383 43114 21392
rect 43062 21349 43071 21383
rect 43071 21349 43105 21383
rect 43105 21349 43114 21383
rect 43062 21340 43114 21349
rect 6344 21238 6396 21290
rect 6408 21238 6460 21290
rect 6472 21238 6524 21290
rect 6536 21238 6588 21290
rect 38312 21238 38364 21290
rect 38376 21238 38428 21290
rect 38440 21238 38492 21290
rect 38504 21238 38556 21290
rect 6078 21136 6130 21188
rect 34138 21136 34190 21188
rect 6906 21111 6958 21120
rect 6906 21077 6915 21111
rect 6915 21077 6949 21111
rect 6949 21077 6958 21111
rect 6906 21068 6958 21077
rect 3410 21000 3462 21052
rect 6722 21000 6774 21052
rect 34506 21000 34558 21052
rect 35334 21136 35386 21188
rect 37450 21136 37502 21188
rect 39658 21136 39710 21188
rect 35426 21068 35478 21120
rect 35886 21111 35938 21120
rect 35886 21077 35895 21111
rect 35895 21077 35929 21111
rect 35929 21077 35938 21111
rect 35886 21068 35938 21077
rect 35334 21043 35386 21052
rect 35334 21009 35343 21043
rect 35343 21009 35377 21043
rect 35377 21009 35386 21043
rect 35334 21000 35386 21009
rect 36622 21000 36674 21052
rect 38094 21000 38146 21052
rect 39474 21000 39526 21052
rect 4974 20932 5026 20984
rect 37450 20932 37502 20984
rect 39658 20932 39710 20984
rect 41498 20839 41550 20848
rect 41498 20805 41507 20839
rect 41507 20805 41541 20839
rect 41541 20805 41550 20839
rect 41498 20796 41550 20805
rect 3680 20694 3732 20746
rect 3744 20694 3796 20746
rect 3808 20694 3860 20746
rect 3872 20694 3924 20746
rect 35648 20694 35700 20746
rect 35712 20694 35764 20746
rect 35776 20694 35828 20746
rect 35840 20694 35892 20746
rect 40976 20694 41028 20746
rect 41040 20694 41092 20746
rect 41104 20694 41156 20746
rect 41168 20694 41220 20746
rect 2398 20635 2450 20644
rect 2398 20601 2407 20635
rect 2407 20601 2441 20635
rect 2441 20601 2450 20635
rect 2398 20592 2450 20601
rect 6170 20592 6222 20644
rect 34690 20592 34742 20644
rect 2766 20431 2818 20440
rect 2766 20397 2775 20431
rect 2775 20397 2809 20431
rect 2809 20397 2818 20431
rect 2766 20388 2818 20397
rect 3318 20431 3370 20440
rect 3318 20397 3327 20431
rect 3327 20397 3361 20431
rect 3361 20397 3370 20431
rect 3318 20388 3370 20397
rect 4238 20388 4290 20440
rect 39658 20592 39710 20644
rect 3594 20320 3646 20372
rect 4054 20320 4106 20372
rect 30274 20320 30326 20372
rect 43062 20456 43114 20508
rect 40946 20431 40998 20440
rect 40946 20397 40955 20431
rect 40955 20397 40989 20431
rect 40989 20397 40998 20431
rect 40946 20388 40998 20397
rect 42326 20363 42378 20372
rect 42326 20329 42335 20363
rect 42335 20329 42369 20363
rect 42369 20329 42378 20363
rect 42326 20320 42378 20329
rect 6814 20252 6866 20304
rect 34414 20295 34466 20304
rect 34414 20261 34423 20295
rect 34423 20261 34457 20295
rect 34457 20261 34466 20295
rect 34414 20252 34466 20261
rect 36438 20295 36490 20304
rect 36438 20261 36447 20295
rect 36447 20261 36481 20295
rect 36481 20261 36490 20295
rect 36438 20252 36490 20261
rect 43062 20295 43114 20304
rect 43062 20261 43071 20295
rect 43071 20261 43105 20295
rect 43105 20261 43114 20295
rect 43062 20252 43114 20261
rect 6344 20150 6396 20202
rect 6408 20150 6460 20202
rect 6472 20150 6524 20202
rect 6536 20150 6588 20202
rect 38312 20150 38364 20202
rect 38376 20150 38428 20202
rect 38440 20150 38492 20202
rect 38504 20150 38556 20202
rect 39290 20048 39342 20100
rect 6814 20023 6866 20032
rect 6814 19989 6823 20023
rect 6823 19989 6857 20023
rect 6857 19989 6866 20023
rect 6814 19980 6866 19989
rect 5066 19912 5118 19964
rect 37634 19912 37686 19964
rect 67166 19980 67218 20032
rect 70478 19980 70530 20032
rect 71306 19980 71358 20032
rect 6722 19844 6774 19896
rect 39198 19887 39250 19896
rect 39198 19853 39207 19887
rect 39207 19853 39241 19887
rect 39241 19853 39250 19887
rect 39198 19844 39250 19853
rect 30826 19776 30878 19828
rect 42326 19912 42378 19964
rect 40946 19844 40998 19896
rect 6722 19708 6774 19760
rect 6998 19751 7050 19760
rect 6998 19717 7007 19751
rect 7007 19717 7041 19751
rect 7041 19717 7050 19751
rect 6998 19708 7050 19717
rect 3680 19606 3732 19658
rect 3744 19606 3796 19658
rect 3808 19606 3860 19658
rect 3872 19606 3924 19658
rect 35648 19606 35700 19658
rect 35712 19606 35764 19658
rect 35776 19606 35828 19658
rect 35840 19606 35892 19658
rect 40976 19606 41028 19658
rect 41040 19606 41092 19658
rect 41104 19606 41156 19658
rect 41168 19606 41220 19658
rect 4238 19547 4290 19556
rect 4238 19513 4247 19547
rect 4247 19513 4281 19547
rect 4281 19513 4290 19547
rect 4238 19504 4290 19513
rect 34506 19504 34558 19556
rect 34966 19504 35018 19556
rect 37450 19504 37502 19556
rect 4054 19368 4106 19420
rect 4146 19343 4198 19352
rect 4146 19309 4155 19343
rect 4155 19309 4189 19343
rect 4189 19309 4198 19343
rect 4146 19300 4198 19309
rect 35426 19343 35478 19352
rect 35426 19309 35435 19343
rect 35435 19309 35469 19343
rect 35469 19309 35478 19343
rect 35426 19300 35478 19309
rect 37634 19343 37686 19352
rect 37634 19309 37643 19343
rect 37643 19309 37677 19343
rect 37677 19309 37686 19343
rect 37634 19300 37686 19309
rect 36438 19232 36490 19284
rect 38922 19300 38974 19352
rect 40578 19300 40630 19352
rect 39382 19232 39434 19284
rect 3502 19207 3554 19216
rect 3502 19173 3511 19207
rect 3511 19173 3545 19207
rect 3545 19173 3554 19207
rect 3502 19164 3554 19173
rect 34414 19207 34466 19216
rect 34414 19173 34423 19207
rect 34423 19173 34457 19207
rect 34457 19173 34466 19207
rect 34414 19164 34466 19173
rect 6344 19062 6396 19114
rect 6408 19062 6460 19114
rect 6472 19062 6524 19114
rect 6536 19062 6588 19114
rect 38312 19062 38364 19114
rect 38376 19062 38428 19114
rect 38440 19062 38492 19114
rect 38504 19062 38556 19114
rect 5986 18960 6038 19012
rect 3594 18824 3646 18876
rect 4330 18892 4382 18944
rect 4422 18867 4474 18876
rect 4422 18833 4431 18867
rect 4431 18833 4465 18867
rect 4465 18833 4474 18867
rect 4422 18824 4474 18833
rect 6906 18867 6958 18876
rect 4606 18731 4658 18740
rect 4606 18697 4615 18731
rect 4615 18697 4649 18731
rect 4649 18697 4658 18731
rect 4606 18688 4658 18697
rect 6906 18833 6915 18867
rect 6915 18833 6949 18867
rect 6949 18833 6958 18867
rect 6906 18824 6958 18833
rect 34414 18867 34466 18876
rect 34414 18833 34423 18867
rect 34423 18833 34457 18867
rect 34457 18833 34466 18867
rect 34414 18824 34466 18833
rect 34598 18867 34650 18876
rect 34598 18833 34626 18867
rect 34626 18833 34650 18867
rect 34598 18824 34650 18833
rect 34966 18824 35018 18876
rect 37634 18824 37686 18876
rect 39658 18960 39710 19012
rect 40578 18960 40630 19012
rect 39382 18867 39434 18876
rect 39382 18833 39391 18867
rect 39391 18833 39425 18867
rect 39425 18833 39434 18867
rect 39382 18824 39434 18833
rect 7090 18731 7142 18740
rect 7090 18697 7099 18731
rect 7099 18697 7133 18731
rect 7133 18697 7142 18731
rect 7090 18688 7142 18697
rect 35518 18731 35570 18740
rect 35518 18697 35527 18731
rect 35527 18697 35561 18731
rect 35561 18697 35570 18731
rect 35518 18688 35570 18697
rect 70386 18824 70438 18876
rect 70846 18824 70898 18876
rect 43338 18620 43390 18672
rect 3680 18518 3732 18570
rect 3744 18518 3796 18570
rect 3808 18518 3860 18570
rect 3872 18518 3924 18570
rect 35648 18518 35700 18570
rect 35712 18518 35764 18570
rect 35776 18518 35828 18570
rect 35840 18518 35892 18570
rect 40976 18518 41028 18570
rect 41040 18518 41092 18570
rect 41104 18518 41156 18570
rect 41168 18518 41220 18570
rect 6906 18416 6958 18468
rect 4606 18280 4658 18332
rect 36714 18416 36766 18468
rect 39658 18416 39710 18468
rect 35518 18280 35570 18332
rect 3502 18212 3554 18264
rect 35426 18212 35478 18264
rect 43522 18280 43574 18332
rect 40762 18255 40814 18264
rect 40762 18221 40771 18255
rect 40771 18221 40805 18255
rect 40805 18221 40814 18255
rect 40762 18212 40814 18221
rect 5066 18119 5118 18128
rect 5066 18085 5075 18119
rect 5075 18085 5109 18119
rect 5109 18085 5118 18119
rect 5066 18076 5118 18085
rect 5526 18119 5578 18128
rect 5526 18085 5535 18119
rect 5535 18085 5569 18119
rect 5569 18085 5578 18119
rect 5526 18076 5578 18085
rect 7274 18076 7326 18128
rect 34414 18119 34466 18128
rect 34414 18085 34423 18119
rect 34423 18085 34457 18119
rect 34457 18085 34466 18119
rect 34414 18076 34466 18085
rect 42050 18119 42102 18128
rect 42050 18085 42059 18119
rect 42059 18085 42093 18119
rect 42093 18085 42102 18119
rect 42050 18076 42102 18085
rect 6344 17974 6396 18026
rect 6408 17974 6460 18026
rect 6472 17974 6524 18026
rect 6536 17974 6588 18026
rect 38312 17974 38364 18026
rect 38376 17974 38428 18026
rect 38440 17974 38492 18026
rect 38504 17974 38556 18026
rect 4422 17872 4474 17924
rect 5066 17736 5118 17788
rect 7090 17736 7142 17788
rect 38094 17736 38146 17788
rect 39198 17779 39250 17788
rect 39198 17745 39207 17779
rect 39207 17745 39241 17779
rect 39241 17745 39250 17779
rect 39198 17736 39250 17745
rect 40670 17779 40722 17788
rect 40670 17745 40679 17779
rect 40679 17745 40713 17779
rect 40713 17745 40722 17779
rect 42050 17872 42102 17924
rect 40670 17736 40722 17745
rect 5526 17668 5578 17720
rect 6078 17668 6130 17720
rect 6998 17668 7050 17720
rect 5066 17575 5118 17584
rect 5066 17541 5075 17575
rect 5075 17541 5109 17575
rect 5109 17541 5118 17575
rect 5066 17532 5118 17541
rect 7274 17575 7326 17584
rect 7274 17541 7283 17575
rect 7283 17541 7317 17575
rect 7317 17541 7326 17575
rect 7274 17532 7326 17541
rect 37542 17532 37594 17584
rect 38002 17532 38054 17584
rect 40762 17668 40814 17720
rect 3680 17430 3732 17482
rect 3744 17430 3796 17482
rect 3808 17430 3860 17482
rect 3872 17430 3924 17482
rect 35648 17430 35700 17482
rect 35712 17430 35764 17482
rect 35776 17430 35828 17482
rect 35840 17430 35892 17482
rect 40976 17430 41028 17482
rect 41040 17430 41092 17482
rect 41104 17430 41156 17482
rect 41168 17430 41220 17482
rect 36714 17260 36766 17312
rect 39750 17260 39802 17312
rect 37358 17192 37410 17244
rect 39198 17192 39250 17244
rect 34414 17031 34466 17040
rect 34414 16997 34423 17031
rect 34423 16997 34457 17031
rect 34457 16997 34466 17031
rect 34414 16988 34466 16997
rect 36346 17124 36398 17176
rect 38738 17167 38790 17176
rect 36438 17056 36490 17108
rect 38738 17133 38747 17167
rect 38747 17133 38781 17167
rect 38781 17133 38790 17167
rect 38738 17124 38790 17133
rect 39842 17167 39894 17176
rect 39842 17133 39851 17167
rect 39851 17133 39885 17167
rect 39885 17133 39894 17167
rect 39842 17124 39894 17133
rect 40762 17167 40814 17176
rect 40762 17133 40771 17167
rect 40771 17133 40805 17167
rect 40805 17133 40814 17167
rect 40762 17124 40814 17133
rect 38830 17099 38882 17108
rect 38830 17065 38839 17099
rect 38839 17065 38873 17099
rect 38873 17065 38882 17099
rect 38830 17056 38882 17065
rect 37726 16988 37778 17040
rect 39842 16988 39894 17040
rect 41038 17031 41090 17040
rect 41038 16997 41047 17031
rect 41047 16997 41081 17031
rect 41081 16997 41090 17031
rect 41038 16988 41090 16997
rect 6344 16886 6396 16938
rect 6408 16886 6460 16938
rect 6472 16886 6524 16938
rect 6536 16886 6588 16938
rect 38312 16886 38364 16938
rect 38376 16886 38428 16938
rect 38440 16886 38492 16938
rect 38504 16886 38556 16938
rect 4698 16784 4750 16836
rect 36346 16784 36398 16836
rect 39750 16784 39802 16836
rect 7182 16648 7234 16700
rect 38646 16648 38698 16700
rect 38738 16648 38790 16700
rect 5710 16623 5762 16632
rect 5710 16589 5719 16623
rect 5719 16589 5753 16623
rect 5753 16589 5762 16623
rect 5710 16580 5762 16589
rect 39750 16580 39802 16632
rect 41038 16648 41090 16700
rect 41682 16623 41734 16632
rect 41682 16589 41691 16623
rect 41691 16589 41725 16623
rect 41725 16589 41734 16623
rect 41682 16580 41734 16589
rect 6722 16555 6774 16564
rect 6722 16521 6731 16555
rect 6731 16521 6765 16555
rect 6765 16521 6774 16555
rect 6722 16512 6774 16521
rect 3680 16342 3732 16394
rect 3744 16342 3796 16394
rect 3808 16342 3860 16394
rect 3872 16342 3924 16394
rect 35648 16342 35700 16394
rect 35712 16342 35764 16394
rect 35776 16342 35828 16394
rect 35840 16342 35892 16394
rect 40976 16342 41028 16394
rect 41040 16342 41092 16394
rect 41104 16342 41156 16394
rect 41168 16342 41220 16394
rect 4698 16240 4750 16292
rect 36346 16283 36398 16292
rect 36346 16249 36355 16283
rect 36355 16249 36389 16283
rect 36389 16249 36398 16283
rect 36346 16240 36398 16249
rect 4882 16172 4934 16224
rect 38002 16240 38054 16292
rect 4698 16079 4750 16088
rect 4698 16045 4707 16079
rect 4707 16045 4741 16079
rect 4741 16045 4750 16079
rect 4698 16036 4750 16045
rect 5250 16011 5302 16020
rect 5250 15977 5259 16011
rect 5259 15977 5293 16011
rect 5293 15977 5302 16011
rect 5250 15968 5302 15977
rect 36438 16036 36490 16088
rect 37174 16079 37226 16088
rect 37174 16045 37183 16079
rect 37183 16045 37217 16079
rect 37217 16045 37226 16079
rect 37174 16036 37226 16045
rect 38922 16036 38974 16088
rect 6998 15900 7050 15952
rect 37726 15943 37778 15952
rect 37726 15909 37735 15943
rect 37735 15909 37769 15943
rect 37769 15909 37778 15943
rect 37726 15900 37778 15909
rect 6344 15798 6396 15850
rect 6408 15798 6460 15850
rect 6472 15798 6524 15850
rect 6536 15798 6588 15850
rect 38312 15798 38364 15850
rect 38376 15798 38428 15850
rect 38440 15798 38492 15850
rect 38504 15798 38556 15850
rect 68362 15832 68414 15884
rect 70478 15832 70530 15884
rect 71490 15832 71542 15884
rect 36714 15696 36766 15748
rect 5250 15560 5302 15612
rect 37082 15603 37134 15612
rect 37082 15569 37091 15603
rect 37091 15569 37125 15603
rect 37125 15569 37134 15603
rect 37082 15560 37134 15569
rect 37358 15603 37410 15612
rect 37358 15569 37367 15603
rect 37367 15569 37401 15603
rect 37401 15569 37410 15603
rect 37358 15560 37410 15569
rect 6078 15492 6130 15544
rect 6998 15399 7050 15408
rect 6998 15365 7007 15399
rect 7007 15365 7041 15399
rect 7041 15365 7050 15399
rect 6998 15356 7050 15365
rect 38646 15399 38698 15408
rect 38646 15365 38655 15399
rect 38655 15365 38689 15399
rect 38689 15365 38698 15399
rect 38646 15356 38698 15365
rect 43522 15356 43574 15408
rect 3680 15254 3732 15306
rect 3744 15254 3796 15306
rect 3808 15254 3860 15306
rect 3872 15254 3924 15306
rect 35648 15254 35700 15306
rect 35712 15254 35764 15306
rect 35776 15254 35828 15306
rect 35840 15254 35892 15306
rect 40976 15254 41028 15306
rect 41040 15254 41092 15306
rect 41104 15254 41156 15306
rect 41168 15254 41220 15306
rect 7182 15195 7234 15204
rect 7182 15161 7191 15195
rect 7191 15161 7225 15195
rect 7225 15161 7234 15195
rect 7182 15152 7234 15161
rect 37082 15195 37134 15204
rect 37082 15161 37091 15195
rect 37091 15161 37125 15195
rect 37125 15161 37134 15195
rect 37082 15152 37134 15161
rect 37726 15016 37778 15068
rect 38922 14923 38974 14932
rect 38922 14889 38931 14923
rect 38931 14889 38965 14923
rect 38965 14889 38974 14923
rect 38922 14880 38974 14889
rect 7366 14855 7418 14864
rect 7366 14821 7375 14855
rect 7375 14821 7409 14855
rect 7409 14821 7418 14855
rect 7366 14812 7418 14821
rect 34414 14855 34466 14864
rect 34414 14821 34423 14855
rect 34423 14821 34457 14855
rect 34457 14821 34466 14855
rect 34414 14812 34466 14821
rect 6344 14710 6396 14762
rect 6408 14710 6460 14762
rect 6472 14710 6524 14762
rect 6536 14710 6588 14762
rect 38312 14710 38364 14762
rect 38376 14710 38428 14762
rect 38440 14710 38492 14762
rect 38504 14710 38556 14762
rect 6078 14608 6130 14660
rect 6722 14472 6774 14524
rect 7366 14515 7418 14524
rect 7366 14481 7375 14515
rect 7375 14481 7409 14515
rect 7409 14481 7418 14515
rect 7366 14472 7418 14481
rect 3680 14166 3732 14218
rect 3744 14166 3796 14218
rect 3808 14166 3860 14218
rect 3872 14166 3924 14218
rect 35648 14166 35700 14218
rect 35712 14166 35764 14218
rect 35776 14166 35828 14218
rect 35840 14166 35892 14218
rect 40976 14166 41028 14218
rect 41040 14166 41092 14218
rect 41104 14166 41156 14218
rect 41168 14166 41220 14218
rect 6344 13622 6396 13674
rect 6408 13622 6460 13674
rect 6472 13622 6524 13674
rect 6536 13622 6588 13674
rect 38312 13622 38364 13674
rect 38376 13622 38428 13674
rect 38440 13622 38492 13674
rect 38504 13622 38556 13674
rect 3680 13078 3732 13130
rect 3744 13078 3796 13130
rect 3808 13078 3860 13130
rect 3872 13078 3924 13130
rect 35648 13078 35700 13130
rect 35712 13078 35764 13130
rect 35776 13078 35828 13130
rect 35840 13078 35892 13130
rect 40976 13078 41028 13130
rect 41040 13078 41092 13130
rect 41104 13078 41156 13130
rect 41168 13078 41220 13130
rect 6344 12534 6396 12586
rect 6408 12534 6460 12586
rect 6472 12534 6524 12586
rect 6536 12534 6588 12586
rect 38312 12534 38364 12586
rect 38376 12534 38428 12586
rect 38440 12534 38492 12586
rect 38504 12534 38556 12586
rect 3680 11990 3732 12042
rect 3744 11990 3796 12042
rect 3808 11990 3860 12042
rect 3872 11990 3924 12042
rect 35648 11990 35700 12042
rect 35712 11990 35764 12042
rect 35776 11990 35828 12042
rect 35840 11990 35892 12042
rect 40976 11990 41028 12042
rect 41040 11990 41092 12042
rect 41104 11990 41156 12042
rect 41168 11990 41220 12042
rect 38922 11616 38974 11668
rect 43522 11616 43574 11668
rect 6344 11446 6396 11498
rect 6408 11446 6460 11498
rect 6472 11446 6524 11498
rect 6536 11446 6588 11498
rect 38312 11446 38364 11498
rect 38376 11446 38428 11498
rect 38440 11446 38492 11498
rect 38504 11446 38556 11498
rect 3680 10902 3732 10954
rect 3744 10902 3796 10954
rect 3808 10902 3860 10954
rect 3872 10902 3924 10954
rect 35648 10902 35700 10954
rect 35712 10902 35764 10954
rect 35776 10902 35828 10954
rect 35840 10902 35892 10954
rect 40976 10902 41028 10954
rect 41040 10902 41092 10954
rect 41104 10902 41156 10954
rect 41168 10902 41220 10954
rect 34414 10503 34466 10512
rect 34414 10469 34423 10503
rect 34423 10469 34457 10503
rect 34457 10469 34466 10503
rect 34414 10460 34466 10469
rect 6344 10358 6396 10410
rect 6408 10358 6460 10410
rect 6472 10358 6524 10410
rect 6536 10358 6588 10410
rect 38312 10358 38364 10410
rect 38376 10358 38428 10410
rect 38440 10358 38492 10410
rect 38504 10358 38556 10410
rect 6078 10120 6130 10172
rect 11138 10188 11190 10240
rect 7090 9959 7142 9968
rect 7090 9925 7099 9959
rect 7099 9925 7133 9959
rect 7133 9925 7142 9959
rect 7090 9916 7142 9925
rect 3680 9814 3732 9866
rect 3744 9814 3796 9866
rect 3808 9814 3860 9866
rect 3872 9814 3924 9866
rect 35648 9814 35700 9866
rect 35712 9814 35764 9866
rect 35776 9814 35828 9866
rect 35840 9814 35892 9866
rect 40976 9814 41028 9866
rect 41040 9814 41092 9866
rect 41104 9814 41156 9866
rect 41168 9814 41220 9866
rect 6344 9270 6396 9322
rect 6408 9270 6460 9322
rect 6472 9270 6524 9322
rect 6536 9270 6588 9322
rect 38312 9270 38364 9322
rect 38376 9270 38428 9322
rect 38440 9270 38492 9322
rect 38504 9270 38556 9322
rect 3680 8726 3732 8778
rect 3744 8726 3796 8778
rect 3808 8726 3860 8778
rect 3872 8726 3924 8778
rect 35648 8726 35700 8778
rect 35712 8726 35764 8778
rect 35776 8726 35828 8778
rect 35840 8726 35892 8778
rect 40976 8726 41028 8778
rect 41040 8726 41092 8778
rect 41104 8726 41156 8778
rect 41168 8726 41220 8778
rect 6344 8182 6396 8234
rect 6408 8182 6460 8234
rect 6472 8182 6524 8234
rect 6536 8182 6588 8234
rect 38312 8182 38364 8234
rect 38376 8182 38428 8234
rect 38440 8182 38492 8234
rect 38504 8182 38556 8234
rect 3680 7638 3732 7690
rect 3744 7638 3796 7690
rect 3808 7638 3860 7690
rect 3872 7638 3924 7690
rect 35648 7638 35700 7690
rect 35712 7638 35764 7690
rect 35776 7638 35828 7690
rect 35840 7638 35892 7690
rect 40976 7638 41028 7690
rect 41040 7638 41092 7690
rect 41104 7638 41156 7690
rect 41168 7638 41220 7690
rect 6344 7094 6396 7146
rect 6408 7094 6460 7146
rect 6472 7094 6524 7146
rect 6536 7094 6588 7146
rect 38312 7094 38364 7146
rect 38376 7094 38428 7146
rect 38440 7094 38492 7146
rect 38504 7094 38556 7146
rect 3680 6550 3732 6602
rect 3744 6550 3796 6602
rect 3808 6550 3860 6602
rect 3872 6550 3924 6602
rect 35648 6550 35700 6602
rect 35712 6550 35764 6602
rect 35776 6550 35828 6602
rect 35840 6550 35892 6602
rect 40976 6550 41028 6602
rect 41040 6550 41092 6602
rect 41104 6550 41156 6602
rect 41168 6550 41220 6602
rect 6344 6006 6396 6058
rect 6408 6006 6460 6058
rect 6472 6006 6524 6058
rect 6536 6006 6588 6058
rect 38312 6006 38364 6058
rect 38376 6006 38428 6058
rect 38440 6006 38492 6058
rect 38504 6006 38556 6058
rect 3680 5462 3732 5514
rect 3744 5462 3796 5514
rect 3808 5462 3860 5514
rect 3872 5462 3924 5514
rect 35648 5462 35700 5514
rect 35712 5462 35764 5514
rect 35776 5462 35828 5514
rect 35840 5462 35892 5514
rect 40976 5462 41028 5514
rect 41040 5462 41092 5514
rect 41104 5462 41156 5514
rect 41168 5462 41220 5514
rect 6344 4918 6396 4970
rect 6408 4918 6460 4970
rect 6472 4918 6524 4970
rect 6536 4918 6588 4970
rect 38312 4918 38364 4970
rect 38376 4918 38428 4970
rect 38440 4918 38492 4970
rect 38504 4918 38556 4970
rect 3680 4374 3732 4426
rect 3744 4374 3796 4426
rect 3808 4374 3860 4426
rect 3872 4374 3924 4426
rect 35648 4374 35700 4426
rect 35712 4374 35764 4426
rect 35776 4374 35828 4426
rect 35840 4374 35892 4426
rect 40976 4374 41028 4426
rect 41040 4374 41092 4426
rect 41104 4374 41156 4426
rect 41168 4374 41220 4426
rect 6344 3830 6396 3882
rect 6408 3830 6460 3882
rect 6472 3830 6524 3882
rect 6536 3830 6588 3882
rect 38312 3830 38364 3882
rect 38376 3830 38428 3882
rect 38440 3830 38492 3882
rect 38504 3830 38556 3882
rect 3680 3286 3732 3338
rect 3744 3286 3796 3338
rect 3808 3286 3860 3338
rect 3872 3286 3924 3338
rect 35648 3286 35700 3338
rect 35712 3286 35764 3338
rect 35776 3286 35828 3338
rect 35840 3286 35892 3338
rect 40976 3286 41028 3338
rect 41040 3286 41092 3338
rect 41104 3286 41156 3338
rect 41168 3286 41220 3338
rect 6344 2742 6396 2794
rect 6408 2742 6460 2794
rect 6472 2742 6524 2794
rect 6536 2742 6588 2794
rect 38312 2742 38364 2794
rect 38376 2742 38428 2794
rect 38440 2742 38492 2794
rect 38504 2742 38556 2794
rect 43246 2640 43298 2692
rect 31378 2300 31430 2352
rect 3680 2198 3732 2250
rect 3744 2198 3796 2250
rect 3808 2198 3860 2250
rect 3872 2198 3924 2250
rect 35648 2198 35700 2250
rect 35712 2198 35764 2250
rect 35776 2198 35828 2250
rect 35840 2198 35892 2250
rect 40976 2198 41028 2250
rect 41040 2198 41092 2250
rect 41104 2198 41156 2250
rect 41168 2198 41220 2250
rect 7090 2096 7142 2148
rect 31378 2096 31430 2148
rect 6344 1654 6396 1706
rect 6408 1654 6460 1706
rect 6472 1654 6524 1706
rect 6536 1654 6588 1706
rect 38312 1654 38364 1706
rect 38376 1654 38428 1706
rect 38440 1654 38492 1706
rect 38504 1654 38556 1706
rect 3680 1110 3732 1162
rect 3744 1110 3796 1162
rect 3808 1110 3860 1162
rect 3872 1110 3924 1162
rect 35648 1110 35700 1162
rect 35712 1110 35764 1162
rect 35776 1110 35828 1162
rect 35840 1110 35892 1162
rect 40976 1110 41028 1162
rect 41040 1110 41092 1162
rect 41104 1110 41156 1162
rect 41168 1110 41220 1162
rect 6344 566 6396 618
rect 6408 566 6460 618
rect 6472 566 6524 618
rect 6536 566 6588 618
rect 38312 566 38364 618
rect 38376 566 38428 618
rect 38440 566 38492 618
rect 38504 566 38556 618
rect 3680 22 3732 74
rect 3744 22 3796 74
rect 3808 22 3860 74
rect 3872 22 3924 74
rect 35648 22 35700 74
rect 35712 22 35764 74
rect 35776 22 35828 74
rect 35840 22 35892 74
rect 40976 22 41028 74
rect 41040 22 41092 74
rect 41104 22 41156 74
rect 41168 22 41220 74
<< metal2 >>
rect 4 43312 60 44112
rect 1200 43312 1256 44112
rect 2396 43312 2452 44112
rect 3592 43312 3648 44112
rect 4880 43312 4936 44112
rect 6076 43312 6132 44112
rect 7272 43312 7328 44112
rect 8468 43312 8524 44112
rect 9756 43312 9812 44112
rect 10952 43312 11008 44112
rect 12148 43312 12204 44112
rect 13436 43312 13492 44112
rect 14632 43312 14688 44112
rect 15828 43312 15884 44112
rect 17024 43312 17080 44112
rect 18312 43312 18368 44112
rect 19508 43312 19564 44112
rect 20704 43312 20760 44112
rect 21992 43312 22048 44112
rect 23188 43312 23244 44112
rect 24384 43312 24440 44112
rect 25580 43312 25636 44112
rect 26868 43312 26924 44112
rect 28064 43312 28120 44112
rect 29260 43312 29316 44112
rect 30548 43312 30604 44112
rect 31744 43312 31800 44112
rect 32940 43312 32996 44112
rect 34136 43312 34192 44112
rect 35424 43312 35480 44112
rect 36620 43312 36676 44112
rect 37816 43312 37872 44112
rect 39104 43312 39160 44112
rect 40300 43312 40356 44112
rect 41496 43312 41552 44112
rect 42692 43312 42748 44112
rect 43980 43312 44036 44112
rect 45176 43312 45232 44112
rect 46372 43312 46428 44112
rect 47660 43312 47716 44112
rect 48856 43312 48912 44112
rect 50052 43312 50108 44112
rect 51248 43312 51304 44112
rect 52536 43312 52592 44112
rect 53732 43312 53788 44112
rect 54928 43312 54984 44112
rect 56124 43312 56180 44112
rect 57412 43312 57468 44112
rect 58608 43312 58664 44112
rect 59804 43312 59860 44112
rect 61092 43312 61148 44112
rect 62288 43312 62344 44112
rect 63484 43312 63540 44112
rect 64680 43312 64736 44112
rect 65968 43312 66024 44112
rect 67164 43312 67220 44112
rect 68360 43312 68416 44112
rect 69648 43312 69704 44112
rect 70844 43312 70900 44112
rect 72040 43312 72096 44112
rect 73236 43312 73292 44112
rect 74524 43312 74580 44112
rect 75720 43312 75776 44112
rect 76916 43312 76972 44112
rect 78204 43312 78260 44112
rect 79400 43312 79456 44112
rect 80596 43312 80652 44112
rect 81792 43312 81848 44112
rect 83080 43312 83136 44112
rect 84276 43312 84332 44112
rect 85472 43312 85528 44112
rect 86760 43312 86816 44112
rect 87956 43312 88012 44112
rect 89152 43312 89208 44112
rect 90348 43312 90404 44112
rect 91636 43312 91692 44112
rect 92832 43312 92888 44112
rect 94028 43312 94084 44112
rect 18 40642 46 43312
rect 1214 43242 1242 43312
rect 846 43214 1242 43242
rect 6 40636 58 40642
rect 6 40578 58 40584
rect 846 31530 874 43214
rect 2410 41322 2438 43312
rect 3606 41610 3634 43312
rect 3606 41582 4094 41610
rect 3502 41520 3554 41526
rect 3502 41462 3554 41468
rect 3514 41322 3542 41462
rect 3654 41420 3950 41440
rect 3710 41418 3734 41420
rect 3790 41418 3814 41420
rect 3870 41418 3894 41420
rect 3732 41366 3734 41418
rect 3796 41366 3808 41418
rect 3870 41366 3872 41418
rect 3710 41364 3734 41366
rect 3790 41364 3814 41366
rect 3870 41364 3894 41366
rect 3654 41344 3950 41364
rect 2398 41316 2450 41322
rect 2398 41258 2450 41264
rect 3502 41316 3554 41322
rect 3502 41258 3554 41264
rect 3502 41112 3554 41118
rect 3502 41054 3554 41060
rect 3514 40778 3542 41054
rect 3502 40772 3554 40778
rect 3502 40714 3554 40720
rect 3514 40642 3542 40714
rect 4066 40642 4094 41582
rect 4606 41112 4658 41118
rect 4606 41054 4658 41060
rect 3502 40636 3554 40642
rect 3502 40578 3554 40584
rect 4054 40636 4106 40642
rect 4054 40578 4106 40584
rect 2490 40432 2542 40438
rect 3514 40386 3542 40578
rect 4618 40506 4646 41054
rect 4894 40574 4922 43312
rect 6090 43242 6118 43312
rect 5446 43214 6118 43242
rect 5066 40636 5118 40642
rect 5066 40578 5118 40584
rect 4882 40568 4934 40574
rect 4882 40510 4934 40516
rect 4606 40500 4658 40506
rect 4606 40442 4658 40448
rect 2490 40374 2542 40380
rect 2502 40234 2530 40374
rect 3422 40358 3542 40386
rect 2490 40228 2542 40234
rect 2490 40170 2542 40176
rect 2490 39004 2542 39010
rect 2490 38946 2542 38952
rect 2214 38936 2266 38942
rect 2214 38878 2266 38884
rect 2226 37854 2254 38878
rect 2502 38602 2530 38946
rect 3422 38942 3450 40358
rect 3654 40332 3950 40352
rect 3710 40330 3734 40332
rect 3790 40330 3814 40332
rect 3870 40330 3894 40332
rect 3732 40278 3734 40330
rect 3796 40278 3808 40330
rect 3870 40278 3872 40330
rect 3710 40276 3734 40278
rect 3790 40276 3814 40278
rect 3870 40276 3894 40278
rect 3654 40256 3950 40276
rect 4618 39690 4646 40442
rect 4606 39684 4658 39690
rect 4606 39626 4658 39632
rect 3502 39480 3554 39486
rect 3502 39422 3554 39428
rect 3514 39010 3542 39422
rect 3654 39244 3950 39264
rect 3710 39242 3734 39244
rect 3790 39242 3814 39244
rect 3870 39242 3894 39244
rect 3732 39190 3734 39242
rect 3796 39190 3808 39242
rect 3870 39190 3872 39242
rect 3710 39188 3734 39190
rect 3790 39188 3814 39190
rect 3870 39188 3894 39190
rect 3654 39168 3950 39188
rect 3502 39004 3554 39010
rect 3502 38946 3554 38952
rect 3410 38936 3462 38942
rect 3410 38878 3462 38884
rect 3422 38806 3450 38878
rect 4330 38868 4382 38874
rect 4330 38810 4382 38816
rect 3410 38800 3462 38806
rect 3410 38742 3462 38748
rect 4054 38800 4106 38806
rect 4054 38742 4106 38748
rect 2490 38596 2542 38602
rect 2490 38538 2542 38544
rect 4066 38398 4094 38742
rect 4342 38466 4370 38810
rect 4330 38460 4382 38466
rect 4330 38402 4382 38408
rect 2398 38392 2450 38398
rect 2398 38334 2450 38340
rect 4054 38392 4106 38398
rect 4054 38334 4106 38340
rect 2410 37854 2438 38334
rect 3654 38156 3950 38176
rect 3710 38154 3734 38156
rect 3790 38154 3814 38156
rect 3870 38154 3894 38156
rect 3732 38102 3734 38154
rect 3796 38102 3808 38154
rect 3870 38102 3872 38154
rect 3710 38100 3734 38102
rect 3790 38100 3814 38102
rect 3870 38100 3894 38102
rect 3654 38080 3950 38100
rect 4066 37938 4094 38334
rect 3974 37910 4094 37938
rect 2214 37848 2266 37854
rect 2214 37790 2266 37796
rect 2398 37848 2450 37854
rect 2398 37790 2450 37796
rect 2410 36970 2438 37790
rect 3974 37718 4002 37910
rect 4422 37780 4474 37786
rect 4422 37722 4474 37728
rect 3962 37712 4014 37718
rect 3962 37654 4014 37660
rect 3974 37514 4002 37654
rect 3134 37508 3186 37514
rect 3134 37450 3186 37456
rect 3962 37508 4014 37514
rect 3962 37450 4014 37456
rect 2398 36964 2450 36970
rect 2398 36906 2450 36912
rect 3146 36834 3174 37450
rect 4434 37378 4462 37722
rect 4422 37372 4474 37378
rect 4422 37314 4474 37320
rect 3654 37068 3950 37088
rect 3710 37066 3734 37068
rect 3790 37066 3814 37068
rect 3870 37066 3894 37068
rect 3732 37014 3734 37066
rect 3796 37014 3808 37066
rect 3870 37014 3872 37066
rect 3710 37012 3734 37014
rect 3790 37012 3814 37014
rect 3870 37012 3894 37014
rect 3654 36992 3950 37012
rect 3134 36828 3186 36834
rect 3134 36770 3186 36776
rect 2490 36760 2542 36766
rect 2490 36702 2542 36708
rect 3410 36760 3462 36766
rect 3410 36702 3462 36708
rect 2502 36426 2530 36702
rect 3422 36426 3450 36702
rect 4974 36624 5026 36630
rect 4974 36566 5026 36572
rect 4986 36426 5014 36566
rect 2490 36420 2542 36426
rect 2490 36362 2542 36368
rect 3410 36420 3462 36426
rect 3410 36362 3462 36368
rect 4974 36420 5026 36426
rect 4974 36362 5026 36368
rect 2674 36216 2726 36222
rect 2674 36158 2726 36164
rect 2686 35746 2714 36158
rect 3654 35980 3950 36000
rect 3710 35978 3734 35980
rect 3790 35978 3814 35980
rect 3870 35978 3894 35980
rect 3732 35926 3734 35978
rect 3796 35926 3808 35978
rect 3870 35926 3872 35978
rect 3710 35924 3734 35926
rect 3790 35924 3814 35926
rect 3870 35924 3894 35926
rect 3654 35904 3950 35924
rect 2674 35740 2726 35746
rect 2674 35682 2726 35688
rect 2686 35338 2714 35682
rect 3962 35536 4014 35542
rect 3962 35478 4014 35484
rect 4238 35536 4290 35542
rect 4238 35478 4290 35484
rect 2674 35332 2726 35338
rect 2674 35274 2726 35280
rect 3974 35202 4002 35478
rect 2582 35196 2634 35202
rect 2582 35138 2634 35144
rect 3962 35196 4014 35202
rect 3962 35138 4014 35144
rect 2594 34590 2622 35138
rect 4250 35134 4278 35478
rect 4238 35128 4290 35134
rect 4238 35070 4290 35076
rect 3654 34892 3950 34912
rect 3710 34890 3734 34892
rect 3790 34890 3814 34892
rect 3870 34890 3894 34892
rect 3732 34838 3734 34890
rect 3796 34838 3808 34890
rect 3870 34838 3872 34890
rect 3710 34836 3734 34838
rect 3790 34836 3814 34838
rect 3870 34836 3894 34838
rect 3654 34816 3950 34836
rect 4250 34794 4278 35070
rect 4238 34788 4290 34794
rect 4238 34730 4290 34736
rect 2582 34584 2634 34590
rect 2582 34526 2634 34532
rect 3226 34584 3278 34590
rect 3226 34526 3278 34532
rect 2594 33706 2622 34526
rect 2582 33700 2634 33706
rect 2582 33642 2634 33648
rect 3238 33434 3266 34526
rect 3870 34448 3922 34454
rect 3870 34390 3922 34396
rect 3882 34114 3910 34390
rect 3870 34108 3922 34114
rect 3870 34050 3922 34056
rect 4698 34040 4750 34046
rect 4698 33982 4750 33988
rect 3654 33804 3950 33824
rect 3710 33802 3734 33804
rect 3790 33802 3814 33804
rect 3870 33802 3894 33804
rect 3732 33750 3734 33802
rect 3796 33750 3808 33802
rect 3870 33750 3872 33802
rect 3710 33748 3734 33750
rect 3790 33748 3814 33750
rect 3870 33748 3894 33750
rect 3654 33728 3950 33748
rect 3502 33496 3554 33502
rect 3502 33438 3554 33444
rect 3226 33428 3278 33434
rect 3226 33370 3278 33376
rect 2766 32408 2818 32414
rect 2766 32350 2818 32356
rect 1662 32340 1714 32346
rect 1662 32282 1714 32288
rect 834 31524 886 31530
rect 834 31466 886 31472
rect 1674 31394 1702 32282
rect 2778 31530 2806 32350
rect 2766 31524 2818 31530
rect 2766 31466 2818 31472
rect 1662 31388 1714 31394
rect 1662 31330 1714 31336
rect 3238 30442 3266 33370
rect 3514 31802 3542 33438
rect 4710 33026 4738 33982
rect 4974 33360 5026 33366
rect 4974 33302 5026 33308
rect 4986 33026 5014 33302
rect 4698 33020 4750 33026
rect 4698 32962 4750 32968
rect 4974 33020 5026 33026
rect 4974 32962 5026 32968
rect 3654 32716 3950 32736
rect 3710 32714 3734 32716
rect 3790 32714 3814 32716
rect 3870 32714 3894 32716
rect 3732 32662 3734 32714
rect 3796 32662 3808 32714
rect 3870 32662 3872 32714
rect 3710 32660 3734 32662
rect 3790 32660 3814 32662
rect 3870 32660 3894 32662
rect 3654 32640 3950 32660
rect 4710 32550 4738 32962
rect 5078 32550 5106 40578
rect 5342 40432 5394 40438
rect 5342 40374 5394 40380
rect 5354 39554 5382 40374
rect 5342 39548 5394 39554
rect 5342 39490 5394 39496
rect 5446 39434 5474 43214
rect 6318 41964 6614 41984
rect 6374 41962 6398 41964
rect 6454 41962 6478 41964
rect 6534 41962 6558 41964
rect 6396 41910 6398 41962
rect 6460 41910 6472 41962
rect 6534 41910 6536 41962
rect 6374 41908 6398 41910
rect 6454 41908 6478 41910
rect 6534 41908 6558 41910
rect 6318 41888 6614 41908
rect 6170 41112 6222 41118
rect 6170 41054 6222 41060
rect 6182 40778 6210 41054
rect 6318 40876 6614 40896
rect 6374 40874 6398 40876
rect 6454 40874 6478 40876
rect 6534 40874 6558 40876
rect 6396 40822 6398 40874
rect 6460 40822 6472 40874
rect 6534 40822 6536 40874
rect 6374 40820 6398 40822
rect 6454 40820 6478 40822
rect 6534 40820 6558 40822
rect 6318 40800 6614 40820
rect 6170 40772 6222 40778
rect 6170 40714 6222 40720
rect 6182 40574 6210 40714
rect 7286 40658 7314 43312
rect 8482 43242 8510 43312
rect 8390 43214 8510 43242
rect 7826 40976 7878 40982
rect 7826 40918 7878 40924
rect 8010 40976 8062 40982
rect 8010 40918 8062 40924
rect 7286 40630 7406 40658
rect 7378 40574 7406 40630
rect 6170 40568 6222 40574
rect 6170 40510 6222 40516
rect 7366 40568 7418 40574
rect 7366 40510 7418 40516
rect 6182 40098 6210 40510
rect 7838 40098 7866 40918
rect 8022 40642 8050 40918
rect 8010 40636 8062 40642
rect 8010 40578 8062 40584
rect 8022 40522 8050 40578
rect 8022 40494 8142 40522
rect 8010 40432 8062 40438
rect 8010 40374 8062 40380
rect 8022 40098 8050 40374
rect 8114 40166 8142 40494
rect 8102 40160 8154 40166
rect 8102 40102 8154 40108
rect 6170 40092 6222 40098
rect 6170 40034 6222 40040
rect 7826 40092 7878 40098
rect 7826 40034 7878 40040
rect 8010 40092 8062 40098
rect 8010 40034 8062 40040
rect 8114 40030 8142 40102
rect 8102 40024 8154 40030
rect 8102 39966 8154 39972
rect 8010 39956 8062 39962
rect 8010 39898 8062 39904
rect 6318 39788 6614 39808
rect 6374 39786 6398 39788
rect 6454 39786 6478 39788
rect 6534 39786 6558 39788
rect 6396 39734 6398 39786
rect 6460 39734 6472 39786
rect 6534 39734 6536 39786
rect 6374 39732 6398 39734
rect 6454 39732 6478 39734
rect 6534 39732 6558 39734
rect 6318 39712 6614 39732
rect 5354 39406 5474 39434
rect 5158 33496 5210 33502
rect 5158 33438 5210 33444
rect 5170 32618 5198 33438
rect 5158 32612 5210 32618
rect 5158 32554 5210 32560
rect 4698 32544 4750 32550
rect 4698 32486 4750 32492
rect 5066 32544 5118 32550
rect 5066 32486 5118 32492
rect 4974 31932 5026 31938
rect 4974 31874 5026 31880
rect 3502 31796 3554 31802
rect 3502 31738 3554 31744
rect 3514 31530 3542 31738
rect 3654 31628 3950 31648
rect 3710 31626 3734 31628
rect 3790 31626 3814 31628
rect 3870 31626 3894 31628
rect 3732 31574 3734 31626
rect 3796 31574 3808 31626
rect 3870 31574 3872 31626
rect 3710 31572 3734 31574
rect 3790 31572 3814 31574
rect 3870 31572 3894 31574
rect 3654 31552 3950 31572
rect 3502 31524 3554 31530
rect 3502 31466 3554 31472
rect 3514 31394 3542 31466
rect 3502 31388 3554 31394
rect 3502 31330 3554 31336
rect 4882 31252 4934 31258
rect 4882 31194 4934 31200
rect 3654 30540 3950 30560
rect 3710 30538 3734 30540
rect 3790 30538 3814 30540
rect 3870 30538 3894 30540
rect 3732 30486 3734 30538
rect 3796 30486 3808 30538
rect 3870 30486 3872 30538
rect 3710 30484 3734 30486
rect 3790 30484 3814 30486
rect 3870 30484 3894 30486
rect 3654 30464 3950 30484
rect 3226 30436 3278 30442
rect 3226 30378 3278 30384
rect 2398 30300 2450 30306
rect 2398 30242 2450 30248
rect 2306 29008 2358 29014
rect 2306 28950 2358 28956
rect 2318 28130 2346 28950
rect 926 28124 978 28130
rect 926 28066 978 28072
rect 2306 28124 2358 28130
rect 2306 28066 2358 28072
rect 938 27586 966 28066
rect 1938 28056 1990 28062
rect 1938 27998 1990 28004
rect 1950 27722 1978 27998
rect 1938 27716 1990 27722
rect 1938 27658 1990 27664
rect 926 27580 978 27586
rect 926 27522 978 27528
rect 2410 20650 2438 30242
rect 3042 30232 3094 30238
rect 3042 30174 3094 30180
rect 2950 30096 3002 30102
rect 2950 30038 3002 30044
rect 2962 29014 2990 30038
rect 3054 29354 3082 30174
rect 4330 29552 4382 29558
rect 4330 29494 4382 29500
rect 3654 29452 3950 29472
rect 3710 29450 3734 29452
rect 3790 29450 3814 29452
rect 3870 29450 3894 29452
rect 3732 29398 3734 29450
rect 3796 29398 3808 29450
rect 3870 29398 3872 29450
rect 3710 29396 3734 29398
rect 3790 29396 3814 29398
rect 3870 29396 3894 29398
rect 3654 29376 3950 29396
rect 3042 29348 3094 29354
rect 3042 29290 3094 29296
rect 3042 29144 3094 29150
rect 3042 29086 3094 29092
rect 2950 29008 3002 29014
rect 2950 28950 3002 28956
rect 3054 28266 3082 29086
rect 3654 28364 3950 28384
rect 3710 28362 3734 28364
rect 3790 28362 3814 28364
rect 3870 28362 3894 28364
rect 3732 28310 3734 28362
rect 3796 28310 3808 28362
rect 3870 28310 3872 28362
rect 3710 28308 3734 28310
rect 3790 28308 3814 28310
rect 3870 28308 3894 28310
rect 3654 28288 3950 28308
rect 3042 28260 3094 28266
rect 3042 28202 3094 28208
rect 4054 27920 4106 27926
rect 4054 27862 4106 27868
rect 2950 27376 3002 27382
rect 2950 27318 3002 27324
rect 2962 27042 2990 27318
rect 3654 27276 3950 27296
rect 3710 27274 3734 27276
rect 3790 27274 3814 27276
rect 3870 27274 3894 27276
rect 3732 27222 3734 27274
rect 3796 27222 3808 27274
rect 3870 27222 3872 27274
rect 3710 27220 3734 27222
rect 3790 27220 3814 27222
rect 3870 27220 3894 27222
rect 3654 27200 3950 27220
rect 4066 27178 4094 27862
rect 4238 27376 4290 27382
rect 4238 27318 4290 27324
rect 4054 27172 4106 27178
rect 3974 27132 4054 27160
rect 2950 27036 3002 27042
rect 2950 26978 3002 26984
rect 3974 26634 4002 27132
rect 4054 27114 4106 27120
rect 4054 26968 4106 26974
rect 4054 26910 4106 26916
rect 3962 26628 4014 26634
rect 3962 26570 4014 26576
rect 3502 26288 3554 26294
rect 3502 26230 3554 26236
rect 3514 25886 3542 26230
rect 3654 26188 3950 26208
rect 3710 26186 3734 26188
rect 3790 26186 3814 26188
rect 3870 26186 3894 26188
rect 3732 26134 3734 26186
rect 3796 26134 3808 26186
rect 3870 26134 3872 26186
rect 3710 26132 3734 26134
rect 3790 26132 3814 26134
rect 3870 26132 3894 26134
rect 3654 26112 3950 26132
rect 4066 26090 4094 26910
rect 4054 26084 4106 26090
rect 4054 26026 4106 26032
rect 4250 26022 4278 27318
rect 4238 26016 4290 26022
rect 4238 25958 4290 25964
rect 2766 25880 2818 25886
rect 2766 25822 2818 25828
rect 3502 25880 3554 25886
rect 3502 25822 3554 25828
rect 2778 25478 2806 25822
rect 2766 25472 2818 25478
rect 2766 25414 2818 25420
rect 4238 25472 4290 25478
rect 4238 25414 4290 25420
rect 2778 25002 2806 25414
rect 4146 25268 4198 25274
rect 4146 25210 4198 25216
rect 4054 25200 4106 25206
rect 4054 25142 4106 25148
rect 3654 25100 3950 25120
rect 3710 25098 3734 25100
rect 3790 25098 3814 25100
rect 3870 25098 3894 25100
rect 3732 25046 3734 25098
rect 3796 25046 3808 25098
rect 3870 25046 3872 25098
rect 3710 25044 3734 25046
rect 3790 25044 3814 25046
rect 3870 25044 3894 25046
rect 3654 25024 3950 25044
rect 2766 24996 2818 25002
rect 2766 24938 2818 24944
rect 3410 24860 3462 24866
rect 3410 24802 3462 24808
rect 2490 24384 2542 24390
rect 2490 24326 2542 24332
rect 2502 23710 2530 24326
rect 2490 23704 2542 23710
rect 2490 23646 2542 23652
rect 2674 23704 2726 23710
rect 2674 23646 2726 23652
rect 2686 22214 2714 23646
rect 3318 23568 3370 23574
rect 3318 23510 3370 23516
rect 3330 22690 3358 23510
rect 3422 23302 3450 24802
rect 4066 24730 4094 25142
rect 4054 24724 4106 24730
rect 4054 24666 4106 24672
rect 3686 24656 3738 24662
rect 3686 24598 3738 24604
rect 3698 24322 3726 24598
rect 4158 24322 4186 25210
rect 4250 24322 4278 25414
rect 3686 24316 3738 24322
rect 3686 24258 3738 24264
rect 4146 24316 4198 24322
rect 4146 24258 4198 24264
rect 4238 24316 4290 24322
rect 4238 24258 4290 24264
rect 3654 24012 3950 24032
rect 3710 24010 3734 24012
rect 3790 24010 3814 24012
rect 3870 24010 3894 24012
rect 3732 23958 3734 24010
rect 3796 23958 3808 24010
rect 3870 23958 3872 24010
rect 3710 23956 3734 23958
rect 3790 23956 3814 23958
rect 3870 23956 3894 23958
rect 3654 23936 3950 23956
rect 3594 23704 3646 23710
rect 3594 23646 3646 23652
rect 3606 23370 3634 23646
rect 3594 23364 3646 23370
rect 3594 23306 3646 23312
rect 3410 23296 3462 23302
rect 3410 23238 3462 23244
rect 3422 22690 3450 23238
rect 3502 23228 3554 23234
rect 3502 23170 3554 23176
rect 3514 23030 3542 23170
rect 3502 23024 3554 23030
rect 3502 22966 3554 22972
rect 3514 22758 3542 22966
rect 3654 22924 3950 22944
rect 3710 22922 3734 22924
rect 3790 22922 3814 22924
rect 3870 22922 3894 22924
rect 3732 22870 3734 22922
rect 3796 22870 3808 22922
rect 3870 22870 3872 22922
rect 3710 22868 3734 22870
rect 3790 22868 3814 22870
rect 3870 22868 3894 22870
rect 3654 22848 3950 22868
rect 3502 22752 3554 22758
rect 3500 22720 3502 22729
rect 3554 22720 3556 22729
rect 3318 22684 3370 22690
rect 3318 22626 3370 22632
rect 3410 22684 3462 22690
rect 3500 22655 3556 22664
rect 3410 22626 3462 22632
rect 3514 22629 3542 22655
rect 2674 22208 2726 22214
rect 2674 22150 2726 22156
rect 2686 21534 2714 22150
rect 2766 22140 2818 22146
rect 2766 22082 2818 22088
rect 2778 21942 2806 22082
rect 2766 21936 2818 21942
rect 2766 21878 2818 21884
rect 2778 21534 2806 21878
rect 2674 21528 2726 21534
rect 2674 21470 2726 21476
rect 2766 21528 2818 21534
rect 2766 21470 2818 21476
rect 2398 20644 2450 20650
rect 2398 20586 2450 20592
rect 2778 20446 2806 21470
rect 3318 21392 3370 21398
rect 3318 21334 3370 21340
rect 3330 20446 3358 21334
rect 3422 21058 3450 22626
rect 3594 22616 3646 22622
rect 3594 22558 3646 22564
rect 3606 22078 3634 22558
rect 3870 22276 3922 22282
rect 3870 22218 3922 22224
rect 3882 22078 3910 22218
rect 3594 22072 3646 22078
rect 3594 22014 3646 22020
rect 3870 22072 3922 22078
rect 3870 22014 3922 22020
rect 3654 21836 3950 21856
rect 3710 21834 3734 21836
rect 3790 21834 3814 21836
rect 3870 21834 3894 21836
rect 3732 21782 3734 21834
rect 3796 21782 3808 21834
rect 3870 21782 3872 21834
rect 3710 21780 3734 21782
rect 3790 21780 3814 21782
rect 3870 21780 3894 21782
rect 3654 21760 3950 21780
rect 3410 21052 3462 21058
rect 3410 20994 3462 21000
rect 3654 20748 3950 20768
rect 3710 20746 3734 20748
rect 3790 20746 3814 20748
rect 3870 20746 3894 20748
rect 3732 20694 3734 20746
rect 3796 20694 3808 20746
rect 3870 20694 3872 20746
rect 3710 20692 3734 20694
rect 3790 20692 3814 20694
rect 3870 20692 3894 20694
rect 3654 20672 3950 20692
rect 2766 20440 2818 20446
rect 2766 20382 2818 20388
rect 3318 20440 3370 20446
rect 3318 20382 3370 20388
rect 4238 20440 4290 20446
rect 4238 20382 4290 20388
rect 3594 20372 3646 20378
rect 3594 20314 3646 20320
rect 4054 20372 4106 20378
rect 4054 20314 4106 20320
rect 3606 19850 3634 20314
rect 3514 19822 3634 19850
rect 3514 19442 3542 19822
rect 3654 19660 3950 19680
rect 3710 19658 3734 19660
rect 3790 19658 3814 19660
rect 3870 19658 3894 19660
rect 3732 19606 3734 19658
rect 3796 19606 3808 19658
rect 3870 19606 3872 19658
rect 3710 19604 3734 19606
rect 3790 19604 3814 19606
rect 3870 19604 3894 19606
rect 3654 19584 3950 19604
rect 3514 19414 3634 19442
rect 4066 19426 4094 20314
rect 4250 19562 4278 20382
rect 4238 19556 4290 19562
rect 4238 19498 4290 19504
rect 3502 19216 3554 19222
rect 3502 19158 3554 19164
rect 3514 18270 3542 19158
rect 3606 18882 3634 19414
rect 4054 19420 4106 19426
rect 4054 19362 4106 19368
rect 4146 19352 4198 19358
rect 4144 19320 4146 19329
rect 4198 19320 4200 19329
rect 4144 19255 4200 19264
rect 4342 18950 4370 29494
rect 4698 29280 4750 29286
rect 4698 29222 4750 29228
rect 4606 27104 4658 27110
rect 4606 27046 4658 27052
rect 4422 26968 4474 26974
rect 4422 26910 4474 26916
rect 4434 22622 4462 26910
rect 4514 26016 4566 26022
rect 4514 25958 4566 25964
rect 4422 22616 4474 22622
rect 4422 22558 4474 22564
rect 4422 22480 4474 22486
rect 4422 22422 4474 22428
rect 4434 22214 4462 22422
rect 4422 22208 4474 22214
rect 4422 22150 4474 22156
rect 4526 21738 4554 25958
rect 4618 25342 4646 27046
rect 4710 26974 4738 29222
rect 4790 27444 4842 27450
rect 4790 27386 4842 27392
rect 4698 26968 4750 26974
rect 4698 26910 4750 26916
rect 4802 26838 4830 27386
rect 4790 26832 4842 26838
rect 4790 26774 4842 26780
rect 4606 25336 4658 25342
rect 4606 25278 4658 25284
rect 4618 22282 4646 25278
rect 4698 24792 4750 24798
rect 4698 24734 4750 24740
rect 4710 24458 4738 24734
rect 4698 24452 4750 24458
rect 4698 24394 4750 24400
rect 4802 24338 4830 26774
rect 4710 24310 4830 24338
rect 4606 22276 4658 22282
rect 4606 22218 4658 22224
rect 4514 21732 4566 21738
rect 4514 21674 4566 21680
rect 4330 18944 4382 18950
rect 4330 18886 4382 18892
rect 3594 18876 3646 18882
rect 3594 18818 3646 18824
rect 4422 18876 4474 18882
rect 4422 18818 4474 18824
rect 3654 18572 3950 18592
rect 3710 18570 3734 18572
rect 3790 18570 3814 18572
rect 3870 18570 3894 18572
rect 3732 18518 3734 18570
rect 3796 18518 3808 18570
rect 3870 18518 3872 18570
rect 3710 18516 3734 18518
rect 3790 18516 3814 18518
rect 3870 18516 3894 18518
rect 3654 18496 3950 18516
rect 3502 18264 3554 18270
rect 3502 18206 3554 18212
rect 4434 17930 4462 18818
rect 4606 18740 4658 18746
rect 4606 18682 4658 18688
rect 4618 18338 4646 18682
rect 4606 18332 4658 18338
rect 4606 18274 4658 18280
rect 4422 17924 4474 17930
rect 4422 17866 4474 17872
rect 3654 17484 3950 17504
rect 3710 17482 3734 17484
rect 3790 17482 3814 17484
rect 3870 17482 3894 17484
rect 3732 17430 3734 17482
rect 3796 17430 3808 17482
rect 3870 17430 3872 17482
rect 3710 17428 3734 17430
rect 3790 17428 3814 17430
rect 3870 17428 3894 17430
rect 3654 17408 3950 17428
rect 4710 16842 4738 24310
rect 4698 16836 4750 16842
rect 4698 16778 4750 16784
rect 3654 16396 3950 16416
rect 3710 16394 3734 16396
rect 3790 16394 3814 16396
rect 3870 16394 3894 16396
rect 3732 16342 3734 16394
rect 3796 16342 3808 16394
rect 3870 16342 3872 16394
rect 3710 16340 3734 16342
rect 3790 16340 3814 16342
rect 3870 16340 3894 16342
rect 3654 16320 3950 16340
rect 4710 16298 4738 16778
rect 4698 16292 4750 16298
rect 4698 16234 4750 16240
rect 4710 16094 4738 16234
rect 4894 16230 4922 31194
rect 4986 30986 5014 31874
rect 5078 31546 5106 32486
rect 5354 32074 5382 39406
rect 8022 39010 8050 39898
rect 8010 39004 8062 39010
rect 8010 38946 8062 38952
rect 8102 38868 8154 38874
rect 8102 38810 8154 38816
rect 6318 38700 6614 38720
rect 6374 38698 6398 38700
rect 6454 38698 6478 38700
rect 6534 38698 6558 38700
rect 6396 38646 6398 38698
rect 6460 38646 6472 38698
rect 6534 38646 6536 38698
rect 6374 38644 6398 38646
rect 6454 38644 6478 38646
rect 6534 38644 6558 38646
rect 6318 38624 6614 38644
rect 7642 38392 7694 38398
rect 7642 38334 7694 38340
rect 5894 38256 5946 38262
rect 5894 38198 5946 38204
rect 5906 37514 5934 38198
rect 7458 37848 7510 37854
rect 7458 37790 7510 37796
rect 6318 37612 6614 37632
rect 6374 37610 6398 37612
rect 6454 37610 6478 37612
rect 6534 37610 6558 37612
rect 6396 37558 6398 37610
rect 6460 37558 6472 37610
rect 6534 37558 6536 37610
rect 6374 37556 6398 37558
rect 6454 37556 6478 37558
rect 6534 37556 6558 37558
rect 6318 37536 6614 37556
rect 7470 37514 7498 37790
rect 5894 37508 5946 37514
rect 5894 37450 5946 37456
rect 7458 37508 7510 37514
rect 7458 37450 7510 37456
rect 5802 36692 5854 36698
rect 5802 36634 5854 36640
rect 5814 36290 5842 36634
rect 6318 36524 6614 36544
rect 6374 36522 6398 36524
rect 6454 36522 6478 36524
rect 6534 36522 6558 36524
rect 6396 36470 6398 36522
rect 6460 36470 6472 36522
rect 6534 36470 6536 36522
rect 6374 36468 6398 36470
rect 6454 36468 6478 36470
rect 6534 36468 6558 36470
rect 6318 36448 6614 36468
rect 7470 36426 7498 37450
rect 7654 37446 7682 38334
rect 8114 37922 8142 38810
rect 8102 37916 8154 37922
rect 8102 37858 8154 37864
rect 7642 37440 7694 37446
rect 7642 37382 7694 37388
rect 7458 36420 7510 36426
rect 7458 36362 7510 36368
rect 5802 36284 5854 36290
rect 5802 36226 5854 36232
rect 6318 35436 6614 35456
rect 6374 35434 6398 35436
rect 6454 35434 6478 35436
rect 6534 35434 6558 35436
rect 6396 35382 6398 35434
rect 6460 35382 6472 35434
rect 6534 35382 6536 35434
rect 6374 35380 6398 35382
rect 6454 35380 6478 35382
rect 6534 35380 6558 35382
rect 6318 35360 6614 35380
rect 8390 34998 8418 43214
rect 8982 41420 9278 41440
rect 9038 41418 9062 41420
rect 9118 41418 9142 41420
rect 9198 41418 9222 41420
rect 9060 41366 9062 41418
rect 9124 41366 9136 41418
rect 9198 41366 9200 41418
rect 9038 41364 9062 41366
rect 9118 41364 9142 41366
rect 9198 41364 9222 41366
rect 8982 41344 9278 41364
rect 9770 40642 9798 43312
rect 9758 40636 9810 40642
rect 9758 40578 9810 40584
rect 8982 40332 9278 40352
rect 9038 40330 9062 40332
rect 9118 40330 9142 40332
rect 9198 40330 9222 40332
rect 9060 40278 9062 40330
rect 9124 40278 9136 40330
rect 9198 40278 9200 40330
rect 9038 40276 9062 40278
rect 9118 40276 9142 40278
rect 9198 40276 9222 40278
rect 8982 40256 9278 40276
rect 10966 39690 10994 43312
rect 11646 41964 11942 41984
rect 11702 41962 11726 41964
rect 11782 41962 11806 41964
rect 11862 41962 11886 41964
rect 11724 41910 11726 41962
rect 11788 41910 11800 41962
rect 11862 41910 11864 41962
rect 11702 41908 11726 41910
rect 11782 41908 11806 41910
rect 11862 41908 11886 41910
rect 11646 41888 11942 41908
rect 11646 40876 11942 40896
rect 11702 40874 11726 40876
rect 11782 40874 11806 40876
rect 11862 40874 11886 40876
rect 11724 40822 11726 40874
rect 11788 40822 11800 40874
rect 11862 40822 11864 40874
rect 11702 40820 11726 40822
rect 11782 40820 11806 40822
rect 11862 40820 11886 40822
rect 11646 40800 11942 40820
rect 11046 40568 11098 40574
rect 11046 40510 11098 40516
rect 11058 40166 11086 40510
rect 12162 40506 12190 43312
rect 12334 41112 12386 41118
rect 12334 41054 12386 41060
rect 13450 41066 13478 43312
rect 14310 41420 14606 41440
rect 14366 41418 14390 41420
rect 14446 41418 14470 41420
rect 14526 41418 14550 41420
rect 14388 41366 14390 41418
rect 14452 41366 14464 41418
rect 14526 41366 14528 41418
rect 14366 41364 14390 41366
rect 14446 41364 14470 41366
rect 14526 41364 14550 41366
rect 14310 41344 14606 41364
rect 12150 40500 12202 40506
rect 12150 40442 12202 40448
rect 12346 40234 12374 41054
rect 13070 41044 13122 41050
rect 13450 41038 13570 41066
rect 13070 40986 13122 40992
rect 13082 40438 13110 40986
rect 13438 40976 13490 40982
rect 13438 40918 13490 40924
rect 13450 40642 13478 40918
rect 13438 40636 13490 40642
rect 13438 40578 13490 40584
rect 13070 40432 13122 40438
rect 13070 40374 13122 40380
rect 11966 40228 12018 40234
rect 11966 40170 12018 40176
rect 12334 40228 12386 40234
rect 12334 40170 12386 40176
rect 11046 40160 11098 40166
rect 11046 40102 11098 40108
rect 11058 40030 11086 40102
rect 11046 40024 11098 40030
rect 11046 39966 11098 39972
rect 11646 39788 11942 39808
rect 11702 39786 11726 39788
rect 11782 39786 11806 39788
rect 11862 39786 11886 39788
rect 11724 39734 11726 39786
rect 11788 39734 11800 39786
rect 11862 39734 11864 39786
rect 11702 39732 11726 39734
rect 11782 39732 11806 39734
rect 11862 39732 11886 39734
rect 11646 39712 11942 39732
rect 10954 39684 11006 39690
rect 10954 39626 11006 39632
rect 11506 39480 11558 39486
rect 11506 39422 11558 39428
rect 8982 39244 9278 39264
rect 9038 39242 9062 39244
rect 9118 39242 9142 39244
rect 9198 39242 9222 39244
rect 9060 39190 9062 39242
rect 9124 39190 9136 39242
rect 9198 39190 9200 39242
rect 9038 39188 9062 39190
rect 9118 39188 9142 39190
rect 9198 39188 9222 39190
rect 8982 39168 9278 39188
rect 8654 39004 8706 39010
rect 8654 38946 8706 38952
rect 8666 37990 8694 38946
rect 9114 38936 9166 38942
rect 9114 38878 9166 38884
rect 9126 38806 9154 38878
rect 9758 38868 9810 38874
rect 9758 38810 9810 38816
rect 9114 38800 9166 38806
rect 9114 38742 9166 38748
rect 9482 38800 9534 38806
rect 9482 38742 9534 38748
rect 9298 38460 9350 38466
rect 9298 38402 9350 38408
rect 8982 38156 9278 38176
rect 9038 38154 9062 38156
rect 9118 38154 9142 38156
rect 9198 38154 9222 38156
rect 9060 38102 9062 38154
rect 9124 38102 9136 38154
rect 9198 38102 9200 38154
rect 9038 38100 9062 38102
rect 9118 38100 9142 38102
rect 9198 38100 9222 38102
rect 8982 38080 9278 38100
rect 9310 38058 9338 38402
rect 9298 38052 9350 38058
rect 9298 37994 9350 38000
rect 8654 37984 8706 37990
rect 9114 37984 9166 37990
rect 8654 37926 8706 37932
rect 9112 37952 9114 37961
rect 9166 37952 9168 37961
rect 9112 37887 9168 37896
rect 8982 37068 9278 37088
rect 9038 37066 9062 37068
rect 9118 37066 9142 37068
rect 9198 37066 9222 37068
rect 9060 37014 9062 37066
rect 9124 37014 9136 37066
rect 9198 37014 9200 37066
rect 9038 37012 9062 37014
rect 9118 37012 9142 37014
rect 9198 37012 9222 37014
rect 8982 36992 9278 37012
rect 9494 36630 9522 38742
rect 9770 38058 9798 38810
rect 10310 38392 10362 38398
rect 10310 38334 10362 38340
rect 9758 38052 9810 38058
rect 9758 37994 9810 38000
rect 9482 36624 9534 36630
rect 9482 36566 9534 36572
rect 8982 35980 9278 36000
rect 9038 35978 9062 35980
rect 9118 35978 9142 35980
rect 9198 35978 9222 35980
rect 9060 35926 9062 35978
rect 9124 35926 9136 35978
rect 9198 35926 9200 35978
rect 9038 35924 9062 35926
rect 9118 35924 9142 35926
rect 9198 35924 9222 35926
rect 8982 35904 9278 35924
rect 7090 34992 7142 34998
rect 7090 34934 7142 34940
rect 8378 34992 8430 34998
rect 8378 34934 8430 34940
rect 6630 34516 6682 34522
rect 6630 34458 6682 34464
rect 6318 34348 6614 34368
rect 6374 34346 6398 34348
rect 6454 34346 6478 34348
rect 6534 34346 6558 34348
rect 6396 34294 6398 34346
rect 6460 34294 6472 34346
rect 6534 34294 6536 34346
rect 6374 34292 6398 34294
rect 6454 34292 6478 34294
rect 6534 34292 6558 34294
rect 6318 34272 6614 34292
rect 6642 34182 6670 34458
rect 6630 34176 6682 34182
rect 6630 34118 6682 34124
rect 6642 33502 6670 34118
rect 7102 33978 7130 34934
rect 7090 33972 7142 33978
rect 7090 33914 7142 33920
rect 7102 33502 7130 33914
rect 6630 33496 6682 33502
rect 6630 33438 6682 33444
rect 7090 33496 7142 33502
rect 7090 33438 7142 33444
rect 6170 33428 6222 33434
rect 6170 33370 6222 33376
rect 6182 33042 6210 33370
rect 6318 33260 6614 33280
rect 6374 33258 6398 33260
rect 6454 33258 6478 33260
rect 6534 33258 6558 33260
rect 6396 33206 6398 33258
rect 6460 33206 6472 33258
rect 6534 33206 6536 33258
rect 6374 33204 6398 33206
rect 6454 33204 6478 33206
rect 6534 33204 6558 33206
rect 6318 33184 6614 33204
rect 7102 33162 7130 33438
rect 7090 33156 7142 33162
rect 7090 33098 7142 33104
rect 6182 33014 6302 33042
rect 6274 32822 6302 33014
rect 6262 32816 6314 32822
rect 6262 32758 6314 32764
rect 6274 32618 6302 32758
rect 6262 32612 6314 32618
rect 6262 32554 6314 32560
rect 7918 32544 7970 32550
rect 7918 32486 7970 32492
rect 6630 32408 6682 32414
rect 6630 32350 6682 32356
rect 6998 32408 7050 32414
rect 6998 32350 7050 32356
rect 6318 32172 6614 32192
rect 6374 32170 6398 32172
rect 6454 32170 6478 32172
rect 6534 32170 6558 32172
rect 6396 32118 6398 32170
rect 6460 32118 6472 32170
rect 6534 32118 6536 32170
rect 6374 32116 6398 32118
rect 6454 32116 6478 32118
rect 6534 32116 6558 32118
rect 6318 32096 6614 32116
rect 5342 32068 5394 32074
rect 5342 32010 5394 32016
rect 6078 32068 6130 32074
rect 6078 32010 6130 32016
rect 6090 31802 6118 32010
rect 6170 32000 6222 32006
rect 6170 31942 6222 31948
rect 6078 31796 6130 31802
rect 6078 31738 6130 31744
rect 6182 31734 6210 31942
rect 6642 31802 6670 32350
rect 7010 31870 7038 32350
rect 6998 31864 7050 31870
rect 6998 31806 7050 31812
rect 6630 31796 6682 31802
rect 6630 31738 6682 31744
rect 6170 31728 6222 31734
rect 6170 31670 6222 31676
rect 5078 31530 5198 31546
rect 5078 31524 5210 31530
rect 5078 31518 5158 31524
rect 5078 30986 5106 31518
rect 5158 31466 5210 31472
rect 6182 31462 6210 31670
rect 6446 31524 6498 31530
rect 6446 31466 6498 31472
rect 6170 31456 6222 31462
rect 6170 31398 6222 31404
rect 6458 31326 6486 31466
rect 6446 31320 6498 31326
rect 6446 31262 6498 31268
rect 6642 31274 6670 31738
rect 7010 31394 7038 31806
rect 6998 31388 7050 31394
rect 6998 31330 7050 31336
rect 6722 31320 6774 31326
rect 6642 31268 6722 31274
rect 6642 31262 6774 31268
rect 6642 31246 6762 31262
rect 6814 31252 6866 31258
rect 6318 31084 6614 31104
rect 6374 31082 6398 31084
rect 6454 31082 6478 31084
rect 6534 31082 6558 31084
rect 6396 31030 6398 31082
rect 6460 31030 6472 31082
rect 6534 31030 6536 31082
rect 6374 31028 6398 31030
rect 6454 31028 6478 31030
rect 6534 31028 6558 31030
rect 6318 31008 6614 31028
rect 4974 30980 5026 30986
rect 4974 30922 5026 30928
rect 5066 30980 5118 30986
rect 5066 30922 5118 30928
rect 6642 30850 6670 31246
rect 6814 31194 6866 31200
rect 6630 30844 6682 30850
rect 6630 30786 6682 30792
rect 6262 30776 6314 30782
rect 6262 30718 6314 30724
rect 5066 30708 5118 30714
rect 5066 30650 5118 30656
rect 5078 30238 5106 30650
rect 5710 30436 5762 30442
rect 5710 30378 5762 30384
rect 5066 30232 5118 30238
rect 5066 30174 5118 30180
rect 5722 29830 5750 30378
rect 6274 30238 6302 30718
rect 6826 30238 6854 31194
rect 6906 30844 6958 30850
rect 6906 30786 6958 30792
rect 6918 30646 6946 30786
rect 6906 30640 6958 30646
rect 6906 30582 6958 30588
rect 7090 30640 7142 30646
rect 7090 30582 7142 30588
rect 6918 30306 6946 30582
rect 7102 30306 7130 30582
rect 6906 30300 6958 30306
rect 6906 30242 6958 30248
rect 7090 30300 7142 30306
rect 7090 30242 7142 30248
rect 6262 30232 6314 30238
rect 6182 30192 6262 30220
rect 5710 29824 5762 29830
rect 5710 29766 5762 29772
rect 6182 29762 6210 30192
rect 6262 30174 6314 30180
rect 6814 30232 6866 30238
rect 6814 30174 6866 30180
rect 6722 30096 6774 30102
rect 6722 30038 6774 30044
rect 6318 29996 6614 30016
rect 6374 29994 6398 29996
rect 6454 29994 6478 29996
rect 6534 29994 6558 29996
rect 6396 29942 6398 29994
rect 6460 29942 6472 29994
rect 6534 29942 6536 29994
rect 6374 29940 6398 29942
rect 6454 29940 6478 29942
rect 6534 29940 6558 29942
rect 6318 29920 6614 29940
rect 6734 29762 6762 30038
rect 6170 29756 6222 29762
rect 6170 29698 6222 29704
rect 6354 29756 6406 29762
rect 6354 29698 6406 29704
rect 6446 29756 6498 29762
rect 6446 29698 6498 29704
rect 6722 29756 6774 29762
rect 6722 29698 6774 29704
rect 6182 28674 6210 29698
rect 6366 29150 6394 29698
rect 6458 29218 6486 29698
rect 6446 29212 6498 29218
rect 6446 29154 6498 29160
rect 6918 29150 6946 30242
rect 7930 30238 7958 32486
rect 8194 31728 8246 31734
rect 8194 31670 8246 31676
rect 8102 31184 8154 31190
rect 8102 31126 8154 31132
rect 8114 30374 8142 31126
rect 8206 30714 8234 31670
rect 8194 30708 8246 30714
rect 8194 30650 8246 30656
rect 8102 30368 8154 30374
rect 8102 30310 8154 30316
rect 7734 30232 7786 30238
rect 7734 30174 7786 30180
rect 7918 30232 7970 30238
rect 7918 30174 7970 30180
rect 7746 29218 7774 30174
rect 8114 29830 8142 30310
rect 8206 30238 8234 30650
rect 8286 30368 8338 30374
rect 8286 30310 8338 30316
rect 8194 30232 8246 30238
rect 8194 30174 8246 30180
rect 8102 29824 8154 29830
rect 8102 29766 8154 29772
rect 8010 29756 8062 29762
rect 8010 29698 8062 29704
rect 8022 29354 8050 29698
rect 8010 29348 8062 29354
rect 8010 29290 8062 29296
rect 7734 29212 7786 29218
rect 7734 29154 7786 29160
rect 8114 29150 8142 29766
rect 8194 29756 8246 29762
rect 8194 29698 8246 29704
rect 8206 29218 8234 29698
rect 8298 29354 8326 30310
rect 8286 29348 8338 29354
rect 8286 29290 8338 29296
rect 8194 29212 8246 29218
rect 8194 29154 8246 29160
rect 6354 29144 6406 29150
rect 6354 29086 6406 29092
rect 6906 29144 6958 29150
rect 6906 29086 6958 29092
rect 8102 29144 8154 29150
rect 8102 29086 8154 29092
rect 6722 29008 6774 29014
rect 6722 28950 6774 28956
rect 6318 28908 6614 28928
rect 6374 28906 6398 28908
rect 6454 28906 6478 28908
rect 6534 28906 6558 28908
rect 6396 28854 6398 28906
rect 6460 28854 6472 28906
rect 6534 28854 6536 28906
rect 6374 28852 6398 28854
rect 6454 28852 6478 28854
rect 6534 28852 6558 28854
rect 6318 28832 6614 28852
rect 6734 28810 6762 28950
rect 6722 28804 6774 28810
rect 6722 28746 6774 28752
rect 8114 28674 8142 29086
rect 6170 28668 6222 28674
rect 6170 28610 6222 28616
rect 8102 28668 8154 28674
rect 8102 28610 8154 28616
rect 5986 28532 6038 28538
rect 5986 28474 6038 28480
rect 5526 26900 5578 26906
rect 5526 26842 5578 26848
rect 5538 26634 5566 26842
rect 5526 26628 5578 26634
rect 5526 26570 5578 26576
rect 5802 26424 5854 26430
rect 5802 26366 5854 26372
rect 5814 25478 5842 26366
rect 5802 25472 5854 25478
rect 5802 25414 5854 25420
rect 5066 24860 5118 24866
rect 5066 24802 5118 24808
rect 5078 24390 5106 24802
rect 5066 24384 5118 24390
rect 5066 24326 5118 24332
rect 4974 21936 5026 21942
rect 4974 21878 5026 21884
rect 4986 20990 5014 21878
rect 5066 21460 5118 21466
rect 5066 21402 5118 21408
rect 4974 20984 5026 20990
rect 4974 20926 5026 20932
rect 5078 19970 5106 21402
rect 5066 19964 5118 19970
rect 5066 19906 5118 19912
rect 5998 19018 6026 28474
rect 8102 28192 8154 28198
rect 8102 28134 8154 28140
rect 6170 28124 6222 28130
rect 6170 28066 6222 28072
rect 6182 26634 6210 28066
rect 7734 28056 7786 28062
rect 7734 27998 7786 28004
rect 6318 27820 6614 27840
rect 6374 27818 6398 27820
rect 6454 27818 6478 27820
rect 6534 27818 6558 27820
rect 6396 27766 6398 27818
rect 6460 27766 6472 27818
rect 6534 27766 6536 27818
rect 6374 27764 6398 27766
rect 6454 27764 6478 27766
rect 6534 27764 6558 27766
rect 6318 27744 6614 27764
rect 7746 27722 7774 27998
rect 8114 27722 8142 28134
rect 7734 27716 7786 27722
rect 7734 27658 7786 27664
rect 8102 27716 8154 27722
rect 8102 27658 8154 27664
rect 8114 27586 8142 27658
rect 8102 27580 8154 27586
rect 8102 27522 8154 27528
rect 7550 27376 7602 27382
rect 7550 27318 7602 27324
rect 6318 26732 6614 26752
rect 6374 26730 6398 26732
rect 6454 26730 6478 26732
rect 6534 26730 6558 26732
rect 6396 26678 6398 26730
rect 6460 26678 6472 26730
rect 6534 26678 6536 26730
rect 6374 26676 6398 26678
rect 6454 26676 6478 26678
rect 6534 26676 6558 26678
rect 6318 26656 6614 26676
rect 6170 26628 6222 26634
rect 6170 26570 6222 26576
rect 6630 26356 6682 26362
rect 6630 26298 6682 26304
rect 6642 26090 6670 26298
rect 6630 26084 6682 26090
rect 6630 26026 6682 26032
rect 6630 25812 6682 25818
rect 6630 25754 6682 25760
rect 6318 25644 6614 25664
rect 6374 25642 6398 25644
rect 6454 25642 6478 25644
rect 6534 25642 6558 25644
rect 6396 25590 6398 25642
rect 6460 25590 6472 25642
rect 6534 25590 6536 25642
rect 6374 25588 6398 25590
rect 6454 25588 6478 25590
rect 6534 25588 6558 25590
rect 6318 25568 6614 25588
rect 6642 25410 6670 25754
rect 6630 25404 6682 25410
rect 6630 25346 6682 25352
rect 7090 24996 7142 25002
rect 7090 24938 7142 24944
rect 7102 24798 7130 24938
rect 7090 24792 7142 24798
rect 7090 24734 7142 24740
rect 6722 24656 6774 24662
rect 6722 24598 6774 24604
rect 6318 24556 6614 24576
rect 6374 24554 6398 24556
rect 6454 24554 6478 24556
rect 6534 24554 6558 24556
rect 6396 24502 6398 24554
rect 6460 24502 6472 24554
rect 6534 24502 6536 24554
rect 6374 24500 6398 24502
rect 6454 24500 6478 24502
rect 6534 24500 6558 24502
rect 6318 24480 6614 24500
rect 6734 24254 6762 24598
rect 7562 24390 7590 27318
rect 7550 24384 7602 24390
rect 7550 24326 7602 24332
rect 7562 24254 7590 24326
rect 6722 24248 6774 24254
rect 6722 24190 6774 24196
rect 7550 24248 7602 24254
rect 7550 24190 7602 24196
rect 6630 23772 6682 23778
rect 6630 23714 6682 23720
rect 6318 23468 6614 23488
rect 6374 23466 6398 23468
rect 6454 23466 6478 23468
rect 6534 23466 6558 23468
rect 6396 23414 6398 23466
rect 6460 23414 6472 23466
rect 6534 23414 6536 23466
rect 6374 23412 6398 23414
rect 6454 23412 6478 23414
rect 6534 23412 6558 23414
rect 6318 23392 6614 23412
rect 6642 23302 6670 23714
rect 6734 23370 6762 24190
rect 7274 24112 7326 24118
rect 7274 24054 7326 24060
rect 7286 23914 7314 24054
rect 7274 23908 7326 23914
rect 7274 23850 7326 23856
rect 6906 23840 6958 23846
rect 6906 23782 6958 23788
rect 6722 23364 6774 23370
rect 6722 23306 6774 23312
rect 6630 23296 6682 23302
rect 6630 23238 6682 23244
rect 6642 22826 6670 23238
rect 6630 22820 6682 22826
rect 6630 22762 6682 22768
rect 6630 22548 6682 22554
rect 6630 22490 6682 22496
rect 6318 22380 6614 22400
rect 6374 22378 6398 22380
rect 6454 22378 6478 22380
rect 6534 22378 6558 22380
rect 6396 22326 6398 22378
rect 6460 22326 6472 22378
rect 6534 22326 6536 22378
rect 6374 22324 6398 22326
rect 6454 22324 6478 22326
rect 6534 22324 6558 22326
rect 6318 22304 6614 22324
rect 6642 22146 6670 22490
rect 6078 22140 6130 22146
rect 6078 22082 6130 22088
rect 6630 22140 6682 22146
rect 6630 22082 6682 22088
rect 6090 21194 6118 22082
rect 6170 21528 6222 21534
rect 6170 21470 6222 21476
rect 6078 21188 6130 21194
rect 6078 21130 6130 21136
rect 6182 20650 6210 21470
rect 6318 21292 6614 21312
rect 6374 21290 6398 21292
rect 6454 21290 6478 21292
rect 6534 21290 6558 21292
rect 6396 21238 6398 21290
rect 6460 21238 6472 21290
rect 6534 21238 6536 21290
rect 6374 21236 6398 21238
rect 6454 21236 6478 21238
rect 6534 21236 6558 21238
rect 6318 21216 6614 21236
rect 6734 21058 6762 23306
rect 6918 21126 6946 23782
rect 7286 23710 7314 23850
rect 7274 23704 7326 23710
rect 7274 23646 7326 23652
rect 7182 23160 7234 23166
rect 7182 23102 7234 23108
rect 7194 22282 7222 23102
rect 7182 22276 7234 22282
rect 7182 22218 7234 22224
rect 8390 22010 8418 34934
rect 8982 34892 9278 34912
rect 9038 34890 9062 34892
rect 9118 34890 9142 34892
rect 9198 34890 9222 34892
rect 9060 34838 9062 34890
rect 9124 34838 9136 34890
rect 9198 34838 9200 34890
rect 9038 34836 9062 34838
rect 9118 34836 9142 34838
rect 9198 34836 9222 34838
rect 8982 34816 9278 34836
rect 9494 34590 9522 36566
rect 9770 36426 9798 37994
rect 10322 37514 10350 38334
rect 10770 38256 10822 38262
rect 10770 38198 10822 38204
rect 10402 38052 10454 38058
rect 10402 37994 10454 38000
rect 10414 37530 10442 37994
rect 10414 37514 10534 37530
rect 10310 37508 10362 37514
rect 10414 37508 10546 37514
rect 10414 37502 10494 37508
rect 10310 37450 10362 37456
rect 10494 37450 10546 37456
rect 10782 37378 10810 38198
rect 11518 37378 11546 39422
rect 11646 38700 11942 38720
rect 11702 38698 11726 38700
rect 11782 38698 11806 38700
rect 11862 38698 11886 38700
rect 11724 38646 11726 38698
rect 11788 38646 11800 38698
rect 11862 38646 11864 38698
rect 11702 38644 11726 38646
rect 11782 38644 11806 38646
rect 11862 38644 11886 38646
rect 11646 38624 11942 38644
rect 11978 38482 12006 40170
rect 13082 40166 13110 40374
rect 13542 40166 13570 41038
rect 14646 40642 14674 43312
rect 14910 40976 14962 40982
rect 14910 40918 14962 40924
rect 14922 40778 14950 40918
rect 14910 40772 14962 40778
rect 14910 40714 14962 40720
rect 14634 40636 14686 40642
rect 14634 40578 14686 40584
rect 14922 40574 14950 40714
rect 14174 40568 14226 40574
rect 14174 40510 14226 40516
rect 14910 40568 14962 40574
rect 14910 40510 14962 40516
rect 14186 40234 14214 40510
rect 14310 40332 14606 40352
rect 14366 40330 14390 40332
rect 14446 40330 14470 40332
rect 14526 40330 14550 40332
rect 14388 40278 14390 40330
rect 14452 40278 14464 40330
rect 14526 40278 14528 40330
rect 14366 40276 14390 40278
rect 14446 40276 14470 40278
rect 14526 40276 14550 40278
rect 14310 40256 14606 40276
rect 14174 40228 14226 40234
rect 14174 40170 14226 40176
rect 13070 40160 13122 40166
rect 13070 40102 13122 40108
rect 13530 40160 13582 40166
rect 13530 40102 13582 40108
rect 12242 39956 12294 39962
rect 12242 39898 12294 39904
rect 12978 39956 13030 39962
rect 12978 39898 13030 39904
rect 12254 39554 12282 39898
rect 12242 39548 12294 39554
rect 12242 39490 12294 39496
rect 12334 39480 12386 39486
rect 11886 38454 12006 38482
rect 12070 39428 12334 39434
rect 12070 39422 12386 39428
rect 12070 39406 12374 39422
rect 11886 37700 11914 38454
rect 11966 38256 12018 38262
rect 11966 38198 12018 38204
rect 11978 37922 12006 38198
rect 11966 37916 12018 37922
rect 11966 37858 12018 37864
rect 11886 37672 12006 37700
rect 11646 37612 11942 37632
rect 11702 37610 11726 37612
rect 11782 37610 11806 37612
rect 11862 37610 11886 37612
rect 11724 37558 11726 37610
rect 11788 37558 11800 37610
rect 11862 37558 11864 37610
rect 11702 37556 11726 37558
rect 11782 37556 11806 37558
rect 11862 37556 11886 37558
rect 11646 37536 11942 37556
rect 10770 37372 10822 37378
rect 10770 37314 10822 37320
rect 11506 37372 11558 37378
rect 11506 37314 11558 37320
rect 10494 36624 10546 36630
rect 10494 36566 10546 36572
rect 9758 36420 9810 36426
rect 9758 36362 9810 36368
rect 10506 36290 10534 36566
rect 11518 36290 11546 37314
rect 11646 36524 11942 36544
rect 11702 36522 11726 36524
rect 11782 36522 11806 36524
rect 11862 36522 11886 36524
rect 11724 36470 11726 36522
rect 11788 36470 11800 36522
rect 11862 36470 11864 36522
rect 11702 36468 11726 36470
rect 11782 36468 11806 36470
rect 11862 36468 11886 36470
rect 11646 36448 11942 36468
rect 10218 36284 10270 36290
rect 10218 36226 10270 36232
rect 10494 36284 10546 36290
rect 10494 36226 10546 36232
rect 11506 36284 11558 36290
rect 11506 36226 11558 36232
rect 10230 35814 10258 36226
rect 10218 35808 10270 35814
rect 10218 35750 10270 35756
rect 10126 35536 10178 35542
rect 10126 35478 10178 35484
rect 10138 35202 10166 35478
rect 10126 35196 10178 35202
rect 10126 35138 10178 35144
rect 9114 34584 9166 34590
rect 9114 34526 9166 34532
rect 9482 34584 9534 34590
rect 9482 34526 9534 34532
rect 9126 34114 9154 34526
rect 10230 34250 10258 35750
rect 10506 35746 10534 36226
rect 10494 35740 10546 35746
rect 10494 35682 10546 35688
rect 10586 35672 10638 35678
rect 10586 35614 10638 35620
rect 11322 35672 11374 35678
rect 11322 35614 11374 35620
rect 10598 35338 10626 35614
rect 10586 35332 10638 35338
rect 10586 35274 10638 35280
rect 11334 35134 11362 35614
rect 11414 35604 11466 35610
rect 11414 35546 11466 35552
rect 11426 35202 11454 35546
rect 11646 35436 11942 35456
rect 11702 35434 11726 35436
rect 11782 35434 11806 35436
rect 11862 35434 11886 35436
rect 11724 35382 11726 35434
rect 11788 35382 11800 35434
rect 11862 35382 11864 35434
rect 11702 35380 11726 35382
rect 11782 35380 11806 35382
rect 11862 35380 11886 35382
rect 11646 35360 11942 35380
rect 11978 35338 12006 37672
rect 12070 37446 12098 39406
rect 12242 39344 12294 39350
rect 12242 39286 12294 39292
rect 12254 39010 12282 39286
rect 12242 39004 12294 39010
rect 12242 38946 12294 38952
rect 12794 37848 12846 37854
rect 12794 37790 12846 37796
rect 12806 37514 12834 37790
rect 12794 37508 12846 37514
rect 12794 37450 12846 37456
rect 12058 37440 12110 37446
rect 12058 37382 12110 37388
rect 12070 36222 12098 37382
rect 12058 36216 12110 36222
rect 12058 36158 12110 36164
rect 12610 36148 12662 36154
rect 12610 36090 12662 36096
rect 12150 36080 12202 36086
rect 12150 36022 12202 36028
rect 12162 35746 12190 36022
rect 12150 35740 12202 35746
rect 12150 35682 12202 35688
rect 12622 35542 12650 36090
rect 12610 35536 12662 35542
rect 12610 35478 12662 35484
rect 11966 35332 12018 35338
rect 11966 35274 12018 35280
rect 11414 35196 11466 35202
rect 11414 35138 11466 35144
rect 11322 35128 11374 35134
rect 11322 35070 11374 35076
rect 11334 34998 11362 35070
rect 11322 34992 11374 34998
rect 11322 34934 11374 34940
rect 10218 34244 10270 34250
rect 10218 34186 10270 34192
rect 9114 34108 9166 34114
rect 9114 34050 9166 34056
rect 10402 33972 10454 33978
rect 10402 33914 10454 33920
rect 9390 33904 9442 33910
rect 9390 33846 9442 33852
rect 8982 33804 9278 33824
rect 9038 33802 9062 33804
rect 9118 33802 9142 33804
rect 9198 33802 9222 33804
rect 9060 33750 9062 33802
rect 9124 33750 9136 33802
rect 9198 33750 9200 33802
rect 9038 33748 9062 33750
rect 9118 33748 9142 33750
rect 9198 33748 9222 33750
rect 8982 33728 9278 33748
rect 9402 33570 9430 33846
rect 9390 33564 9442 33570
rect 9390 33506 9442 33512
rect 10034 33496 10086 33502
rect 10034 33438 10086 33444
rect 10046 33026 10074 33438
rect 10414 33434 10442 33914
rect 10402 33428 10454 33434
rect 10402 33370 10454 33376
rect 10034 33020 10086 33026
rect 10034 32962 10086 32968
rect 10414 32822 10442 33370
rect 11334 33026 11362 34934
rect 11322 33020 11374 33026
rect 11322 32962 11374 32968
rect 10402 32816 10454 32822
rect 10402 32758 10454 32764
rect 11230 32816 11282 32822
rect 11230 32758 11282 32764
rect 8982 32716 9278 32736
rect 9038 32714 9062 32716
rect 9118 32714 9142 32716
rect 9198 32714 9222 32716
rect 9060 32662 9062 32714
rect 9124 32662 9136 32714
rect 9198 32662 9200 32714
rect 9038 32660 9062 32662
rect 9118 32660 9142 32662
rect 9198 32660 9222 32662
rect 8982 32640 9278 32660
rect 11242 31938 11270 32758
rect 8470 31932 8522 31938
rect 8470 31874 8522 31880
rect 11046 31932 11098 31938
rect 11046 31874 11098 31880
rect 11230 31932 11282 31938
rect 11230 31874 11282 31880
rect 8482 29558 8510 31874
rect 8982 31628 9278 31648
rect 9038 31626 9062 31628
rect 9118 31626 9142 31628
rect 9198 31626 9222 31628
rect 9060 31574 9062 31626
rect 9124 31574 9136 31626
rect 9198 31574 9200 31626
rect 9038 31572 9062 31574
rect 9118 31572 9142 31574
rect 9198 31572 9222 31574
rect 8982 31552 9278 31572
rect 11058 31530 11086 31874
rect 11046 31524 11098 31530
rect 11046 31466 11098 31472
rect 9298 31320 9350 31326
rect 9298 31262 9350 31268
rect 8982 30540 9278 30560
rect 9038 30538 9062 30540
rect 9118 30538 9142 30540
rect 9198 30538 9222 30540
rect 9060 30486 9062 30538
rect 9124 30486 9136 30538
rect 9198 30486 9200 30538
rect 9038 30484 9062 30486
rect 9118 30484 9142 30486
rect 9198 30484 9222 30486
rect 8982 30464 9278 30484
rect 9310 30306 9338 31262
rect 10310 30844 10362 30850
rect 10310 30786 10362 30792
rect 10402 30844 10454 30850
rect 10402 30786 10454 30792
rect 9482 30776 9534 30782
rect 9482 30718 9534 30724
rect 10126 30776 10178 30782
rect 10126 30718 10178 30724
rect 9298 30300 9350 30306
rect 9298 30242 9350 30248
rect 9494 30238 9522 30718
rect 9482 30232 9534 30238
rect 9482 30174 9534 30180
rect 9482 29824 9534 29830
rect 9482 29766 9534 29772
rect 9390 29756 9442 29762
rect 9390 29698 9442 29704
rect 9298 29620 9350 29626
rect 9298 29562 9350 29568
rect 8470 29552 8522 29558
rect 8470 29494 8522 29500
rect 8982 29452 9278 29472
rect 9038 29450 9062 29452
rect 9118 29450 9142 29452
rect 9198 29450 9222 29452
rect 9060 29398 9062 29450
rect 9124 29398 9136 29450
rect 9198 29398 9200 29450
rect 9038 29396 9062 29398
rect 9118 29396 9142 29398
rect 9198 29396 9222 29398
rect 8982 29376 9278 29396
rect 9310 28810 9338 29562
rect 9402 29354 9430 29698
rect 9494 29558 9522 29766
rect 9850 29688 9902 29694
rect 9850 29630 9902 29636
rect 9482 29552 9534 29558
rect 9482 29494 9534 29500
rect 9390 29348 9442 29354
rect 9390 29290 9442 29296
rect 9298 28804 9350 28810
rect 9298 28746 9350 28752
rect 9402 28674 9430 29290
rect 9494 29082 9522 29494
rect 9482 29076 9534 29082
rect 9482 29018 9534 29024
rect 9482 28736 9534 28742
rect 9482 28678 9534 28684
rect 9390 28668 9442 28674
rect 9390 28610 9442 28616
rect 8982 28364 9278 28384
rect 9038 28362 9062 28364
rect 9118 28362 9142 28364
rect 9198 28362 9222 28364
rect 9060 28310 9062 28362
rect 9124 28310 9136 28362
rect 9198 28310 9200 28362
rect 9038 28308 9062 28310
rect 9118 28308 9142 28310
rect 9198 28308 9222 28310
rect 8982 28288 9278 28308
rect 8562 28124 8614 28130
rect 8562 28066 8614 28072
rect 8574 27926 8602 28066
rect 9494 28062 9522 28678
rect 9482 28056 9534 28062
rect 9482 27998 9534 28004
rect 8562 27920 8614 27926
rect 8562 27862 8614 27868
rect 9298 27920 9350 27926
rect 9298 27862 9350 27868
rect 8574 27654 8602 27862
rect 8562 27648 8614 27654
rect 8562 27590 8614 27596
rect 9310 27450 9338 27862
rect 9298 27444 9350 27450
rect 9298 27386 9350 27392
rect 8982 27276 9278 27296
rect 9038 27274 9062 27276
rect 9118 27274 9142 27276
rect 9198 27274 9222 27276
rect 9060 27222 9062 27274
rect 9124 27222 9136 27274
rect 9198 27222 9200 27274
rect 9038 27220 9062 27222
rect 9118 27220 9142 27222
rect 9198 27220 9222 27222
rect 8982 27200 9278 27220
rect 9310 27178 9338 27386
rect 9298 27172 9350 27178
rect 9298 27114 9350 27120
rect 9310 26974 9338 27114
rect 9298 26968 9350 26974
rect 9298 26910 9350 26916
rect 9022 26900 9074 26906
rect 9022 26842 9074 26848
rect 9034 23574 9062 26842
rect 9862 24662 9890 29630
rect 10138 29626 10166 30718
rect 10322 29830 10350 30786
rect 10310 29824 10362 29830
rect 10310 29766 10362 29772
rect 10126 29620 10178 29626
rect 10126 29562 10178 29568
rect 10138 29218 10166 29562
rect 10414 29354 10442 30786
rect 10402 29348 10454 29354
rect 10402 29290 10454 29296
rect 10126 29212 10178 29218
rect 10126 29154 10178 29160
rect 10954 29076 11006 29082
rect 10954 29018 11006 29024
rect 10966 28742 10994 29018
rect 10954 28736 11006 28742
rect 10954 28678 11006 28684
rect 10954 28600 11006 28606
rect 10954 28542 11006 28548
rect 10966 28062 10994 28542
rect 10954 28056 11006 28062
rect 10954 27998 11006 28004
rect 10310 27512 10362 27518
rect 10124 27480 10180 27489
rect 10310 27454 10362 27460
rect 10124 27415 10180 27424
rect 10138 26974 10166 27415
rect 10322 26974 10350 27454
rect 10586 27376 10638 27382
rect 10586 27318 10638 27324
rect 10598 27110 10626 27318
rect 10586 27104 10638 27110
rect 10586 27046 10638 27052
rect 10126 26968 10178 26974
rect 10126 26910 10178 26916
rect 10310 26968 10362 26974
rect 10310 26910 10362 26916
rect 10678 26900 10730 26906
rect 10678 26842 10730 26848
rect 9850 24656 9902 24662
rect 9850 24598 9902 24604
rect 10690 24322 10718 26842
rect 10678 24316 10730 24322
rect 10678 24258 10730 24264
rect 9022 23568 9074 23574
rect 9022 23510 9074 23516
rect 8378 22004 8430 22010
rect 8378 21946 8430 21952
rect 6906 21120 6958 21126
rect 6906 21062 6958 21068
rect 6722 21052 6774 21058
rect 6722 20994 6774 21000
rect 6170 20644 6222 20650
rect 6170 20586 6222 20592
rect 6318 20204 6614 20224
rect 6374 20202 6398 20204
rect 6454 20202 6478 20204
rect 6534 20202 6558 20204
rect 6396 20150 6398 20202
rect 6460 20150 6472 20202
rect 6534 20150 6536 20202
rect 6374 20148 6398 20150
rect 6454 20148 6478 20150
rect 6534 20148 6558 20150
rect 6318 20128 6614 20148
rect 6734 19902 6762 20994
rect 6814 20304 6866 20310
rect 6814 20246 6866 20252
rect 6826 20038 6854 20246
rect 6814 20032 6866 20038
rect 6812 20000 6814 20009
rect 6866 20000 6868 20009
rect 6812 19935 6868 19944
rect 6722 19896 6774 19902
rect 6722 19838 6774 19844
rect 6734 19766 6762 19838
rect 6722 19760 6774 19766
rect 6722 19702 6774 19708
rect 6998 19760 7050 19766
rect 6998 19702 7050 19708
rect 6318 19116 6614 19136
rect 6374 19114 6398 19116
rect 6454 19114 6478 19116
rect 6534 19114 6558 19116
rect 6396 19062 6398 19114
rect 6460 19062 6472 19114
rect 6534 19062 6536 19114
rect 6374 19060 6398 19062
rect 6454 19060 6478 19062
rect 6534 19060 6558 19062
rect 6318 19040 6614 19060
rect 5986 19012 6038 19018
rect 5986 18954 6038 18960
rect 6906 18876 6958 18882
rect 6906 18818 6958 18824
rect 6918 18474 6946 18818
rect 6906 18468 6958 18474
rect 6906 18410 6958 18416
rect 5066 18128 5118 18134
rect 5066 18070 5118 18076
rect 5526 18128 5578 18134
rect 5526 18070 5578 18076
rect 5078 17794 5106 18070
rect 5066 17788 5118 17794
rect 5066 17730 5118 17736
rect 5078 17590 5106 17730
rect 5538 17726 5566 18070
rect 6318 18028 6614 18048
rect 6374 18026 6398 18028
rect 6454 18026 6478 18028
rect 6534 18026 6558 18028
rect 6396 17974 6398 18026
rect 6460 17974 6472 18026
rect 6534 17974 6536 18026
rect 6374 17972 6398 17974
rect 6454 17972 6478 17974
rect 6534 17972 6558 17974
rect 6318 17952 6614 17972
rect 7010 17726 7038 19702
rect 7090 18740 7142 18746
rect 7090 18682 7142 18688
rect 7102 17794 7130 18682
rect 7274 18128 7326 18134
rect 7274 18070 7326 18076
rect 7090 17788 7142 17794
rect 7090 17730 7142 17736
rect 5526 17720 5578 17726
rect 5526 17662 5578 17668
rect 6078 17720 6130 17726
rect 6078 17662 6130 17668
rect 6998 17720 7050 17726
rect 6998 17662 7050 17668
rect 5066 17584 5118 17590
rect 5066 17526 5118 17532
rect 5078 17289 5106 17526
rect 5064 17280 5120 17289
rect 5064 17215 5120 17224
rect 5710 16632 5762 16638
rect 5708 16600 5710 16609
rect 5762 16600 5764 16609
rect 5708 16535 5764 16544
rect 4882 16224 4934 16230
rect 4882 16166 4934 16172
rect 4698 16088 4750 16094
rect 4698 16030 4750 16036
rect 5250 16020 5302 16026
rect 5250 15962 5302 15968
rect 5262 15618 5290 15962
rect 5250 15612 5302 15618
rect 5250 15554 5302 15560
rect 6090 15550 6118 17662
rect 7286 17590 7314 18070
rect 7274 17584 7326 17590
rect 7272 17552 7274 17561
rect 7326 17552 7328 17561
rect 7272 17487 7328 17496
rect 6318 16940 6614 16960
rect 6374 16938 6398 16940
rect 6454 16938 6478 16940
rect 6534 16938 6558 16940
rect 6396 16886 6398 16938
rect 6460 16886 6472 16938
rect 6534 16886 6536 16938
rect 6374 16884 6398 16886
rect 6454 16884 6478 16886
rect 6534 16884 6558 16886
rect 6318 16864 6614 16884
rect 7182 16700 7234 16706
rect 7182 16642 7234 16648
rect 6722 16564 6774 16570
rect 6722 16506 6774 16512
rect 6318 15852 6614 15872
rect 6374 15850 6398 15852
rect 6454 15850 6478 15852
rect 6534 15850 6558 15852
rect 6396 15798 6398 15850
rect 6460 15798 6472 15850
rect 6534 15798 6536 15850
rect 6374 15796 6398 15798
rect 6454 15796 6478 15798
rect 6534 15796 6558 15798
rect 6318 15776 6614 15796
rect 6078 15544 6130 15550
rect 6078 15486 6130 15492
rect 3654 15308 3950 15328
rect 3710 15306 3734 15308
rect 3790 15306 3814 15308
rect 3870 15306 3894 15308
rect 3732 15254 3734 15306
rect 3796 15254 3808 15306
rect 3870 15254 3872 15306
rect 3710 15252 3734 15254
rect 3790 15252 3814 15254
rect 3870 15252 3894 15254
rect 3654 15232 3950 15252
rect 6090 14666 6118 15486
rect 6318 14764 6614 14784
rect 6374 14762 6398 14764
rect 6454 14762 6478 14764
rect 6534 14762 6558 14764
rect 6396 14710 6398 14762
rect 6460 14710 6472 14762
rect 6534 14710 6536 14762
rect 6374 14708 6398 14710
rect 6454 14708 6478 14710
rect 6534 14708 6558 14710
rect 6318 14688 6614 14708
rect 6078 14660 6130 14666
rect 6078 14602 6130 14608
rect 3654 14220 3950 14240
rect 3710 14218 3734 14220
rect 3790 14218 3814 14220
rect 3870 14218 3894 14220
rect 3732 14166 3734 14218
rect 3796 14166 3808 14218
rect 3870 14166 3872 14218
rect 3710 14164 3734 14166
rect 3790 14164 3814 14166
rect 3870 14164 3894 14166
rect 3654 14144 3950 14164
rect 3654 13132 3950 13152
rect 3710 13130 3734 13132
rect 3790 13130 3814 13132
rect 3870 13130 3894 13132
rect 3732 13078 3734 13130
rect 3796 13078 3808 13130
rect 3870 13078 3872 13130
rect 3710 13076 3734 13078
rect 3790 13076 3814 13078
rect 3870 13076 3894 13078
rect 3654 13056 3950 13076
rect 3654 12044 3950 12064
rect 3710 12042 3734 12044
rect 3790 12042 3814 12044
rect 3870 12042 3894 12044
rect 3732 11990 3734 12042
rect 3796 11990 3808 12042
rect 3870 11990 3872 12042
rect 3710 11988 3734 11990
rect 3790 11988 3814 11990
rect 3870 11988 3894 11990
rect 3654 11968 3950 11988
rect 3654 10956 3950 10976
rect 3710 10954 3734 10956
rect 3790 10954 3814 10956
rect 3870 10954 3894 10956
rect 3732 10902 3734 10954
rect 3796 10902 3808 10954
rect 3870 10902 3872 10954
rect 3710 10900 3734 10902
rect 3790 10900 3814 10902
rect 3870 10900 3894 10902
rect 3654 10880 3950 10900
rect 6090 10178 6118 14602
rect 6734 14530 6762 16506
rect 6998 15952 7050 15958
rect 6998 15894 7050 15900
rect 7010 15414 7038 15894
rect 6998 15408 7050 15414
rect 6998 15350 7050 15356
rect 7010 15249 7038 15350
rect 6996 15240 7052 15249
rect 7194 15210 7222 16642
rect 6996 15175 7052 15184
rect 7182 15204 7234 15210
rect 7182 15146 7234 15152
rect 7366 14864 7418 14870
rect 7366 14806 7418 14812
rect 7378 14569 7406 14806
rect 7364 14560 7420 14569
rect 6722 14524 6774 14530
rect 7364 14495 7366 14504
rect 6722 14466 6774 14472
rect 7418 14495 7420 14504
rect 7366 14466 7418 14472
rect 6318 13676 6614 13696
rect 6374 13674 6398 13676
rect 6454 13674 6478 13676
rect 6534 13674 6558 13676
rect 6396 13622 6398 13674
rect 6460 13622 6472 13674
rect 6534 13622 6536 13674
rect 6374 13620 6398 13622
rect 6454 13620 6478 13622
rect 6534 13620 6558 13622
rect 6318 13600 6614 13620
rect 6318 12588 6614 12608
rect 6374 12586 6398 12588
rect 6454 12586 6478 12588
rect 6534 12586 6558 12588
rect 6396 12534 6398 12586
rect 6460 12534 6472 12586
rect 6534 12534 6536 12586
rect 6374 12532 6398 12534
rect 6454 12532 6478 12534
rect 6534 12532 6558 12534
rect 6318 12512 6614 12532
rect 6318 11500 6614 11520
rect 6374 11498 6398 11500
rect 6454 11498 6478 11500
rect 6534 11498 6558 11500
rect 6396 11446 6398 11498
rect 6460 11446 6472 11498
rect 6534 11446 6536 11498
rect 6374 11444 6398 11446
rect 6454 11444 6478 11446
rect 6534 11444 6558 11446
rect 6318 11424 6614 11444
rect 6318 10412 6614 10432
rect 6374 10410 6398 10412
rect 6454 10410 6478 10412
rect 6534 10410 6558 10412
rect 6396 10358 6398 10410
rect 6460 10358 6472 10410
rect 6534 10358 6536 10410
rect 6374 10356 6398 10358
rect 6454 10356 6478 10358
rect 6534 10356 6558 10358
rect 6318 10336 6614 10356
rect 11138 10240 11190 10246
rect 11242 10194 11270 31874
rect 11426 30850 11454 35138
rect 11646 34348 11942 34368
rect 11702 34346 11726 34348
rect 11782 34346 11806 34348
rect 11862 34346 11886 34348
rect 11724 34294 11726 34346
rect 11788 34294 11800 34346
rect 11862 34294 11864 34346
rect 11702 34292 11726 34294
rect 11782 34292 11806 34294
rect 11862 34292 11886 34294
rect 11646 34272 11942 34292
rect 12518 33496 12570 33502
rect 12518 33438 12570 33444
rect 12426 33428 12478 33434
rect 12426 33370 12478 33376
rect 11506 33360 11558 33366
rect 11506 33302 11558 33308
rect 11518 31938 11546 33302
rect 11646 33260 11942 33280
rect 11702 33258 11726 33260
rect 11782 33258 11806 33260
rect 11862 33258 11886 33260
rect 11724 33206 11726 33258
rect 11788 33206 11800 33258
rect 11862 33206 11864 33258
rect 11702 33204 11726 33206
rect 11782 33204 11806 33206
rect 11862 33204 11886 33206
rect 11646 33184 11942 33204
rect 12438 33026 12466 33370
rect 12426 33020 12478 33026
rect 12426 32962 12478 32968
rect 11646 32172 11942 32192
rect 11702 32170 11726 32172
rect 11782 32170 11806 32172
rect 11862 32170 11886 32172
rect 11724 32118 11726 32170
rect 11788 32118 11800 32170
rect 11862 32118 11864 32170
rect 11702 32116 11726 32118
rect 11782 32116 11806 32118
rect 11862 32116 11886 32118
rect 11646 32096 11942 32116
rect 12530 32006 12558 33438
rect 12518 32000 12570 32006
rect 12518 31942 12570 31948
rect 11506 31932 11558 31938
rect 11506 31874 11558 31880
rect 11518 30918 11546 31874
rect 12622 31852 12650 35478
rect 12794 35332 12846 35338
rect 12794 35274 12846 35280
rect 12806 34794 12834 35274
rect 12794 34788 12846 34794
rect 12794 34730 12846 34736
rect 12806 34590 12834 34730
rect 12794 34584 12846 34590
rect 12794 34526 12846 34532
rect 12886 32408 12938 32414
rect 12886 32350 12938 32356
rect 12898 32074 12926 32350
rect 12886 32068 12938 32074
rect 12886 32010 12938 32016
rect 12530 31824 12650 31852
rect 12334 31388 12386 31394
rect 12334 31330 12386 31336
rect 12150 31184 12202 31190
rect 12150 31126 12202 31132
rect 11646 31084 11942 31104
rect 11702 31082 11726 31084
rect 11782 31082 11806 31084
rect 11862 31082 11886 31084
rect 11724 31030 11726 31082
rect 11788 31030 11800 31082
rect 11862 31030 11864 31082
rect 11702 31028 11726 31030
rect 11782 31028 11806 31030
rect 11862 31028 11886 31030
rect 11646 31008 11942 31028
rect 11506 30912 11558 30918
rect 11506 30854 11558 30860
rect 11414 30844 11466 30850
rect 11414 30786 11466 30792
rect 11506 30776 11558 30782
rect 11506 30718 11558 30724
rect 11414 30164 11466 30170
rect 11414 30106 11466 30112
rect 11426 29898 11454 30106
rect 11414 29892 11466 29898
rect 11414 29834 11466 29840
rect 11322 29008 11374 29014
rect 11322 28950 11374 28956
rect 11334 28538 11362 28950
rect 11518 28674 11546 30718
rect 11966 30164 12018 30170
rect 11966 30106 12018 30112
rect 11646 29996 11942 30016
rect 11702 29994 11726 29996
rect 11782 29994 11806 29996
rect 11862 29994 11886 29996
rect 11724 29942 11726 29994
rect 11788 29942 11800 29994
rect 11862 29942 11864 29994
rect 11702 29940 11726 29942
rect 11782 29940 11806 29942
rect 11862 29940 11886 29942
rect 11646 29920 11942 29940
rect 11646 28908 11942 28928
rect 11702 28906 11726 28908
rect 11782 28906 11806 28908
rect 11862 28906 11886 28908
rect 11724 28854 11726 28906
rect 11788 28854 11800 28906
rect 11862 28854 11864 28906
rect 11702 28852 11726 28854
rect 11782 28852 11806 28854
rect 11862 28852 11886 28854
rect 11646 28832 11942 28852
rect 11506 28668 11558 28674
rect 11506 28610 11558 28616
rect 11322 28532 11374 28538
rect 11322 28474 11374 28480
rect 11506 28532 11558 28538
rect 11506 28474 11558 28480
rect 11518 26362 11546 28474
rect 11978 28130 12006 30106
rect 12058 28668 12110 28674
rect 12058 28610 12110 28616
rect 11966 28124 12018 28130
rect 11966 28066 12018 28072
rect 11646 27820 11942 27840
rect 11702 27818 11726 27820
rect 11782 27818 11806 27820
rect 11862 27818 11886 27820
rect 11724 27766 11726 27818
rect 11788 27766 11800 27818
rect 11862 27766 11864 27818
rect 11702 27764 11726 27766
rect 11782 27764 11806 27766
rect 11862 27764 11886 27766
rect 11646 27744 11942 27764
rect 11874 27580 11926 27586
rect 11874 27522 11926 27528
rect 11886 27382 11914 27522
rect 11874 27376 11926 27382
rect 11874 27318 11926 27324
rect 12070 27042 12098 28610
rect 12162 27382 12190 31126
rect 12346 30850 12374 31330
rect 12426 31320 12478 31326
rect 12426 31262 12478 31268
rect 12438 30850 12466 31262
rect 12334 30844 12386 30850
rect 12334 30786 12386 30792
rect 12426 30844 12478 30850
rect 12426 30786 12478 30792
rect 12346 30306 12374 30786
rect 12334 30300 12386 30306
rect 12334 30242 12386 30248
rect 12530 30238 12558 31824
rect 12794 30844 12846 30850
rect 12794 30786 12846 30792
rect 12610 30368 12662 30374
rect 12610 30310 12662 30316
rect 12518 30232 12570 30238
rect 12518 30174 12570 30180
rect 12242 28056 12294 28062
rect 12242 27998 12294 28004
rect 12254 27586 12282 27998
rect 12622 27625 12650 30310
rect 12806 30238 12834 30786
rect 12794 30232 12846 30238
rect 12794 30174 12846 30180
rect 12806 29762 12834 30174
rect 12794 29756 12846 29762
rect 12794 29698 12846 29704
rect 12886 29552 12938 29558
rect 12886 29494 12938 29500
rect 12898 29354 12926 29494
rect 12886 29348 12938 29354
rect 12886 29290 12938 29296
rect 12990 28742 13018 39898
rect 13082 38602 13110 40102
rect 13254 40024 13306 40030
rect 13254 39966 13306 39972
rect 13898 40024 13950 40030
rect 13898 39966 13950 39972
rect 13070 38596 13122 38602
rect 13070 38538 13122 38544
rect 13070 34448 13122 34454
rect 13070 34390 13122 34396
rect 13082 33638 13110 34390
rect 13070 33632 13122 33638
rect 13070 33574 13122 33580
rect 13162 33020 13214 33026
rect 13162 32962 13214 32968
rect 13070 31932 13122 31938
rect 13070 31874 13122 31880
rect 13082 31258 13110 31874
rect 13070 31252 13122 31258
rect 13070 31194 13122 31200
rect 13174 30646 13202 32962
rect 13162 30640 13214 30646
rect 13162 30582 13214 30588
rect 13162 30096 13214 30102
rect 13162 30038 13214 30044
rect 13174 29762 13202 30038
rect 13162 29756 13214 29762
rect 13162 29698 13214 29704
rect 12978 28736 13030 28742
rect 12978 28678 13030 28684
rect 12886 28260 12938 28266
rect 12886 28202 12938 28208
rect 12700 28160 12756 28169
rect 12700 28095 12756 28104
rect 12714 28062 12742 28095
rect 12898 28062 12926 28202
rect 13266 28198 13294 39966
rect 13910 39622 13938 39966
rect 13622 39616 13674 39622
rect 13622 39558 13674 39564
rect 13898 39616 13950 39622
rect 13898 39558 13950 39564
rect 13634 38942 13662 39558
rect 14310 39244 14606 39264
rect 14366 39242 14390 39244
rect 14446 39242 14470 39244
rect 14526 39242 14550 39244
rect 14388 39190 14390 39242
rect 14452 39190 14464 39242
rect 14526 39190 14528 39242
rect 14366 39188 14390 39190
rect 14446 39188 14470 39190
rect 14526 39188 14550 39190
rect 14310 39168 14606 39188
rect 13622 38936 13674 38942
rect 13622 38878 13674 38884
rect 14082 38800 14134 38806
rect 14082 38742 14134 38748
rect 14094 37718 14122 38742
rect 14310 38156 14606 38176
rect 14366 38154 14390 38156
rect 14446 38154 14470 38156
rect 14526 38154 14550 38156
rect 14388 38102 14390 38154
rect 14452 38102 14464 38154
rect 14526 38102 14528 38154
rect 14366 38100 14390 38102
rect 14446 38100 14470 38102
rect 14526 38100 14550 38102
rect 14310 38080 14606 38100
rect 14174 37780 14226 37786
rect 14174 37722 14226 37728
rect 14082 37712 14134 37718
rect 14082 37654 14134 37660
rect 14094 35542 14122 37654
rect 14186 37446 14214 37722
rect 14174 37440 14226 37446
rect 14174 37382 14226 37388
rect 14310 37068 14606 37088
rect 14366 37066 14390 37068
rect 14446 37066 14470 37068
rect 14526 37066 14550 37068
rect 14388 37014 14390 37066
rect 14452 37014 14464 37066
rect 14526 37014 14528 37066
rect 14366 37012 14390 37014
rect 14446 37012 14470 37014
rect 14526 37012 14550 37014
rect 14310 36992 14606 37012
rect 14922 36426 14950 40510
rect 15738 38256 15790 38262
rect 15738 38198 15790 38204
rect 14910 36420 14962 36426
rect 14910 36362 14962 36368
rect 15554 36080 15606 36086
rect 15554 36022 15606 36028
rect 14310 35980 14606 36000
rect 14366 35978 14390 35980
rect 14446 35978 14470 35980
rect 14526 35978 14550 35980
rect 14388 35926 14390 35978
rect 14452 35926 14464 35978
rect 14526 35926 14528 35978
rect 14366 35924 14390 35926
rect 14446 35924 14470 35926
rect 14526 35924 14550 35926
rect 14310 35904 14606 35924
rect 15566 35542 15594 36022
rect 14082 35536 14134 35542
rect 14082 35478 14134 35484
rect 15554 35536 15606 35542
rect 15554 35478 15606 35484
rect 15566 35338 15594 35478
rect 15554 35332 15606 35338
rect 15554 35274 15606 35280
rect 15094 35264 15146 35270
rect 14724 35232 14780 35241
rect 14724 35167 14726 35176
rect 14778 35167 14780 35176
rect 15092 35232 15094 35241
rect 15146 35232 15148 35241
rect 15092 35167 15148 35176
rect 14726 35138 14778 35144
rect 13530 34992 13582 34998
rect 13530 34934 13582 34940
rect 13346 32408 13398 32414
rect 13346 32350 13398 32356
rect 13358 31394 13386 32350
rect 13542 31870 13570 34934
rect 14310 34892 14606 34912
rect 14366 34890 14390 34892
rect 14446 34890 14470 34892
rect 14526 34890 14550 34892
rect 14388 34838 14390 34890
rect 14452 34838 14464 34890
rect 14526 34838 14528 34890
rect 14366 34836 14390 34838
rect 14446 34836 14470 34838
rect 14526 34836 14550 34838
rect 14310 34816 14606 34836
rect 14310 33804 14606 33824
rect 14366 33802 14390 33804
rect 14446 33802 14470 33804
rect 14526 33802 14550 33804
rect 14388 33750 14390 33802
rect 14452 33750 14464 33802
rect 14526 33750 14528 33802
rect 14366 33748 14390 33750
rect 14446 33748 14470 33750
rect 14526 33748 14550 33750
rect 14310 33728 14606 33748
rect 13898 33496 13950 33502
rect 13896 33464 13898 33473
rect 13950 33464 13952 33473
rect 13896 33399 13952 33408
rect 14174 32884 14226 32890
rect 14174 32826 14226 32832
rect 13622 32816 13674 32822
rect 13622 32758 13674 32764
rect 13634 32346 13662 32758
rect 14186 32414 14214 32826
rect 14310 32716 14606 32736
rect 14366 32714 14390 32716
rect 14446 32714 14470 32716
rect 14526 32714 14550 32716
rect 14388 32662 14390 32714
rect 14452 32662 14464 32714
rect 14526 32662 14528 32714
rect 14366 32660 14390 32662
rect 14446 32660 14470 32662
rect 14526 32660 14550 32662
rect 14310 32640 14606 32660
rect 14174 32408 14226 32414
rect 14174 32350 14226 32356
rect 14266 32408 14318 32414
rect 14266 32350 14318 32356
rect 13622 32340 13674 32346
rect 13622 32282 13674 32288
rect 14278 31938 14306 32350
rect 14266 31932 14318 31938
rect 14266 31874 14318 31880
rect 13530 31864 13582 31870
rect 13530 31806 13582 31812
rect 13346 31388 13398 31394
rect 13346 31330 13398 31336
rect 13542 29354 13570 31806
rect 14310 31628 14606 31648
rect 14366 31626 14390 31628
rect 14446 31626 14470 31628
rect 14526 31626 14550 31628
rect 14388 31574 14390 31626
rect 14452 31574 14464 31626
rect 14526 31574 14528 31626
rect 14366 31572 14390 31574
rect 14446 31572 14470 31574
rect 14526 31572 14550 31574
rect 14310 31552 14606 31572
rect 14738 30986 14766 35138
rect 15566 35134 15594 35274
rect 15554 35128 15606 35134
rect 15554 35070 15606 35076
rect 15094 33156 15146 33162
rect 15094 33098 15146 33104
rect 14726 30980 14778 30986
rect 14726 30922 14778 30928
rect 14818 30844 14870 30850
rect 14818 30786 14870 30792
rect 14310 30540 14606 30560
rect 14366 30538 14390 30540
rect 14446 30538 14470 30540
rect 14526 30538 14550 30540
rect 14388 30486 14390 30538
rect 14452 30486 14464 30538
rect 14526 30486 14528 30538
rect 14366 30484 14390 30486
rect 14446 30484 14470 30486
rect 14526 30484 14550 30486
rect 14310 30464 14606 30484
rect 14726 30164 14778 30170
rect 14726 30106 14778 30112
rect 14310 29452 14606 29472
rect 14366 29450 14390 29452
rect 14446 29450 14470 29452
rect 14526 29450 14550 29452
rect 14388 29398 14390 29450
rect 14452 29398 14464 29450
rect 14526 29398 14528 29450
rect 14366 29396 14390 29398
rect 14446 29396 14470 29398
rect 14526 29396 14550 29398
rect 14310 29376 14606 29396
rect 13530 29348 13582 29354
rect 13530 29290 13582 29296
rect 13530 28804 13582 28810
rect 13530 28746 13582 28752
rect 13542 28266 13570 28746
rect 14738 28674 14766 30106
rect 14726 28668 14778 28674
rect 14726 28610 14778 28616
rect 14310 28364 14606 28384
rect 14366 28362 14390 28364
rect 14446 28362 14470 28364
rect 14526 28362 14550 28364
rect 14388 28310 14390 28362
rect 14452 28310 14464 28362
rect 14526 28310 14528 28362
rect 14366 28308 14390 28310
rect 14446 28308 14470 28310
rect 14526 28308 14550 28310
rect 14310 28288 14606 28308
rect 13530 28260 13582 28266
rect 13530 28202 13582 28208
rect 13254 28192 13306 28198
rect 13254 28134 13306 28140
rect 12702 28056 12754 28062
rect 12702 27998 12754 28004
rect 12886 28056 12938 28062
rect 12886 27998 12938 28004
rect 14830 27926 14858 30786
rect 15106 28470 15134 33098
rect 15566 32550 15594 35070
rect 15750 34250 15778 38198
rect 15842 37938 15870 43312
rect 17038 42154 17066 43312
rect 17038 42126 17342 42154
rect 16974 41964 17270 41984
rect 17030 41962 17054 41964
rect 17110 41962 17134 41964
rect 17190 41962 17214 41964
rect 17052 41910 17054 41962
rect 17116 41910 17128 41962
rect 17190 41910 17192 41962
rect 17030 41908 17054 41910
rect 17110 41908 17134 41910
rect 17190 41908 17214 41910
rect 16974 41888 17270 41908
rect 17314 41338 17342 42126
rect 18326 41338 18354 43312
rect 17314 41322 17434 41338
rect 17314 41316 17446 41322
rect 17314 41310 17394 41316
rect 17394 41258 17446 41264
rect 17590 41310 18354 41338
rect 17394 40976 17446 40982
rect 17394 40918 17446 40924
rect 16974 40876 17270 40896
rect 17030 40874 17054 40876
rect 17110 40874 17134 40876
rect 17190 40874 17214 40876
rect 17052 40822 17054 40874
rect 17116 40822 17128 40874
rect 17190 40822 17192 40874
rect 17030 40820 17054 40822
rect 17110 40820 17134 40822
rect 17190 40820 17214 40822
rect 16974 40800 17270 40820
rect 17406 40710 17434 40918
rect 17394 40704 17446 40710
rect 17394 40646 17446 40652
rect 17406 40574 17434 40646
rect 17394 40568 17446 40574
rect 17394 40510 17446 40516
rect 16658 40160 16710 40166
rect 16658 40102 16710 40108
rect 15922 39684 15974 39690
rect 15922 39626 15974 39632
rect 15934 38262 15962 39626
rect 16014 38868 16066 38874
rect 16014 38810 16066 38816
rect 16026 38466 16054 38810
rect 16014 38460 16066 38466
rect 16014 38402 16066 38408
rect 16382 38460 16434 38466
rect 16382 38402 16434 38408
rect 15922 38256 15974 38262
rect 15922 38198 15974 38204
rect 15842 37910 15962 37938
rect 15830 37780 15882 37786
rect 15830 37722 15882 37728
rect 15842 37378 15870 37722
rect 15830 37372 15882 37378
rect 15830 37314 15882 37320
rect 15830 36828 15882 36834
rect 15830 36770 15882 36776
rect 15738 34244 15790 34250
rect 15738 34186 15790 34192
rect 15842 33162 15870 36770
rect 15830 33156 15882 33162
rect 15830 33098 15882 33104
rect 15554 32544 15606 32550
rect 15554 32486 15606 32492
rect 15934 30986 15962 37910
rect 16026 37786 16054 38402
rect 16394 37961 16422 38402
rect 16380 37952 16436 37961
rect 16380 37887 16436 37896
rect 16014 37780 16066 37786
rect 16014 37722 16066 37728
rect 16026 37446 16054 37722
rect 16014 37440 16066 37446
rect 16014 37382 16066 37388
rect 16026 36970 16054 37382
rect 16474 37304 16526 37310
rect 16474 37246 16526 37252
rect 16014 36964 16066 36970
rect 16014 36906 16066 36912
rect 16198 36624 16250 36630
rect 16198 36566 16250 36572
rect 16106 36284 16158 36290
rect 16106 36226 16158 36232
rect 16118 35678 16146 36226
rect 16106 35672 16158 35678
rect 16106 35614 16158 35620
rect 16014 35128 16066 35134
rect 16014 35070 16066 35076
rect 16026 34250 16054 35070
rect 16118 34794 16146 35614
rect 16106 34788 16158 34794
rect 16106 34730 16158 34736
rect 16014 34244 16066 34250
rect 16014 34186 16066 34192
rect 16014 34108 16066 34114
rect 16014 34050 16066 34056
rect 16026 32006 16054 34050
rect 16106 32816 16158 32822
rect 16106 32758 16158 32764
rect 16118 32618 16146 32758
rect 16106 32612 16158 32618
rect 16106 32554 16158 32560
rect 16210 32498 16238 36566
rect 16486 32618 16514 37246
rect 16474 32612 16526 32618
rect 16474 32554 16526 32560
rect 16118 32470 16238 32498
rect 16014 32000 16066 32006
rect 16014 31942 16066 31948
rect 15922 30980 15974 30986
rect 15922 30922 15974 30928
rect 15934 30850 15962 30922
rect 15922 30844 15974 30850
rect 15922 30786 15974 30792
rect 15922 30096 15974 30102
rect 15922 30038 15974 30044
rect 15934 29762 15962 30038
rect 15922 29756 15974 29762
rect 15922 29698 15974 29704
rect 15830 29552 15882 29558
rect 15830 29494 15882 29500
rect 15094 28464 15146 28470
rect 15094 28406 15146 28412
rect 15106 28266 15134 28406
rect 15094 28260 15146 28266
rect 15094 28202 15146 28208
rect 15186 28192 15238 28198
rect 15186 28134 15238 28140
rect 14818 27920 14870 27926
rect 14818 27862 14870 27868
rect 12608 27616 12664 27625
rect 12242 27580 12294 27586
rect 12608 27551 12610 27560
rect 12242 27522 12294 27528
rect 12662 27551 12664 27560
rect 12610 27522 12662 27528
rect 12622 27491 12650 27522
rect 15198 27450 15226 28134
rect 15738 28056 15790 28062
rect 15738 27998 15790 28004
rect 15370 27920 15422 27926
rect 15370 27862 15422 27868
rect 15382 27722 15410 27862
rect 15370 27716 15422 27722
rect 15370 27658 15422 27664
rect 15750 27654 15778 27998
rect 15842 27722 15870 29494
rect 15922 28668 15974 28674
rect 15922 28610 15974 28616
rect 15934 28266 15962 28610
rect 15922 28260 15974 28266
rect 15922 28202 15974 28208
rect 15830 27716 15882 27722
rect 15830 27658 15882 27664
rect 15738 27648 15790 27654
rect 15738 27590 15790 27596
rect 15646 27580 15698 27586
rect 15646 27522 15698 27528
rect 16026 27568 16054 31942
rect 16118 31734 16146 32470
rect 16290 32408 16342 32414
rect 16290 32350 16342 32356
rect 16198 32340 16250 32346
rect 16198 32282 16250 32288
rect 16106 31728 16158 31734
rect 16106 31670 16158 31676
rect 16118 29218 16146 31670
rect 16106 29212 16158 29218
rect 16106 29154 16158 29160
rect 16106 28464 16158 28470
rect 16106 28406 16158 28412
rect 16118 28062 16146 28406
rect 16210 28130 16238 32282
rect 16302 28470 16330 32350
rect 16670 31394 16698 40102
rect 17406 40098 17434 40510
rect 17394 40092 17446 40098
rect 17394 40034 17446 40040
rect 16974 39788 17270 39808
rect 17030 39786 17054 39788
rect 17110 39786 17134 39788
rect 17190 39786 17214 39788
rect 17052 39734 17054 39786
rect 17116 39734 17128 39786
rect 17190 39734 17192 39786
rect 17030 39732 17054 39734
rect 17110 39732 17134 39734
rect 17190 39732 17214 39734
rect 16974 39712 17270 39732
rect 17486 39548 17538 39554
rect 17486 39490 17538 39496
rect 17394 39412 17446 39418
rect 17394 39354 17446 39360
rect 16750 38868 16802 38874
rect 16750 38810 16802 38816
rect 16762 38534 16790 38810
rect 16974 38700 17270 38720
rect 17030 38698 17054 38700
rect 17110 38698 17134 38700
rect 17190 38698 17214 38700
rect 17052 38646 17054 38698
rect 17116 38646 17128 38698
rect 17190 38646 17192 38698
rect 17030 38644 17054 38646
rect 17110 38644 17134 38646
rect 17190 38644 17214 38646
rect 16974 38624 17270 38644
rect 16750 38528 16802 38534
rect 16750 38470 16802 38476
rect 16974 37612 17270 37632
rect 17030 37610 17054 37612
rect 17110 37610 17134 37612
rect 17190 37610 17214 37612
rect 17052 37558 17054 37610
rect 17116 37558 17128 37610
rect 17190 37558 17192 37610
rect 17030 37556 17054 37558
rect 17110 37556 17134 37558
rect 17190 37556 17214 37558
rect 16974 37536 17270 37556
rect 17210 37372 17262 37378
rect 17210 37314 17262 37320
rect 17222 36970 17250 37314
rect 17406 37174 17434 39354
rect 17498 39010 17526 39490
rect 17486 39004 17538 39010
rect 17486 38946 17538 38952
rect 17590 38346 17618 41310
rect 17762 41112 17814 41118
rect 17762 41054 17814 41060
rect 17670 40568 17722 40574
rect 17670 40510 17722 40516
rect 17498 38318 17618 38346
rect 17394 37168 17446 37174
rect 17394 37110 17446 37116
rect 17210 36964 17262 36970
rect 17210 36906 17262 36912
rect 16974 36524 17270 36544
rect 17030 36522 17054 36524
rect 17110 36522 17134 36524
rect 17190 36522 17214 36524
rect 17052 36470 17054 36522
rect 17116 36470 17128 36522
rect 17190 36470 17192 36522
rect 17030 36468 17054 36470
rect 17110 36468 17134 36470
rect 17190 36468 17214 36470
rect 16974 36448 17270 36468
rect 16750 36216 16802 36222
rect 16750 36158 16802 36164
rect 16762 35882 16790 36158
rect 16750 35876 16802 35882
rect 16750 35818 16802 35824
rect 16842 35536 16894 35542
rect 16842 35478 16894 35484
rect 16854 34658 16882 35478
rect 16974 35436 17270 35456
rect 17030 35434 17054 35436
rect 17110 35434 17134 35436
rect 17190 35434 17214 35436
rect 17052 35382 17054 35434
rect 17116 35382 17128 35434
rect 17190 35382 17192 35434
rect 17030 35380 17054 35382
rect 17110 35380 17134 35382
rect 17190 35380 17214 35382
rect 16974 35360 17270 35380
rect 17498 35218 17526 38318
rect 17682 38262 17710 40510
rect 17774 39350 17802 41054
rect 17854 40432 17906 40438
rect 17854 40374 17906 40380
rect 17866 39978 17894 40374
rect 19522 40234 19550 43312
rect 20614 41520 20666 41526
rect 20614 41462 20666 41468
rect 19638 41420 19934 41440
rect 19694 41418 19718 41420
rect 19774 41418 19798 41420
rect 19854 41418 19878 41420
rect 19716 41366 19718 41418
rect 19780 41366 19792 41418
rect 19854 41366 19856 41418
rect 19694 41364 19718 41366
rect 19774 41364 19798 41366
rect 19854 41364 19878 41366
rect 19638 41344 19934 41364
rect 19638 40332 19934 40352
rect 19694 40330 19718 40332
rect 19774 40330 19798 40332
rect 19854 40330 19878 40332
rect 19716 40278 19718 40330
rect 19780 40278 19792 40330
rect 19854 40278 19856 40330
rect 19694 40276 19718 40278
rect 19774 40276 19798 40278
rect 19854 40276 19878 40278
rect 19638 40256 19934 40276
rect 19510 40228 19562 40234
rect 19510 40170 19562 40176
rect 19050 40024 19102 40030
rect 17866 39950 17986 39978
rect 19050 39966 19102 39972
rect 17762 39344 17814 39350
rect 17762 39286 17814 39292
rect 17762 38460 17814 38466
rect 17762 38402 17814 38408
rect 17578 38256 17630 38262
rect 17578 38198 17630 38204
rect 17670 38256 17722 38262
rect 17670 38198 17722 38204
rect 17590 38058 17618 38198
rect 17578 38052 17630 38058
rect 17578 37994 17630 38000
rect 17590 37242 17618 37994
rect 17774 37990 17802 38402
rect 17762 37984 17814 37990
rect 17762 37926 17814 37932
rect 17958 37922 17986 39950
rect 18774 39616 18826 39622
rect 18774 39558 18826 39564
rect 18314 39344 18366 39350
rect 18314 39286 18366 39292
rect 17946 37916 17998 37922
rect 17946 37858 17998 37864
rect 17670 37780 17722 37786
rect 17670 37722 17722 37728
rect 17946 37780 17998 37786
rect 17946 37722 17998 37728
rect 17682 37446 17710 37722
rect 17670 37440 17722 37446
rect 17670 37382 17722 37388
rect 17578 37236 17630 37242
rect 17578 37178 17630 37184
rect 17670 36760 17722 36766
rect 17670 36702 17722 36708
rect 17682 36426 17710 36702
rect 17670 36420 17722 36426
rect 17670 36362 17722 36368
rect 17578 35672 17630 35678
rect 17578 35614 17630 35620
rect 17590 35270 17618 35614
rect 17406 35190 17526 35218
rect 17578 35264 17630 35270
rect 17578 35206 17630 35212
rect 17302 34992 17354 34998
rect 17302 34934 17354 34940
rect 16842 34652 16894 34658
rect 16842 34594 16894 34600
rect 16854 34454 16882 34594
rect 16842 34448 16894 34454
rect 16842 34390 16894 34396
rect 16974 34348 17270 34368
rect 17030 34346 17054 34348
rect 17110 34346 17134 34348
rect 17190 34346 17214 34348
rect 17052 34294 17054 34346
rect 17116 34294 17128 34346
rect 17190 34294 17192 34346
rect 17030 34292 17054 34294
rect 17110 34292 17134 34294
rect 17190 34292 17214 34294
rect 16974 34272 17270 34292
rect 17314 33502 17342 34934
rect 17302 33496 17354 33502
rect 17302 33438 17354 33444
rect 16974 33260 17270 33280
rect 17030 33258 17054 33260
rect 17110 33258 17134 33260
rect 17190 33258 17214 33260
rect 17052 33206 17054 33258
rect 17116 33206 17128 33258
rect 17190 33206 17192 33258
rect 17030 33204 17054 33206
rect 17110 33204 17134 33206
rect 17190 33204 17214 33206
rect 16974 33184 17270 33204
rect 17314 32958 17342 33438
rect 17302 32952 17354 32958
rect 17302 32894 17354 32900
rect 16974 32172 17270 32192
rect 17030 32170 17054 32172
rect 17110 32170 17134 32172
rect 17190 32170 17214 32172
rect 17052 32118 17054 32170
rect 17116 32118 17128 32170
rect 17190 32118 17192 32170
rect 17030 32116 17054 32118
rect 17110 32116 17134 32118
rect 17190 32116 17214 32118
rect 16974 32096 17270 32116
rect 17302 31864 17354 31870
rect 17300 31832 17302 31841
rect 17354 31832 17356 31841
rect 17300 31767 17356 31776
rect 16658 31388 16710 31394
rect 16658 31330 16710 31336
rect 16382 30708 16434 30714
rect 16382 30650 16434 30656
rect 16394 29762 16422 30650
rect 16382 29756 16434 29762
rect 16382 29698 16434 29704
rect 16670 28742 16698 31330
rect 16974 31084 17270 31104
rect 17030 31082 17054 31084
rect 17110 31082 17134 31084
rect 17190 31082 17214 31084
rect 17052 31030 17054 31082
rect 17116 31030 17128 31082
rect 17190 31030 17192 31082
rect 17030 31028 17054 31030
rect 17110 31028 17134 31030
rect 17190 31028 17214 31030
rect 16974 31008 17270 31028
rect 16748 30880 16804 30889
rect 16748 30815 16750 30824
rect 16802 30815 16804 30824
rect 16750 30786 16802 30792
rect 17406 30102 17434 35190
rect 17670 34448 17722 34454
rect 17670 34390 17722 34396
rect 17578 34244 17630 34250
rect 17578 34186 17630 34192
rect 17590 34114 17618 34186
rect 17578 34108 17630 34114
rect 17578 34050 17630 34056
rect 17486 34040 17538 34046
rect 17486 33982 17538 33988
rect 17498 32414 17526 33982
rect 17590 33706 17618 34050
rect 17682 33910 17710 34390
rect 17762 34176 17814 34182
rect 17762 34118 17814 34124
rect 17670 33904 17722 33910
rect 17670 33846 17722 33852
rect 17578 33700 17630 33706
rect 17578 33642 17630 33648
rect 17486 32408 17538 32414
rect 17486 32350 17538 32356
rect 17774 31326 17802 34118
rect 17854 31932 17906 31938
rect 17854 31874 17906 31880
rect 17866 31802 17894 31874
rect 17854 31796 17906 31802
rect 17854 31738 17906 31744
rect 17762 31320 17814 31326
rect 17762 31262 17814 31268
rect 17670 30980 17722 30986
rect 17670 30922 17722 30928
rect 17578 30844 17630 30850
rect 17578 30786 17630 30792
rect 17590 30646 17618 30786
rect 17578 30640 17630 30646
rect 17578 30582 17630 30588
rect 17486 30232 17538 30238
rect 17486 30174 17538 30180
rect 17394 30096 17446 30102
rect 17394 30038 17446 30044
rect 16974 29996 17270 30016
rect 17030 29994 17054 29996
rect 17110 29994 17134 29996
rect 17190 29994 17214 29996
rect 17052 29942 17054 29994
rect 17116 29942 17128 29994
rect 17190 29942 17192 29994
rect 17030 29940 17054 29942
rect 17110 29940 17134 29942
rect 17190 29940 17214 29942
rect 16974 29920 17270 29940
rect 17498 29898 17526 30174
rect 17486 29892 17538 29898
rect 17486 29834 17538 29840
rect 17302 29620 17354 29626
rect 17302 29562 17354 29568
rect 16974 28908 17270 28928
rect 17030 28906 17054 28908
rect 17110 28906 17134 28908
rect 17190 28906 17214 28908
rect 17052 28854 17054 28906
rect 17116 28854 17128 28906
rect 17190 28854 17192 28906
rect 17030 28852 17054 28854
rect 17110 28852 17134 28854
rect 17190 28852 17214 28854
rect 16974 28832 17270 28852
rect 17314 28810 17342 29562
rect 17498 29150 17526 29834
rect 17486 29144 17538 29150
rect 17486 29086 17538 29092
rect 17590 29014 17618 30582
rect 17682 29694 17710 30922
rect 17774 30889 17802 31262
rect 17760 30880 17816 30889
rect 17760 30815 17816 30824
rect 17762 30164 17814 30170
rect 17762 30106 17814 30112
rect 17670 29688 17722 29694
rect 17670 29630 17722 29636
rect 17578 29008 17630 29014
rect 17578 28950 17630 28956
rect 17302 28804 17354 28810
rect 17302 28746 17354 28752
rect 16658 28736 16710 28742
rect 16658 28678 16710 28684
rect 17302 28668 17354 28674
rect 17302 28610 17354 28616
rect 16750 28600 16802 28606
rect 16750 28542 16802 28548
rect 16290 28464 16342 28470
rect 16290 28406 16342 28412
rect 16198 28124 16250 28130
rect 16198 28066 16250 28072
rect 16658 28124 16710 28130
rect 16658 28066 16710 28072
rect 16106 28056 16158 28062
rect 16106 27998 16158 28004
rect 16670 27722 16698 28066
rect 16658 27716 16710 27722
rect 16658 27658 16710 27664
rect 16106 27580 16158 27586
rect 16026 27540 16106 27568
rect 12426 27444 12478 27450
rect 12426 27386 12478 27392
rect 13162 27444 13214 27450
rect 13162 27386 13214 27392
rect 15186 27444 15238 27450
rect 15186 27386 15238 27392
rect 12150 27376 12202 27382
rect 12150 27318 12202 27324
rect 12162 27178 12190 27318
rect 12150 27172 12202 27178
rect 12150 27114 12202 27120
rect 12058 27036 12110 27042
rect 12058 26978 12110 26984
rect 12438 26974 12466 27386
rect 13174 27178 13202 27386
rect 15278 27376 15330 27382
rect 15278 27318 15330 27324
rect 14310 27276 14606 27296
rect 14366 27274 14390 27276
rect 14446 27274 14470 27276
rect 14526 27274 14550 27276
rect 14388 27222 14390 27274
rect 14452 27222 14464 27274
rect 14526 27222 14528 27274
rect 14366 27220 14390 27222
rect 14446 27220 14470 27222
rect 14526 27220 14550 27222
rect 14310 27200 14606 27220
rect 12702 27172 12754 27178
rect 12702 27114 12754 27120
rect 13162 27172 13214 27178
rect 13162 27114 13214 27120
rect 12714 26974 12742 27114
rect 12426 26968 12478 26974
rect 12426 26910 12478 26916
rect 12702 26968 12754 26974
rect 12702 26910 12754 26916
rect 11646 26732 11942 26752
rect 11702 26730 11726 26732
rect 11782 26730 11806 26732
rect 11862 26730 11886 26732
rect 11724 26678 11726 26730
rect 11788 26678 11800 26730
rect 11862 26678 11864 26730
rect 11702 26676 11726 26678
rect 11782 26676 11806 26678
rect 11862 26676 11886 26678
rect 11646 26656 11942 26676
rect 11506 26356 11558 26362
rect 11506 26298 11558 26304
rect 15290 24390 15318 27318
rect 15658 27042 15686 27522
rect 16026 27382 16054 27540
rect 16106 27522 16158 27528
rect 16474 27580 16526 27586
rect 16474 27522 16526 27528
rect 16566 27580 16618 27586
rect 16566 27522 16618 27528
rect 16014 27376 16066 27382
rect 16014 27318 16066 27324
rect 16486 27178 16514 27522
rect 16578 27489 16606 27522
rect 16564 27480 16620 27489
rect 16564 27415 16620 27424
rect 16474 27172 16526 27178
rect 16474 27114 16526 27120
rect 16566 27172 16618 27178
rect 16566 27114 16618 27120
rect 15646 27036 15698 27042
rect 15646 26978 15698 26984
rect 16578 26974 16606 27114
rect 16566 26968 16618 26974
rect 16566 26910 16618 26916
rect 16762 25546 16790 28542
rect 17314 27926 17342 28610
rect 17670 28600 17722 28606
rect 17670 28542 17722 28548
rect 17394 28192 17446 28198
rect 17394 28134 17446 28140
rect 17406 27926 17434 28134
rect 17302 27920 17354 27926
rect 17302 27862 17354 27868
rect 17394 27920 17446 27926
rect 17394 27862 17446 27868
rect 16974 27820 17270 27840
rect 17030 27818 17054 27820
rect 17110 27818 17134 27820
rect 17190 27818 17214 27820
rect 17052 27766 17054 27818
rect 17116 27766 17128 27818
rect 17190 27766 17192 27818
rect 17030 27764 17054 27766
rect 17110 27764 17134 27766
rect 17190 27764 17214 27766
rect 16974 27744 17270 27764
rect 17682 27722 17710 28542
rect 17774 28130 17802 30106
rect 17958 30050 17986 37722
rect 18222 32408 18274 32414
rect 18222 32350 18274 32356
rect 18234 32006 18262 32350
rect 18222 32000 18274 32006
rect 18222 31942 18274 31948
rect 18130 31864 18182 31870
rect 18130 31806 18182 31812
rect 18142 31190 18170 31806
rect 18130 31184 18182 31190
rect 18130 31126 18182 31132
rect 18038 30776 18090 30782
rect 18038 30718 18090 30724
rect 18050 30238 18078 30718
rect 18038 30232 18090 30238
rect 18038 30174 18090 30180
rect 17866 30022 17986 30050
rect 17866 28810 17894 30022
rect 18326 29558 18354 39286
rect 18786 39078 18814 39558
rect 19062 39146 19090 39966
rect 20246 39888 20298 39894
rect 20246 39830 20298 39836
rect 19638 39244 19934 39264
rect 19694 39242 19718 39244
rect 19774 39242 19798 39244
rect 19854 39242 19878 39244
rect 19716 39190 19718 39242
rect 19780 39190 19792 39242
rect 19854 39190 19856 39242
rect 19694 39188 19718 39190
rect 19774 39188 19798 39190
rect 19854 39188 19878 39190
rect 19638 39168 19934 39188
rect 19050 39140 19102 39146
rect 19050 39082 19102 39088
rect 18774 39072 18826 39078
rect 18774 39014 18826 39020
rect 20258 38942 20286 39830
rect 19050 38936 19102 38942
rect 19050 38878 19102 38884
rect 20246 38936 20298 38942
rect 20246 38878 20298 38884
rect 18590 38256 18642 38262
rect 18590 38198 18642 38204
rect 18498 35808 18550 35814
rect 18498 35750 18550 35756
rect 18510 35542 18538 35750
rect 18498 35536 18550 35542
rect 18498 35478 18550 35484
rect 18406 34448 18458 34454
rect 18406 34390 18458 34396
rect 18418 34182 18446 34390
rect 18406 34176 18458 34182
rect 18406 34118 18458 34124
rect 18510 33065 18538 35478
rect 18496 33056 18552 33065
rect 18496 32991 18552 33000
rect 18314 29552 18366 29558
rect 18314 29494 18366 29500
rect 17854 28804 17906 28810
rect 17854 28746 17906 28752
rect 18602 28742 18630 38198
rect 18958 35332 19010 35338
rect 18958 35274 19010 35280
rect 18970 35202 18998 35274
rect 18958 35196 19010 35202
rect 18958 35138 19010 35144
rect 18774 33496 18826 33502
rect 18774 33438 18826 33444
rect 18682 33428 18734 33434
rect 18682 33370 18734 33376
rect 18694 33162 18722 33370
rect 18682 33156 18734 33162
rect 18682 33098 18734 33104
rect 18694 33026 18722 33098
rect 18682 33020 18734 33026
rect 18682 32962 18734 32968
rect 18694 32006 18722 32962
rect 18786 32618 18814 33438
rect 18970 33094 18998 35138
rect 18958 33088 19010 33094
rect 18958 33030 19010 33036
rect 18866 32884 18918 32890
rect 18866 32826 18918 32832
rect 18774 32612 18826 32618
rect 18774 32554 18826 32560
rect 18682 32000 18734 32006
rect 18682 31942 18734 31948
rect 18694 31802 18722 31942
rect 18682 31796 18734 31802
rect 18682 31738 18734 31744
rect 18878 31394 18906 32826
rect 18956 31968 19012 31977
rect 18956 31903 18958 31912
rect 19010 31903 19012 31912
rect 18958 31874 19010 31880
rect 18866 31388 18918 31394
rect 18866 31330 18918 31336
rect 18682 31184 18734 31190
rect 18682 31126 18734 31132
rect 18694 30306 18722 31126
rect 18878 30850 18906 31330
rect 18958 31320 19010 31326
rect 18958 31262 19010 31268
rect 18970 31190 18998 31262
rect 18958 31184 19010 31190
rect 18958 31126 19010 31132
rect 18866 30844 18918 30850
rect 18866 30786 18918 30792
rect 18866 30640 18918 30646
rect 18866 30582 18918 30588
rect 18878 30442 18906 30582
rect 18866 30436 18918 30442
rect 18866 30378 18918 30384
rect 18682 30300 18734 30306
rect 18682 30242 18734 30248
rect 18970 29898 18998 31126
rect 18958 29892 19010 29898
rect 18958 29834 19010 29840
rect 18774 29280 18826 29286
rect 18774 29222 18826 29228
rect 18958 29280 19010 29286
rect 18958 29222 19010 29228
rect 18786 29150 18814 29222
rect 18774 29144 18826 29150
rect 18774 29086 18826 29092
rect 18590 28736 18642 28742
rect 18590 28678 18642 28684
rect 18970 28674 18998 29222
rect 18958 28668 19010 28674
rect 18958 28610 19010 28616
rect 18222 28532 18274 28538
rect 18222 28474 18274 28480
rect 18234 28130 18262 28474
rect 17762 28124 17814 28130
rect 17762 28066 17814 28072
rect 18222 28124 18274 28130
rect 18222 28066 18274 28072
rect 17670 27716 17722 27722
rect 17670 27658 17722 27664
rect 17578 27648 17630 27654
rect 17116 27616 17172 27625
rect 17578 27590 17630 27596
rect 17116 27551 17172 27560
rect 17130 27382 17158 27551
rect 17026 27376 17078 27382
rect 17026 27318 17078 27324
rect 17118 27376 17170 27382
rect 17118 27318 17170 27324
rect 17038 27042 17066 27318
rect 17590 27110 17618 27590
rect 17682 27518 17710 27658
rect 17670 27512 17722 27518
rect 17670 27454 17722 27460
rect 17578 27104 17630 27110
rect 17578 27046 17630 27052
rect 17026 27036 17078 27042
rect 17026 26978 17078 26984
rect 17682 26974 17710 27454
rect 17774 27110 17802 28066
rect 18866 28056 18918 28062
rect 18864 28024 18866 28033
rect 18918 28024 18920 28033
rect 19062 27994 19090 38878
rect 19638 38156 19934 38176
rect 19694 38154 19718 38156
rect 19774 38154 19798 38156
rect 19854 38154 19878 38156
rect 19716 38102 19718 38154
rect 19780 38102 19792 38154
rect 19854 38102 19856 38154
rect 19694 38100 19718 38102
rect 19774 38100 19798 38102
rect 19854 38100 19878 38102
rect 19638 38080 19934 38100
rect 20258 38058 20286 38878
rect 20246 38052 20298 38058
rect 20246 37994 20298 38000
rect 20626 37922 20654 41462
rect 20614 37916 20666 37922
rect 20614 37858 20666 37864
rect 20430 37848 20482 37854
rect 20430 37790 20482 37796
rect 20338 37780 20390 37786
rect 20338 37722 20390 37728
rect 19418 37508 19470 37514
rect 19418 37450 19470 37456
rect 19430 35338 19458 37450
rect 19638 37068 19934 37088
rect 19694 37066 19718 37068
rect 19774 37066 19798 37068
rect 19854 37066 19878 37068
rect 19716 37014 19718 37066
rect 19780 37014 19792 37066
rect 19854 37014 19856 37066
rect 19694 37012 19718 37014
rect 19774 37012 19798 37014
rect 19854 37012 19878 37014
rect 19638 36992 19934 37012
rect 20350 36834 20378 37722
rect 20338 36828 20390 36834
rect 20338 36770 20390 36776
rect 20154 36080 20206 36086
rect 20154 36022 20206 36028
rect 19638 35980 19934 36000
rect 19694 35978 19718 35980
rect 19774 35978 19798 35980
rect 19854 35978 19878 35980
rect 19716 35926 19718 35978
rect 19780 35926 19792 35978
rect 19854 35926 19856 35978
rect 19694 35924 19718 35926
rect 19774 35924 19798 35926
rect 19854 35924 19878 35926
rect 19638 35904 19934 35924
rect 19418 35332 19470 35338
rect 19418 35274 19470 35280
rect 20166 35270 20194 36022
rect 20154 35264 20206 35270
rect 20154 35206 20206 35212
rect 19638 34892 19934 34912
rect 19694 34890 19718 34892
rect 19774 34890 19798 34892
rect 19854 34890 19878 34892
rect 19716 34838 19718 34890
rect 19780 34838 19792 34890
rect 19854 34838 19856 34890
rect 19694 34836 19718 34838
rect 19774 34836 19798 34838
rect 19854 34836 19878 34838
rect 19638 34816 19934 34836
rect 20166 34114 20194 35206
rect 20154 34108 20206 34114
rect 20154 34050 20206 34056
rect 19638 33804 19934 33824
rect 19694 33802 19718 33804
rect 19774 33802 19798 33804
rect 19854 33802 19878 33804
rect 19716 33750 19718 33802
rect 19780 33750 19792 33802
rect 19854 33750 19856 33802
rect 19694 33748 19718 33750
rect 19774 33748 19798 33750
rect 19854 33748 19878 33750
rect 19638 33728 19934 33748
rect 19326 33088 19378 33094
rect 19326 33030 19378 33036
rect 19142 32272 19194 32278
rect 19142 32214 19194 32220
rect 19154 31938 19182 32214
rect 19142 31932 19194 31938
rect 19142 31874 19194 31880
rect 19154 31530 19182 31874
rect 19338 31734 19366 33030
rect 19638 32716 19934 32736
rect 19694 32714 19718 32716
rect 19774 32714 19798 32716
rect 19854 32714 19878 32716
rect 19716 32662 19718 32714
rect 19780 32662 19792 32714
rect 19854 32662 19856 32714
rect 19694 32660 19718 32662
rect 19774 32660 19798 32662
rect 19854 32660 19878 32662
rect 19638 32640 19934 32660
rect 20442 32618 20470 37790
rect 20522 35604 20574 35610
rect 20522 35546 20574 35552
rect 20534 34590 20562 35546
rect 20522 34584 20574 34590
rect 20522 34526 20574 34532
rect 20614 34584 20666 34590
rect 20614 34526 20666 34532
rect 20626 34454 20654 34526
rect 20614 34448 20666 34454
rect 20614 34390 20666 34396
rect 20430 32612 20482 32618
rect 20430 32554 20482 32560
rect 19418 31864 19470 31870
rect 19416 31832 19418 31841
rect 19470 31832 19472 31841
rect 19416 31767 19472 31776
rect 19326 31728 19378 31734
rect 19326 31670 19378 31676
rect 19638 31628 19934 31648
rect 19694 31626 19718 31628
rect 19774 31626 19798 31628
rect 19854 31626 19878 31628
rect 19716 31574 19718 31626
rect 19780 31574 19792 31626
rect 19854 31574 19856 31626
rect 19694 31572 19718 31574
rect 19774 31572 19798 31574
rect 19854 31572 19878 31574
rect 19638 31552 19934 31572
rect 19142 31524 19194 31530
rect 19142 31466 19194 31472
rect 20718 31258 20746 43312
rect 20890 40976 20942 40982
rect 20890 40918 20942 40924
rect 20902 40438 20930 40918
rect 22006 40574 22034 43312
rect 22302 41964 22598 41984
rect 22358 41962 22382 41964
rect 22438 41962 22462 41964
rect 22518 41962 22542 41964
rect 22380 41910 22382 41962
rect 22444 41910 22456 41962
rect 22518 41910 22520 41962
rect 22358 41908 22382 41910
rect 22438 41908 22462 41910
rect 22518 41908 22542 41910
rect 22302 41888 22598 41908
rect 22302 40876 22598 40896
rect 22358 40874 22382 40876
rect 22438 40874 22462 40876
rect 22518 40874 22542 40876
rect 22380 40822 22382 40874
rect 22444 40822 22456 40874
rect 22518 40822 22520 40874
rect 22358 40820 22382 40822
rect 22438 40820 22462 40822
rect 22518 40820 22542 40822
rect 22302 40800 22598 40820
rect 21258 40568 21310 40574
rect 21258 40510 21310 40516
rect 21994 40568 22046 40574
rect 21994 40510 22046 40516
rect 20890 40432 20942 40438
rect 20890 40374 20942 40380
rect 20902 40098 20930 40374
rect 20890 40092 20942 40098
rect 20890 40034 20942 40040
rect 20902 37938 20930 40034
rect 21270 39622 21298 40510
rect 22302 39788 22598 39808
rect 22358 39786 22382 39788
rect 22438 39786 22462 39788
rect 22518 39786 22542 39788
rect 22380 39734 22382 39786
rect 22444 39734 22456 39786
rect 22518 39734 22520 39786
rect 22358 39732 22382 39734
rect 22438 39732 22462 39734
rect 22518 39732 22542 39734
rect 22302 39712 22598 39732
rect 21258 39616 21310 39622
rect 21258 39558 21310 39564
rect 21074 39480 21126 39486
rect 21074 39422 21126 39428
rect 21086 39146 21114 39422
rect 21074 39140 21126 39146
rect 21074 39082 21126 39088
rect 22302 38700 22598 38720
rect 22358 38698 22382 38700
rect 22438 38698 22462 38700
rect 22518 38698 22542 38700
rect 22380 38646 22382 38698
rect 22444 38646 22456 38698
rect 22518 38646 22520 38698
rect 22358 38644 22382 38646
rect 22438 38644 22462 38646
rect 22518 38644 22542 38646
rect 22302 38624 22598 38644
rect 20902 37922 21114 37938
rect 20902 37916 21126 37922
rect 20902 37910 21074 37916
rect 20902 37378 20930 37910
rect 21074 37858 21126 37864
rect 22302 37612 22598 37632
rect 22358 37610 22382 37612
rect 22438 37610 22462 37612
rect 22518 37610 22542 37612
rect 22380 37558 22382 37610
rect 22444 37558 22456 37610
rect 22518 37558 22520 37610
rect 22358 37556 22382 37558
rect 22438 37556 22462 37558
rect 22518 37556 22542 37558
rect 22302 37536 22598 37556
rect 20890 37372 20942 37378
rect 20890 37314 20942 37320
rect 21350 37304 21402 37310
rect 21350 37246 21402 37252
rect 21362 36970 21390 37246
rect 21534 37168 21586 37174
rect 21534 37110 21586 37116
rect 21350 36964 21402 36970
rect 21350 36906 21402 36912
rect 21258 36760 21310 36766
rect 21258 36702 21310 36708
rect 21074 35672 21126 35678
rect 21074 35614 21126 35620
rect 21086 35202 21114 35614
rect 21166 35332 21218 35338
rect 21166 35274 21218 35280
rect 21074 35196 21126 35202
rect 21074 35138 21126 35144
rect 21178 34794 21206 35274
rect 21166 34788 21218 34794
rect 21166 34730 21218 34736
rect 21270 34658 21298 36702
rect 21546 36698 21574 37110
rect 22822 36896 22874 36902
rect 22822 36838 22874 36844
rect 21534 36692 21586 36698
rect 21534 36634 21586 36640
rect 21546 36290 21574 36634
rect 22302 36524 22598 36544
rect 22358 36522 22382 36524
rect 22438 36522 22462 36524
rect 22518 36522 22542 36524
rect 22380 36470 22382 36522
rect 22444 36470 22456 36522
rect 22518 36470 22520 36522
rect 22358 36468 22382 36470
rect 22438 36468 22462 36470
rect 22518 36468 22542 36470
rect 22302 36448 22598 36468
rect 21534 36284 21586 36290
rect 21534 36226 21586 36232
rect 21534 36080 21586 36086
rect 21534 36022 21586 36028
rect 21546 35610 21574 36022
rect 22834 35882 22862 36838
rect 21626 35876 21678 35882
rect 21626 35818 21678 35824
rect 22822 35876 22874 35882
rect 22822 35818 22874 35824
rect 21534 35604 21586 35610
rect 21534 35546 21586 35552
rect 21258 34652 21310 34658
rect 21258 34594 21310 34600
rect 20798 33496 20850 33502
rect 20798 33438 20850 33444
rect 20810 33366 20838 33438
rect 21638 33366 21666 35818
rect 22822 35604 22874 35610
rect 22822 35546 22874 35552
rect 22302 35436 22598 35456
rect 22358 35434 22382 35436
rect 22438 35434 22462 35436
rect 22518 35434 22542 35436
rect 22380 35382 22382 35434
rect 22444 35382 22456 35434
rect 22518 35382 22520 35434
rect 22358 35380 22382 35382
rect 22438 35380 22462 35382
rect 22518 35380 22542 35382
rect 22302 35360 22598 35380
rect 21718 35196 21770 35202
rect 21718 35138 21770 35144
rect 21730 33978 21758 35138
rect 22730 35060 22782 35066
rect 22730 35002 22782 35008
rect 22302 34348 22598 34368
rect 22358 34346 22382 34348
rect 22438 34346 22462 34348
rect 22518 34346 22542 34348
rect 22380 34294 22382 34346
rect 22444 34294 22456 34346
rect 22518 34294 22520 34346
rect 22358 34292 22382 34294
rect 22438 34292 22462 34294
rect 22518 34292 22542 34294
rect 22302 34272 22598 34292
rect 22742 34114 22770 35002
rect 22834 34794 22862 35546
rect 22822 34788 22874 34794
rect 22822 34730 22874 34736
rect 23006 34448 23058 34454
rect 23006 34390 23058 34396
rect 23018 34182 23046 34390
rect 23006 34176 23058 34182
rect 23006 34118 23058 34124
rect 22730 34108 22782 34114
rect 22730 34050 22782 34056
rect 21718 33972 21770 33978
rect 21718 33914 21770 33920
rect 20798 33360 20850 33366
rect 20798 33302 20850 33308
rect 21626 33360 21678 33366
rect 21626 33302 21678 33308
rect 20810 31802 20838 33302
rect 21638 33162 21666 33302
rect 22302 33260 22598 33280
rect 22358 33258 22382 33260
rect 22438 33258 22462 33260
rect 22518 33258 22542 33260
rect 22380 33206 22382 33258
rect 22444 33206 22456 33258
rect 22518 33206 22520 33258
rect 22358 33204 22382 33206
rect 22438 33204 22462 33206
rect 22518 33204 22542 33206
rect 22302 33184 22598 33204
rect 21626 33156 21678 33162
rect 21626 33098 21678 33104
rect 21074 32816 21126 32822
rect 21074 32758 21126 32764
rect 21086 32482 21114 32758
rect 22086 32544 22138 32550
rect 22086 32486 22138 32492
rect 21074 32476 21126 32482
rect 21074 32418 21126 32424
rect 21350 32408 21402 32414
rect 21350 32350 21402 32356
rect 20798 31796 20850 31802
rect 20798 31738 20850 31744
rect 20706 31252 20758 31258
rect 20706 31194 20758 31200
rect 19878 31184 19930 31190
rect 19878 31126 19930 31132
rect 19890 30918 19918 31126
rect 19878 30912 19930 30918
rect 19878 30854 19930 30860
rect 19510 30708 19562 30714
rect 19510 30650 19562 30656
rect 19522 30322 19550 30650
rect 19890 30628 19918 30854
rect 19890 30600 20010 30628
rect 19638 30540 19934 30560
rect 19694 30538 19718 30540
rect 19774 30538 19798 30540
rect 19854 30538 19878 30540
rect 19716 30486 19718 30538
rect 19780 30486 19792 30538
rect 19854 30486 19856 30538
rect 19694 30484 19718 30486
rect 19774 30484 19798 30486
rect 19854 30484 19878 30486
rect 19638 30464 19934 30484
rect 19600 30336 19656 30345
rect 19522 30294 19600 30322
rect 19600 30271 19602 30280
rect 19654 30271 19656 30280
rect 19602 30242 19654 30248
rect 19614 29762 19642 30242
rect 19602 29756 19654 29762
rect 19602 29698 19654 29704
rect 19638 29452 19934 29472
rect 19694 29450 19718 29452
rect 19774 29450 19798 29452
rect 19854 29450 19878 29452
rect 19716 29398 19718 29450
rect 19780 29398 19792 29450
rect 19854 29398 19856 29450
rect 19694 29396 19718 29398
rect 19774 29396 19798 29398
rect 19854 29396 19878 29398
rect 19638 29376 19934 29396
rect 19982 29354 20010 30600
rect 19326 29348 19378 29354
rect 19326 29290 19378 29296
rect 19970 29348 20022 29354
rect 19970 29290 20022 29296
rect 19338 29014 19366 29290
rect 19326 29008 19378 29014
rect 19326 28950 19378 28956
rect 19338 28130 19366 28950
rect 20982 28532 21034 28538
rect 20982 28474 21034 28480
rect 19638 28364 19934 28384
rect 19694 28362 19718 28364
rect 19774 28362 19798 28364
rect 19854 28362 19878 28364
rect 19716 28310 19718 28362
rect 19780 28310 19792 28362
rect 19854 28310 19856 28362
rect 19694 28308 19718 28310
rect 19774 28308 19798 28310
rect 19854 28308 19878 28310
rect 19638 28288 19934 28308
rect 20994 28266 21022 28474
rect 20982 28260 21034 28266
rect 20982 28202 21034 28208
rect 19326 28124 19378 28130
rect 19326 28066 19378 28072
rect 20994 28062 21022 28202
rect 21362 28062 21390 32350
rect 21810 31932 21862 31938
rect 21810 31874 21862 31880
rect 21534 31864 21586 31870
rect 21534 31806 21586 31812
rect 21546 31734 21574 31806
rect 21822 31734 21850 31874
rect 21534 31728 21586 31734
rect 21534 31670 21586 31676
rect 21810 31728 21862 31734
rect 21810 31670 21862 31676
rect 21822 29694 21850 31670
rect 22098 31530 22126 32486
rect 22302 32172 22598 32192
rect 22358 32170 22382 32172
rect 22438 32170 22462 32172
rect 22518 32170 22542 32172
rect 22380 32118 22382 32170
rect 22444 32118 22456 32170
rect 22518 32118 22520 32170
rect 22358 32116 22382 32118
rect 22438 32116 22462 32118
rect 22518 32116 22542 32118
rect 22302 32096 22598 32116
rect 22086 31524 22138 31530
rect 22086 31466 22138 31472
rect 22914 31184 22966 31190
rect 22914 31126 22966 31132
rect 22302 31084 22598 31104
rect 22358 31082 22382 31084
rect 22438 31082 22462 31084
rect 22518 31082 22542 31084
rect 22380 31030 22382 31082
rect 22444 31030 22456 31082
rect 22518 31030 22520 31082
rect 22358 31028 22382 31030
rect 22438 31028 22462 31030
rect 22518 31028 22542 31030
rect 22302 31008 22598 31028
rect 22822 30164 22874 30170
rect 22822 30106 22874 30112
rect 22302 29996 22598 30016
rect 22358 29994 22382 29996
rect 22438 29994 22462 29996
rect 22518 29994 22542 29996
rect 22380 29942 22382 29994
rect 22444 29942 22456 29994
rect 22518 29942 22520 29994
rect 22358 29940 22382 29942
rect 22438 29940 22462 29942
rect 22518 29940 22542 29942
rect 22302 29920 22598 29940
rect 22728 29928 22784 29937
rect 22728 29863 22730 29872
rect 22782 29863 22784 29872
rect 22730 29834 22782 29840
rect 22834 29830 22862 30106
rect 22822 29824 22874 29830
rect 22822 29766 22874 29772
rect 21810 29688 21862 29694
rect 21810 29630 21862 29636
rect 22822 29620 22874 29626
rect 22822 29562 22874 29568
rect 22730 29212 22782 29218
rect 22730 29154 22782 29160
rect 22302 28908 22598 28928
rect 22358 28906 22382 28908
rect 22438 28906 22462 28908
rect 22518 28906 22542 28908
rect 22380 28854 22382 28906
rect 22444 28854 22456 28906
rect 22518 28854 22520 28906
rect 22358 28852 22382 28854
rect 22438 28852 22462 28854
rect 22518 28852 22542 28854
rect 22302 28832 22598 28852
rect 22742 28674 22770 29154
rect 22730 28668 22782 28674
rect 22730 28610 22782 28616
rect 22834 28577 22862 29562
rect 22820 28568 22876 28577
rect 22820 28503 22876 28512
rect 22638 28464 22690 28470
rect 22638 28406 22690 28412
rect 20982 28056 21034 28062
rect 20982 27998 21034 28004
rect 21350 28056 21402 28062
rect 21350 27998 21402 28004
rect 18864 27959 18920 27968
rect 19050 27988 19102 27994
rect 19050 27930 19102 27936
rect 20890 27920 20942 27926
rect 20890 27862 20942 27868
rect 18590 27580 18642 27586
rect 18774 27580 18826 27586
rect 18642 27540 18774 27568
rect 18590 27522 18642 27528
rect 18774 27522 18826 27528
rect 17762 27104 17814 27110
rect 17762 27046 17814 27052
rect 17774 26974 17802 27046
rect 17670 26968 17722 26974
rect 17670 26910 17722 26916
rect 17762 26968 17814 26974
rect 17762 26910 17814 26916
rect 18786 26838 18814 27522
rect 20902 27518 20930 27862
rect 22302 27820 22598 27840
rect 22358 27818 22382 27820
rect 22438 27818 22462 27820
rect 22518 27818 22542 27820
rect 22380 27766 22382 27818
rect 22444 27766 22456 27818
rect 22518 27766 22520 27818
rect 22358 27764 22382 27766
rect 22438 27764 22462 27766
rect 22518 27764 22542 27766
rect 22302 27744 22598 27764
rect 22650 27586 22678 28406
rect 22546 27580 22598 27586
rect 22546 27522 22598 27528
rect 22638 27580 22690 27586
rect 22638 27522 22690 27528
rect 20890 27512 20942 27518
rect 20890 27454 20942 27460
rect 19142 27444 19194 27450
rect 19142 27386 19194 27392
rect 19154 26974 19182 27386
rect 19638 27276 19934 27296
rect 19694 27274 19718 27276
rect 19774 27274 19798 27276
rect 19854 27274 19878 27276
rect 19716 27222 19718 27274
rect 19780 27222 19792 27274
rect 19854 27222 19856 27274
rect 19694 27220 19718 27222
rect 19774 27220 19798 27222
rect 19854 27220 19878 27222
rect 19638 27200 19934 27220
rect 22558 27042 22586 27522
rect 22926 27382 22954 31126
rect 23098 30776 23150 30782
rect 23098 30718 23150 30724
rect 23110 30306 23138 30718
rect 23098 30300 23150 30306
rect 23098 30242 23150 30248
rect 23006 30096 23058 30102
rect 23006 30038 23058 30044
rect 23018 29354 23046 30038
rect 23202 29626 23230 43312
rect 24398 41322 24426 43312
rect 24966 41420 25262 41440
rect 25022 41418 25046 41420
rect 25102 41418 25126 41420
rect 25182 41418 25206 41420
rect 25044 41366 25046 41418
rect 25108 41366 25120 41418
rect 25182 41366 25184 41418
rect 25022 41364 25046 41366
rect 25102 41364 25126 41366
rect 25182 41364 25206 41366
rect 24966 41344 25262 41364
rect 24386 41316 24438 41322
rect 24386 41258 24438 41264
rect 24966 40332 25262 40352
rect 25022 40330 25046 40332
rect 25102 40330 25126 40332
rect 25182 40330 25206 40332
rect 25044 40278 25046 40330
rect 25108 40278 25120 40330
rect 25182 40278 25184 40330
rect 25022 40276 25046 40278
rect 25102 40276 25126 40278
rect 25182 40276 25206 40278
rect 24966 40256 25262 40276
rect 25594 39894 25622 43312
rect 26882 42154 26910 43312
rect 28078 43242 28106 43312
rect 28078 43214 28198 43242
rect 26882 42126 27002 42154
rect 26974 42018 27002 42126
rect 26974 41990 27094 42018
rect 27066 41322 27094 41990
rect 27630 41964 27926 41984
rect 27686 41962 27710 41964
rect 27766 41962 27790 41964
rect 27846 41962 27870 41964
rect 27708 41910 27710 41962
rect 27772 41910 27784 41962
rect 27846 41910 27848 41962
rect 27686 41908 27710 41910
rect 27766 41908 27790 41910
rect 27846 41908 27870 41910
rect 27630 41888 27926 41908
rect 27054 41316 27106 41322
rect 27054 41258 27106 41264
rect 25674 41112 25726 41118
rect 25674 41054 25726 41060
rect 25686 40642 25714 41054
rect 26778 40976 26830 40982
rect 26778 40918 26830 40924
rect 26790 40642 26818 40918
rect 27630 40876 27926 40896
rect 27686 40874 27710 40876
rect 27766 40874 27790 40876
rect 27846 40874 27870 40876
rect 27708 40822 27710 40874
rect 27772 40822 27784 40874
rect 27846 40822 27848 40874
rect 27686 40820 27710 40822
rect 27766 40820 27790 40822
rect 27846 40820 27870 40822
rect 27630 40800 27926 40820
rect 25674 40636 25726 40642
rect 25674 40578 25726 40584
rect 26778 40636 26830 40642
rect 26778 40578 26830 40584
rect 27054 40568 27106 40574
rect 27054 40510 27106 40516
rect 27066 40098 27094 40510
rect 27054 40092 27106 40098
rect 27054 40034 27106 40040
rect 27146 40024 27198 40030
rect 27422 40024 27474 40030
rect 27198 39984 27278 40012
rect 27146 39966 27198 39972
rect 25582 39888 25634 39894
rect 25582 39830 25634 39836
rect 27146 39888 27198 39894
rect 27146 39830 27198 39836
rect 24202 39412 24254 39418
rect 24202 39354 24254 39360
rect 27054 39412 27106 39418
rect 27054 39354 27106 39360
rect 24018 36284 24070 36290
rect 24018 36226 24070 36232
rect 23374 36080 23426 36086
rect 23374 36022 23426 36028
rect 23386 35746 23414 36022
rect 23374 35740 23426 35746
rect 23374 35682 23426 35688
rect 23834 35536 23886 35542
rect 23834 35478 23886 35484
rect 23846 35338 23874 35478
rect 24030 35338 24058 36226
rect 23834 35332 23886 35338
rect 23834 35274 23886 35280
rect 24018 35332 24070 35338
rect 24018 35274 24070 35280
rect 23846 35202 23874 35274
rect 23282 35196 23334 35202
rect 23282 35138 23334 35144
rect 23834 35196 23886 35202
rect 23834 35138 23886 35144
rect 23294 34590 23322 35138
rect 23282 34584 23334 34590
rect 23282 34526 23334 34532
rect 23294 33706 23322 34526
rect 23374 34108 23426 34114
rect 23374 34050 23426 34056
rect 23282 33700 23334 33706
rect 23282 33642 23334 33648
rect 23386 33502 23414 34050
rect 23374 33496 23426 33502
rect 23374 33438 23426 33444
rect 24018 33496 24070 33502
rect 24018 33438 24070 33444
rect 23386 32958 23414 33438
rect 23374 32952 23426 32958
rect 23374 32894 23426 32900
rect 23834 32340 23886 32346
rect 23834 32282 23886 32288
rect 23742 31932 23794 31938
rect 23742 31874 23794 31880
rect 23754 31734 23782 31874
rect 23742 31728 23794 31734
rect 23742 31670 23794 31676
rect 23282 31320 23334 31326
rect 23282 31262 23334 31268
rect 23190 29620 23242 29626
rect 23190 29562 23242 29568
rect 23202 29370 23230 29562
rect 23294 29506 23322 31262
rect 23754 30714 23782 31670
rect 23846 31326 23874 32282
rect 24030 31977 24058 33438
rect 24016 31968 24072 31977
rect 24016 31903 24072 31912
rect 24030 31734 24058 31903
rect 24018 31728 24070 31734
rect 24018 31670 24070 31676
rect 23834 31320 23886 31326
rect 23834 31262 23886 31268
rect 24110 31320 24162 31326
rect 24110 31262 24162 31268
rect 24122 31190 24150 31262
rect 24110 31184 24162 31190
rect 24110 31126 24162 31132
rect 23926 30844 23978 30850
rect 23926 30786 23978 30792
rect 23742 30708 23794 30714
rect 23742 30650 23794 30656
rect 23650 30640 23702 30646
rect 23650 30582 23702 30588
rect 23662 30374 23690 30582
rect 23650 30368 23702 30374
rect 23650 30310 23702 30316
rect 23650 30232 23702 30238
rect 23650 30174 23702 30180
rect 23294 29478 23598 29506
rect 23006 29348 23058 29354
rect 23006 29290 23058 29296
rect 23110 29342 23230 29370
rect 23466 29348 23518 29354
rect 23006 29144 23058 29150
rect 23110 29132 23138 29342
rect 23466 29290 23518 29296
rect 23374 29212 23426 29218
rect 23294 29172 23374 29200
rect 23058 29104 23138 29132
rect 23190 29144 23242 29150
rect 23006 29086 23058 29092
rect 23294 29098 23322 29172
rect 23374 29154 23426 29160
rect 23242 29092 23322 29098
rect 23190 29086 23322 29092
rect 23202 29070 23322 29086
rect 23478 28674 23506 29290
rect 23466 28668 23518 28674
rect 23466 28610 23518 28616
rect 23098 28600 23150 28606
rect 23098 28542 23150 28548
rect 23110 27722 23138 28542
rect 23570 28062 23598 29478
rect 23558 28056 23610 28062
rect 23294 27994 23506 28010
rect 23558 27998 23610 28004
rect 23294 27988 23518 27994
rect 23294 27982 23466 27988
rect 23294 27926 23322 27982
rect 23466 27930 23518 27936
rect 23282 27920 23334 27926
rect 23282 27862 23334 27868
rect 23662 27722 23690 30174
rect 23754 29762 23782 30650
rect 23834 30436 23886 30442
rect 23834 30378 23886 30384
rect 23846 30238 23874 30378
rect 23834 30232 23886 30238
rect 23834 30174 23886 30180
rect 23742 29756 23794 29762
rect 23742 29698 23794 29704
rect 23754 29354 23782 29698
rect 23742 29348 23794 29354
rect 23742 29290 23794 29296
rect 23754 29150 23782 29290
rect 23742 29144 23794 29150
rect 23742 29086 23794 29092
rect 23832 28704 23888 28713
rect 23832 28639 23834 28648
rect 23886 28639 23888 28648
rect 23834 28610 23886 28616
rect 23742 28600 23794 28606
rect 23742 28542 23794 28548
rect 23754 28470 23782 28542
rect 23742 28464 23794 28470
rect 23742 28406 23794 28412
rect 23938 28198 23966 30786
rect 24018 30368 24070 30374
rect 24018 30310 24070 30316
rect 24030 29218 24058 30310
rect 24110 29688 24162 29694
rect 24110 29630 24162 29636
rect 24018 29212 24070 29218
rect 24018 29154 24070 29160
rect 23926 28192 23978 28198
rect 23926 28134 23978 28140
rect 24018 28056 24070 28062
rect 24018 27998 24070 28004
rect 23098 27716 23150 27722
rect 23098 27658 23150 27664
rect 23650 27716 23702 27722
rect 23650 27658 23702 27664
rect 23662 27518 23690 27658
rect 23926 27648 23978 27654
rect 23926 27590 23978 27596
rect 23374 27512 23426 27518
rect 23374 27454 23426 27460
rect 23650 27512 23702 27518
rect 23834 27512 23886 27518
rect 23650 27454 23702 27460
rect 23740 27480 23796 27489
rect 23386 27382 23414 27454
rect 23834 27454 23886 27460
rect 23740 27415 23796 27424
rect 22914 27376 22966 27382
rect 22914 27318 22966 27324
rect 23374 27376 23426 27382
rect 23374 27318 23426 27324
rect 22546 27036 22598 27042
rect 22546 26978 22598 26984
rect 22926 26974 22954 27318
rect 23754 27110 23782 27415
rect 23742 27104 23794 27110
rect 23742 27046 23794 27052
rect 19142 26968 19194 26974
rect 19142 26910 19194 26916
rect 22914 26968 22966 26974
rect 22914 26910 22966 26916
rect 23650 26900 23702 26906
rect 23650 26842 23702 26848
rect 18774 26832 18826 26838
rect 18774 26774 18826 26780
rect 16974 26732 17270 26752
rect 17030 26730 17054 26732
rect 17110 26730 17134 26732
rect 17190 26730 17214 26732
rect 17052 26678 17054 26730
rect 17116 26678 17128 26730
rect 17190 26678 17192 26730
rect 17030 26676 17054 26678
rect 17110 26676 17134 26678
rect 17190 26676 17214 26678
rect 16974 26656 17270 26676
rect 22302 26732 22598 26752
rect 22358 26730 22382 26732
rect 22438 26730 22462 26732
rect 22518 26730 22542 26732
rect 22380 26678 22382 26730
rect 22444 26678 22456 26730
rect 22518 26678 22520 26730
rect 22358 26676 22382 26678
rect 22438 26676 22462 26678
rect 22518 26676 22542 26678
rect 22302 26656 22598 26676
rect 23662 26634 23690 26842
rect 23650 26628 23702 26634
rect 23650 26570 23702 26576
rect 16750 25540 16802 25546
rect 16750 25482 16802 25488
rect 16762 24730 16790 25482
rect 23846 25206 23874 27454
rect 23938 26906 23966 27590
rect 24030 26974 24058 27998
rect 24122 27994 24150 29630
rect 24214 29218 24242 39354
rect 24966 39244 25262 39264
rect 25022 39242 25046 39244
rect 25102 39242 25126 39244
rect 25182 39242 25206 39244
rect 25044 39190 25046 39242
rect 25108 39190 25120 39242
rect 25182 39190 25184 39242
rect 25022 39188 25046 39190
rect 25102 39188 25126 39190
rect 25182 39188 25206 39190
rect 24966 39168 25262 39188
rect 25674 38936 25726 38942
rect 25674 38878 25726 38884
rect 25686 38466 25714 38878
rect 27066 38534 27094 39354
rect 27054 38528 27106 38534
rect 27054 38470 27106 38476
rect 25674 38460 25726 38466
rect 25674 38402 25726 38408
rect 24662 38324 24714 38330
rect 24662 38266 24714 38272
rect 24674 37922 24702 38266
rect 24966 38156 25262 38176
rect 25022 38154 25046 38156
rect 25102 38154 25126 38156
rect 25182 38154 25206 38156
rect 25044 38102 25046 38154
rect 25108 38102 25120 38154
rect 25182 38102 25184 38154
rect 25022 38100 25046 38102
rect 25102 38100 25126 38102
rect 25182 38100 25206 38102
rect 24966 38080 25262 38100
rect 25686 37922 25714 38402
rect 24662 37916 24714 37922
rect 24662 37858 24714 37864
rect 25674 37916 25726 37922
rect 25674 37858 25726 37864
rect 25582 37848 25634 37854
rect 25580 37816 25582 37825
rect 25634 37816 25636 37825
rect 25580 37751 25636 37760
rect 27054 37780 27106 37786
rect 27054 37722 27106 37728
rect 27066 37514 27094 37722
rect 27054 37508 27106 37514
rect 27054 37450 27106 37456
rect 24966 37068 25262 37088
rect 25022 37066 25046 37068
rect 25102 37066 25126 37068
rect 25182 37066 25206 37068
rect 25044 37014 25046 37066
rect 25108 37014 25120 37066
rect 25182 37014 25184 37066
rect 25022 37012 25046 37014
rect 25102 37012 25126 37014
rect 25182 37012 25206 37014
rect 24966 36992 25262 37012
rect 25674 36284 25726 36290
rect 25674 36226 25726 36232
rect 24570 36080 24622 36086
rect 24570 36022 24622 36028
rect 24582 35270 24610 36022
rect 24966 35980 25262 36000
rect 25022 35978 25046 35980
rect 25102 35978 25126 35980
rect 25182 35978 25206 35980
rect 25044 35926 25046 35978
rect 25108 35926 25120 35978
rect 25182 35926 25184 35978
rect 25022 35924 25046 35926
rect 25102 35924 25126 35926
rect 25182 35924 25206 35926
rect 24966 35904 25262 35924
rect 25686 35678 25714 36226
rect 27054 36148 27106 36154
rect 27054 36090 27106 36096
rect 27066 35814 27094 36090
rect 27054 35808 27106 35814
rect 27054 35750 27106 35756
rect 25674 35672 25726 35678
rect 25674 35614 25726 35620
rect 24570 35264 24622 35270
rect 24570 35206 24622 35212
rect 27066 35202 27094 35750
rect 27054 35196 27106 35202
rect 27054 35138 27106 35144
rect 24294 34992 24346 34998
rect 24294 34934 24346 34940
rect 24306 33570 24334 34934
rect 24966 34892 25262 34912
rect 25022 34890 25046 34892
rect 25102 34890 25126 34892
rect 25182 34890 25206 34892
rect 25044 34838 25046 34890
rect 25108 34838 25120 34890
rect 25182 34838 25184 34890
rect 25022 34836 25046 34838
rect 25102 34836 25126 34838
rect 25182 34836 25206 34838
rect 24966 34816 25262 34836
rect 25858 34652 25910 34658
rect 25858 34594 25910 34600
rect 26226 34652 26278 34658
rect 26226 34594 26278 34600
rect 26870 34652 26922 34658
rect 26870 34594 26922 34600
rect 25490 34584 25542 34590
rect 25490 34526 25542 34532
rect 24938 34516 24990 34522
rect 24938 34458 24990 34464
rect 24950 33978 24978 34458
rect 25502 34114 25530 34526
rect 25870 34454 25898 34594
rect 25766 34448 25818 34454
rect 25766 34390 25818 34396
rect 25858 34448 25910 34454
rect 25858 34390 25910 34396
rect 25490 34108 25542 34114
rect 25490 34050 25542 34056
rect 24938 33972 24990 33978
rect 24938 33914 24990 33920
rect 25398 33904 25450 33910
rect 25398 33846 25450 33852
rect 24966 33804 25262 33824
rect 25022 33802 25046 33804
rect 25102 33802 25126 33804
rect 25182 33802 25206 33804
rect 25044 33750 25046 33802
rect 25108 33750 25120 33802
rect 25182 33750 25184 33802
rect 25022 33748 25046 33750
rect 25102 33748 25126 33750
rect 25182 33748 25206 33750
rect 24966 33728 25262 33748
rect 25410 33706 25438 33846
rect 25398 33700 25450 33706
rect 25398 33642 25450 33648
rect 24294 33564 24346 33570
rect 24294 33506 24346 33512
rect 24306 33162 24334 33506
rect 24294 33156 24346 33162
rect 24294 33098 24346 33104
rect 25410 32890 25438 33642
rect 25490 33360 25542 33366
rect 25490 33302 25542 33308
rect 25398 32884 25450 32890
rect 25398 32826 25450 32832
rect 24966 32716 25262 32736
rect 25022 32714 25046 32716
rect 25102 32714 25126 32716
rect 25182 32714 25206 32716
rect 25044 32662 25046 32714
rect 25108 32662 25120 32714
rect 25182 32662 25184 32714
rect 25022 32660 25046 32662
rect 25102 32660 25126 32662
rect 25182 32660 25206 32662
rect 24966 32640 25262 32660
rect 25502 32482 25530 33302
rect 25778 33026 25806 34390
rect 25950 34108 26002 34114
rect 25950 34050 26002 34056
rect 25962 33094 25990 34050
rect 26238 33910 26266 34594
rect 26778 34448 26830 34454
rect 26778 34390 26830 34396
rect 26226 33904 26278 33910
rect 26226 33846 26278 33852
rect 26134 33496 26186 33502
rect 26134 33438 26186 33444
rect 25950 33088 26002 33094
rect 25950 33030 26002 33036
rect 25766 33020 25818 33026
rect 25766 32962 25818 32968
rect 26146 32958 26174 33438
rect 26790 33026 26818 34390
rect 26882 34250 26910 34594
rect 27054 34448 27106 34454
rect 27054 34390 27106 34396
rect 27066 34250 27094 34390
rect 26870 34244 26922 34250
rect 26870 34186 26922 34192
rect 27054 34244 27106 34250
rect 27054 34186 27106 34192
rect 26868 34008 26924 34017
rect 26868 33943 26870 33952
rect 26922 33943 26924 33952
rect 26870 33914 26922 33920
rect 26778 33020 26830 33026
rect 26778 32962 26830 32968
rect 26134 32952 26186 32958
rect 26134 32894 26186 32900
rect 26870 32952 26922 32958
rect 26870 32894 26922 32900
rect 25766 32816 25818 32822
rect 25766 32758 25818 32764
rect 25490 32476 25542 32482
rect 25490 32418 25542 32424
rect 24846 32272 24898 32278
rect 24846 32214 24898 32220
rect 24570 32000 24622 32006
rect 24570 31942 24622 31948
rect 24478 31864 24530 31870
rect 24478 31806 24530 31812
rect 24490 30238 24518 31806
rect 24582 31530 24610 31942
rect 24570 31524 24622 31530
rect 24570 31466 24622 31472
rect 24582 31326 24610 31466
rect 24570 31320 24622 31326
rect 24570 31262 24622 31268
rect 24858 30850 24886 32214
rect 24966 31628 25262 31648
rect 25022 31626 25046 31628
rect 25102 31626 25126 31628
rect 25182 31626 25206 31628
rect 25044 31574 25046 31626
rect 25108 31574 25120 31626
rect 25182 31574 25184 31626
rect 25022 31572 25046 31574
rect 25102 31572 25126 31574
rect 25182 31572 25206 31574
rect 24966 31552 25262 31572
rect 24846 30844 24898 30850
rect 24846 30786 24898 30792
rect 24966 30540 25262 30560
rect 25022 30538 25046 30540
rect 25102 30538 25126 30540
rect 25182 30538 25206 30540
rect 25044 30486 25046 30538
rect 25108 30486 25120 30538
rect 25182 30486 25184 30538
rect 25022 30484 25046 30486
rect 25102 30484 25126 30486
rect 25182 30484 25206 30486
rect 24966 30464 25262 30484
rect 24294 30232 24346 30238
rect 24294 30174 24346 30180
rect 24478 30232 24530 30238
rect 24478 30174 24530 30180
rect 24306 29830 24334 30174
rect 24294 29824 24346 29830
rect 24294 29766 24346 29772
rect 24490 29762 24518 30174
rect 24478 29756 24530 29762
rect 24478 29698 24530 29704
rect 24662 29620 24714 29626
rect 24662 29562 24714 29568
rect 24202 29212 24254 29218
rect 24202 29154 24254 29160
rect 24674 29150 24702 29562
rect 24966 29452 25262 29472
rect 25022 29450 25046 29452
rect 25102 29450 25126 29452
rect 25182 29450 25206 29452
rect 25044 29398 25046 29450
rect 25108 29398 25120 29450
rect 25182 29398 25184 29450
rect 25022 29396 25046 29398
rect 25102 29396 25126 29398
rect 25182 29396 25206 29398
rect 24966 29376 25262 29396
rect 24846 29348 24898 29354
rect 24846 29290 24898 29296
rect 24662 29144 24714 29150
rect 24662 29086 24714 29092
rect 24662 29008 24714 29014
rect 24662 28950 24714 28956
rect 24754 29008 24806 29014
rect 24754 28950 24806 28956
rect 24674 28810 24702 28950
rect 24662 28804 24714 28810
rect 24662 28746 24714 28752
rect 24766 28146 24794 28950
rect 24858 28713 24886 29290
rect 25778 28742 25806 32758
rect 25858 31864 25910 31870
rect 25858 31806 25910 31812
rect 25870 31462 25898 31806
rect 26146 31734 26174 32894
rect 26778 32816 26830 32822
rect 26778 32758 26830 32764
rect 26318 32272 26370 32278
rect 26318 32214 26370 32220
rect 26330 32074 26358 32214
rect 26318 32068 26370 32074
rect 26318 32010 26370 32016
rect 26134 31728 26186 31734
rect 26134 31670 26186 31676
rect 25858 31456 25910 31462
rect 25858 31398 25910 31404
rect 25870 29626 25898 31398
rect 26146 31394 26174 31670
rect 26134 31388 26186 31394
rect 26134 31330 26186 31336
rect 26790 31258 26818 32758
rect 26882 32618 26910 32894
rect 26870 32612 26922 32618
rect 26870 32554 26922 32560
rect 26882 31938 26910 32554
rect 26962 32340 27014 32346
rect 26962 32282 27014 32288
rect 26870 31932 26922 31938
rect 26870 31874 26922 31880
rect 26974 31462 27002 32282
rect 27158 31870 27186 39830
rect 27250 37514 27278 39984
rect 27422 39966 27474 39972
rect 27434 39146 27462 39966
rect 27630 39788 27926 39808
rect 27686 39786 27710 39788
rect 27766 39786 27790 39788
rect 27846 39786 27870 39788
rect 27708 39734 27710 39786
rect 27772 39734 27784 39786
rect 27846 39734 27848 39786
rect 27686 39732 27710 39734
rect 27766 39732 27790 39734
rect 27846 39732 27870 39734
rect 27630 39712 27926 39732
rect 27974 39548 28026 39554
rect 27974 39490 28026 39496
rect 27422 39140 27474 39146
rect 27422 39082 27474 39088
rect 27986 38942 28014 39490
rect 27422 38936 27474 38942
rect 27422 38878 27474 38884
rect 27514 38936 27566 38942
rect 27514 38878 27566 38884
rect 27974 38936 28026 38942
rect 27974 38878 28026 38884
rect 27434 38058 27462 38878
rect 27422 38052 27474 38058
rect 27422 37994 27474 38000
rect 27330 37848 27382 37854
rect 27330 37790 27382 37796
rect 27342 37718 27370 37790
rect 27330 37712 27382 37718
rect 27330 37654 27382 37660
rect 27238 37508 27290 37514
rect 27238 37450 27290 37456
rect 27342 36902 27370 37654
rect 27434 37378 27462 37994
rect 27526 37446 27554 38878
rect 27630 38700 27926 38720
rect 27686 38698 27710 38700
rect 27766 38698 27790 38700
rect 27846 38698 27870 38700
rect 27708 38646 27710 38698
rect 27772 38646 27784 38698
rect 27846 38646 27848 38698
rect 27686 38644 27710 38646
rect 27766 38644 27790 38646
rect 27846 38644 27870 38646
rect 27630 38624 27926 38644
rect 27986 37922 28014 38878
rect 27974 37916 28026 37922
rect 27974 37858 28026 37864
rect 27630 37612 27926 37632
rect 27686 37610 27710 37612
rect 27766 37610 27790 37612
rect 27846 37610 27870 37612
rect 27708 37558 27710 37610
rect 27772 37558 27784 37610
rect 27846 37558 27848 37610
rect 27686 37556 27710 37558
rect 27766 37556 27790 37558
rect 27846 37556 27870 37558
rect 27630 37536 27926 37556
rect 27514 37440 27566 37446
rect 27514 37382 27566 37388
rect 27422 37372 27474 37378
rect 27422 37314 27474 37320
rect 27698 37304 27750 37310
rect 27698 37246 27750 37252
rect 27710 36970 27738 37246
rect 27698 36964 27750 36970
rect 27698 36906 27750 36912
rect 27330 36896 27382 36902
rect 27330 36838 27382 36844
rect 27630 36524 27926 36544
rect 27686 36522 27710 36524
rect 27766 36522 27790 36524
rect 27846 36522 27870 36524
rect 27708 36470 27710 36522
rect 27772 36470 27784 36522
rect 27846 36470 27848 36522
rect 27686 36468 27710 36470
rect 27766 36468 27790 36470
rect 27846 36468 27870 36470
rect 27630 36448 27926 36468
rect 28066 36216 28118 36222
rect 28066 36158 28118 36164
rect 27630 35436 27926 35456
rect 27686 35434 27710 35436
rect 27766 35434 27790 35436
rect 27846 35434 27870 35436
rect 27708 35382 27710 35434
rect 27772 35382 27784 35434
rect 27846 35382 27848 35434
rect 27686 35380 27710 35382
rect 27766 35380 27790 35382
rect 27846 35380 27870 35382
rect 27630 35360 27926 35380
rect 28078 35338 28106 36158
rect 28066 35332 28118 35338
rect 28066 35274 28118 35280
rect 27630 34348 27926 34368
rect 27686 34346 27710 34348
rect 27766 34346 27790 34348
rect 27846 34346 27870 34348
rect 27708 34294 27710 34346
rect 27772 34294 27784 34346
rect 27846 34294 27848 34346
rect 27686 34292 27710 34294
rect 27766 34292 27790 34294
rect 27846 34292 27870 34294
rect 27630 34272 27926 34292
rect 27630 33260 27926 33280
rect 27686 33258 27710 33260
rect 27766 33258 27790 33260
rect 27846 33258 27870 33260
rect 27708 33206 27710 33258
rect 27772 33206 27784 33258
rect 27846 33206 27848 33258
rect 27686 33204 27710 33206
rect 27766 33204 27790 33206
rect 27846 33204 27870 33206
rect 27630 33184 27926 33204
rect 27514 32816 27566 32822
rect 27514 32758 27566 32764
rect 27526 32346 27554 32758
rect 27514 32340 27566 32346
rect 27514 32282 27566 32288
rect 27630 32172 27926 32192
rect 27686 32170 27710 32172
rect 27766 32170 27790 32172
rect 27846 32170 27870 32172
rect 27708 32118 27710 32170
rect 27772 32118 27784 32170
rect 27846 32118 27848 32170
rect 27686 32116 27710 32118
rect 27766 32116 27790 32118
rect 27846 32116 27870 32118
rect 27630 32096 27926 32116
rect 28170 31938 28198 43214
rect 28434 41112 28486 41118
rect 28434 41054 28486 41060
rect 28802 41112 28854 41118
rect 28802 41054 28854 41060
rect 28446 39894 28474 41054
rect 28526 40976 28578 40982
rect 28526 40918 28578 40924
rect 28538 40710 28566 40918
rect 28526 40704 28578 40710
rect 28526 40646 28578 40652
rect 28814 40098 28842 41054
rect 29274 40778 29302 43312
rect 30562 41610 30590 43312
rect 30562 41582 30682 41610
rect 30294 41420 30590 41440
rect 30350 41418 30374 41420
rect 30430 41418 30454 41420
rect 30510 41418 30534 41420
rect 30372 41366 30374 41418
rect 30436 41366 30448 41418
rect 30510 41366 30512 41418
rect 30350 41364 30374 41366
rect 30430 41364 30454 41366
rect 30510 41364 30534 41366
rect 30294 41344 30590 41364
rect 29354 40976 29406 40982
rect 29354 40918 29406 40924
rect 30458 40976 30510 40982
rect 30458 40918 30510 40924
rect 29262 40772 29314 40778
rect 29262 40714 29314 40720
rect 28802 40092 28854 40098
rect 28802 40034 28854 40040
rect 28434 39888 28486 39894
rect 28434 39830 28486 39836
rect 28250 39412 28302 39418
rect 28250 39354 28302 39360
rect 28262 38466 28290 39354
rect 29366 38602 29394 40918
rect 30470 40642 30498 40918
rect 30458 40636 30510 40642
rect 30458 40578 30510 40584
rect 30294 40332 30590 40352
rect 30350 40330 30374 40332
rect 30430 40330 30454 40332
rect 30510 40330 30534 40332
rect 30372 40278 30374 40330
rect 30436 40278 30448 40330
rect 30510 40278 30512 40330
rect 30350 40276 30374 40278
rect 30430 40276 30454 40278
rect 30510 40276 30534 40278
rect 30294 40256 30590 40276
rect 30654 39350 30682 41582
rect 31758 41322 31786 43312
rect 32954 42154 32982 43312
rect 32862 42126 32982 42154
rect 31746 41316 31798 41322
rect 31746 41258 31798 41264
rect 32758 41112 32810 41118
rect 32758 41054 32810 41060
rect 32770 40982 32798 41054
rect 31562 40976 31614 40982
rect 31562 40918 31614 40924
rect 32758 40976 32810 40982
rect 32758 40918 32810 40924
rect 31378 40024 31430 40030
rect 31378 39966 31430 39972
rect 30642 39344 30694 39350
rect 30642 39286 30694 39292
rect 30294 39244 30590 39264
rect 30350 39242 30374 39244
rect 30430 39242 30454 39244
rect 30510 39242 30534 39244
rect 30372 39190 30374 39242
rect 30436 39190 30448 39242
rect 30510 39190 30512 39242
rect 30350 39188 30374 39190
rect 30430 39188 30454 39190
rect 30510 39188 30534 39190
rect 30294 39168 30590 39188
rect 29354 38596 29406 38602
rect 29354 38538 29406 38544
rect 28250 38460 28302 38466
rect 28250 38402 28302 38408
rect 28894 37712 28946 37718
rect 28894 37654 28946 37660
rect 28906 37514 28934 37654
rect 28894 37508 28946 37514
rect 28894 37450 28946 37456
rect 28802 37372 28854 37378
rect 28802 37314 28854 37320
rect 28250 36964 28302 36970
rect 28250 36906 28302 36912
rect 28262 35678 28290 36906
rect 28814 36630 28842 37314
rect 28986 36760 29038 36766
rect 28986 36702 29038 36708
rect 28802 36624 28854 36630
rect 28802 36566 28854 36572
rect 28342 36216 28394 36222
rect 28342 36158 28394 36164
rect 28250 35672 28302 35678
rect 28250 35614 28302 35620
rect 28354 33706 28382 36158
rect 28814 35202 28842 36566
rect 28998 36086 29026 36702
rect 29366 36426 29394 38538
rect 29722 38392 29774 38398
rect 29722 38334 29774 38340
rect 29630 38256 29682 38262
rect 29630 38198 29682 38204
rect 29642 37990 29670 38198
rect 29630 37984 29682 37990
rect 29630 37926 29682 37932
rect 29642 37174 29670 37926
rect 29734 37854 29762 38334
rect 30294 38156 30590 38176
rect 30350 38154 30374 38156
rect 30430 38154 30454 38156
rect 30510 38154 30534 38156
rect 30372 38102 30374 38154
rect 30436 38102 30448 38154
rect 30510 38102 30512 38154
rect 30350 38100 30374 38102
rect 30430 38100 30454 38102
rect 30510 38100 30534 38102
rect 30294 38080 30590 38100
rect 29722 37848 29774 37854
rect 29722 37790 29774 37796
rect 29734 37718 29762 37790
rect 29722 37712 29774 37718
rect 29722 37654 29774 37660
rect 29630 37168 29682 37174
rect 29630 37110 29682 37116
rect 29734 36970 29762 37654
rect 29814 37304 29866 37310
rect 29814 37246 29866 37252
rect 29826 37174 29854 37246
rect 29814 37168 29866 37174
rect 29814 37110 29866 37116
rect 29722 36964 29774 36970
rect 29722 36906 29774 36912
rect 29354 36420 29406 36426
rect 29354 36362 29406 36368
rect 29078 36352 29130 36358
rect 29078 36294 29130 36300
rect 28986 36080 29038 36086
rect 28986 36022 29038 36028
rect 28998 35270 29026 36022
rect 29090 35542 29118 36294
rect 29262 36080 29314 36086
rect 29262 36022 29314 36028
rect 29078 35536 29130 35542
rect 29078 35478 29130 35484
rect 28986 35264 29038 35270
rect 28986 35206 29038 35212
rect 28802 35196 28854 35202
rect 28802 35138 28854 35144
rect 28894 34108 28946 34114
rect 28894 34050 28946 34056
rect 28342 33700 28394 33706
rect 28342 33642 28394 33648
rect 28906 33502 28934 34050
rect 29090 33978 29118 35478
rect 29274 35338 29302 36022
rect 29354 35672 29406 35678
rect 29354 35614 29406 35620
rect 29366 35542 29394 35614
rect 29354 35536 29406 35542
rect 29354 35478 29406 35484
rect 29262 35332 29314 35338
rect 29262 35274 29314 35280
rect 29826 34726 29854 37110
rect 30294 37068 30590 37088
rect 30350 37066 30374 37068
rect 30430 37066 30454 37068
rect 30510 37066 30534 37068
rect 30372 37014 30374 37066
rect 30436 37014 30448 37066
rect 30510 37014 30512 37066
rect 30350 37012 30374 37014
rect 30430 37012 30454 37014
rect 30510 37012 30534 37014
rect 30294 36992 30590 37012
rect 31390 36834 31418 39966
rect 31574 39962 31602 40918
rect 32298 40568 32350 40574
rect 32298 40510 32350 40516
rect 32114 40024 32166 40030
rect 32114 39966 32166 39972
rect 31562 39956 31614 39962
rect 31562 39898 31614 39904
rect 31574 39554 31602 39898
rect 31562 39548 31614 39554
rect 31562 39490 31614 39496
rect 32022 39548 32074 39554
rect 32022 39490 32074 39496
rect 31930 39480 31982 39486
rect 31930 39422 31982 39428
rect 31838 39344 31890 39350
rect 31838 39286 31890 39292
rect 31378 36828 31430 36834
rect 31378 36770 31430 36776
rect 29906 36420 29958 36426
rect 29906 36362 29958 36368
rect 29918 36154 29946 36362
rect 29906 36148 29958 36154
rect 29906 36090 29958 36096
rect 29918 34726 29946 36090
rect 30294 35980 30590 36000
rect 30350 35978 30374 35980
rect 30430 35978 30454 35980
rect 30510 35978 30534 35980
rect 30372 35926 30374 35978
rect 30436 35926 30448 35978
rect 30510 35926 30512 35978
rect 30350 35924 30374 35926
rect 30430 35924 30454 35926
rect 30510 35924 30534 35926
rect 30294 35904 30590 35924
rect 30458 35808 30510 35814
rect 30458 35750 30510 35756
rect 30274 35672 30326 35678
rect 30274 35614 30326 35620
rect 30090 35536 30142 35542
rect 30090 35478 30142 35484
rect 30102 35134 30130 35478
rect 30286 35202 30314 35614
rect 30470 35270 30498 35750
rect 30458 35264 30510 35270
rect 30458 35206 30510 35212
rect 30274 35196 30326 35202
rect 30194 35156 30274 35184
rect 30090 35128 30142 35134
rect 30090 35070 30142 35076
rect 29814 34720 29866 34726
rect 29814 34662 29866 34668
rect 29906 34720 29958 34726
rect 29906 34662 29958 34668
rect 29826 34590 29854 34662
rect 29814 34584 29866 34590
rect 29814 34526 29866 34532
rect 29826 34114 29854 34526
rect 29814 34108 29866 34114
rect 29814 34050 29866 34056
rect 29078 33972 29130 33978
rect 29078 33914 29130 33920
rect 29826 33858 29854 34050
rect 29734 33830 29854 33858
rect 29734 33706 29762 33830
rect 30194 33706 30222 35156
rect 30274 35138 30326 35144
rect 30734 35128 30786 35134
rect 30734 35070 30786 35076
rect 30642 34992 30694 34998
rect 30642 34934 30694 34940
rect 30294 34892 30590 34912
rect 30350 34890 30374 34892
rect 30430 34890 30454 34892
rect 30510 34890 30534 34892
rect 30372 34838 30374 34890
rect 30436 34838 30448 34890
rect 30510 34838 30512 34890
rect 30350 34836 30374 34838
rect 30430 34836 30454 34838
rect 30510 34836 30534 34838
rect 30294 34816 30590 34836
rect 30654 34794 30682 34934
rect 30642 34788 30694 34794
rect 30642 34730 30694 34736
rect 30294 33804 30590 33824
rect 30350 33802 30374 33804
rect 30430 33802 30454 33804
rect 30510 33802 30534 33804
rect 30372 33750 30374 33802
rect 30436 33750 30448 33802
rect 30510 33750 30512 33802
rect 30350 33748 30374 33750
rect 30430 33748 30454 33750
rect 30510 33748 30534 33750
rect 30294 33728 30590 33748
rect 29722 33700 29774 33706
rect 29722 33642 29774 33648
rect 30182 33700 30234 33706
rect 30182 33642 30234 33648
rect 30194 33502 30222 33642
rect 30746 33609 30774 35070
rect 31850 34454 31878 39286
rect 31942 37922 31970 39422
rect 32034 39146 32062 39490
rect 32022 39140 32074 39146
rect 32022 39082 32074 39088
rect 31930 37916 31982 37922
rect 31930 37858 31982 37864
rect 32126 37514 32154 39966
rect 32310 39622 32338 40510
rect 32770 40166 32798 40918
rect 32758 40160 32810 40166
rect 32758 40102 32810 40108
rect 32770 39622 32798 40102
rect 32298 39616 32350 39622
rect 32298 39558 32350 39564
rect 32758 39616 32810 39622
rect 32758 39558 32810 39564
rect 32758 38936 32810 38942
rect 32758 38878 32810 38884
rect 32666 38868 32718 38874
rect 32666 38810 32718 38816
rect 32298 37780 32350 37786
rect 32298 37722 32350 37728
rect 32114 37508 32166 37514
rect 32114 37450 32166 37456
rect 31930 37372 31982 37378
rect 31930 37314 31982 37320
rect 31942 36766 31970 37314
rect 32310 36834 32338 37722
rect 32678 37378 32706 38810
rect 32770 37446 32798 38878
rect 32758 37440 32810 37446
rect 32758 37382 32810 37388
rect 32666 37372 32718 37378
rect 32666 37314 32718 37320
rect 32770 37258 32798 37382
rect 32678 37242 32798 37258
rect 32666 37236 32798 37242
rect 32718 37230 32798 37236
rect 32666 37178 32718 37184
rect 32114 36828 32166 36834
rect 32114 36770 32166 36776
rect 32298 36828 32350 36834
rect 32298 36770 32350 36776
rect 31930 36760 31982 36766
rect 31930 36702 31982 36708
rect 32126 36630 32154 36770
rect 32482 36760 32534 36766
rect 32770 36748 32798 37230
rect 32534 36720 32798 36748
rect 32482 36702 32534 36708
rect 32206 36692 32258 36698
rect 32206 36634 32258 36640
rect 32022 36624 32074 36630
rect 32022 36566 32074 36572
rect 32114 36624 32166 36630
rect 32114 36566 32166 36572
rect 32034 36442 32062 36566
rect 32218 36442 32246 36634
rect 32758 36624 32810 36630
rect 32758 36566 32810 36572
rect 32034 36414 32246 36442
rect 32114 36284 32166 36290
rect 32114 36226 32166 36232
rect 32126 35678 32154 36226
rect 32770 35678 32798 36566
rect 32862 36222 32890 42126
rect 32958 41964 33254 41984
rect 33014 41962 33038 41964
rect 33094 41962 33118 41964
rect 33174 41962 33198 41964
rect 33036 41910 33038 41962
rect 33100 41910 33112 41962
rect 33174 41910 33176 41962
rect 33014 41908 33038 41910
rect 33094 41908 33118 41910
rect 33174 41908 33198 41910
rect 32958 41888 33254 41908
rect 32958 40876 33254 40896
rect 33014 40874 33038 40876
rect 33094 40874 33118 40876
rect 33174 40874 33198 40876
rect 33036 40822 33038 40874
rect 33100 40822 33112 40874
rect 33174 40822 33176 40874
rect 33014 40820 33038 40822
rect 33094 40820 33118 40822
rect 33174 40820 33198 40822
rect 32958 40800 33254 40820
rect 34150 40642 34178 43312
rect 34138 40636 34190 40642
rect 34138 40578 34190 40584
rect 34598 40568 34650 40574
rect 34598 40510 34650 40516
rect 34610 40098 34638 40510
rect 34690 40432 34742 40438
rect 34690 40374 34742 40380
rect 34598 40092 34650 40098
rect 34598 40034 34650 40040
rect 34230 39956 34282 39962
rect 34230 39898 34282 39904
rect 33310 39888 33362 39894
rect 33310 39830 33362 39836
rect 32958 39788 33254 39808
rect 33014 39786 33038 39788
rect 33094 39786 33118 39788
rect 33174 39786 33198 39788
rect 33036 39734 33038 39786
rect 33100 39734 33112 39786
rect 33174 39734 33176 39786
rect 33014 39732 33038 39734
rect 33094 39732 33118 39734
rect 33174 39732 33198 39734
rect 32958 39712 33254 39732
rect 33322 39486 33350 39830
rect 34046 39548 34098 39554
rect 34046 39490 34098 39496
rect 33310 39480 33362 39486
rect 33310 39422 33362 39428
rect 33402 38800 33454 38806
rect 33402 38742 33454 38748
rect 32958 38700 33254 38720
rect 33014 38698 33038 38700
rect 33094 38698 33118 38700
rect 33174 38698 33198 38700
rect 33036 38646 33038 38698
rect 33100 38646 33112 38698
rect 33174 38646 33176 38698
rect 33014 38644 33038 38646
rect 33094 38644 33118 38646
rect 33174 38644 33198 38646
rect 32958 38624 33254 38644
rect 33414 37854 33442 38742
rect 33586 38392 33638 38398
rect 33586 38334 33638 38340
rect 33598 38058 33626 38334
rect 33954 38256 34006 38262
rect 33954 38198 34006 38204
rect 33586 38052 33638 38058
rect 33586 37994 33638 38000
rect 33402 37848 33454 37854
rect 33402 37790 33454 37796
rect 33586 37848 33638 37854
rect 33586 37790 33638 37796
rect 33598 37718 33626 37790
rect 33586 37712 33638 37718
rect 33586 37654 33638 37660
rect 32958 37612 33254 37632
rect 33014 37610 33038 37612
rect 33094 37610 33118 37612
rect 33174 37610 33198 37612
rect 33036 37558 33038 37610
rect 33100 37558 33112 37610
rect 33174 37558 33176 37610
rect 33014 37556 33038 37558
rect 33094 37556 33118 37558
rect 33174 37556 33198 37558
rect 32958 37536 33254 37556
rect 33598 36766 33626 37654
rect 33494 36760 33546 36766
rect 33494 36702 33546 36708
rect 33586 36760 33638 36766
rect 33586 36702 33638 36708
rect 33506 36578 33534 36702
rect 33506 36550 33626 36578
rect 32958 36524 33254 36544
rect 33014 36522 33038 36524
rect 33094 36522 33118 36524
rect 33174 36522 33198 36524
rect 33036 36470 33038 36522
rect 33100 36470 33112 36522
rect 33174 36470 33176 36522
rect 33014 36468 33038 36470
rect 33094 36468 33118 36470
rect 33174 36468 33198 36470
rect 32958 36448 33254 36468
rect 33598 36290 33626 36550
rect 33586 36284 33638 36290
rect 33586 36226 33638 36232
rect 32850 36216 32902 36222
rect 32850 36158 32902 36164
rect 32862 35814 32890 36158
rect 33966 36086 33994 38198
rect 34058 37922 34086 39490
rect 34046 37916 34098 37922
rect 34046 37858 34098 37864
rect 33954 36080 34006 36086
rect 33954 36022 34006 36028
rect 34138 36080 34190 36086
rect 34138 36022 34190 36028
rect 32850 35808 32902 35814
rect 32850 35750 32902 35756
rect 34046 35808 34098 35814
rect 34046 35750 34098 35756
rect 32114 35672 32166 35678
rect 32114 35614 32166 35620
rect 32758 35672 32810 35678
rect 32758 35614 32810 35620
rect 32022 35604 32074 35610
rect 32022 35546 32074 35552
rect 32034 35202 32062 35546
rect 32022 35196 32074 35202
rect 32022 35138 32074 35144
rect 31838 34448 31890 34454
rect 31838 34390 31890 34396
rect 31470 33904 31522 33910
rect 31470 33846 31522 33852
rect 30364 33600 30420 33609
rect 30364 33535 30366 33544
rect 30418 33535 30420 33544
rect 30732 33600 30788 33609
rect 30732 33535 30788 33544
rect 30366 33506 30418 33512
rect 31482 33502 31510 33846
rect 31850 33502 31878 34390
rect 32126 33502 32154 35614
rect 33310 35604 33362 35610
rect 33310 35546 33362 35552
rect 32958 35436 33254 35456
rect 33014 35434 33038 35436
rect 33094 35434 33118 35436
rect 33174 35434 33198 35436
rect 33036 35382 33038 35434
rect 33100 35382 33112 35434
rect 33174 35382 33176 35434
rect 33014 35380 33038 35382
rect 33094 35380 33118 35382
rect 33174 35380 33198 35382
rect 32958 35360 33254 35380
rect 33126 35196 33178 35202
rect 33322 35184 33350 35546
rect 33402 35196 33454 35202
rect 33322 35156 33402 35184
rect 33126 35138 33178 35144
rect 33402 35138 33454 35144
rect 33138 34794 33166 35138
rect 33126 34788 33178 34794
rect 33126 34730 33178 34736
rect 33402 34788 33454 34794
rect 33402 34730 33454 34736
rect 32482 34448 32534 34454
rect 32482 34390 32534 34396
rect 32494 34114 32522 34390
rect 32958 34348 33254 34368
rect 33014 34346 33038 34348
rect 33094 34346 33118 34348
rect 33174 34346 33198 34348
rect 33036 34294 33038 34346
rect 33100 34294 33112 34346
rect 33174 34294 33176 34346
rect 33014 34292 33038 34294
rect 33094 34292 33118 34294
rect 33174 34292 33198 34294
rect 32958 34272 33254 34292
rect 32482 34108 32534 34114
rect 32482 34050 32534 34056
rect 28894 33496 28946 33502
rect 28894 33438 28946 33444
rect 30182 33496 30234 33502
rect 30182 33438 30234 33444
rect 31470 33496 31522 33502
rect 31470 33438 31522 33444
rect 31838 33496 31890 33502
rect 31838 33438 31890 33444
rect 32114 33496 32166 33502
rect 32114 33438 32166 33444
rect 32574 33496 32626 33502
rect 32574 33438 32626 33444
rect 28906 33162 28934 33438
rect 28802 33156 28854 33162
rect 28802 33098 28854 33104
rect 28894 33156 28946 33162
rect 28894 33098 28946 33104
rect 28814 32550 28842 33098
rect 29170 33020 29222 33026
rect 29170 32962 29222 32968
rect 28802 32544 28854 32550
rect 28802 32486 28854 32492
rect 28618 32068 28670 32074
rect 28618 32010 28670 32016
rect 28894 32068 28946 32074
rect 28894 32010 28946 32016
rect 28158 31932 28210 31938
rect 28158 31874 28210 31880
rect 27146 31864 27198 31870
rect 27146 31806 27198 31812
rect 28170 31734 28198 31874
rect 28526 31864 28578 31870
rect 28524 31832 28526 31841
rect 28578 31832 28580 31841
rect 28524 31767 28580 31776
rect 27698 31728 27750 31734
rect 27698 31670 27750 31676
rect 28158 31728 28210 31734
rect 28158 31670 28210 31676
rect 27710 31462 27738 31670
rect 26962 31456 27014 31462
rect 26962 31398 27014 31404
rect 27698 31456 27750 31462
rect 27698 31398 27750 31404
rect 28158 31456 28210 31462
rect 28434 31456 28486 31462
rect 28158 31398 28210 31404
rect 28432 31424 28434 31433
rect 28486 31424 28488 31433
rect 26778 31252 26830 31258
rect 26778 31194 26830 31200
rect 27630 31084 27926 31104
rect 27686 31082 27710 31084
rect 27766 31082 27790 31084
rect 27846 31082 27870 31084
rect 27708 31030 27710 31082
rect 27772 31030 27784 31082
rect 27846 31030 27848 31082
rect 27686 31028 27710 31030
rect 27766 31028 27790 31030
rect 27846 31028 27870 31030
rect 27630 31008 27926 31028
rect 27514 30776 27566 30782
rect 27514 30718 27566 30724
rect 27698 30776 27750 30782
rect 27698 30718 27750 30724
rect 27330 30708 27382 30714
rect 27330 30650 27382 30656
rect 27146 30436 27198 30442
rect 27146 30378 27198 30384
rect 27054 30232 27106 30238
rect 27054 30174 27106 30180
rect 27066 29694 27094 30174
rect 27054 29688 27106 29694
rect 27054 29630 27106 29636
rect 25858 29620 25910 29626
rect 25858 29562 25910 29568
rect 25490 28736 25542 28742
rect 24844 28704 24900 28713
rect 25766 28736 25818 28742
rect 25490 28678 25542 28684
rect 25764 28704 25766 28713
rect 26502 28736 26554 28742
rect 25818 28704 25820 28713
rect 24844 28639 24846 28648
rect 24898 28639 24900 28648
rect 24846 28610 24898 28616
rect 24858 28579 24886 28610
rect 25502 28470 25530 28678
rect 26502 28678 26554 28684
rect 25764 28639 25820 28648
rect 26514 28538 26542 28678
rect 27158 28674 27186 30378
rect 27342 30238 27370 30650
rect 27330 30232 27382 30238
rect 27330 30174 27382 30180
rect 27422 30164 27474 30170
rect 27422 30106 27474 30112
rect 27434 29937 27462 30106
rect 27420 29928 27476 29937
rect 27420 29863 27476 29872
rect 27526 29830 27554 30718
rect 27710 30374 27738 30718
rect 27974 30436 28026 30442
rect 27974 30378 28026 30384
rect 27698 30368 27750 30374
rect 27698 30310 27750 30316
rect 27630 29996 27926 30016
rect 27686 29994 27710 29996
rect 27766 29994 27790 29996
rect 27846 29994 27870 29996
rect 27708 29942 27710 29994
rect 27772 29942 27784 29994
rect 27846 29942 27848 29994
rect 27686 29940 27710 29942
rect 27766 29940 27790 29942
rect 27846 29940 27870 29942
rect 27630 29920 27926 29940
rect 27514 29824 27566 29830
rect 27514 29766 27566 29772
rect 27606 29824 27658 29830
rect 27606 29766 27658 29772
rect 27618 29694 27646 29766
rect 27986 29762 28014 30378
rect 28170 29762 28198 31398
rect 28432 31359 28488 31368
rect 28526 31388 28578 31394
rect 28526 31330 28578 31336
rect 28538 31297 28566 31330
rect 28524 31288 28580 31297
rect 28524 31223 28580 31232
rect 28342 30368 28394 30374
rect 28340 30336 28342 30345
rect 28394 30336 28396 30345
rect 28340 30271 28396 30280
rect 28630 29830 28658 32010
rect 28906 31938 28934 32010
rect 28710 31932 28762 31938
rect 28710 31874 28762 31880
rect 28894 31932 28946 31938
rect 28894 31874 28946 31880
rect 28722 31433 28750 31874
rect 29182 31870 29210 32962
rect 30294 32716 30590 32736
rect 30350 32714 30374 32716
rect 30430 32714 30454 32716
rect 30510 32714 30534 32716
rect 30372 32662 30374 32714
rect 30436 32662 30448 32714
rect 30510 32662 30512 32714
rect 30350 32660 30374 32662
rect 30430 32660 30454 32662
rect 30510 32660 30534 32662
rect 30294 32640 30590 32660
rect 30090 31932 30142 31938
rect 30090 31874 30142 31880
rect 29170 31864 29222 31870
rect 28984 31832 29040 31841
rect 29170 31806 29222 31812
rect 28984 31767 29040 31776
rect 28708 31424 28764 31433
rect 28998 31394 29026 31767
rect 28708 31359 28764 31368
rect 28986 31388 29038 31394
rect 28986 31330 29038 31336
rect 28802 31184 28854 31190
rect 28802 31126 28854 31132
rect 28814 30850 28842 31126
rect 28802 30844 28854 30850
rect 28802 30786 28854 30792
rect 28710 30640 28762 30646
rect 28710 30582 28762 30588
rect 28618 29824 28670 29830
rect 28618 29766 28670 29772
rect 28722 29762 28750 30582
rect 27974 29756 28026 29762
rect 27974 29698 28026 29704
rect 28158 29756 28210 29762
rect 28158 29698 28210 29704
rect 28710 29756 28762 29762
rect 28710 29698 28762 29704
rect 27606 29688 27658 29694
rect 27606 29630 27658 29636
rect 27986 29626 28014 29698
rect 27974 29620 28026 29626
rect 27974 29562 28026 29568
rect 28158 29620 28210 29626
rect 28158 29562 28210 29568
rect 28170 29286 28198 29562
rect 28158 29280 28210 29286
rect 28158 29222 28210 29228
rect 28710 29212 28762 29218
rect 28710 29154 28762 29160
rect 28526 29144 28578 29150
rect 28526 29086 28578 29092
rect 27630 28908 27926 28928
rect 27686 28906 27710 28908
rect 27766 28906 27790 28908
rect 27846 28906 27870 28908
rect 27708 28854 27710 28906
rect 27772 28854 27784 28906
rect 27846 28854 27848 28906
rect 27686 28852 27710 28854
rect 27766 28852 27790 28854
rect 27846 28852 27870 28854
rect 27630 28832 27926 28852
rect 28538 28810 28566 29086
rect 28526 28804 28578 28810
rect 28526 28746 28578 28752
rect 27422 28736 27474 28742
rect 28342 28736 28394 28742
rect 27474 28696 27922 28724
rect 27422 28678 27474 28684
rect 27146 28668 27198 28674
rect 27146 28610 27198 28616
rect 27894 28606 27922 28696
rect 27972 28704 28028 28713
rect 28342 28678 28394 28684
rect 27972 28639 28028 28648
rect 27698 28600 27750 28606
rect 27698 28542 27750 28548
rect 27882 28600 27934 28606
rect 27882 28542 27934 28548
rect 26502 28532 26554 28538
rect 26502 28474 26554 28480
rect 25398 28464 25450 28470
rect 25398 28406 25450 28412
rect 25490 28464 25542 28470
rect 25490 28406 25542 28412
rect 24966 28364 25262 28384
rect 25022 28362 25046 28364
rect 25102 28362 25126 28364
rect 25182 28362 25206 28364
rect 25044 28310 25046 28362
rect 25108 28310 25120 28362
rect 25182 28310 25184 28362
rect 25022 28308 25046 28310
rect 25102 28308 25126 28310
rect 25182 28308 25206 28310
rect 24966 28288 25262 28308
rect 24386 28124 24438 28130
rect 24386 28066 24438 28072
rect 24674 28118 24794 28146
rect 24398 28033 24426 28066
rect 24384 28024 24440 28033
rect 24110 27988 24162 27994
rect 24384 27959 24440 27968
rect 24110 27930 24162 27936
rect 24122 27738 24150 27930
rect 24122 27710 24242 27738
rect 24110 27580 24162 27586
rect 24110 27522 24162 27528
rect 24122 27042 24150 27522
rect 24214 27330 24242 27710
rect 24570 27716 24622 27722
rect 24570 27658 24622 27664
rect 24582 27602 24610 27658
rect 24674 27602 24702 28118
rect 24754 28056 24806 28062
rect 24754 27998 24806 28004
rect 24766 27722 24794 27998
rect 24754 27716 24806 27722
rect 24754 27658 24806 27664
rect 25214 27648 25266 27654
rect 24582 27574 24794 27602
rect 25214 27590 25266 27596
rect 24766 27518 24794 27574
rect 24754 27512 24806 27518
rect 25226 27489 25254 27590
rect 24754 27454 24806 27460
rect 25212 27480 25268 27489
rect 24846 27444 24898 27450
rect 25212 27415 25268 27424
rect 24846 27386 24898 27392
rect 24858 27330 24886 27386
rect 24214 27302 24886 27330
rect 24966 27276 25262 27296
rect 25022 27274 25046 27276
rect 25102 27274 25126 27276
rect 25182 27274 25206 27276
rect 25044 27222 25046 27274
rect 25108 27222 25120 27274
rect 25182 27222 25184 27274
rect 25022 27220 25046 27222
rect 25102 27220 25126 27222
rect 25182 27220 25206 27222
rect 24966 27200 25262 27220
rect 24662 27172 24714 27178
rect 24662 27114 24714 27120
rect 24478 27104 24530 27110
rect 24674 27058 24702 27114
rect 24530 27052 24702 27058
rect 24478 27046 24702 27052
rect 24110 27036 24162 27042
rect 24490 27030 24702 27046
rect 24110 26978 24162 26984
rect 24674 26974 24702 27030
rect 24018 26968 24070 26974
rect 24018 26910 24070 26916
rect 24662 26968 24714 26974
rect 24662 26910 24714 26916
rect 23926 26900 23978 26906
rect 23926 26842 23978 26848
rect 25410 26634 25438 28406
rect 27710 28198 27738 28542
rect 27986 28538 28014 28639
rect 27974 28532 28026 28538
rect 27974 28474 28026 28480
rect 28354 28470 28382 28678
rect 28722 28674 28750 29154
rect 28710 28668 28762 28674
rect 28710 28610 28762 28616
rect 28524 28568 28580 28577
rect 28524 28503 28580 28512
rect 28538 28470 28566 28503
rect 28342 28464 28394 28470
rect 28342 28406 28394 28412
rect 28526 28464 28578 28470
rect 28526 28406 28578 28412
rect 28354 28266 28382 28406
rect 28342 28260 28394 28266
rect 28342 28202 28394 28208
rect 27698 28192 27750 28198
rect 27698 28134 27750 28140
rect 25858 28056 25910 28062
rect 25858 27998 25910 28004
rect 25870 27926 25898 27998
rect 25858 27920 25910 27926
rect 25858 27862 25910 27868
rect 25870 27110 25898 27862
rect 27630 27820 27926 27840
rect 27686 27818 27710 27820
rect 27766 27818 27790 27820
rect 27846 27818 27870 27820
rect 27708 27766 27710 27818
rect 27772 27766 27784 27818
rect 27846 27766 27848 27818
rect 27686 27764 27710 27766
rect 27766 27764 27790 27766
rect 27846 27764 27870 27766
rect 27630 27744 27926 27764
rect 27066 27710 27462 27738
rect 27066 27518 27094 27710
rect 27146 27648 27198 27654
rect 27198 27608 27278 27636
rect 27146 27590 27198 27596
rect 27250 27518 27278 27608
rect 27434 27586 27462 27710
rect 28814 27586 28842 30786
rect 28894 30096 28946 30102
rect 28894 30038 28946 30044
rect 28906 29898 28934 30038
rect 28894 29892 28946 29898
rect 28894 29834 28946 29840
rect 28906 29286 28934 29834
rect 29078 29756 29130 29762
rect 29078 29698 29130 29704
rect 29090 29558 29118 29698
rect 29182 29694 29210 31806
rect 30102 31462 30130 31874
rect 30294 31628 30590 31648
rect 30350 31626 30374 31628
rect 30430 31626 30454 31628
rect 30510 31626 30534 31628
rect 30372 31574 30374 31626
rect 30436 31574 30448 31626
rect 30510 31574 30512 31626
rect 30350 31572 30374 31574
rect 30430 31572 30454 31574
rect 30510 31572 30534 31574
rect 30294 31552 30590 31572
rect 30090 31456 30142 31462
rect 30090 31398 30142 31404
rect 29262 31184 29314 31190
rect 29262 31126 29314 31132
rect 29274 30986 29302 31126
rect 29262 30980 29314 30986
rect 29262 30922 29314 30928
rect 29354 30980 29406 30986
rect 29354 30922 29406 30928
rect 29366 30374 29394 30922
rect 30102 30374 30130 31398
rect 31482 31326 31510 33438
rect 32586 33366 32614 33438
rect 31838 33360 31890 33366
rect 31838 33302 31890 33308
rect 32574 33360 32626 33366
rect 32574 33302 32626 33308
rect 31850 33026 31878 33302
rect 31838 33020 31890 33026
rect 31838 32962 31890 32968
rect 32586 32618 32614 33302
rect 32958 33260 33254 33280
rect 33014 33258 33038 33260
rect 33094 33258 33118 33260
rect 33174 33258 33198 33260
rect 33036 33206 33038 33258
rect 33100 33206 33112 33258
rect 33174 33206 33176 33258
rect 33014 33204 33038 33206
rect 33094 33204 33118 33206
rect 33174 33204 33198 33206
rect 32958 33184 33254 33204
rect 33414 33162 33442 34730
rect 34058 34114 34086 35750
rect 34150 34590 34178 36022
rect 34242 35202 34270 39898
rect 34506 39344 34558 39350
rect 34506 39286 34558 39292
rect 34518 39010 34546 39286
rect 34702 39146 34730 40374
rect 35438 39962 35466 43312
rect 35622 41420 35918 41440
rect 35678 41418 35702 41420
rect 35758 41418 35782 41420
rect 35838 41418 35862 41420
rect 35700 41366 35702 41418
rect 35764 41366 35776 41418
rect 35838 41366 35840 41418
rect 35678 41364 35702 41366
rect 35758 41364 35782 41366
rect 35838 41364 35862 41366
rect 35622 41344 35918 41364
rect 36346 41112 36398 41118
rect 36346 41054 36398 41060
rect 35622 40332 35918 40352
rect 35678 40330 35702 40332
rect 35758 40330 35782 40332
rect 35838 40330 35862 40332
rect 35700 40278 35702 40330
rect 35764 40278 35776 40330
rect 35838 40278 35840 40330
rect 35678 40276 35702 40278
rect 35758 40276 35782 40278
rect 35838 40276 35862 40278
rect 35622 40256 35918 40276
rect 35426 39956 35478 39962
rect 35426 39898 35478 39904
rect 36358 39554 36386 41054
rect 36634 40642 36662 43312
rect 37082 41180 37134 41186
rect 37082 41122 37134 41128
rect 36622 40636 36674 40642
rect 36622 40578 36674 40584
rect 37094 39894 37122 41122
rect 37542 40976 37594 40982
rect 37542 40918 37594 40924
rect 37554 40642 37582 40918
rect 37542 40636 37594 40642
rect 37542 40578 37594 40584
rect 37082 39888 37134 39894
rect 37082 39830 37134 39836
rect 34874 39548 34926 39554
rect 34874 39490 34926 39496
rect 36346 39548 36398 39554
rect 36346 39490 36398 39496
rect 34886 39350 34914 39490
rect 37830 39418 37858 43312
rect 38286 41964 38582 41984
rect 38342 41962 38366 41964
rect 38422 41962 38446 41964
rect 38502 41962 38526 41964
rect 38364 41910 38366 41962
rect 38428 41910 38440 41962
rect 38502 41910 38504 41962
rect 38342 41908 38366 41910
rect 38422 41908 38446 41910
rect 38502 41908 38526 41910
rect 38286 41888 38582 41908
rect 38286 40876 38582 40896
rect 38342 40874 38366 40876
rect 38422 40874 38446 40876
rect 38502 40874 38526 40876
rect 38364 40822 38366 40874
rect 38428 40822 38440 40874
rect 38502 40822 38504 40874
rect 38342 40820 38366 40822
rect 38422 40820 38446 40822
rect 38502 40820 38526 40822
rect 38286 40800 38582 40820
rect 39118 40642 39146 43312
rect 39106 40636 39158 40642
rect 39106 40578 39158 40584
rect 39658 40568 39710 40574
rect 39658 40510 39710 40516
rect 39934 40568 39986 40574
rect 39934 40510 39986 40516
rect 39670 40234 39698 40510
rect 39658 40228 39710 40234
rect 39658 40170 39710 40176
rect 38094 40092 38146 40098
rect 38094 40034 38146 40040
rect 38106 39894 38134 40034
rect 39198 40024 39250 40030
rect 39198 39966 39250 39972
rect 38094 39888 38146 39894
rect 38094 39830 38146 39836
rect 38106 39690 38134 39830
rect 38286 39788 38582 39808
rect 38342 39786 38366 39788
rect 38422 39786 38446 39788
rect 38502 39786 38526 39788
rect 38364 39734 38366 39786
rect 38428 39734 38440 39786
rect 38502 39734 38504 39786
rect 38342 39732 38366 39734
rect 38422 39732 38446 39734
rect 38502 39732 38526 39734
rect 38286 39712 38582 39732
rect 38094 39684 38146 39690
rect 38094 39626 38146 39632
rect 37818 39412 37870 39418
rect 37818 39354 37870 39360
rect 34874 39344 34926 39350
rect 34874 39286 34926 39292
rect 34690 39140 34742 39146
rect 34690 39082 34742 39088
rect 34506 39004 34558 39010
rect 34506 38946 34558 38952
rect 34702 38942 34730 39082
rect 34886 39078 34914 39286
rect 35622 39244 35918 39264
rect 35678 39242 35702 39244
rect 35758 39242 35782 39244
rect 35838 39242 35862 39244
rect 35700 39190 35702 39242
rect 35764 39190 35776 39242
rect 35838 39190 35840 39242
rect 35678 39188 35702 39190
rect 35758 39188 35782 39190
rect 35838 39188 35862 39190
rect 35622 39168 35918 39188
rect 34874 39072 34926 39078
rect 34874 39014 34926 39020
rect 34690 38936 34742 38942
rect 34690 38878 34742 38884
rect 34702 38602 34730 38878
rect 34690 38596 34742 38602
rect 34690 38538 34742 38544
rect 34886 38534 34914 39014
rect 38286 38700 38582 38720
rect 38342 38698 38366 38700
rect 38422 38698 38446 38700
rect 38502 38698 38526 38700
rect 38364 38646 38366 38698
rect 38428 38646 38440 38698
rect 38502 38646 38504 38698
rect 38342 38644 38366 38646
rect 38422 38644 38446 38646
rect 38502 38644 38526 38646
rect 38286 38624 38582 38644
rect 34874 38528 34926 38534
rect 34874 38470 34926 38476
rect 34874 38256 34926 38262
rect 34874 38198 34926 38204
rect 34886 37990 34914 38198
rect 35622 38156 35918 38176
rect 35678 38154 35702 38156
rect 35758 38154 35782 38156
rect 35838 38154 35862 38156
rect 35700 38102 35702 38154
rect 35764 38102 35776 38154
rect 35838 38102 35840 38154
rect 35678 38100 35702 38102
rect 35758 38100 35782 38102
rect 35838 38100 35862 38102
rect 35622 38080 35918 38100
rect 34874 37984 34926 37990
rect 34874 37926 34926 37932
rect 37738 37922 37858 37938
rect 34966 37916 35018 37922
rect 34966 37858 35018 37864
rect 36622 37916 36674 37922
rect 36622 37858 36674 37864
rect 37738 37916 37870 37922
rect 37738 37910 37818 37916
rect 34978 37718 35006 37858
rect 35150 37848 35202 37854
rect 35150 37790 35202 37796
rect 34966 37712 35018 37718
rect 34966 37654 35018 37660
rect 35058 37712 35110 37718
rect 35058 37654 35110 37660
rect 34978 37378 35006 37654
rect 35070 37514 35098 37654
rect 35162 37514 35190 37790
rect 35058 37508 35110 37514
rect 35058 37450 35110 37456
rect 35150 37508 35202 37514
rect 35150 37450 35202 37456
rect 34966 37372 35018 37378
rect 34966 37314 35018 37320
rect 34782 36624 34834 36630
rect 34782 36566 34834 36572
rect 34506 36148 34558 36154
rect 34506 36090 34558 36096
rect 34518 35814 34546 36090
rect 34794 35814 34822 36566
rect 35058 36216 35110 36222
rect 35058 36158 35110 36164
rect 34506 35808 34558 35814
rect 34506 35750 34558 35756
rect 34782 35808 34834 35814
rect 34782 35750 34834 35756
rect 34794 35678 34822 35750
rect 34782 35672 34834 35678
rect 34782 35614 34834 35620
rect 34230 35196 34282 35202
rect 34230 35138 34282 35144
rect 34598 35060 34650 35066
rect 34598 35002 34650 35008
rect 34610 34794 34638 35002
rect 34598 34788 34650 34794
rect 34598 34730 34650 34736
rect 34610 34590 34638 34730
rect 34138 34584 34190 34590
rect 34138 34526 34190 34532
rect 34598 34584 34650 34590
rect 34598 34526 34650 34532
rect 34046 34108 34098 34114
rect 34046 34050 34098 34056
rect 33954 33972 34006 33978
rect 33954 33914 34006 33920
rect 34414 33972 34466 33978
rect 34414 33914 34466 33920
rect 33966 33570 33994 33914
rect 33954 33564 34006 33570
rect 33954 33506 34006 33512
rect 33402 33156 33454 33162
rect 33402 33098 33454 33104
rect 34426 33026 34454 33914
rect 34414 33020 34466 33026
rect 34414 32962 34466 32968
rect 34794 32906 34822 35614
rect 35070 34590 35098 36158
rect 35058 34584 35110 34590
rect 35058 34526 35110 34532
rect 35058 33904 35110 33910
rect 35058 33846 35110 33852
rect 35070 33570 35098 33846
rect 35058 33564 35110 33570
rect 35058 33506 35110 33512
rect 34794 32878 35006 32906
rect 33034 32816 33086 32822
rect 33034 32758 33086 32764
rect 32574 32612 32626 32618
rect 32574 32554 32626 32560
rect 33046 32414 33074 32758
rect 34874 32544 34926 32550
rect 34874 32486 34926 32492
rect 33034 32408 33086 32414
rect 33034 32350 33086 32356
rect 34690 32408 34742 32414
rect 34690 32350 34742 32356
rect 34322 32272 34374 32278
rect 34322 32214 34374 32220
rect 32958 32172 33254 32192
rect 33014 32170 33038 32172
rect 33094 32170 33118 32172
rect 33174 32170 33198 32172
rect 33036 32118 33038 32170
rect 33100 32118 33112 32170
rect 33174 32118 33176 32170
rect 33014 32116 33038 32118
rect 33094 32116 33118 32118
rect 33174 32116 33198 32118
rect 32958 32096 33254 32116
rect 32482 31796 32534 31802
rect 32482 31738 32534 31744
rect 32574 31796 32626 31802
rect 32574 31738 32626 31744
rect 32494 31530 32522 31738
rect 32298 31524 32350 31530
rect 32298 31466 32350 31472
rect 32482 31524 32534 31530
rect 32482 31466 32534 31472
rect 32310 31326 32338 31466
rect 32586 31433 32614 31738
rect 32572 31424 32628 31433
rect 32572 31359 32628 31368
rect 33138 31348 33534 31376
rect 31470 31320 31522 31326
rect 31470 31262 31522 31268
rect 32206 31320 32258 31326
rect 32206 31262 32258 31268
rect 32298 31320 32350 31326
rect 32298 31262 32350 31268
rect 32666 31320 32718 31326
rect 32666 31262 32718 31268
rect 32218 31190 32246 31262
rect 32206 31184 32258 31190
rect 32206 31126 32258 31132
rect 30918 30912 30970 30918
rect 30918 30854 30970 30860
rect 30294 30540 30590 30560
rect 30350 30538 30374 30540
rect 30430 30538 30454 30540
rect 30510 30538 30534 30540
rect 30372 30486 30374 30538
rect 30436 30486 30448 30538
rect 30510 30486 30512 30538
rect 30350 30484 30374 30486
rect 30430 30484 30454 30486
rect 30510 30484 30534 30486
rect 30294 30464 30590 30484
rect 29354 30368 29406 30374
rect 29354 30310 29406 30316
rect 30090 30368 30142 30374
rect 30090 30310 30142 30316
rect 30102 29830 30130 30310
rect 30090 29824 30142 29830
rect 30090 29766 30142 29772
rect 30826 29824 30878 29830
rect 30826 29766 30878 29772
rect 29170 29688 29222 29694
rect 29170 29630 29222 29636
rect 30090 29688 30142 29694
rect 30090 29630 30142 29636
rect 28986 29552 29038 29558
rect 28986 29494 29038 29500
rect 29078 29552 29130 29558
rect 29078 29494 29130 29500
rect 28998 29286 29026 29494
rect 28894 29280 28946 29286
rect 28894 29222 28946 29228
rect 28986 29280 29038 29286
rect 28986 29222 29038 29228
rect 29090 29150 29118 29494
rect 29538 29212 29590 29218
rect 29538 29154 29590 29160
rect 29078 29144 29130 29150
rect 29078 29086 29130 29092
rect 29550 28606 29578 29154
rect 29998 29144 30050 29150
rect 29998 29086 30050 29092
rect 29814 28668 29866 28674
rect 29814 28610 29866 28616
rect 29538 28600 29590 28606
rect 29538 28542 29590 28548
rect 29722 28600 29774 28606
rect 29722 28542 29774 28548
rect 29550 28062 29578 28542
rect 29734 28470 29762 28542
rect 29722 28464 29774 28470
rect 29722 28406 29774 28412
rect 29734 28062 29762 28406
rect 29446 28056 29498 28062
rect 29446 27998 29498 28004
rect 29538 28056 29590 28062
rect 29538 27998 29590 28004
rect 29722 28056 29774 28062
rect 29722 27998 29774 28004
rect 27422 27580 27474 27586
rect 27422 27522 27474 27528
rect 28802 27580 28854 27586
rect 28802 27522 28854 27528
rect 27054 27512 27106 27518
rect 27054 27454 27106 27460
rect 27238 27512 27290 27518
rect 27238 27454 27290 27460
rect 26962 27444 27014 27450
rect 26962 27386 27014 27392
rect 28618 27444 28670 27450
rect 28618 27386 28670 27392
rect 26974 27110 27002 27386
rect 28630 27110 28658 27386
rect 25858 27104 25910 27110
rect 25858 27046 25910 27052
rect 26962 27104 27014 27110
rect 27974 27104 28026 27110
rect 26962 27046 27014 27052
rect 27618 27052 27974 27058
rect 27618 27046 28026 27052
rect 28618 27104 28670 27110
rect 28618 27046 28670 27052
rect 25870 26974 25898 27046
rect 27618 27030 28014 27046
rect 29458 27042 29486 27998
rect 29826 27722 29854 28610
rect 30010 28062 30038 29086
rect 30102 28674 30130 29630
rect 30294 29452 30590 29472
rect 30350 29450 30374 29452
rect 30430 29450 30454 29452
rect 30510 29450 30534 29452
rect 30372 29398 30374 29450
rect 30436 29398 30448 29450
rect 30510 29398 30512 29450
rect 30350 29396 30374 29398
rect 30430 29396 30454 29398
rect 30510 29396 30534 29398
rect 30294 29376 30590 29396
rect 30182 29212 30234 29218
rect 30182 29154 30234 29160
rect 30090 28668 30142 28674
rect 30090 28610 30142 28616
rect 30194 28062 30222 29154
rect 30838 29150 30866 29766
rect 30458 29144 30510 29150
rect 30458 29086 30510 29092
rect 30826 29144 30878 29150
rect 30826 29086 30878 29092
rect 30274 29008 30326 29014
rect 30274 28950 30326 28956
rect 30366 29008 30418 29014
rect 30366 28950 30418 28956
rect 30286 28606 30314 28950
rect 30378 28810 30406 28950
rect 30470 28810 30498 29086
rect 30366 28804 30418 28810
rect 30366 28746 30418 28752
rect 30458 28804 30510 28810
rect 30458 28746 30510 28752
rect 30274 28600 30326 28606
rect 30274 28542 30326 28548
rect 30826 28464 30878 28470
rect 30826 28406 30878 28412
rect 30294 28364 30590 28384
rect 30350 28362 30374 28364
rect 30430 28362 30454 28364
rect 30510 28362 30534 28364
rect 30372 28310 30374 28362
rect 30436 28310 30448 28362
rect 30510 28310 30512 28362
rect 30350 28308 30374 28310
rect 30430 28308 30454 28310
rect 30510 28308 30534 28310
rect 30294 28288 30590 28308
rect 30734 28192 30786 28198
rect 30734 28134 30786 28140
rect 30642 28124 30694 28130
rect 30642 28066 30694 28072
rect 29906 28056 29958 28062
rect 29906 27998 29958 28004
rect 29998 28056 30050 28062
rect 29998 27998 30050 28004
rect 30182 28056 30234 28062
rect 30182 27998 30234 28004
rect 30364 28024 30420 28033
rect 29918 27761 29946 27998
rect 30364 27959 30420 27968
rect 29904 27752 29960 27761
rect 29814 27716 29866 27722
rect 29904 27687 29960 27696
rect 29814 27658 29866 27664
rect 30378 27654 30406 27959
rect 30654 27722 30682 28066
rect 30642 27716 30694 27722
rect 30642 27658 30694 27664
rect 30366 27648 30418 27654
rect 29812 27616 29868 27625
rect 29722 27580 29774 27586
rect 30366 27590 30418 27596
rect 29812 27551 29868 27560
rect 29722 27522 29774 27528
rect 29734 27081 29762 27522
rect 29720 27072 29776 27081
rect 29446 27036 29498 27042
rect 27618 26974 27646 27030
rect 29720 27007 29776 27016
rect 29446 26978 29498 26984
rect 29826 26974 29854 27551
rect 30180 27480 30236 27489
rect 30180 27415 30236 27424
rect 30194 27092 30222 27415
rect 30294 27276 30590 27296
rect 30350 27274 30374 27276
rect 30430 27274 30454 27276
rect 30510 27274 30534 27276
rect 30372 27222 30374 27274
rect 30436 27222 30448 27274
rect 30510 27222 30512 27274
rect 30350 27220 30374 27222
rect 30430 27220 30454 27222
rect 30510 27220 30534 27222
rect 30294 27200 30590 27220
rect 30746 27178 30774 28134
rect 30838 28062 30866 28406
rect 30826 28056 30878 28062
rect 30826 27998 30878 28004
rect 30734 27172 30786 27178
rect 30734 27114 30786 27120
rect 30826 27104 30878 27110
rect 30194 27064 30314 27092
rect 30286 26974 30314 27064
rect 30826 27046 30878 27052
rect 25858 26968 25910 26974
rect 25858 26910 25910 26916
rect 27606 26968 27658 26974
rect 29814 26968 29866 26974
rect 27606 26910 27658 26916
rect 29352 26936 29408 26945
rect 29814 26910 29866 26916
rect 30274 26968 30326 26974
rect 30734 26968 30786 26974
rect 30274 26910 30326 26916
rect 30364 26936 30420 26945
rect 29352 26871 29354 26880
rect 29406 26871 29408 26880
rect 30364 26871 30420 26880
rect 30732 26936 30734 26945
rect 30786 26936 30788 26945
rect 30732 26871 30788 26880
rect 29354 26842 29406 26848
rect 27630 26732 27926 26752
rect 27686 26730 27710 26732
rect 27766 26730 27790 26732
rect 27846 26730 27870 26732
rect 27708 26678 27710 26730
rect 27772 26678 27784 26730
rect 27846 26678 27848 26730
rect 27686 26676 27710 26678
rect 27766 26676 27790 26678
rect 27846 26676 27870 26678
rect 27630 26656 27926 26676
rect 25398 26628 25450 26634
rect 25398 26570 25450 26576
rect 23834 25200 23886 25206
rect 23834 25142 23886 25148
rect 25410 24730 25438 26570
rect 16750 24724 16802 24730
rect 16750 24666 16802 24672
rect 25398 24724 25450 24730
rect 25398 24666 25450 24672
rect 15278 24384 15330 24390
rect 15278 24326 15330 24332
rect 30274 24112 30326 24118
rect 30274 24054 30326 24060
rect 30286 20378 30314 24054
rect 30378 22690 30406 26871
rect 30366 22684 30418 22690
rect 30366 22626 30418 22632
rect 30274 20372 30326 20378
rect 30274 20314 30326 20320
rect 30838 19834 30866 27046
rect 30930 22622 30958 30854
rect 32310 29286 32338 31262
rect 32678 31190 32706 31262
rect 33138 31258 33166 31348
rect 33126 31252 33178 31258
rect 33126 31194 33178 31200
rect 33310 31252 33362 31258
rect 33310 31194 33362 31200
rect 32666 31184 32718 31190
rect 32666 31126 32718 31132
rect 32958 31084 33254 31104
rect 33014 31082 33038 31084
rect 33094 31082 33118 31084
rect 33174 31082 33198 31084
rect 33036 31030 33038 31082
rect 33100 31030 33112 31082
rect 33174 31030 33176 31082
rect 33014 31028 33038 31030
rect 33094 31028 33118 31030
rect 33174 31028 33198 31030
rect 32958 31008 33254 31028
rect 33322 30850 33350 31194
rect 33506 31190 33534 31348
rect 33494 31184 33546 31190
rect 33494 31126 33546 31132
rect 33310 30844 33362 30850
rect 33310 30786 33362 30792
rect 34230 30708 34282 30714
rect 34230 30650 34282 30656
rect 34046 30640 34098 30646
rect 34046 30582 34098 30588
rect 34058 30306 34086 30582
rect 34046 30300 34098 30306
rect 34046 30242 34098 30248
rect 34242 30238 34270 30650
rect 34230 30232 34282 30238
rect 34230 30174 34282 30180
rect 32958 29996 33254 30016
rect 33014 29994 33038 29996
rect 33094 29994 33118 29996
rect 33174 29994 33198 29996
rect 33036 29942 33038 29994
rect 33100 29942 33112 29994
rect 33174 29942 33176 29994
rect 33014 29940 33038 29942
rect 33094 29940 33118 29942
rect 33174 29940 33198 29942
rect 32958 29920 33254 29940
rect 34230 29892 34282 29898
rect 34230 29834 34282 29840
rect 32298 29280 32350 29286
rect 32298 29222 32350 29228
rect 34138 29280 34190 29286
rect 34138 29222 34190 29228
rect 32022 29212 32074 29218
rect 32022 29154 32074 29160
rect 31286 29144 31338 29150
rect 31206 29104 31286 29132
rect 31206 29098 31234 29104
rect 31022 29070 31234 29098
rect 31286 29086 31338 29092
rect 31022 28470 31050 29070
rect 32034 28674 32062 29154
rect 33954 29144 34006 29150
rect 33216 29112 33272 29121
rect 33954 29086 34006 29092
rect 33216 29047 33218 29056
rect 33270 29047 33272 29056
rect 33218 29018 33270 29024
rect 32958 28908 33254 28928
rect 33014 28906 33038 28908
rect 33094 28906 33118 28908
rect 33174 28906 33198 28908
rect 33036 28854 33038 28906
rect 33100 28854 33112 28906
rect 33174 28854 33176 28906
rect 33014 28852 33038 28854
rect 33094 28852 33118 28854
rect 33174 28852 33198 28854
rect 32958 28832 33254 28852
rect 31562 28668 31614 28674
rect 31562 28610 31614 28616
rect 32022 28668 32074 28674
rect 32022 28610 32074 28616
rect 31102 28532 31154 28538
rect 31154 28492 31234 28520
rect 31102 28474 31154 28480
rect 31010 28464 31062 28470
rect 31010 28406 31062 28412
rect 31102 28056 31154 28062
rect 31022 28016 31102 28044
rect 31022 27518 31050 28016
rect 31102 27998 31154 28004
rect 31206 27994 31234 28492
rect 31378 28056 31430 28062
rect 31376 28024 31378 28033
rect 31430 28024 31432 28033
rect 31194 27988 31246 27994
rect 31376 27959 31432 27968
rect 31194 27930 31246 27936
rect 31286 27920 31338 27926
rect 31284 27888 31286 27897
rect 31378 27920 31430 27926
rect 31338 27888 31340 27897
rect 31378 27862 31430 27868
rect 31284 27823 31340 27832
rect 31192 27616 31248 27625
rect 31192 27551 31248 27560
rect 31010 27512 31062 27518
rect 31010 27454 31062 27460
rect 31206 26974 31234 27551
rect 31286 27512 31338 27518
rect 31286 27454 31338 27460
rect 31298 27042 31326 27454
rect 31390 27450 31418 27862
rect 31468 27752 31524 27761
rect 31468 27687 31524 27696
rect 31378 27444 31430 27450
rect 31378 27386 31430 27392
rect 31482 27110 31510 27687
rect 31574 27654 31602 28610
rect 33966 28606 33994 29086
rect 34046 29008 34098 29014
rect 34046 28950 34098 28956
rect 34058 28810 34086 28950
rect 34046 28804 34098 28810
rect 34046 28746 34098 28752
rect 33954 28600 34006 28606
rect 33954 28542 34006 28548
rect 34046 28124 34098 28130
rect 34046 28066 34098 28072
rect 33954 28056 34006 28062
rect 33954 27998 34006 28004
rect 32958 27820 33254 27840
rect 33014 27818 33038 27820
rect 33094 27818 33118 27820
rect 33174 27818 33198 27820
rect 33036 27766 33038 27818
rect 33100 27766 33112 27818
rect 33174 27766 33176 27818
rect 33014 27764 33038 27766
rect 33094 27764 33118 27766
rect 33174 27764 33198 27766
rect 32958 27744 33254 27764
rect 31562 27648 31614 27654
rect 31562 27590 31614 27596
rect 33770 27648 33822 27654
rect 33770 27590 33822 27596
rect 31838 27580 31890 27586
rect 31838 27522 31890 27528
rect 33126 27580 33178 27586
rect 33126 27522 33178 27528
rect 31744 27480 31800 27489
rect 31744 27415 31800 27424
rect 31758 27382 31786 27415
rect 31746 27376 31798 27382
rect 31746 27318 31798 27324
rect 31470 27104 31522 27110
rect 31654 27104 31706 27110
rect 31470 27046 31522 27052
rect 31652 27072 31654 27081
rect 31706 27072 31708 27081
rect 31286 27036 31338 27042
rect 31652 27007 31708 27016
rect 31286 26978 31338 26984
rect 31194 26968 31246 26974
rect 31194 26910 31246 26916
rect 31376 26936 31432 26945
rect 31376 26871 31432 26880
rect 31390 26566 31418 26871
rect 31378 26560 31430 26566
rect 31378 26502 31430 26508
rect 31850 25954 31878 27522
rect 33138 27382 33166 27522
rect 33126 27376 33178 27382
rect 33126 27318 33178 27324
rect 33138 27110 33166 27318
rect 33782 27178 33810 27590
rect 33966 27178 33994 27998
rect 33770 27172 33822 27178
rect 33770 27114 33822 27120
rect 33954 27172 34006 27178
rect 33954 27114 34006 27120
rect 33126 27104 33178 27110
rect 33126 27046 33178 27052
rect 32958 26732 33254 26752
rect 33014 26730 33038 26732
rect 33094 26730 33118 26732
rect 33174 26730 33198 26732
rect 33036 26678 33038 26730
rect 33100 26678 33112 26730
rect 33174 26678 33176 26730
rect 33014 26676 33038 26678
rect 33094 26676 33118 26678
rect 33174 26676 33198 26678
rect 32958 26656 33254 26676
rect 33966 26430 33994 27114
rect 33954 26424 34006 26430
rect 33954 26366 34006 26372
rect 31838 25948 31890 25954
rect 31838 25890 31890 25896
rect 34058 23914 34086 28066
rect 34150 27178 34178 29222
rect 34242 28062 34270 29834
rect 34230 28056 34282 28062
rect 34230 27998 34282 28004
rect 34138 27172 34190 27178
rect 34138 27114 34190 27120
rect 34150 26498 34178 27114
rect 34138 26492 34190 26498
rect 34138 26434 34190 26440
rect 33954 23908 34006 23914
rect 33954 23850 34006 23856
rect 34046 23908 34098 23914
rect 34046 23850 34098 23856
rect 31378 23772 31430 23778
rect 31378 23714 31430 23720
rect 31390 23069 31418 23714
rect 31376 23060 31432 23069
rect 31376 22995 31432 23004
rect 30918 22616 30970 22622
rect 30918 22558 30970 22564
rect 33966 21369 33994 23850
rect 33952 21360 34008 21369
rect 33952 21295 34008 21304
rect 34150 21194 34178 26434
rect 34334 23545 34362 32214
rect 34414 31184 34466 31190
rect 34414 31126 34466 31132
rect 34426 30102 34454 31126
rect 34506 30776 34558 30782
rect 34506 30718 34558 30724
rect 34414 30096 34466 30102
rect 34414 30038 34466 30044
rect 34426 29830 34454 30038
rect 34414 29824 34466 29830
rect 34414 29766 34466 29772
rect 34518 29694 34546 30718
rect 34702 30714 34730 32350
rect 34690 30708 34742 30714
rect 34690 30650 34742 30656
rect 34506 29688 34558 29694
rect 34506 29630 34558 29636
rect 34506 28804 34558 28810
rect 34506 28746 34558 28752
rect 34414 28600 34466 28606
rect 34414 28542 34466 28548
rect 34426 27382 34454 28542
rect 34518 28146 34546 28746
rect 34518 28130 34638 28146
rect 34518 28124 34650 28130
rect 34518 28118 34598 28124
rect 34598 28066 34650 28072
rect 34414 27376 34466 27382
rect 34414 27318 34466 27324
rect 34426 26838 34454 27318
rect 34414 26832 34466 26838
rect 34414 26774 34466 26780
rect 34426 25886 34454 26774
rect 34690 26288 34742 26294
rect 34690 26230 34742 26236
rect 34702 25954 34730 26230
rect 34690 25948 34742 25954
rect 34690 25890 34742 25896
rect 34414 25880 34466 25886
rect 34414 25822 34466 25828
rect 34426 25478 34454 25822
rect 34414 25472 34466 25478
rect 34414 25414 34466 25420
rect 34886 24934 34914 32486
rect 34978 30730 35006 32878
rect 35070 32550 35098 33506
rect 35162 32618 35190 37450
rect 36634 37446 36662 37858
rect 37634 37780 37686 37786
rect 37634 37722 37686 37728
rect 36622 37440 36674 37446
rect 36622 37382 36674 37388
rect 35622 37068 35918 37088
rect 35678 37066 35702 37068
rect 35758 37066 35782 37068
rect 35838 37066 35862 37068
rect 35700 37014 35702 37066
rect 35764 37014 35776 37066
rect 35838 37014 35840 37066
rect 35678 37012 35702 37014
rect 35758 37012 35782 37014
rect 35838 37012 35862 37014
rect 35622 36992 35918 37012
rect 37540 36864 37596 36873
rect 37540 36799 37596 36808
rect 37554 36766 37582 36799
rect 37542 36760 37594 36766
rect 37542 36702 37594 36708
rect 37450 36692 37502 36698
rect 37450 36634 37502 36640
rect 37462 36193 37490 36634
rect 37448 36184 37504 36193
rect 37646 36154 37674 37722
rect 37738 37514 37766 37910
rect 37818 37858 37870 37864
rect 37818 37780 37870 37786
rect 37818 37722 37870 37728
rect 37726 37508 37778 37514
rect 37726 37450 37778 37456
rect 37724 36728 37780 36737
rect 37724 36663 37780 36672
rect 37738 36630 37766 36663
rect 37726 36624 37778 36630
rect 37726 36566 37778 36572
rect 37448 36119 37504 36128
rect 37634 36148 37686 36154
rect 37634 36090 37686 36096
rect 35622 35980 35918 36000
rect 35678 35978 35702 35980
rect 35758 35978 35782 35980
rect 35838 35978 35862 35980
rect 35700 35926 35702 35978
rect 35764 35926 35776 35978
rect 35838 35926 35840 35978
rect 35678 35924 35702 35926
rect 35758 35924 35782 35926
rect 35838 35924 35862 35926
rect 35622 35904 35918 35924
rect 37174 35672 37226 35678
rect 37174 35614 37226 35620
rect 35518 35604 35570 35610
rect 35518 35546 35570 35552
rect 35530 35338 35558 35546
rect 37186 35542 37214 35614
rect 36070 35536 36122 35542
rect 36070 35478 36122 35484
rect 37174 35536 37226 35542
rect 37174 35478 37226 35484
rect 35518 35332 35570 35338
rect 35518 35274 35570 35280
rect 36082 35202 36110 35478
rect 36070 35196 36122 35202
rect 36070 35138 36122 35144
rect 35622 34892 35918 34912
rect 35678 34890 35702 34892
rect 35758 34890 35782 34892
rect 35838 34890 35862 34892
rect 35700 34838 35702 34890
rect 35764 34838 35776 34890
rect 35838 34838 35840 34890
rect 35678 34836 35702 34838
rect 35758 34836 35782 34838
rect 35838 34836 35862 34838
rect 35622 34816 35918 34836
rect 35518 34788 35570 34794
rect 35518 34730 35570 34736
rect 35530 34114 35558 34730
rect 35518 34108 35570 34114
rect 35518 34050 35570 34056
rect 35240 33600 35296 33609
rect 35240 33535 35242 33544
rect 35294 33535 35296 33544
rect 35242 33506 35294 33512
rect 35530 33502 35558 34050
rect 35622 33804 35918 33824
rect 35678 33802 35702 33804
rect 35758 33802 35782 33804
rect 35838 33802 35862 33804
rect 35700 33750 35702 33802
rect 35764 33750 35776 33802
rect 35838 33750 35840 33802
rect 35678 33748 35702 33750
rect 35758 33748 35782 33750
rect 35838 33748 35862 33750
rect 35622 33728 35918 33748
rect 35426 33496 35478 33502
rect 35426 33438 35478 33444
rect 35518 33496 35570 33502
rect 35518 33438 35570 33444
rect 35438 33162 35466 33438
rect 35426 33156 35478 33162
rect 35426 33098 35478 33104
rect 35622 32716 35918 32736
rect 35678 32714 35702 32716
rect 35758 32714 35782 32716
rect 35838 32714 35862 32716
rect 35700 32662 35702 32714
rect 35764 32662 35776 32714
rect 35838 32662 35840 32714
rect 35678 32660 35702 32662
rect 35758 32660 35782 32662
rect 35838 32660 35862 32662
rect 35622 32640 35918 32660
rect 35150 32612 35202 32618
rect 35150 32554 35202 32560
rect 35058 32544 35110 32550
rect 35058 32486 35110 32492
rect 35162 32414 35190 32554
rect 35150 32408 35202 32414
rect 35150 32350 35202 32356
rect 36082 32074 36110 35138
rect 37186 35066 37214 35478
rect 37830 35202 37858 37722
rect 38286 37612 38582 37632
rect 38342 37610 38366 37612
rect 38422 37610 38446 37612
rect 38502 37610 38526 37612
rect 38364 37558 38366 37610
rect 38428 37558 38440 37610
rect 38502 37558 38504 37610
rect 38342 37556 38366 37558
rect 38422 37556 38446 37558
rect 38502 37556 38526 37558
rect 38286 37536 38582 37556
rect 38002 37440 38054 37446
rect 38002 37382 38054 37388
rect 37910 37372 37962 37378
rect 37910 37314 37962 37320
rect 37922 36630 37950 37314
rect 38014 37242 38042 37382
rect 39104 37272 39160 37281
rect 38002 37236 38054 37242
rect 38002 37178 38054 37184
rect 38094 37236 38146 37242
rect 39104 37207 39160 37216
rect 38094 37178 38146 37184
rect 37910 36624 37962 36630
rect 37910 36566 37962 36572
rect 38106 35746 38134 37178
rect 39118 37174 39146 37207
rect 39106 37168 39158 37174
rect 39106 37110 39158 37116
rect 38286 36524 38582 36544
rect 38342 36522 38366 36524
rect 38422 36522 38446 36524
rect 38502 36522 38526 36524
rect 38364 36470 38366 36522
rect 38428 36470 38440 36522
rect 38502 36470 38504 36522
rect 38342 36468 38366 36470
rect 38422 36468 38446 36470
rect 38502 36468 38526 36470
rect 38286 36448 38582 36468
rect 39210 36358 39238 39966
rect 39474 39684 39526 39690
rect 39474 39626 39526 39632
rect 39486 39078 39514 39626
rect 39474 39072 39526 39078
rect 39474 39014 39526 39020
rect 39486 38466 39514 39014
rect 39474 38460 39526 38466
rect 39474 38402 39526 38408
rect 39946 38330 39974 40510
rect 40314 39962 40342 43312
rect 40950 41420 41246 41440
rect 41006 41418 41030 41420
rect 41086 41418 41110 41420
rect 41166 41418 41190 41420
rect 41028 41366 41030 41418
rect 41092 41366 41104 41418
rect 41166 41366 41168 41418
rect 41006 41364 41030 41366
rect 41086 41364 41110 41366
rect 41166 41364 41190 41366
rect 40950 41344 41246 41364
rect 40854 41112 40906 41118
rect 40854 41054 40906 41060
rect 40302 39956 40354 39962
rect 40302 39898 40354 39904
rect 40394 39548 40446 39554
rect 40394 39490 40446 39496
rect 40026 38460 40078 38466
rect 40026 38402 40078 38408
rect 39934 38324 39986 38330
rect 39934 38266 39986 38272
rect 40038 38058 40066 38402
rect 40302 38392 40354 38398
rect 40302 38334 40354 38340
rect 40026 38052 40078 38058
rect 40026 37994 40078 38000
rect 39566 37712 39618 37718
rect 39288 37680 39344 37689
rect 39566 37654 39618 37660
rect 39842 37712 39894 37718
rect 39842 37654 39894 37660
rect 39288 37615 39344 37624
rect 39302 37378 39330 37615
rect 39290 37372 39342 37378
rect 39290 37314 39342 37320
rect 39302 37174 39330 37314
rect 39474 37236 39526 37242
rect 39474 37178 39526 37184
rect 39290 37168 39342 37174
rect 39290 37110 39342 37116
rect 39302 36902 39330 37110
rect 39290 36896 39342 36902
rect 39290 36838 39342 36844
rect 39198 36352 39250 36358
rect 39198 36294 39250 36300
rect 38186 36216 38238 36222
rect 38186 36158 38238 36164
rect 38094 35740 38146 35746
rect 38094 35682 38146 35688
rect 37818 35196 37870 35202
rect 37818 35138 37870 35144
rect 37174 35060 37226 35066
rect 37174 35002 37226 35008
rect 38198 34454 38226 36158
rect 38286 35436 38582 35456
rect 38342 35434 38366 35436
rect 38422 35434 38446 35436
rect 38502 35434 38526 35436
rect 38364 35382 38366 35434
rect 38428 35382 38440 35434
rect 38502 35382 38504 35434
rect 38342 35380 38366 35382
rect 38422 35380 38446 35382
rect 38502 35380 38526 35382
rect 38286 35360 38582 35380
rect 39486 34998 39514 37178
rect 39578 35814 39606 37654
rect 39750 37372 39802 37378
rect 39750 37314 39802 37320
rect 39658 36216 39710 36222
rect 39658 36158 39710 36164
rect 39566 35808 39618 35814
rect 39566 35750 39618 35756
rect 39474 34992 39526 34998
rect 39474 34934 39526 34940
rect 39382 34720 39434 34726
rect 39380 34688 39382 34697
rect 39434 34688 39436 34697
rect 39380 34623 39436 34632
rect 38186 34448 38238 34454
rect 38186 34390 38238 34396
rect 38286 34348 38582 34368
rect 38342 34346 38366 34348
rect 38422 34346 38446 34348
rect 38502 34346 38526 34348
rect 38364 34294 38366 34346
rect 38428 34294 38440 34346
rect 38502 34294 38504 34346
rect 38342 34292 38366 34294
rect 38422 34292 38446 34294
rect 38502 34292 38526 34294
rect 38286 34272 38582 34292
rect 39670 33706 39698 36158
rect 39762 35082 39790 37314
rect 39854 37174 39882 37654
rect 40314 37446 40342 38334
rect 40406 37854 40434 39490
rect 40866 39010 40894 41054
rect 41510 40642 41538 43312
rect 41498 40636 41550 40642
rect 41498 40578 41550 40584
rect 41590 40568 41642 40574
rect 41590 40510 41642 40516
rect 41406 40500 41458 40506
rect 41406 40442 41458 40448
rect 40950 40332 41246 40352
rect 41006 40330 41030 40332
rect 41086 40330 41110 40332
rect 41166 40330 41190 40332
rect 41028 40278 41030 40330
rect 41092 40278 41104 40330
rect 41166 40278 41168 40330
rect 41006 40276 41030 40278
rect 41086 40276 41110 40278
rect 41166 40276 41190 40278
rect 40950 40256 41246 40276
rect 41314 39548 41366 39554
rect 41314 39490 41366 39496
rect 40950 39244 41246 39264
rect 41006 39242 41030 39244
rect 41086 39242 41110 39244
rect 41166 39242 41190 39244
rect 41028 39190 41030 39242
rect 41092 39190 41104 39242
rect 41166 39190 41168 39242
rect 41006 39188 41030 39190
rect 41086 39188 41110 39190
rect 41166 39188 41190 39190
rect 40950 39168 41246 39188
rect 41326 39010 41354 39490
rect 40854 39004 40906 39010
rect 40854 38946 40906 38952
rect 41314 39004 41366 39010
rect 41314 38946 41366 38952
rect 41314 38868 41366 38874
rect 41314 38810 41366 38816
rect 41326 38262 41354 38810
rect 40854 38256 40906 38262
rect 40854 38198 40906 38204
rect 41314 38256 41366 38262
rect 41314 38198 41366 38204
rect 40578 37916 40630 37922
rect 40578 37858 40630 37864
rect 40394 37848 40446 37854
rect 40394 37790 40446 37796
rect 40302 37440 40354 37446
rect 40302 37382 40354 37388
rect 40406 37174 40434 37790
rect 40590 37786 40618 37858
rect 40578 37780 40630 37786
rect 40578 37722 40630 37728
rect 40486 37712 40538 37718
rect 40486 37654 40538 37660
rect 40498 37514 40526 37654
rect 40486 37508 40538 37514
rect 40486 37450 40538 37456
rect 40486 37304 40538 37310
rect 40486 37246 40538 37252
rect 39842 37168 39894 37174
rect 39842 37110 39894 37116
rect 40394 37168 40446 37174
rect 40394 37110 40446 37116
rect 39854 36290 39882 37110
rect 40498 36902 40526 37246
rect 40486 36896 40538 36902
rect 40486 36838 40538 36844
rect 40498 36358 40526 36838
rect 40866 36766 40894 38198
rect 40950 38156 41246 38176
rect 41006 38154 41030 38156
rect 41086 38154 41110 38156
rect 41166 38154 41190 38156
rect 41028 38102 41030 38154
rect 41092 38102 41104 38154
rect 41166 38102 41168 38154
rect 41006 38100 41030 38102
rect 41086 38100 41110 38102
rect 41166 38100 41190 38102
rect 40950 38080 41246 38100
rect 41418 37938 41446 40442
rect 41602 40234 41630 40510
rect 42706 40506 42734 43312
rect 43614 41964 43910 41984
rect 43670 41962 43694 41964
rect 43750 41962 43774 41964
rect 43830 41962 43854 41964
rect 43692 41910 43694 41962
rect 43756 41910 43768 41962
rect 43830 41910 43832 41962
rect 43670 41908 43694 41910
rect 43750 41908 43774 41910
rect 43830 41908 43854 41910
rect 43614 41888 43910 41908
rect 43614 40876 43910 40896
rect 43670 40874 43694 40876
rect 43750 40874 43774 40876
rect 43830 40874 43854 40876
rect 43692 40822 43694 40874
rect 43756 40822 43768 40874
rect 43830 40822 43832 40874
rect 43670 40820 43694 40822
rect 43750 40820 43774 40822
rect 43830 40820 43854 40822
rect 43614 40800 43910 40820
rect 43994 40574 44022 43312
rect 44074 41044 44126 41050
rect 44074 40986 44126 40992
rect 44086 40642 44114 40986
rect 44074 40636 44126 40642
rect 44074 40578 44126 40584
rect 43982 40568 44034 40574
rect 43982 40510 44034 40516
rect 42694 40500 42746 40506
rect 42694 40442 42746 40448
rect 41590 40228 41642 40234
rect 41590 40170 41642 40176
rect 41958 40024 42010 40030
rect 41958 39966 42010 39972
rect 41970 39690 41998 39966
rect 43062 39888 43114 39894
rect 43062 39830 43114 39836
rect 41958 39684 42010 39690
rect 41958 39626 42010 39632
rect 42878 39684 42930 39690
rect 42878 39626 42930 39632
rect 41774 39140 41826 39146
rect 41774 39082 41826 39088
rect 41786 38942 41814 39082
rect 41774 38936 41826 38942
rect 41774 38878 41826 38884
rect 41786 38602 41814 38878
rect 42326 38800 42378 38806
rect 42326 38742 42378 38748
rect 42338 38602 42366 38742
rect 41774 38596 41826 38602
rect 41774 38538 41826 38544
rect 42326 38596 42378 38602
rect 42326 38538 42378 38544
rect 42338 38058 42366 38538
rect 42326 38052 42378 38058
rect 42326 37994 42378 38000
rect 41050 37910 41446 37938
rect 41050 37718 41078 37910
rect 41222 37848 41274 37854
rect 41222 37790 41274 37796
rect 41774 37848 41826 37854
rect 41774 37790 41826 37796
rect 41234 37718 41262 37790
rect 41786 37718 41814 37790
rect 41038 37712 41090 37718
rect 41038 37654 41090 37660
rect 41222 37712 41274 37718
rect 41774 37712 41826 37718
rect 41222 37654 41274 37660
rect 41772 37680 41774 37689
rect 41826 37680 41828 37689
rect 41234 37417 41262 37654
rect 41772 37615 41828 37624
rect 41220 37408 41276 37417
rect 41220 37343 41276 37352
rect 42142 37372 42194 37378
rect 42142 37314 42194 37320
rect 42154 37174 42182 37314
rect 42890 37310 42918 39626
rect 43074 39554 43102 39830
rect 43614 39788 43910 39808
rect 43670 39786 43694 39788
rect 43750 39786 43774 39788
rect 43830 39786 43854 39788
rect 43692 39734 43694 39786
rect 43756 39734 43768 39786
rect 43830 39734 43832 39786
rect 43670 39732 43694 39734
rect 43750 39732 43774 39734
rect 43830 39732 43854 39734
rect 43614 39712 43910 39732
rect 43062 39548 43114 39554
rect 43062 39490 43114 39496
rect 45190 39350 45218 43312
rect 46386 41610 46414 43312
rect 46386 41582 46690 41610
rect 46278 41420 46574 41440
rect 46334 41418 46358 41420
rect 46414 41418 46438 41420
rect 46494 41418 46518 41420
rect 46356 41366 46358 41418
rect 46420 41366 46432 41418
rect 46494 41366 46496 41418
rect 46334 41364 46358 41366
rect 46414 41364 46438 41366
rect 46494 41364 46518 41366
rect 46278 41344 46574 41364
rect 46662 40574 46690 41582
rect 47110 41112 47162 41118
rect 47110 41054 47162 41060
rect 47386 41112 47438 41118
rect 47386 41054 47438 41060
rect 47122 40982 47150 41054
rect 46742 40976 46794 40982
rect 46742 40918 46794 40924
rect 47110 40976 47162 40982
rect 47110 40918 47162 40924
rect 45730 40568 45782 40574
rect 45730 40510 45782 40516
rect 46650 40568 46702 40574
rect 46650 40510 46702 40516
rect 45742 40098 45770 40510
rect 46278 40332 46574 40352
rect 46334 40330 46358 40332
rect 46414 40330 46438 40332
rect 46494 40330 46518 40332
rect 46356 40278 46358 40330
rect 46420 40278 46432 40330
rect 46494 40278 46496 40330
rect 46334 40276 46358 40278
rect 46414 40276 46438 40278
rect 46494 40276 46518 40278
rect 46278 40256 46574 40276
rect 46754 40234 46782 40918
rect 47122 40778 47150 40918
rect 47110 40772 47162 40778
rect 47110 40714 47162 40720
rect 46742 40228 46794 40234
rect 46742 40170 46794 40176
rect 45730 40092 45782 40098
rect 45730 40034 45782 40040
rect 46754 40030 46782 40170
rect 46742 40024 46794 40030
rect 46742 39966 46794 39972
rect 43062 39344 43114 39350
rect 43062 39286 43114 39292
rect 45178 39344 45230 39350
rect 45178 39286 45230 39292
rect 43074 39010 43102 39286
rect 46278 39244 46574 39264
rect 46334 39242 46358 39244
rect 46414 39242 46438 39244
rect 46494 39242 46518 39244
rect 46356 39190 46358 39242
rect 46420 39190 46432 39242
rect 46494 39190 46496 39242
rect 46334 39188 46358 39190
rect 46414 39188 46438 39190
rect 46494 39188 46518 39190
rect 46278 39168 46574 39188
rect 44810 39140 44862 39146
rect 44810 39082 44862 39088
rect 43062 39004 43114 39010
rect 43062 38946 43114 38952
rect 43154 38936 43206 38942
rect 43154 38878 43206 38884
rect 43166 37530 43194 38878
rect 44822 38874 44850 39082
rect 47202 39072 47254 39078
rect 47202 39014 47254 39020
rect 46006 38936 46058 38942
rect 47214 38924 47242 39014
rect 47294 38936 47346 38942
rect 47214 38896 47294 38924
rect 46006 38878 46058 38884
rect 47294 38878 47346 38884
rect 44718 38868 44770 38874
rect 44718 38810 44770 38816
rect 44810 38868 44862 38874
rect 44810 38810 44862 38816
rect 43614 38700 43910 38720
rect 43670 38698 43694 38700
rect 43750 38698 43774 38700
rect 43830 38698 43854 38700
rect 43692 38646 43694 38698
rect 43756 38646 43768 38698
rect 43830 38646 43832 38698
rect 43670 38644 43694 38646
rect 43750 38644 43774 38646
rect 43830 38644 43854 38646
rect 43614 38624 43910 38644
rect 43522 38528 43574 38534
rect 43522 38470 43574 38476
rect 43534 37854 43562 38470
rect 44730 38466 44758 38810
rect 44718 38460 44770 38466
rect 44718 38402 44770 38408
rect 46018 38262 46046 38878
rect 47398 38806 47426 41054
rect 47674 39690 47702 43312
rect 48870 41322 48898 43312
rect 48942 41964 49238 41984
rect 48998 41962 49022 41964
rect 49078 41962 49102 41964
rect 49158 41962 49182 41964
rect 49020 41910 49022 41962
rect 49084 41910 49096 41962
rect 49158 41910 49160 41962
rect 48998 41908 49022 41910
rect 49078 41908 49102 41910
rect 49158 41908 49182 41910
rect 48942 41888 49238 41908
rect 48858 41316 48910 41322
rect 48858 41258 48910 41264
rect 49502 40976 49554 40982
rect 49502 40918 49554 40924
rect 48942 40876 49238 40896
rect 48998 40874 49022 40876
rect 49078 40874 49102 40876
rect 49158 40874 49182 40876
rect 49020 40822 49022 40874
rect 49084 40822 49096 40874
rect 49158 40822 49160 40874
rect 48998 40820 49022 40822
rect 49078 40820 49102 40822
rect 49158 40820 49182 40822
rect 48942 40800 49238 40820
rect 49514 40642 49542 40918
rect 49502 40636 49554 40642
rect 49502 40578 49554 40584
rect 49778 40568 49830 40574
rect 49778 40510 49830 40516
rect 49502 40024 49554 40030
rect 49502 39966 49554 39972
rect 48942 39788 49238 39808
rect 48998 39786 49022 39788
rect 49078 39786 49102 39788
rect 49158 39786 49182 39788
rect 49020 39734 49022 39786
rect 49084 39734 49096 39786
rect 49158 39734 49160 39786
rect 48998 39732 49022 39734
rect 49078 39732 49102 39734
rect 49158 39732 49182 39734
rect 48942 39712 49238 39732
rect 49514 39690 49542 39966
rect 49790 39690 49818 40510
rect 50066 40166 50094 43312
rect 50790 41180 50842 41186
rect 50790 41122 50842 41128
rect 50054 40160 50106 40166
rect 50054 40102 50106 40108
rect 49870 39956 49922 39962
rect 49870 39898 49922 39904
rect 49882 39690 49910 39898
rect 47662 39684 47714 39690
rect 47662 39626 47714 39632
rect 49502 39684 49554 39690
rect 49502 39626 49554 39632
rect 49778 39684 49830 39690
rect 49778 39626 49830 39632
rect 49870 39684 49922 39690
rect 49870 39626 49922 39632
rect 49514 39554 49542 39626
rect 49502 39548 49554 39554
rect 49502 39490 49554 39496
rect 50330 39140 50382 39146
rect 50514 39140 50566 39146
rect 50330 39082 50382 39088
rect 50434 39100 50514 39128
rect 50342 39049 50370 39082
rect 50328 39040 50384 39049
rect 47478 39004 47530 39010
rect 50328 38975 50384 38984
rect 47478 38946 47530 38952
rect 47386 38800 47438 38806
rect 47386 38742 47438 38748
rect 45454 38256 45506 38262
rect 45454 38198 45506 38204
rect 46006 38256 46058 38262
rect 46006 38198 46058 38204
rect 46098 38256 46150 38262
rect 46098 38198 46150 38204
rect 45362 37984 45414 37990
rect 45362 37926 45414 37932
rect 43522 37848 43574 37854
rect 43522 37790 43574 37796
rect 43614 37612 43910 37632
rect 43670 37610 43694 37612
rect 43750 37610 43774 37612
rect 43830 37610 43854 37612
rect 43692 37558 43694 37610
rect 43756 37558 43768 37610
rect 43830 37558 43832 37610
rect 43670 37556 43694 37558
rect 43750 37556 43774 37558
rect 43830 37556 43854 37558
rect 43614 37536 43910 37556
rect 43166 37502 43286 37530
rect 42878 37304 42930 37310
rect 42878 37246 42930 37252
rect 42142 37168 42194 37174
rect 42142 37110 42194 37116
rect 40950 37068 41246 37088
rect 41006 37066 41030 37068
rect 41086 37066 41110 37068
rect 41166 37066 41190 37068
rect 41028 37014 41030 37066
rect 41092 37014 41104 37066
rect 41166 37014 41168 37066
rect 41006 37012 41030 37014
rect 41086 37012 41110 37014
rect 41166 37012 41190 37014
rect 40950 36992 41246 37012
rect 42890 36766 42918 37246
rect 43062 37236 43114 37242
rect 43062 37178 43114 37184
rect 43074 36902 43102 37178
rect 43062 36896 43114 36902
rect 43062 36838 43114 36844
rect 43074 36766 43102 36838
rect 43258 36766 43286 37502
rect 43612 37408 43668 37417
rect 45374 37378 45402 37926
rect 45466 37854 45494 38198
rect 45454 37848 45506 37854
rect 45454 37790 45506 37796
rect 45546 37712 45598 37718
rect 45546 37654 45598 37660
rect 43612 37343 43614 37352
rect 43666 37343 43668 37352
rect 45086 37372 45138 37378
rect 43614 37314 43666 37320
rect 45086 37314 45138 37320
rect 45362 37372 45414 37378
rect 45362 37314 45414 37320
rect 44166 37168 44218 37174
rect 44166 37110 44218 37116
rect 43982 36896 44034 36902
rect 43982 36838 44034 36844
rect 43706 36828 43758 36834
rect 43706 36770 43758 36776
rect 40854 36760 40906 36766
rect 40854 36702 40906 36708
rect 42694 36760 42746 36766
rect 42694 36702 42746 36708
rect 42878 36760 42930 36766
rect 42878 36702 42930 36708
rect 43062 36760 43114 36766
rect 43062 36702 43114 36708
rect 43246 36760 43298 36766
rect 43718 36737 43746 36770
rect 43246 36702 43298 36708
rect 43704 36728 43760 36737
rect 42706 36630 42734 36702
rect 43258 36630 43286 36702
rect 43704 36663 43760 36672
rect 42694 36624 42746 36630
rect 42694 36566 42746 36572
rect 43246 36624 43298 36630
rect 43246 36566 43298 36572
rect 43614 36524 43910 36544
rect 43670 36522 43694 36524
rect 43750 36522 43774 36524
rect 43830 36522 43854 36524
rect 43692 36470 43694 36522
rect 43756 36470 43768 36522
rect 43830 36470 43832 36522
rect 43670 36468 43694 36470
rect 43750 36468 43774 36470
rect 43830 36468 43854 36470
rect 43614 36448 43910 36468
rect 40486 36352 40538 36358
rect 40486 36294 40538 36300
rect 40578 36352 40630 36358
rect 40578 36294 40630 36300
rect 39842 36284 39894 36290
rect 39842 36226 39894 36232
rect 39854 36086 39882 36226
rect 40118 36216 40170 36222
rect 40118 36158 40170 36164
rect 39842 36080 39894 36086
rect 39842 36022 39894 36028
rect 40026 35672 40078 35678
rect 40026 35614 40078 35620
rect 39842 35604 39894 35610
rect 39842 35546 39894 35552
rect 39854 35202 39882 35546
rect 40038 35338 40066 35614
rect 40026 35332 40078 35338
rect 40026 35274 40078 35280
rect 39842 35196 39894 35202
rect 39894 35156 39974 35184
rect 39842 35138 39894 35144
rect 39762 35054 39882 35082
rect 39290 33700 39342 33706
rect 39290 33642 39342 33648
rect 39658 33700 39710 33706
rect 39658 33642 39710 33648
rect 38286 33260 38582 33280
rect 38342 33258 38366 33260
rect 38422 33258 38446 33260
rect 38502 33258 38526 33260
rect 38364 33206 38366 33258
rect 38428 33206 38440 33258
rect 38502 33206 38504 33258
rect 38342 33204 38366 33206
rect 38422 33204 38446 33206
rect 38502 33204 38526 33206
rect 38286 33184 38582 33204
rect 39302 33162 39330 33642
rect 39670 33434 39698 33642
rect 39658 33428 39710 33434
rect 39658 33370 39710 33376
rect 39566 33360 39618 33366
rect 39566 33302 39618 33308
rect 39290 33156 39342 33162
rect 39290 33098 39342 33104
rect 37818 33020 37870 33026
rect 37818 32962 37870 32968
rect 37830 32890 37858 32962
rect 37818 32884 37870 32890
rect 37818 32826 37870 32832
rect 37726 32816 37778 32822
rect 37726 32758 37778 32764
rect 36070 32068 36122 32074
rect 36070 32010 36122 32016
rect 35334 32000 35386 32006
rect 35334 31942 35386 31948
rect 34978 30714 35098 30730
rect 34978 30708 35110 30714
rect 34978 30702 35058 30708
rect 34978 29898 35006 30702
rect 35058 30650 35110 30656
rect 34966 29892 35018 29898
rect 34966 29834 35018 29840
rect 35150 28260 35202 28266
rect 35150 28202 35202 28208
rect 35162 27058 35190 28202
rect 35242 28056 35294 28062
rect 35346 28044 35374 31942
rect 37542 31728 37594 31734
rect 37542 31670 37594 31676
rect 35622 31628 35918 31648
rect 35678 31626 35702 31628
rect 35758 31626 35782 31628
rect 35838 31626 35862 31628
rect 35700 31574 35702 31626
rect 35764 31574 35776 31626
rect 35838 31574 35840 31626
rect 35678 31572 35702 31574
rect 35758 31572 35782 31574
rect 35838 31572 35862 31574
rect 35622 31552 35918 31572
rect 37358 31320 37410 31326
rect 37358 31262 37410 31268
rect 36990 31252 37042 31258
rect 36990 31194 37042 31200
rect 35426 31184 35478 31190
rect 35426 31126 35478 31132
rect 35438 29014 35466 31126
rect 37002 30850 37030 31194
rect 36990 30844 37042 30850
rect 36990 30786 37042 30792
rect 36990 30640 37042 30646
rect 36910 30588 36990 30594
rect 36910 30582 37042 30588
rect 36910 30566 37030 30582
rect 35622 30540 35918 30560
rect 35678 30538 35702 30540
rect 35758 30538 35782 30540
rect 35838 30538 35862 30540
rect 35700 30486 35702 30538
rect 35764 30486 35776 30538
rect 35838 30486 35840 30538
rect 35678 30484 35702 30486
rect 35758 30484 35782 30486
rect 35838 30484 35862 30486
rect 35622 30464 35918 30484
rect 36806 30436 36858 30442
rect 36806 30378 36858 30384
rect 36346 29620 36398 29626
rect 36346 29562 36398 29568
rect 35622 29452 35918 29472
rect 35678 29450 35702 29452
rect 35758 29450 35782 29452
rect 35838 29450 35862 29452
rect 35700 29398 35702 29450
rect 35764 29398 35776 29450
rect 35838 29398 35840 29450
rect 35678 29396 35702 29398
rect 35758 29396 35782 29398
rect 35838 29396 35862 29398
rect 35622 29376 35918 29396
rect 36358 29354 36386 29562
rect 36346 29348 36398 29354
rect 36346 29290 36398 29296
rect 36254 29280 36306 29286
rect 36254 29222 36306 29228
rect 35886 29144 35938 29150
rect 35886 29086 35938 29092
rect 36162 29144 36214 29150
rect 36162 29086 36214 29092
rect 35426 29008 35478 29014
rect 35426 28950 35478 28956
rect 35438 28690 35466 28950
rect 35438 28662 35558 28690
rect 35530 28606 35558 28662
rect 35426 28600 35478 28606
rect 35426 28542 35478 28548
rect 35518 28600 35570 28606
rect 35518 28542 35570 28548
rect 35438 28198 35466 28542
rect 35898 28538 35926 29086
rect 36174 28742 36202 29086
rect 36266 28742 36294 29222
rect 36714 29144 36766 29150
rect 36714 29086 36766 29092
rect 36726 29014 36754 29086
rect 36714 29008 36766 29014
rect 36714 28950 36766 28956
rect 36162 28736 36214 28742
rect 36162 28678 36214 28684
rect 36254 28736 36306 28742
rect 36254 28678 36306 28684
rect 35886 28532 35938 28538
rect 35886 28474 35938 28480
rect 35622 28364 35918 28384
rect 35678 28362 35702 28364
rect 35758 28362 35782 28364
rect 35838 28362 35862 28364
rect 35700 28310 35702 28362
rect 35764 28310 35776 28362
rect 35838 28310 35840 28362
rect 35678 28308 35702 28310
rect 35758 28308 35782 28310
rect 35838 28308 35862 28310
rect 35622 28288 35918 28308
rect 35426 28192 35478 28198
rect 35426 28134 35478 28140
rect 36174 28062 36202 28678
rect 36162 28056 36214 28062
rect 35346 28016 35558 28044
rect 35242 27998 35294 28004
rect 35254 27586 35282 27998
rect 35242 27580 35294 27586
rect 35242 27522 35294 27528
rect 35242 27444 35294 27450
rect 35242 27386 35294 27392
rect 35254 27178 35282 27386
rect 35242 27172 35294 27178
rect 35242 27114 35294 27120
rect 35162 27030 35282 27058
rect 35254 27024 35282 27030
rect 35254 26996 35466 27024
rect 35150 26968 35202 26974
rect 35150 26910 35202 26916
rect 34966 26900 35018 26906
rect 34966 26842 35018 26848
rect 34874 24928 34926 24934
rect 34874 24870 34926 24876
rect 34414 24792 34466 24798
rect 34414 24734 34466 24740
rect 34320 23536 34376 23545
rect 34320 23471 34376 23480
rect 34426 23234 34454 24734
rect 34886 23914 34914 24870
rect 34874 23908 34926 23914
rect 34874 23850 34926 23856
rect 34598 23704 34650 23710
rect 34598 23646 34650 23652
rect 34414 23228 34466 23234
rect 34414 23170 34466 23176
rect 34610 22826 34638 23646
rect 34598 22820 34650 22826
rect 34598 22762 34650 22768
rect 34610 21618 34638 22762
rect 34782 22480 34834 22486
rect 34780 22448 34782 22457
rect 34834 22448 34836 22457
rect 34780 22383 34836 22392
rect 34610 21590 34730 21618
rect 34598 21392 34650 21398
rect 34598 21334 34650 21340
rect 34138 21188 34190 21194
rect 34138 21130 34190 21136
rect 34506 21052 34558 21058
rect 34506 20994 34558 21000
rect 34414 20304 34466 20310
rect 34412 20272 34414 20281
rect 34466 20272 34468 20281
rect 34412 20207 34468 20216
rect 30826 19828 30878 19834
rect 30826 19770 30878 19776
rect 34518 19562 34546 20994
rect 34506 19556 34558 19562
rect 34506 19498 34558 19504
rect 34414 19216 34466 19222
rect 34412 19184 34414 19193
rect 34466 19184 34468 19193
rect 34412 19119 34468 19128
rect 34414 18876 34466 18882
rect 34518 18864 34546 19498
rect 34610 18882 34638 21334
rect 34702 20650 34730 21590
rect 34782 21392 34834 21398
rect 34780 21360 34782 21369
rect 34834 21360 34836 21369
rect 34780 21295 34836 21304
rect 34690 20644 34742 20650
rect 34690 20586 34742 20592
rect 34978 19562 35006 26842
rect 35162 25002 35190 26910
rect 35150 24996 35202 25002
rect 35150 24938 35202 24944
rect 35162 24322 35190 24938
rect 35150 24316 35202 24322
rect 35150 24258 35202 24264
rect 35334 23024 35386 23030
rect 35334 22966 35386 22972
rect 35346 21194 35374 22966
rect 35438 22146 35466 26996
rect 35530 23794 35558 28016
rect 36162 27998 36214 28004
rect 36712 28024 36768 28033
rect 35794 27988 35846 27994
rect 36712 27959 36714 27968
rect 35794 27930 35846 27936
rect 36766 27959 36768 27968
rect 36714 27930 36766 27936
rect 35806 27450 35834 27930
rect 36162 27580 36214 27586
rect 36162 27522 36214 27528
rect 35794 27444 35846 27450
rect 35794 27386 35846 27392
rect 36174 27382 36202 27522
rect 36162 27376 36214 27382
rect 36162 27318 36214 27324
rect 35622 27276 35918 27296
rect 35678 27274 35702 27276
rect 35758 27274 35782 27276
rect 35838 27274 35862 27276
rect 35700 27222 35702 27274
rect 35764 27222 35776 27274
rect 35838 27222 35840 27274
rect 35678 27220 35702 27222
rect 35758 27220 35782 27222
rect 35838 27220 35862 27222
rect 35622 27200 35918 27220
rect 36174 27110 36202 27318
rect 35610 27104 35662 27110
rect 35610 27046 35662 27052
rect 36162 27104 36214 27110
rect 36162 27046 36214 27052
rect 35622 26906 35650 27046
rect 36346 26968 36398 26974
rect 36346 26910 36398 26916
rect 36530 26968 36582 26974
rect 36530 26910 36582 26916
rect 36714 26968 36766 26974
rect 36714 26910 36766 26916
rect 35610 26900 35662 26906
rect 35610 26842 35662 26848
rect 35978 26492 36030 26498
rect 35978 26434 36030 26440
rect 35622 26188 35918 26208
rect 35678 26186 35702 26188
rect 35758 26186 35782 26188
rect 35838 26186 35862 26188
rect 35700 26134 35702 26186
rect 35764 26134 35776 26186
rect 35838 26134 35840 26186
rect 35678 26132 35702 26134
rect 35758 26132 35782 26134
rect 35838 26132 35862 26134
rect 35622 26112 35918 26132
rect 35990 26090 36018 26434
rect 35978 26084 36030 26090
rect 35978 26026 36030 26032
rect 35622 25100 35918 25120
rect 35678 25098 35702 25100
rect 35758 25098 35782 25100
rect 35838 25098 35862 25100
rect 35700 25046 35702 25098
rect 35764 25046 35776 25098
rect 35838 25046 35840 25098
rect 35678 25044 35702 25046
rect 35758 25044 35782 25046
rect 35838 25044 35862 25046
rect 35622 25024 35918 25044
rect 35622 24012 35918 24032
rect 35678 24010 35702 24012
rect 35758 24010 35782 24012
rect 35838 24010 35862 24012
rect 35700 23958 35702 24010
rect 35764 23958 35776 24010
rect 35838 23958 35840 24010
rect 35678 23956 35702 23958
rect 35758 23956 35782 23958
rect 35838 23956 35862 23958
rect 35622 23936 35918 23956
rect 35530 23766 35650 23794
rect 35622 23710 35650 23766
rect 35610 23704 35662 23710
rect 35610 23646 35662 23652
rect 35622 22924 35918 22944
rect 35678 22922 35702 22924
rect 35758 22922 35782 22924
rect 35838 22922 35862 22924
rect 35700 22870 35702 22922
rect 35764 22870 35776 22922
rect 35838 22870 35840 22922
rect 35678 22868 35702 22870
rect 35758 22868 35782 22870
rect 35838 22868 35862 22870
rect 35622 22848 35918 22868
rect 35426 22140 35478 22146
rect 35426 22082 35478 22088
rect 35426 21936 35478 21942
rect 35426 21878 35478 21884
rect 35334 21188 35386 21194
rect 35334 21130 35386 21136
rect 35346 21058 35374 21130
rect 35438 21126 35466 21878
rect 35622 21836 35918 21856
rect 35678 21834 35702 21836
rect 35758 21834 35782 21836
rect 35838 21834 35862 21836
rect 35700 21782 35702 21834
rect 35764 21782 35776 21834
rect 35838 21782 35840 21834
rect 35678 21780 35702 21782
rect 35758 21780 35782 21782
rect 35838 21780 35862 21782
rect 35622 21760 35918 21780
rect 35886 21528 35938 21534
rect 35886 21470 35938 21476
rect 35898 21126 35926 21470
rect 35426 21120 35478 21126
rect 35426 21062 35478 21068
rect 35886 21120 35938 21126
rect 35886 21062 35938 21068
rect 35334 21052 35386 21058
rect 35334 20994 35386 21000
rect 35622 20748 35918 20768
rect 35678 20746 35702 20748
rect 35758 20746 35782 20748
rect 35838 20746 35862 20748
rect 35700 20694 35702 20746
rect 35764 20694 35776 20746
rect 35838 20694 35840 20746
rect 35678 20692 35702 20694
rect 35758 20692 35782 20694
rect 35838 20692 35862 20694
rect 35622 20672 35918 20692
rect 35622 19660 35918 19680
rect 35678 19658 35702 19660
rect 35758 19658 35782 19660
rect 35838 19658 35862 19660
rect 35700 19606 35702 19658
rect 35764 19606 35776 19658
rect 35838 19606 35840 19658
rect 35678 19604 35702 19606
rect 35758 19604 35782 19606
rect 35838 19604 35862 19606
rect 35622 19584 35918 19604
rect 34966 19556 35018 19562
rect 34966 19498 35018 19504
rect 34978 18882 35006 19498
rect 35426 19352 35478 19358
rect 35426 19294 35478 19300
rect 34466 18836 34546 18864
rect 34598 18876 34650 18882
rect 34414 18818 34466 18824
rect 34598 18818 34650 18824
rect 34966 18876 35018 18882
rect 34966 18818 35018 18824
rect 35438 18270 35466 19294
rect 35518 18740 35570 18746
rect 35518 18682 35570 18688
rect 35530 18338 35558 18682
rect 35622 18572 35918 18592
rect 35678 18570 35702 18572
rect 35758 18570 35782 18572
rect 35838 18570 35862 18572
rect 35700 18518 35702 18570
rect 35764 18518 35776 18570
rect 35838 18518 35840 18570
rect 35678 18516 35702 18518
rect 35758 18516 35782 18518
rect 35838 18516 35862 18518
rect 35622 18496 35918 18516
rect 35518 18332 35570 18338
rect 35518 18274 35570 18280
rect 35426 18264 35478 18270
rect 35426 18206 35478 18212
rect 34414 18128 34466 18134
rect 34412 18096 34414 18105
rect 34466 18096 34468 18105
rect 34412 18031 34468 18040
rect 35622 17484 35918 17504
rect 35678 17482 35702 17484
rect 35758 17482 35782 17484
rect 35838 17482 35862 17484
rect 35700 17430 35702 17482
rect 35764 17430 35776 17482
rect 35838 17430 35840 17482
rect 35678 17428 35702 17430
rect 35758 17428 35782 17430
rect 35838 17428 35862 17430
rect 35622 17408 35918 17428
rect 36358 17182 36386 26910
rect 36542 26090 36570 26910
rect 36530 26084 36582 26090
rect 36530 26026 36582 26032
rect 36726 25954 36754 26910
rect 36818 26294 36846 30378
rect 36910 30238 36938 30566
rect 36898 30232 36950 30238
rect 36898 30174 36950 30180
rect 36910 29762 36938 30174
rect 37370 29898 37398 31262
rect 37358 29892 37410 29898
rect 37358 29834 37410 29840
rect 37370 29762 37398 29834
rect 36898 29756 36950 29762
rect 36898 29698 36950 29704
rect 37358 29756 37410 29762
rect 37358 29698 37410 29704
rect 37266 29280 37318 29286
rect 37266 29222 37318 29228
rect 37278 29150 37306 29222
rect 37266 29144 37318 29150
rect 37266 29086 37318 29092
rect 37450 28600 37502 28606
rect 37450 28542 37502 28548
rect 36898 28532 36950 28538
rect 36898 28474 36950 28480
rect 36910 28266 36938 28474
rect 36898 28260 36950 28266
rect 36898 28202 36950 28208
rect 36990 27648 37042 27654
rect 36990 27590 37042 27596
rect 36806 26288 36858 26294
rect 36806 26230 36858 26236
rect 36714 25948 36766 25954
rect 36714 25890 36766 25896
rect 36806 25472 36858 25478
rect 36806 25414 36858 25420
rect 36714 24656 36766 24662
rect 36714 24598 36766 24604
rect 36726 24186 36754 24598
rect 36714 24180 36766 24186
rect 36714 24122 36766 24128
rect 36530 23636 36582 23642
rect 36530 23578 36582 23584
rect 36542 22554 36570 23578
rect 36726 23030 36754 24122
rect 36818 23914 36846 25414
rect 36898 24792 36950 24798
rect 36898 24734 36950 24740
rect 36806 23908 36858 23914
rect 36806 23850 36858 23856
rect 36818 23710 36846 23850
rect 36806 23704 36858 23710
rect 36806 23646 36858 23652
rect 36714 23024 36766 23030
rect 36714 22966 36766 22972
rect 36530 22548 36582 22554
rect 36530 22490 36582 22496
rect 36530 22140 36582 22146
rect 36530 22082 36582 22088
rect 36622 22140 36674 22146
rect 36622 22082 36674 22088
rect 36542 21602 36570 22082
rect 36530 21596 36582 21602
rect 36530 21538 36582 21544
rect 36634 21058 36662 22082
rect 36726 21738 36754 22966
rect 36910 22622 36938 24734
rect 37002 24322 37030 27590
rect 37174 25812 37226 25818
rect 37174 25754 37226 25760
rect 37082 24792 37134 24798
rect 37082 24734 37134 24740
rect 37094 24458 37122 24734
rect 37082 24452 37134 24458
rect 37082 24394 37134 24400
rect 36990 24316 37042 24322
rect 36990 24258 37042 24264
rect 36898 22616 36950 22622
rect 36898 22558 36950 22564
rect 36714 21732 36766 21738
rect 36714 21674 36766 21680
rect 36622 21052 36674 21058
rect 36622 20994 36674 21000
rect 36438 20304 36490 20310
rect 36438 20246 36490 20252
rect 36450 19290 36478 20246
rect 36438 19284 36490 19290
rect 36438 19226 36490 19232
rect 36346 17176 36398 17182
rect 36346 17118 36398 17124
rect 34414 17040 34466 17046
rect 34412 17008 34414 17017
rect 34466 17008 34468 17017
rect 34412 16943 34468 16952
rect 36358 16842 36386 17118
rect 36450 17114 36478 19226
rect 36726 18474 36754 21674
rect 36990 21596 37042 21602
rect 36990 21538 37042 21544
rect 37002 21505 37030 21538
rect 36988 21496 37044 21505
rect 36988 21431 37044 21440
rect 36714 18468 36766 18474
rect 36714 18410 36766 18416
rect 36726 17318 36754 18410
rect 36714 17312 36766 17318
rect 36714 17254 36766 17260
rect 36438 17108 36490 17114
rect 36438 17050 36490 17056
rect 36346 16836 36398 16842
rect 36346 16778 36398 16784
rect 36344 16600 36400 16609
rect 36344 16535 36400 16544
rect 35622 16396 35918 16416
rect 35678 16394 35702 16396
rect 35758 16394 35782 16396
rect 35838 16394 35862 16396
rect 35700 16342 35702 16394
rect 35764 16342 35776 16394
rect 35838 16342 35840 16394
rect 35678 16340 35702 16342
rect 35758 16340 35782 16342
rect 35838 16340 35862 16342
rect 35622 16320 35918 16340
rect 36358 16298 36386 16535
rect 36346 16292 36398 16298
rect 36346 16234 36398 16240
rect 36450 16094 36478 17050
rect 36438 16088 36490 16094
rect 36438 16030 36490 16036
rect 36726 15754 36754 17254
rect 37186 16094 37214 25754
rect 37462 21194 37490 28542
rect 37554 25342 37582 31670
rect 37738 29354 37766 32758
rect 37830 30782 37858 32826
rect 38094 32544 38146 32550
rect 38094 32486 38146 32492
rect 37818 30776 37870 30782
rect 37818 30718 37870 30724
rect 37818 29552 37870 29558
rect 37818 29494 37870 29500
rect 37830 29354 37858 29494
rect 37726 29348 37778 29354
rect 37726 29290 37778 29296
rect 37818 29348 37870 29354
rect 37818 29290 37870 29296
rect 37818 29212 37870 29218
rect 37818 29154 37870 29160
rect 37830 29121 37858 29154
rect 37816 29112 37872 29121
rect 37726 29076 37778 29082
rect 37816 29047 37872 29056
rect 37726 29018 37778 29024
rect 37738 28810 37766 29018
rect 37726 28804 37778 28810
rect 37726 28746 37778 28752
rect 38106 26634 38134 32486
rect 39302 32482 39330 33098
rect 39290 32476 39342 32482
rect 39290 32418 39342 32424
rect 39474 32408 39526 32414
rect 39474 32350 39526 32356
rect 38286 32172 38582 32192
rect 38342 32170 38366 32172
rect 38422 32170 38446 32172
rect 38502 32170 38526 32172
rect 38364 32118 38366 32170
rect 38428 32118 38440 32170
rect 38502 32118 38504 32170
rect 38342 32116 38366 32118
rect 38422 32116 38446 32118
rect 38502 32116 38526 32118
rect 38286 32096 38582 32116
rect 39486 32006 39514 32350
rect 39474 32000 39526 32006
rect 39474 31942 39526 31948
rect 39578 31938 39606 33302
rect 39750 32952 39802 32958
rect 39750 32894 39802 32900
rect 39566 31932 39618 31938
rect 39566 31874 39618 31880
rect 39762 31734 39790 32894
rect 39750 31728 39802 31734
rect 39750 31670 39802 31676
rect 39854 31530 39882 35054
rect 39946 34114 39974 35156
rect 40038 34658 40066 35274
rect 40130 35134 40158 36158
rect 40590 35882 40618 36294
rect 42878 36080 42930 36086
rect 42878 36022 42930 36028
rect 40950 35980 41246 36000
rect 41006 35978 41030 35980
rect 41086 35978 41110 35980
rect 41166 35978 41190 35980
rect 41028 35926 41030 35978
rect 41092 35926 41104 35978
rect 41166 35926 41168 35978
rect 41006 35924 41030 35926
rect 41086 35924 41110 35926
rect 41166 35924 41190 35926
rect 40950 35904 41246 35924
rect 40578 35876 40630 35882
rect 40578 35818 40630 35824
rect 42890 35746 42918 36022
rect 42878 35740 42930 35746
rect 42878 35682 42930 35688
rect 43994 35542 44022 36838
rect 44074 36692 44126 36698
rect 44074 36634 44126 36640
rect 44086 35746 44114 36634
rect 44074 35740 44126 35746
rect 44074 35682 44126 35688
rect 40762 35536 40814 35542
rect 40762 35478 40814 35484
rect 43062 35536 43114 35542
rect 43062 35478 43114 35484
rect 43982 35536 44034 35542
rect 43982 35478 44034 35484
rect 40578 35264 40630 35270
rect 40578 35206 40630 35212
rect 40118 35128 40170 35134
rect 40118 35070 40170 35076
rect 40130 34794 40158 35070
rect 40118 34788 40170 34794
rect 40118 34730 40170 34736
rect 40210 34788 40262 34794
rect 40210 34730 40262 34736
rect 40026 34652 40078 34658
rect 40026 34594 40078 34600
rect 40118 34584 40170 34590
rect 40118 34526 40170 34532
rect 40130 34182 40158 34526
rect 40222 34454 40250 34730
rect 40590 34590 40618 35206
rect 40578 34584 40630 34590
rect 40578 34526 40630 34532
rect 40670 34584 40722 34590
rect 40670 34526 40722 34532
rect 40302 34516 40354 34522
rect 40302 34458 40354 34464
rect 40210 34448 40262 34454
rect 40210 34390 40262 34396
rect 40118 34176 40170 34182
rect 40118 34118 40170 34124
rect 39934 34108 39986 34114
rect 39934 34050 39986 34056
rect 39934 33428 39986 33434
rect 39934 33370 39986 33376
rect 39946 32618 39974 33370
rect 40026 33020 40078 33026
rect 40026 32962 40078 32968
rect 39934 32612 39986 32618
rect 39934 32554 39986 32560
rect 39842 31524 39894 31530
rect 39842 31466 39894 31472
rect 39946 31326 39974 32554
rect 40038 32482 40066 32962
rect 40130 32929 40158 34118
rect 40314 34114 40342 34458
rect 40682 34182 40710 34526
rect 40670 34176 40722 34182
rect 40670 34118 40722 34124
rect 40302 34108 40354 34114
rect 40302 34050 40354 34056
rect 40394 34108 40446 34114
rect 40394 34050 40446 34056
rect 40116 32920 40172 32929
rect 40116 32855 40172 32864
rect 40026 32476 40078 32482
rect 40026 32418 40078 32424
rect 40038 31530 40066 32418
rect 40406 32414 40434 34050
rect 40670 33700 40722 33706
rect 40670 33642 40722 33648
rect 40682 33502 40710 33642
rect 40578 33496 40630 33502
rect 40578 33438 40630 33444
rect 40670 33496 40722 33502
rect 40670 33438 40722 33444
rect 40590 32618 40618 33438
rect 40774 33042 40802 35478
rect 43074 35338 43102 35478
rect 43614 35436 43910 35456
rect 43670 35434 43694 35436
rect 43750 35434 43774 35436
rect 43830 35434 43854 35436
rect 43692 35382 43694 35434
rect 43756 35382 43768 35434
rect 43830 35382 43832 35434
rect 43670 35380 43694 35382
rect 43750 35380 43774 35382
rect 43830 35380 43854 35382
rect 43614 35360 43910 35380
rect 43062 35332 43114 35338
rect 43062 35274 43114 35280
rect 44178 35202 44206 37110
rect 44256 36728 44312 36737
rect 44256 36663 44312 36672
rect 44270 36193 44298 36663
rect 45098 36222 45126 37314
rect 45374 36290 45402 37314
rect 45454 37168 45506 37174
rect 45454 37110 45506 37116
rect 45466 36873 45494 37110
rect 45558 36902 45586 37654
rect 45546 36896 45598 36902
rect 45452 36864 45508 36873
rect 45546 36838 45598 36844
rect 45452 36799 45508 36808
rect 45362 36284 45414 36290
rect 45466 36272 45494 36799
rect 45558 36766 45586 36838
rect 45546 36760 45598 36766
rect 45546 36702 45598 36708
rect 45638 36284 45690 36290
rect 45466 36244 45638 36272
rect 45362 36226 45414 36232
rect 45638 36226 45690 36232
rect 45086 36216 45138 36222
rect 44256 36184 44312 36193
rect 45086 36158 45138 36164
rect 44256 36119 44312 36128
rect 44626 35604 44678 35610
rect 44626 35546 44678 35552
rect 44166 35196 44218 35202
rect 44166 35138 44218 35144
rect 43430 35128 43482 35134
rect 43430 35070 43482 35076
rect 41314 34992 41366 34998
rect 41314 34934 41366 34940
rect 40950 34892 41246 34912
rect 41006 34890 41030 34892
rect 41086 34890 41110 34892
rect 41166 34890 41190 34892
rect 41028 34838 41030 34890
rect 41092 34838 41104 34890
rect 41166 34838 41168 34890
rect 41006 34836 41030 34838
rect 41086 34836 41110 34838
rect 41166 34836 41190 34838
rect 40950 34816 41246 34836
rect 41326 34658 41354 34934
rect 41314 34652 41366 34658
rect 41314 34594 41366 34600
rect 43338 33904 43390 33910
rect 43338 33846 43390 33852
rect 40950 33804 41246 33824
rect 41006 33802 41030 33804
rect 41086 33802 41110 33804
rect 41166 33802 41190 33804
rect 41028 33750 41030 33802
rect 41092 33750 41104 33802
rect 41166 33750 41168 33802
rect 41006 33748 41030 33750
rect 41086 33748 41110 33750
rect 41166 33748 41190 33750
rect 40950 33728 41246 33748
rect 40682 33014 40802 33042
rect 41130 33020 41182 33026
rect 40682 32958 40710 33014
rect 41130 32962 41182 32968
rect 40670 32952 40722 32958
rect 40670 32894 40722 32900
rect 40762 32952 40814 32958
rect 40762 32894 40814 32900
rect 40578 32612 40630 32618
rect 40578 32554 40630 32560
rect 40682 32550 40710 32894
rect 40670 32544 40722 32550
rect 40670 32486 40722 32492
rect 40394 32408 40446 32414
rect 40394 32350 40446 32356
rect 40670 32408 40722 32414
rect 40774 32396 40802 32894
rect 41142 32890 41170 32962
rect 41130 32884 41182 32890
rect 41130 32826 41182 32832
rect 41774 32884 41826 32890
rect 41774 32826 41826 32832
rect 42326 32884 42378 32890
rect 42326 32826 42378 32832
rect 40854 32816 40906 32822
rect 40854 32758 40906 32764
rect 40722 32368 40802 32396
rect 40670 32350 40722 32356
rect 40762 32068 40814 32074
rect 40762 32010 40814 32016
rect 40774 31870 40802 32010
rect 40866 31938 40894 32758
rect 40950 32716 41246 32736
rect 41006 32714 41030 32716
rect 41086 32714 41110 32716
rect 41166 32714 41190 32716
rect 41028 32662 41030 32714
rect 41092 32662 41104 32714
rect 41166 32662 41168 32714
rect 41006 32660 41030 32662
rect 41086 32660 41110 32662
rect 41166 32660 41190 32662
rect 40950 32640 41246 32660
rect 41682 32408 41734 32414
rect 41786 32385 41814 32826
rect 42338 32482 42366 32826
rect 42326 32476 42378 32482
rect 42326 32418 42378 32424
rect 41682 32350 41734 32356
rect 41772 32376 41828 32385
rect 41694 32074 41722 32350
rect 41772 32311 41828 32320
rect 41682 32068 41734 32074
rect 41682 32010 41734 32016
rect 40854 31932 40906 31938
rect 40854 31874 40906 31880
rect 40762 31864 40814 31870
rect 40762 31806 40814 31812
rect 40950 31628 41246 31648
rect 41006 31626 41030 31628
rect 41086 31626 41110 31628
rect 41166 31626 41190 31628
rect 41028 31574 41030 31626
rect 41092 31574 41104 31626
rect 41166 31574 41168 31626
rect 41006 31572 41030 31574
rect 41086 31572 41110 31574
rect 41166 31572 41190 31574
rect 40950 31552 41246 31572
rect 40026 31524 40078 31530
rect 40026 31466 40078 31472
rect 39934 31320 39986 31326
rect 40854 31320 40906 31326
rect 39934 31262 39986 31268
rect 40852 31288 40854 31297
rect 40906 31288 40908 31297
rect 40852 31223 40908 31232
rect 38286 31084 38582 31104
rect 38342 31082 38366 31084
rect 38422 31082 38446 31084
rect 38502 31082 38526 31084
rect 38364 31030 38366 31082
rect 38428 31030 38440 31082
rect 38502 31030 38504 31082
rect 38342 31028 38366 31030
rect 38422 31028 38446 31030
rect 38502 31028 38526 31030
rect 38286 31008 38582 31028
rect 38646 30980 38698 30986
rect 38646 30922 38698 30928
rect 38658 30442 38686 30922
rect 42878 30776 42930 30782
rect 42878 30718 42930 30724
rect 40950 30540 41246 30560
rect 41006 30538 41030 30540
rect 41086 30538 41110 30540
rect 41166 30538 41190 30540
rect 41028 30486 41030 30538
rect 41092 30486 41104 30538
rect 41166 30486 41168 30538
rect 41006 30484 41030 30486
rect 41086 30484 41110 30486
rect 41166 30484 41190 30486
rect 40950 30464 41246 30484
rect 38646 30436 38698 30442
rect 38646 30378 38698 30384
rect 42786 30436 42838 30442
rect 42786 30378 42838 30384
rect 40946 30368 40998 30374
rect 40946 30310 40998 30316
rect 38186 30096 38238 30102
rect 38186 30038 38238 30044
rect 38646 30096 38698 30102
rect 38646 30038 38698 30044
rect 39750 30096 39802 30102
rect 39750 30038 39802 30044
rect 38198 29014 38226 30038
rect 38286 29996 38582 30016
rect 38342 29994 38366 29996
rect 38422 29994 38446 29996
rect 38502 29994 38526 29996
rect 38364 29942 38366 29994
rect 38428 29942 38440 29994
rect 38502 29942 38504 29994
rect 38342 29940 38366 29942
rect 38422 29940 38446 29942
rect 38502 29940 38526 29942
rect 38286 29920 38582 29940
rect 38658 29286 38686 30038
rect 38830 29756 38882 29762
rect 38830 29698 38882 29704
rect 39198 29756 39250 29762
rect 39198 29698 39250 29704
rect 39474 29756 39526 29762
rect 39474 29698 39526 29704
rect 38646 29280 38698 29286
rect 38646 29222 38698 29228
rect 38842 29150 38870 29698
rect 39210 29558 39238 29698
rect 39198 29552 39250 29558
rect 39198 29494 39250 29500
rect 38830 29144 38882 29150
rect 38276 29112 38332 29121
rect 38830 29086 38882 29092
rect 38276 29047 38278 29056
rect 38330 29047 38332 29056
rect 38278 29018 38330 29024
rect 38186 29008 38238 29014
rect 38186 28950 38238 28956
rect 38286 28908 38582 28928
rect 38342 28906 38366 28908
rect 38422 28906 38446 28908
rect 38502 28906 38526 28908
rect 38364 28854 38366 28906
rect 38428 28854 38440 28906
rect 38502 28854 38504 28906
rect 38342 28852 38366 28854
rect 38422 28852 38446 28854
rect 38502 28852 38526 28854
rect 38286 28832 38582 28852
rect 38842 28674 38870 29086
rect 39014 29008 39066 29014
rect 39014 28950 39066 28956
rect 38830 28668 38882 28674
rect 38830 28610 38882 28616
rect 38554 28600 38606 28606
rect 38554 28542 38606 28548
rect 38370 28464 38422 28470
rect 38370 28406 38422 28412
rect 38186 28192 38238 28198
rect 38186 28134 38238 28140
rect 38094 26628 38146 26634
rect 38094 26570 38146 26576
rect 38106 26498 38134 26570
rect 38094 26492 38146 26498
rect 38094 26434 38146 26440
rect 37726 26288 37778 26294
rect 37726 26230 37778 26236
rect 37542 25336 37594 25342
rect 37542 25278 37594 25284
rect 37450 21188 37502 21194
rect 37450 21130 37502 21136
rect 37462 20990 37490 21130
rect 37450 20984 37502 20990
rect 37450 20926 37502 20932
rect 37462 19562 37490 20926
rect 37450 19556 37502 19562
rect 37450 19498 37502 19504
rect 37554 17590 37582 25278
rect 37634 19964 37686 19970
rect 37634 19906 37686 19912
rect 37646 19358 37674 19906
rect 37634 19352 37686 19358
rect 37634 19294 37686 19300
rect 37646 18882 37674 19294
rect 37634 18876 37686 18882
rect 37634 18818 37686 18824
rect 37542 17584 37594 17590
rect 37542 17526 37594 17532
rect 37358 17244 37410 17250
rect 37358 17186 37410 17192
rect 37174 16088 37226 16094
rect 37174 16030 37226 16036
rect 36714 15748 36766 15754
rect 36714 15690 36766 15696
rect 37370 15618 37398 17186
rect 37738 17046 37766 26230
rect 38106 25410 38134 26434
rect 38094 25404 38146 25410
rect 38094 25346 38146 25352
rect 38198 24866 38226 28134
rect 38382 27994 38410 28406
rect 38566 28062 38594 28542
rect 38554 28056 38606 28062
rect 38554 27998 38606 28004
rect 38370 27988 38422 27994
rect 38370 27930 38422 27936
rect 38646 27988 38698 27994
rect 38646 27930 38698 27936
rect 38286 27820 38582 27840
rect 38342 27818 38366 27820
rect 38422 27818 38446 27820
rect 38502 27818 38526 27820
rect 38364 27766 38366 27818
rect 38428 27766 38440 27818
rect 38502 27766 38504 27818
rect 38342 27764 38366 27766
rect 38422 27764 38446 27766
rect 38502 27764 38526 27766
rect 38286 27744 38582 27764
rect 38658 27722 38686 27930
rect 38738 27920 38790 27926
rect 38738 27862 38790 27868
rect 38646 27716 38698 27722
rect 38646 27658 38698 27664
rect 38286 26732 38582 26752
rect 38342 26730 38366 26732
rect 38422 26730 38446 26732
rect 38502 26730 38526 26732
rect 38364 26678 38366 26730
rect 38428 26678 38440 26730
rect 38502 26678 38504 26730
rect 38342 26676 38366 26678
rect 38422 26676 38446 26678
rect 38502 26676 38526 26678
rect 38286 26656 38582 26676
rect 38554 26424 38606 26430
rect 38554 26366 38606 26372
rect 38566 26294 38594 26366
rect 38554 26288 38606 26294
rect 38554 26230 38606 26236
rect 38286 25644 38582 25664
rect 38342 25642 38366 25644
rect 38422 25642 38446 25644
rect 38502 25642 38526 25644
rect 38364 25590 38366 25642
rect 38428 25590 38440 25642
rect 38502 25590 38504 25642
rect 38342 25588 38366 25590
rect 38422 25588 38446 25590
rect 38502 25588 38526 25590
rect 38286 25568 38582 25588
rect 38186 24860 38238 24866
rect 38186 24802 38238 24808
rect 38186 24724 38238 24730
rect 38186 24666 38238 24672
rect 38198 23234 38226 24666
rect 38286 24556 38582 24576
rect 38342 24554 38366 24556
rect 38422 24554 38446 24556
rect 38502 24554 38526 24556
rect 38364 24502 38366 24554
rect 38428 24502 38440 24554
rect 38502 24502 38504 24554
rect 38342 24500 38366 24502
rect 38422 24500 38446 24502
rect 38502 24500 38526 24502
rect 38286 24480 38582 24500
rect 38646 23568 38698 23574
rect 38646 23510 38698 23516
rect 38286 23468 38582 23488
rect 38342 23466 38366 23468
rect 38422 23466 38446 23468
rect 38502 23466 38526 23468
rect 38364 23414 38366 23466
rect 38428 23414 38440 23466
rect 38502 23414 38504 23466
rect 38342 23412 38366 23414
rect 38422 23412 38446 23414
rect 38502 23412 38526 23414
rect 38286 23392 38582 23412
rect 38186 23228 38238 23234
rect 38186 23170 38238 23176
rect 38658 22622 38686 23510
rect 38646 22616 38698 22622
rect 38646 22558 38698 22564
rect 38094 22480 38146 22486
rect 38094 22422 38146 22428
rect 38106 21058 38134 22422
rect 38286 22380 38582 22400
rect 38342 22378 38366 22380
rect 38422 22378 38446 22380
rect 38502 22378 38526 22380
rect 38364 22326 38366 22378
rect 38428 22326 38440 22378
rect 38502 22326 38504 22378
rect 38342 22324 38366 22326
rect 38422 22324 38446 22326
rect 38502 22324 38526 22326
rect 38286 22304 38582 22324
rect 38750 21670 38778 27862
rect 38842 27722 38870 28610
rect 38830 27716 38882 27722
rect 38830 27658 38882 27664
rect 38830 27580 38882 27586
rect 38830 27522 38882 27528
rect 38842 27466 38870 27522
rect 38842 27438 38962 27466
rect 38830 25744 38882 25750
rect 38830 25686 38882 25692
rect 38842 25410 38870 25686
rect 38830 25404 38882 25410
rect 38830 25346 38882 25352
rect 38830 24860 38882 24866
rect 38830 24802 38882 24808
rect 38738 21664 38790 21670
rect 38738 21606 38790 21612
rect 38842 21516 38870 24802
rect 38750 21488 38870 21516
rect 38286 21292 38582 21312
rect 38342 21290 38366 21292
rect 38422 21290 38446 21292
rect 38502 21290 38526 21292
rect 38364 21238 38366 21290
rect 38428 21238 38440 21290
rect 38502 21238 38504 21290
rect 38342 21236 38366 21238
rect 38422 21236 38446 21238
rect 38502 21236 38526 21238
rect 38286 21216 38582 21236
rect 38094 21052 38146 21058
rect 38094 20994 38146 21000
rect 38106 17794 38134 20994
rect 38286 20204 38582 20224
rect 38342 20202 38366 20204
rect 38422 20202 38446 20204
rect 38502 20202 38526 20204
rect 38364 20150 38366 20202
rect 38428 20150 38440 20202
rect 38502 20150 38504 20202
rect 38342 20148 38366 20150
rect 38422 20148 38446 20150
rect 38502 20148 38526 20150
rect 38286 20128 38582 20148
rect 38286 19116 38582 19136
rect 38342 19114 38366 19116
rect 38422 19114 38446 19116
rect 38502 19114 38526 19116
rect 38364 19062 38366 19114
rect 38428 19062 38440 19114
rect 38502 19062 38504 19114
rect 38342 19060 38366 19062
rect 38422 19060 38446 19062
rect 38502 19060 38526 19062
rect 38286 19040 38582 19060
rect 38286 18028 38582 18048
rect 38342 18026 38366 18028
rect 38422 18026 38446 18028
rect 38502 18026 38526 18028
rect 38364 17974 38366 18026
rect 38428 17974 38440 18026
rect 38502 17974 38504 18026
rect 38342 17972 38366 17974
rect 38422 17972 38446 17974
rect 38502 17972 38526 17974
rect 38286 17952 38582 17972
rect 38094 17788 38146 17794
rect 38094 17730 38146 17736
rect 38002 17584 38054 17590
rect 38002 17526 38054 17532
rect 37726 17040 37778 17046
rect 37726 16982 37778 16988
rect 38014 16298 38042 17526
rect 38750 17182 38778 21488
rect 38934 19358 38962 27438
rect 39026 27042 39054 28950
rect 39486 28674 39514 29698
rect 39762 29626 39790 30038
rect 40958 29898 40986 30310
rect 40946 29892 40998 29898
rect 40946 29834 40998 29840
rect 42798 29762 42826 30378
rect 42786 29756 42838 29762
rect 42786 29698 42838 29704
rect 39750 29620 39802 29626
rect 39750 29562 39802 29568
rect 40950 29452 41246 29472
rect 41006 29450 41030 29452
rect 41086 29450 41110 29452
rect 41166 29450 41190 29452
rect 41028 29398 41030 29450
rect 41092 29398 41104 29450
rect 41166 29398 41168 29450
rect 41006 29396 41030 29398
rect 41086 29396 41110 29398
rect 41166 29396 41190 29398
rect 40950 29376 41246 29396
rect 42234 29348 42286 29354
rect 42234 29290 42286 29296
rect 42246 29150 42274 29290
rect 41774 29144 41826 29150
rect 41774 29086 41826 29092
rect 42234 29144 42286 29150
rect 42234 29086 42286 29092
rect 42326 29144 42378 29150
rect 42326 29086 42378 29092
rect 39566 28736 39618 28742
rect 39566 28678 39618 28684
rect 39198 28668 39250 28674
rect 39198 28610 39250 28616
rect 39474 28668 39526 28674
rect 39474 28610 39526 28616
rect 39210 28470 39238 28610
rect 39198 28464 39250 28470
rect 39198 28406 39250 28412
rect 39210 28198 39238 28406
rect 39198 28192 39250 28198
rect 39198 28134 39250 28140
rect 39014 27036 39066 27042
rect 39014 26978 39066 26984
rect 39290 26968 39342 26974
rect 39290 26910 39342 26916
rect 39302 26498 39330 26910
rect 39382 26628 39434 26634
rect 39382 26570 39434 26576
rect 39394 26498 39422 26570
rect 39290 26492 39342 26498
rect 39290 26434 39342 26440
rect 39382 26492 39434 26498
rect 39382 26434 39434 26440
rect 39302 26090 39330 26434
rect 39290 26084 39342 26090
rect 39290 26026 39342 26032
rect 39290 25200 39342 25206
rect 39290 25142 39342 25148
rect 39302 22282 39330 25142
rect 39474 24316 39526 24322
rect 39474 24258 39526 24264
rect 39486 24186 39514 24258
rect 39474 24180 39526 24186
rect 39474 24122 39526 24128
rect 39486 23370 39514 24122
rect 39474 23364 39526 23370
rect 39474 23306 39526 23312
rect 39578 23302 39606 28678
rect 40670 28668 40722 28674
rect 40670 28610 40722 28616
rect 39842 28532 39894 28538
rect 39842 28474 39894 28480
rect 39750 28464 39802 28470
rect 39750 28406 39802 28412
rect 39762 27654 39790 28406
rect 39750 27648 39802 27654
rect 39750 27590 39802 27596
rect 39566 23296 39618 23302
rect 39566 23238 39618 23244
rect 39658 22480 39710 22486
rect 39658 22422 39710 22428
rect 39290 22276 39342 22282
rect 39290 22218 39342 22224
rect 39302 22078 39330 22218
rect 39290 22072 39342 22078
rect 39290 22014 39342 22020
rect 39302 20106 39330 22014
rect 39670 21738 39698 22422
rect 39658 21732 39710 21738
rect 39658 21674 39710 21680
rect 39474 21392 39526 21398
rect 39474 21334 39526 21340
rect 39486 21058 39514 21334
rect 39670 21194 39698 21674
rect 39854 21534 39882 28474
rect 40578 28260 40630 28266
rect 40578 28202 40630 28208
rect 39842 21528 39894 21534
rect 39842 21470 39894 21476
rect 39658 21188 39710 21194
rect 39658 21130 39710 21136
rect 39474 21052 39526 21058
rect 39474 20994 39526 21000
rect 39670 20990 39698 21130
rect 39658 20984 39710 20990
rect 39658 20926 39710 20932
rect 39670 20650 39698 20926
rect 39658 20644 39710 20650
rect 39658 20586 39710 20592
rect 39290 20100 39342 20106
rect 39290 20042 39342 20048
rect 39302 19986 39330 20042
rect 39210 19958 39330 19986
rect 39210 19902 39238 19958
rect 39198 19896 39250 19902
rect 39198 19838 39250 19844
rect 38922 19352 38974 19358
rect 38922 19294 38974 19300
rect 39382 19284 39434 19290
rect 39382 19226 39434 19232
rect 39394 18882 39422 19226
rect 39670 19018 39698 20586
rect 40590 19442 40618 28202
rect 40682 28062 40710 28610
rect 40950 28364 41246 28384
rect 41006 28362 41030 28364
rect 41086 28362 41110 28364
rect 41166 28362 41190 28364
rect 41028 28310 41030 28362
rect 41092 28310 41104 28362
rect 41166 28310 41168 28362
rect 41006 28308 41030 28310
rect 41086 28308 41110 28310
rect 41166 28308 41190 28310
rect 40950 28288 41246 28308
rect 41786 28062 41814 29086
rect 42338 29014 42366 29086
rect 42326 29008 42378 29014
rect 42326 28950 42378 28956
rect 42890 28810 42918 30718
rect 43062 30096 43114 30102
rect 43062 30038 43114 30044
rect 43074 29898 43102 30038
rect 43062 29892 43114 29898
rect 43062 29834 43114 29840
rect 43062 29756 43114 29762
rect 43062 29698 43114 29704
rect 42970 29144 43022 29150
rect 42970 29086 43022 29092
rect 42878 28804 42930 28810
rect 42878 28746 42930 28752
rect 42878 28464 42930 28470
rect 42878 28406 42930 28412
rect 40670 28056 40722 28062
rect 40670 27998 40722 28004
rect 41774 28056 41826 28062
rect 41774 27998 41826 28004
rect 42510 27988 42562 27994
rect 42510 27930 42562 27936
rect 42522 27722 42550 27930
rect 42890 27926 42918 28406
rect 42982 28130 43010 29086
rect 43074 28742 43102 29698
rect 43062 28736 43114 28742
rect 43062 28678 43114 28684
rect 42970 28124 43022 28130
rect 42970 28066 43022 28072
rect 42878 27920 42930 27926
rect 42878 27862 42930 27868
rect 42510 27716 42562 27722
rect 42510 27658 42562 27664
rect 42786 27716 42838 27722
rect 42786 27658 42838 27664
rect 42798 27586 42826 27658
rect 42786 27580 42838 27586
rect 42786 27522 42838 27528
rect 42234 27512 42286 27518
rect 42234 27454 42286 27460
rect 40950 27276 41246 27296
rect 41006 27274 41030 27276
rect 41086 27274 41110 27276
rect 41166 27274 41190 27276
rect 41028 27222 41030 27274
rect 41092 27222 41104 27274
rect 41166 27222 41168 27274
rect 41006 27220 41030 27222
rect 41086 27220 41110 27222
rect 41166 27220 41190 27222
rect 40950 27200 41246 27220
rect 40854 26288 40906 26294
rect 40854 26230 40906 26236
rect 40866 24866 40894 26230
rect 40950 26188 41246 26208
rect 41006 26186 41030 26188
rect 41086 26186 41110 26188
rect 41166 26186 41190 26188
rect 41028 26134 41030 26186
rect 41092 26134 41104 26186
rect 41166 26134 41168 26186
rect 41006 26132 41030 26134
rect 41086 26132 41110 26134
rect 41166 26132 41190 26134
rect 40950 26112 41246 26132
rect 42246 25886 42274 27454
rect 42510 26968 42562 26974
rect 42510 26910 42562 26916
rect 42522 25954 42550 26910
rect 42890 26566 42918 27862
rect 42982 27586 43010 28066
rect 43062 28056 43114 28062
rect 43062 27998 43114 28004
rect 43074 27586 43102 27998
rect 43246 27920 43298 27926
rect 43246 27862 43298 27868
rect 42970 27580 43022 27586
rect 42970 27522 43022 27528
rect 43062 27580 43114 27586
rect 43062 27522 43114 27528
rect 42982 27382 43010 27522
rect 42970 27376 43022 27382
rect 42970 27318 43022 27324
rect 43258 27178 43286 27862
rect 43246 27172 43298 27178
rect 43246 27114 43298 27120
rect 42878 26560 42930 26566
rect 42878 26502 42930 26508
rect 42510 25948 42562 25954
rect 42510 25890 42562 25896
rect 42234 25880 42286 25886
rect 42234 25822 42286 25828
rect 40950 25100 41246 25120
rect 41006 25098 41030 25100
rect 41086 25098 41110 25100
rect 41166 25098 41190 25100
rect 41028 25046 41030 25098
rect 41092 25046 41104 25098
rect 41166 25046 41168 25098
rect 41006 25044 41030 25046
rect 41086 25044 41110 25046
rect 41166 25044 41190 25046
rect 40950 25024 41246 25044
rect 42246 25002 42274 25822
rect 42522 25478 42550 25890
rect 42510 25472 42562 25478
rect 42510 25414 42562 25420
rect 42234 24996 42286 25002
rect 42234 24938 42286 24944
rect 40854 24860 40906 24866
rect 40854 24802 40906 24808
rect 40950 24012 41246 24032
rect 41006 24010 41030 24012
rect 41086 24010 41110 24012
rect 41166 24010 41190 24012
rect 41028 23958 41030 24010
rect 41092 23958 41104 24010
rect 41166 23958 41168 24010
rect 41006 23956 41030 23958
rect 41086 23956 41110 23958
rect 41166 23956 41190 23958
rect 40950 23936 41246 23956
rect 42326 23772 42378 23778
rect 42326 23714 42378 23720
rect 42338 23166 42366 23714
rect 42326 23160 42378 23166
rect 42326 23102 42378 23108
rect 40670 23024 40722 23030
rect 40670 22966 40722 22972
rect 40682 22146 40710 22966
rect 40950 22924 41246 22944
rect 41006 22922 41030 22924
rect 41086 22922 41110 22924
rect 41166 22922 41190 22924
rect 41028 22870 41030 22922
rect 41092 22870 41104 22922
rect 41166 22870 41168 22922
rect 41006 22868 41030 22870
rect 41086 22868 41110 22870
rect 41166 22868 41190 22870
rect 40950 22848 41246 22868
rect 42338 22690 42366 23102
rect 42326 22684 42378 22690
rect 42326 22626 42378 22632
rect 40946 22616 40998 22622
rect 40946 22558 40998 22564
rect 40958 22282 40986 22558
rect 43062 22480 43114 22486
rect 43060 22448 43062 22457
rect 43114 22448 43116 22457
rect 43060 22383 43116 22392
rect 40946 22276 40998 22282
rect 40946 22218 40998 22224
rect 40670 22140 40722 22146
rect 40670 22082 40722 22088
rect 40950 21836 41246 21856
rect 41006 21834 41030 21836
rect 41086 21834 41110 21836
rect 41166 21834 41190 21836
rect 41028 21782 41030 21834
rect 41092 21782 41104 21834
rect 41166 21782 41168 21834
rect 41006 21780 41030 21782
rect 41086 21780 41110 21782
rect 41166 21780 41190 21782
rect 40950 21760 41246 21780
rect 43062 21664 43114 21670
rect 43062 21606 43114 21612
rect 41498 21528 41550 21534
rect 41498 21470 41550 21476
rect 41510 20854 41538 21470
rect 43074 21398 43102 21606
rect 43062 21392 43114 21398
rect 43060 21360 43062 21369
rect 43114 21360 43116 21369
rect 43060 21295 43116 21304
rect 41498 20848 41550 20854
rect 41498 20790 41550 20796
rect 40950 20748 41246 20768
rect 41006 20746 41030 20748
rect 41086 20746 41110 20748
rect 41166 20746 41190 20748
rect 41028 20694 41030 20746
rect 41092 20694 41104 20746
rect 41166 20694 41168 20746
rect 41006 20692 41030 20694
rect 41086 20692 41110 20694
rect 41166 20692 41190 20694
rect 40950 20672 41246 20692
rect 40946 20440 40998 20446
rect 40946 20382 40998 20388
rect 40958 19902 40986 20382
rect 41510 20009 41538 20790
rect 43062 20508 43114 20514
rect 43062 20450 43114 20456
rect 42326 20372 42378 20378
rect 42326 20314 42378 20320
rect 41496 20000 41552 20009
rect 42338 19970 42366 20314
rect 43074 20310 43102 20450
rect 43062 20304 43114 20310
rect 43060 20272 43062 20281
rect 43114 20272 43116 20281
rect 43060 20207 43116 20216
rect 41496 19935 41552 19944
rect 42326 19964 42378 19970
rect 42326 19906 42378 19912
rect 40946 19896 40998 19902
rect 40946 19838 40998 19844
rect 40950 19660 41246 19680
rect 41006 19658 41030 19660
rect 41086 19658 41110 19660
rect 41166 19658 41190 19660
rect 41028 19606 41030 19658
rect 41092 19606 41104 19658
rect 41166 19606 41168 19658
rect 41006 19604 41030 19606
rect 41086 19604 41110 19606
rect 41166 19604 41190 19606
rect 40950 19584 41246 19604
rect 40590 19414 40710 19442
rect 40578 19352 40630 19358
rect 40578 19294 40630 19300
rect 40590 19018 40618 19294
rect 39658 19012 39710 19018
rect 39658 18954 39710 18960
rect 40578 19012 40630 19018
rect 40578 18954 40630 18960
rect 39382 18876 39434 18882
rect 39382 18818 39434 18824
rect 39670 18474 39698 18954
rect 39658 18468 39710 18474
rect 39658 18410 39710 18416
rect 40682 17794 40710 19414
rect 42338 19193 42366 19906
rect 42324 19184 42380 19193
rect 42324 19119 42380 19128
rect 43350 18762 43378 33846
rect 43442 30782 43470 35070
rect 44442 34516 44494 34522
rect 44442 34458 44494 34464
rect 43522 34448 43574 34454
rect 43522 34390 43574 34396
rect 43534 33910 43562 34390
rect 43614 34348 43910 34368
rect 43670 34346 43694 34348
rect 43750 34346 43774 34348
rect 43830 34346 43854 34348
rect 43692 34294 43694 34346
rect 43756 34294 43768 34346
rect 43830 34294 43832 34346
rect 43670 34292 43694 34294
rect 43750 34292 43774 34294
rect 43830 34292 43854 34294
rect 43614 34272 43910 34292
rect 43522 33904 43574 33910
rect 43522 33846 43574 33852
rect 44454 33638 44482 34458
rect 44442 33632 44494 33638
rect 44442 33574 44494 33580
rect 43522 33496 43574 33502
rect 43522 33438 43574 33444
rect 43982 33496 44034 33502
rect 43982 33438 44034 33444
rect 43534 31938 43562 33438
rect 43994 33366 44022 33438
rect 43982 33360 44034 33366
rect 43982 33302 44034 33308
rect 43614 33260 43910 33280
rect 43670 33258 43694 33260
rect 43750 33258 43774 33260
rect 43830 33258 43854 33260
rect 43692 33206 43694 33258
rect 43756 33206 43768 33258
rect 43830 33206 43832 33258
rect 43670 33204 43694 33206
rect 43750 33204 43774 33206
rect 43830 33204 43854 33206
rect 43614 33184 43910 33204
rect 43994 33162 44022 33302
rect 43982 33156 44034 33162
rect 43982 33098 44034 33104
rect 43994 32346 44022 33098
rect 44074 33088 44126 33094
rect 44074 33030 44126 33036
rect 44086 32414 44114 33030
rect 44442 33020 44494 33026
rect 44442 32962 44494 32968
rect 44454 32822 44482 32962
rect 44166 32816 44218 32822
rect 44166 32758 44218 32764
rect 44442 32816 44494 32822
rect 44442 32758 44494 32764
rect 44178 32618 44206 32758
rect 44166 32612 44218 32618
rect 44166 32554 44218 32560
rect 44454 32550 44482 32758
rect 44442 32544 44494 32550
rect 44442 32486 44494 32492
rect 44074 32408 44126 32414
rect 44074 32350 44126 32356
rect 43982 32340 44034 32346
rect 43982 32282 44034 32288
rect 43614 32172 43910 32192
rect 43670 32170 43694 32172
rect 43750 32170 43774 32172
rect 43830 32170 43854 32172
rect 43692 32118 43694 32170
rect 43756 32118 43768 32170
rect 43830 32118 43832 32170
rect 43670 32116 43694 32118
rect 43750 32116 43774 32118
rect 43830 32116 43854 32118
rect 43614 32096 43910 32116
rect 43522 31932 43574 31938
rect 43522 31874 43574 31880
rect 43430 30776 43482 30782
rect 43430 30718 43482 30724
rect 43534 30186 43562 31874
rect 44442 31456 44494 31462
rect 44442 31398 44494 31404
rect 43614 31084 43910 31104
rect 43670 31082 43694 31084
rect 43750 31082 43774 31084
rect 43830 31082 43854 31084
rect 43692 31030 43694 31082
rect 43756 31030 43768 31082
rect 43830 31030 43832 31082
rect 43670 31028 43694 31030
rect 43750 31028 43774 31030
rect 43830 31028 43854 31030
rect 43614 31008 43910 31028
rect 44454 30850 44482 31398
rect 44638 30850 44666 35546
rect 45098 34182 45126 36158
rect 45178 35196 45230 35202
rect 45178 35138 45230 35144
rect 45086 34176 45138 34182
rect 45086 34118 45138 34124
rect 45190 34114 45218 35138
rect 45178 34108 45230 34114
rect 45178 34050 45230 34056
rect 44718 33360 44770 33366
rect 44718 33302 44770 33308
rect 44992 33328 45048 33337
rect 44730 33026 44758 33302
rect 44992 33263 45048 33272
rect 44718 33020 44770 33026
rect 44718 32962 44770 32968
rect 45006 32958 45034 33263
rect 44994 32952 45046 32958
rect 44900 32920 44956 32929
rect 44994 32894 45046 32900
rect 44900 32855 44902 32864
rect 44954 32855 44956 32864
rect 44902 32826 44954 32832
rect 44810 32816 44862 32822
rect 44810 32758 44862 32764
rect 44822 32006 44850 32758
rect 44810 32000 44862 32006
rect 44810 31942 44862 31948
rect 45190 31938 45218 34050
rect 46018 33706 46046 38198
rect 46110 35338 46138 38198
rect 46278 38156 46574 38176
rect 46334 38154 46358 38156
rect 46414 38154 46438 38156
rect 46494 38154 46518 38156
rect 46356 38102 46358 38154
rect 46420 38102 46432 38154
rect 46494 38102 46496 38154
rect 46334 38100 46358 38102
rect 46414 38100 46438 38102
rect 46494 38100 46518 38102
rect 46278 38080 46574 38100
rect 47386 37984 47438 37990
rect 47386 37926 47438 37932
rect 46834 37848 46886 37854
rect 46834 37790 46886 37796
rect 46558 37372 46610 37378
rect 46558 37314 46610 37320
rect 46742 37372 46794 37378
rect 46742 37314 46794 37320
rect 46570 37224 46598 37314
rect 46570 37196 46690 37224
rect 46278 37068 46574 37088
rect 46334 37066 46358 37068
rect 46414 37066 46438 37068
rect 46494 37066 46518 37068
rect 46356 37014 46358 37066
rect 46420 37014 46432 37066
rect 46494 37014 46496 37066
rect 46334 37012 46358 37014
rect 46414 37012 46438 37014
rect 46494 37012 46518 37014
rect 46278 36992 46574 37012
rect 46558 36760 46610 36766
rect 46662 36714 46690 37196
rect 46754 36766 46782 37314
rect 46846 36766 46874 37790
rect 47398 37786 47426 37926
rect 47490 37922 47518 38946
rect 50434 38942 50462 39100
rect 50514 39082 50566 39088
rect 48030 38936 48082 38942
rect 48030 38878 48082 38884
rect 50422 38936 50474 38942
rect 50422 38878 50474 38884
rect 47570 38800 47622 38806
rect 47570 38742 47622 38748
rect 47582 38602 47610 38742
rect 48042 38602 48070 38878
rect 50802 38874 50830 41122
rect 51066 41112 51118 41118
rect 51066 41054 51118 41060
rect 51078 40710 51106 41054
rect 51066 40704 51118 40710
rect 51066 40646 51118 40652
rect 51262 40642 51290 43312
rect 51606 41420 51902 41440
rect 51662 41418 51686 41420
rect 51742 41418 51766 41420
rect 51822 41418 51846 41420
rect 51684 41366 51686 41418
rect 51748 41366 51760 41418
rect 51822 41366 51824 41418
rect 51662 41364 51686 41366
rect 51742 41364 51766 41366
rect 51822 41364 51846 41366
rect 51606 41344 51902 41364
rect 52550 41186 52578 43312
rect 53746 41322 53774 43312
rect 54270 41964 54566 41984
rect 54326 41962 54350 41964
rect 54406 41962 54430 41964
rect 54486 41962 54510 41964
rect 54348 41910 54350 41962
rect 54412 41910 54424 41962
rect 54486 41910 54488 41962
rect 54326 41908 54350 41910
rect 54406 41908 54430 41910
rect 54486 41908 54510 41910
rect 54270 41888 54566 41908
rect 53734 41316 53786 41322
rect 53734 41258 53786 41264
rect 52538 41180 52590 41186
rect 52538 41122 52590 41128
rect 51434 41112 51486 41118
rect 51434 41054 51486 41060
rect 54654 41112 54706 41118
rect 54654 41054 54706 41060
rect 51250 40636 51302 40642
rect 51250 40578 51302 40584
rect 51342 40432 51394 40438
rect 51342 40374 51394 40380
rect 51158 40024 51210 40030
rect 51158 39966 51210 39972
rect 51170 39010 51198 39966
rect 51158 39004 51210 39010
rect 51158 38946 51210 38952
rect 50790 38868 50842 38874
rect 50790 38810 50842 38816
rect 48942 38700 49238 38720
rect 48998 38698 49022 38700
rect 49078 38698 49102 38700
rect 49158 38698 49182 38700
rect 49020 38646 49022 38698
rect 49084 38646 49096 38698
rect 49158 38646 49160 38698
rect 48998 38644 49022 38646
rect 49078 38644 49102 38646
rect 49158 38644 49182 38646
rect 48942 38624 49238 38644
rect 51354 38602 51382 40374
rect 51446 40098 51474 41054
rect 54270 40876 54566 40896
rect 54326 40874 54350 40876
rect 54406 40874 54430 40876
rect 54486 40874 54510 40876
rect 54348 40822 54350 40874
rect 54412 40822 54424 40874
rect 54486 40822 54488 40874
rect 54326 40820 54350 40822
rect 54406 40820 54430 40822
rect 54486 40820 54510 40822
rect 54270 40800 54566 40820
rect 51606 40332 51902 40352
rect 51662 40330 51686 40332
rect 51742 40330 51766 40332
rect 51822 40330 51846 40332
rect 51684 40278 51686 40330
rect 51748 40278 51760 40330
rect 51822 40278 51824 40330
rect 51662 40276 51686 40278
rect 51742 40276 51766 40278
rect 51822 40276 51846 40278
rect 51606 40256 51902 40276
rect 51434 40092 51486 40098
rect 51434 40034 51486 40040
rect 54666 40030 54694 41054
rect 54942 40250 54970 43312
rect 56034 41112 56086 41118
rect 55954 41072 56034 41100
rect 55574 40976 55626 40982
rect 55574 40918 55626 40924
rect 55850 40976 55902 40982
rect 55954 40964 55982 41072
rect 56034 41054 56086 41060
rect 55902 40936 55982 40964
rect 55850 40918 55902 40924
rect 55586 40642 55614 40918
rect 56138 40642 56166 43312
rect 56934 41420 57230 41440
rect 56990 41418 57014 41420
rect 57070 41418 57094 41420
rect 57150 41418 57174 41420
rect 57012 41366 57014 41418
rect 57076 41366 57088 41418
rect 57150 41366 57152 41418
rect 56990 41364 57014 41366
rect 57070 41364 57094 41366
rect 57150 41364 57174 41366
rect 56934 41344 57230 41364
rect 56770 41112 56822 41118
rect 56770 41054 56822 41060
rect 56678 40976 56730 40982
rect 56678 40918 56730 40924
rect 55574 40636 55626 40642
rect 55574 40578 55626 40584
rect 56126 40636 56178 40642
rect 56126 40578 56178 40584
rect 56690 40574 56718 40918
rect 56782 40710 56810 41054
rect 56770 40704 56822 40710
rect 56770 40646 56822 40652
rect 55850 40568 55902 40574
rect 55850 40510 55902 40516
rect 56678 40568 56730 40574
rect 56678 40510 56730 40516
rect 54850 40222 54970 40250
rect 55862 40234 55890 40510
rect 55850 40228 55902 40234
rect 54654 40024 54706 40030
rect 54654 39966 54706 39972
rect 54270 39788 54566 39808
rect 54326 39786 54350 39788
rect 54406 39786 54430 39788
rect 54486 39786 54510 39788
rect 54348 39734 54350 39786
rect 54412 39734 54424 39786
rect 54486 39734 54488 39786
rect 54326 39732 54350 39734
rect 54406 39732 54430 39734
rect 54486 39732 54510 39734
rect 54270 39712 54566 39732
rect 53918 39548 53970 39554
rect 53918 39490 53970 39496
rect 51606 39244 51902 39264
rect 51662 39242 51686 39244
rect 51742 39242 51766 39244
rect 51822 39242 51846 39244
rect 51684 39190 51686 39242
rect 51748 39190 51760 39242
rect 51822 39190 51824 39242
rect 51662 39188 51686 39190
rect 51742 39188 51766 39190
rect 51822 39188 51846 39190
rect 51606 39168 51902 39188
rect 52170 39140 52222 39146
rect 52170 39082 52222 39088
rect 52182 38942 52210 39082
rect 53930 39010 53958 39490
rect 54654 39480 54706 39486
rect 54654 39422 54706 39428
rect 54194 39344 54246 39350
rect 54194 39286 54246 39292
rect 54206 39146 54234 39286
rect 54194 39140 54246 39146
rect 54194 39082 54246 39088
rect 53918 39004 53970 39010
rect 53918 38946 53970 38952
rect 51710 38936 51762 38942
rect 52170 38936 52222 38942
rect 51762 38884 51934 38890
rect 51710 38878 51934 38884
rect 52170 38878 52222 38884
rect 52262 38936 52314 38942
rect 52262 38878 52314 38884
rect 51722 38862 51934 38878
rect 47570 38596 47622 38602
rect 47570 38538 47622 38544
rect 48030 38596 48082 38602
rect 48030 38538 48082 38544
rect 51342 38596 51394 38602
rect 51342 38538 51394 38544
rect 48122 38460 48174 38466
rect 48122 38402 48174 38408
rect 48134 38262 48162 38402
rect 51354 38346 51382 38538
rect 51906 38482 51934 38862
rect 51906 38466 52026 38482
rect 51906 38460 52038 38466
rect 51906 38454 51986 38460
rect 51986 38402 52038 38408
rect 51262 38318 51382 38346
rect 48122 38256 48174 38262
rect 48122 38198 48174 38204
rect 47478 37916 47530 37922
rect 47478 37858 47530 37864
rect 47386 37780 47438 37786
rect 47386 37722 47438 37728
rect 47398 37514 47426 37722
rect 47386 37508 47438 37514
rect 47386 37450 47438 37456
rect 46926 37440 46978 37446
rect 46926 37382 46978 37388
rect 46938 37281 46966 37382
rect 46924 37272 46980 37281
rect 48134 37242 48162 38198
rect 51262 37922 51290 38318
rect 51606 38156 51902 38176
rect 51662 38154 51686 38156
rect 51742 38154 51766 38156
rect 51822 38154 51846 38156
rect 51684 38102 51686 38154
rect 51748 38102 51760 38154
rect 51822 38102 51824 38154
rect 51662 38100 51686 38102
rect 51742 38100 51766 38102
rect 51822 38100 51846 38102
rect 51606 38080 51902 38100
rect 51250 37916 51302 37922
rect 51250 37858 51302 37864
rect 48490 37848 48542 37854
rect 48490 37790 48542 37796
rect 51894 37848 51946 37854
rect 51894 37790 51946 37796
rect 48502 37514 48530 37790
rect 48942 37612 49238 37632
rect 48998 37610 49022 37612
rect 49078 37610 49102 37612
rect 49158 37610 49182 37612
rect 49020 37558 49022 37610
rect 49084 37558 49096 37610
rect 49158 37558 49160 37610
rect 48998 37556 49022 37558
rect 49078 37556 49102 37558
rect 49158 37556 49182 37558
rect 48942 37536 49238 37556
rect 48490 37508 48542 37514
rect 48490 37450 48542 37456
rect 51906 37446 51934 37790
rect 51894 37440 51946 37446
rect 51894 37382 51946 37388
rect 48214 37304 48266 37310
rect 50606 37304 50658 37310
rect 48214 37246 48266 37252
rect 50420 37272 50476 37281
rect 46924 37207 46980 37216
rect 48122 37236 48174 37242
rect 48122 37178 48174 37184
rect 47478 37168 47530 37174
rect 47478 37110 47530 37116
rect 46610 36708 46690 36714
rect 46558 36702 46690 36708
rect 46742 36760 46794 36766
rect 46742 36702 46794 36708
rect 46834 36760 46886 36766
rect 46834 36702 46886 36708
rect 46570 36686 46690 36702
rect 46278 35980 46574 36000
rect 46334 35978 46358 35980
rect 46414 35978 46438 35980
rect 46494 35978 46518 35980
rect 46356 35926 46358 35978
rect 46420 35926 46432 35978
rect 46494 35926 46496 35978
rect 46334 35924 46358 35926
rect 46414 35924 46438 35926
rect 46494 35924 46518 35926
rect 46278 35904 46574 35924
rect 46662 35542 46690 36686
rect 46754 35678 46782 36702
rect 46742 35672 46794 35678
rect 46742 35614 46794 35620
rect 46650 35536 46702 35542
rect 46650 35478 46702 35484
rect 46098 35332 46150 35338
rect 46098 35274 46150 35280
rect 46110 35134 46138 35274
rect 46098 35128 46150 35134
rect 46098 35070 46150 35076
rect 46110 34590 46138 35070
rect 46278 34892 46574 34912
rect 46334 34890 46358 34892
rect 46414 34890 46438 34892
rect 46494 34890 46518 34892
rect 46356 34838 46358 34890
rect 46420 34838 46432 34890
rect 46494 34838 46496 34890
rect 46334 34836 46358 34838
rect 46414 34836 46438 34838
rect 46494 34836 46518 34838
rect 46278 34816 46574 34836
rect 46098 34584 46150 34590
rect 46098 34526 46150 34532
rect 46754 34266 46782 35614
rect 47110 35536 47162 35542
rect 47110 35478 47162 35484
rect 46926 34992 46978 34998
rect 46926 34934 46978 34940
rect 46834 34584 46886 34590
rect 46834 34526 46886 34532
rect 46570 34238 46782 34266
rect 46570 34114 46598 34238
rect 46650 34176 46702 34182
rect 46650 34118 46702 34124
rect 46558 34108 46610 34114
rect 46558 34050 46610 34056
rect 46278 33804 46574 33824
rect 46334 33802 46358 33804
rect 46414 33802 46438 33804
rect 46494 33802 46518 33804
rect 46356 33750 46358 33802
rect 46420 33750 46432 33802
rect 46494 33750 46496 33802
rect 46334 33748 46358 33750
rect 46414 33748 46438 33750
rect 46494 33748 46518 33750
rect 46278 33728 46574 33748
rect 46006 33700 46058 33706
rect 46006 33642 46058 33648
rect 46662 33366 46690 34118
rect 46650 33360 46702 33366
rect 46650 33302 46702 33308
rect 46846 32822 46874 34526
rect 46938 34454 46966 34934
rect 47016 34688 47072 34697
rect 47016 34623 47072 34632
rect 46926 34448 46978 34454
rect 46926 34390 46978 34396
rect 47030 34114 47058 34623
rect 47018 34108 47070 34114
rect 47018 34050 47070 34056
rect 47122 33502 47150 35478
rect 47490 35270 47518 37110
rect 47662 36760 47714 36766
rect 47660 36728 47662 36737
rect 47714 36728 47716 36737
rect 47660 36663 47716 36672
rect 47662 36624 47714 36630
rect 47662 36566 47714 36572
rect 47674 35746 47702 36566
rect 47662 35740 47714 35746
rect 47662 35682 47714 35688
rect 48226 35338 48254 37246
rect 50606 37246 50658 37252
rect 50420 37207 50422 37216
rect 50474 37207 50476 37216
rect 50422 37178 50474 37184
rect 50618 36698 50646 37246
rect 51998 37122 52026 38402
rect 52274 37854 52302 38878
rect 53930 38602 53958 38946
rect 53918 38596 53970 38602
rect 53918 38538 53970 38544
rect 54206 38534 54234 39082
rect 54270 38700 54566 38720
rect 54326 38698 54350 38700
rect 54406 38698 54430 38700
rect 54486 38698 54510 38700
rect 54348 38646 54350 38698
rect 54412 38646 54424 38698
rect 54486 38646 54488 38698
rect 54326 38644 54350 38646
rect 54406 38644 54430 38646
rect 54486 38644 54510 38646
rect 54270 38624 54566 38644
rect 54666 38534 54694 39422
rect 54194 38528 54246 38534
rect 54194 38470 54246 38476
rect 54654 38528 54706 38534
rect 54654 38470 54706 38476
rect 52446 38324 52498 38330
rect 52446 38266 52498 38272
rect 52262 37848 52314 37854
rect 52262 37790 52314 37796
rect 52170 37168 52222 37174
rect 51998 37094 52118 37122
rect 52170 37110 52222 37116
rect 51606 37068 51902 37088
rect 51662 37066 51686 37068
rect 51742 37066 51766 37068
rect 51822 37066 51846 37068
rect 51684 37014 51686 37066
rect 51748 37014 51760 37066
rect 51822 37014 51824 37066
rect 51662 37012 51686 37014
rect 51742 37012 51766 37014
rect 51822 37012 51846 37014
rect 51606 36992 51902 37012
rect 51434 36964 51486 36970
rect 51986 36964 52038 36970
rect 51434 36906 51486 36912
rect 51906 36924 51986 36952
rect 51342 36896 51394 36902
rect 51342 36838 51394 36844
rect 50422 36692 50474 36698
rect 50422 36634 50474 36640
rect 50606 36692 50658 36698
rect 50606 36634 50658 36640
rect 50434 36601 50462 36634
rect 50420 36592 50476 36601
rect 48942 36524 49238 36544
rect 50420 36527 50476 36536
rect 48998 36522 49022 36524
rect 49078 36522 49102 36524
rect 49158 36522 49182 36524
rect 49020 36470 49022 36522
rect 49084 36470 49096 36522
rect 49158 36470 49160 36522
rect 48998 36468 49022 36470
rect 49078 36468 49102 36470
rect 49158 36468 49182 36470
rect 48942 36448 49238 36468
rect 51354 36358 51382 36838
rect 51446 36737 51474 36906
rect 51800 36864 51856 36873
rect 51800 36799 51856 36808
rect 51814 36766 51842 36799
rect 51802 36760 51854 36766
rect 51432 36728 51488 36737
rect 51802 36702 51854 36708
rect 51432 36663 51488 36672
rect 51802 36624 51854 36630
rect 51906 36612 51934 36924
rect 51986 36906 52038 36912
rect 51854 36584 51934 36612
rect 51802 36566 51854 36572
rect 49318 36352 49370 36358
rect 49318 36294 49370 36300
rect 51342 36352 51394 36358
rect 51342 36294 51394 36300
rect 48858 36216 48910 36222
rect 48858 36158 48910 36164
rect 48398 36080 48450 36086
rect 48398 36022 48450 36028
rect 48410 35882 48438 36022
rect 48398 35876 48450 35882
rect 48398 35818 48450 35824
rect 48410 35678 48438 35818
rect 48870 35678 48898 36158
rect 48398 35672 48450 35678
rect 48398 35614 48450 35620
rect 48858 35672 48910 35678
rect 48858 35614 48910 35620
rect 48942 35436 49238 35456
rect 48998 35434 49022 35436
rect 49078 35434 49102 35436
rect 49158 35434 49182 35436
rect 49020 35382 49022 35434
rect 49084 35382 49096 35434
rect 49158 35382 49160 35434
rect 48998 35380 49022 35382
rect 49078 35380 49102 35382
rect 49158 35380 49182 35382
rect 48942 35360 49238 35380
rect 49330 35338 49358 36294
rect 51354 36222 51382 36294
rect 51618 36284 51670 36290
rect 51618 36226 51670 36232
rect 51342 36216 51394 36222
rect 51342 36158 51394 36164
rect 51630 36154 51658 36226
rect 51906 36222 51934 36584
rect 52090 36222 52118 37094
rect 52182 36970 52210 37110
rect 52170 36964 52222 36970
rect 52170 36906 52222 36912
rect 52274 36358 52302 37790
rect 52354 37712 52406 37718
rect 52354 37654 52406 37660
rect 52366 37378 52394 37654
rect 52354 37372 52406 37378
rect 52354 37314 52406 37320
rect 52354 37168 52406 37174
rect 52354 37110 52406 37116
rect 52366 36970 52394 37110
rect 52354 36964 52406 36970
rect 52354 36906 52406 36912
rect 52366 36873 52394 36906
rect 52352 36864 52408 36873
rect 52458 36834 52486 38266
rect 53918 38256 53970 38262
rect 53918 38198 53970 38204
rect 53930 37990 53958 38198
rect 53918 37984 53970 37990
rect 53918 37926 53970 37932
rect 54746 37848 54798 37854
rect 54746 37790 54798 37796
rect 54270 37612 54566 37632
rect 54326 37610 54350 37612
rect 54406 37610 54430 37612
rect 54486 37610 54510 37612
rect 54348 37558 54350 37610
rect 54412 37558 54424 37610
rect 54486 37558 54488 37610
rect 54326 37556 54350 37558
rect 54406 37556 54430 37558
rect 54486 37556 54510 37558
rect 54270 37536 54566 37556
rect 54758 37310 54786 37790
rect 54850 37310 54878 40222
rect 55850 40170 55902 40176
rect 55206 40024 55258 40030
rect 55034 39984 55206 40012
rect 55034 39894 55062 39984
rect 55206 39966 55258 39972
rect 55390 40024 55442 40030
rect 55390 39966 55442 39972
rect 55402 39894 55430 39966
rect 55022 39888 55074 39894
rect 55022 39830 55074 39836
rect 55390 39888 55442 39894
rect 55390 39830 55442 39836
rect 55850 39888 55902 39894
rect 55850 39830 55902 39836
rect 55034 37718 55062 39830
rect 55298 39684 55350 39690
rect 55298 39626 55350 39632
rect 55206 39480 55258 39486
rect 55310 39468 55338 39626
rect 55390 39548 55442 39554
rect 55390 39490 55442 39496
rect 55258 39440 55338 39468
rect 55206 39422 55258 39428
rect 55114 39140 55166 39146
rect 55114 39082 55166 39088
rect 55126 39010 55154 39082
rect 55402 39078 55430 39490
rect 55862 39146 55890 39830
rect 56690 39690 56718 40510
rect 56678 39684 56730 39690
rect 56678 39626 56730 39632
rect 56782 39418 56810 40646
rect 57322 40636 57374 40642
rect 57322 40578 57374 40584
rect 56862 40432 56914 40438
rect 56862 40374 56914 40380
rect 56874 40030 56902 40374
rect 56934 40332 57230 40352
rect 56990 40330 57014 40332
rect 57070 40330 57094 40332
rect 57150 40330 57174 40332
rect 57012 40278 57014 40330
rect 57076 40278 57088 40330
rect 57150 40278 57152 40330
rect 56990 40276 57014 40278
rect 57070 40276 57094 40278
rect 57150 40276 57174 40278
rect 56934 40256 57230 40276
rect 57334 40166 57362 40578
rect 57322 40160 57374 40166
rect 57322 40102 57374 40108
rect 56862 40024 56914 40030
rect 56862 39966 56914 39972
rect 57426 39978 57454 43312
rect 58058 40976 58110 40982
rect 58058 40918 58110 40924
rect 58070 40642 58098 40918
rect 58058 40636 58110 40642
rect 58058 40578 58110 40584
rect 57426 39950 57730 39978
rect 57322 39684 57374 39690
rect 57322 39626 57374 39632
rect 56862 39548 56914 39554
rect 56862 39490 56914 39496
rect 56586 39412 56638 39418
rect 56586 39354 56638 39360
rect 56770 39412 56822 39418
rect 56770 39354 56822 39360
rect 55850 39140 55902 39146
rect 55850 39082 55902 39088
rect 55390 39072 55442 39078
rect 55482 39072 55534 39078
rect 55390 39014 55442 39020
rect 55480 39040 55482 39049
rect 55534 39040 55536 39049
rect 55114 39004 55166 39010
rect 55114 38946 55166 38952
rect 55402 38534 55430 39014
rect 55480 38975 55536 38984
rect 55390 38528 55442 38534
rect 55390 38470 55442 38476
rect 55206 38460 55258 38466
rect 55206 38402 55258 38408
rect 55218 37938 55246 38402
rect 55218 37910 55614 37938
rect 55206 37848 55258 37854
rect 55206 37790 55258 37796
rect 55022 37712 55074 37718
rect 55022 37654 55074 37660
rect 54930 37440 54982 37446
rect 54930 37382 54982 37388
rect 54746 37304 54798 37310
rect 52536 37272 52592 37281
rect 54746 37246 54798 37252
rect 54838 37304 54890 37310
rect 54838 37246 54890 37252
rect 52536 37207 52592 37216
rect 52550 37174 52578 37207
rect 52538 37168 52590 37174
rect 52538 37110 52590 37116
rect 54942 36970 54970 37382
rect 55034 37378 55062 37654
rect 55218 37446 55246 37790
rect 55298 37780 55350 37786
rect 55298 37722 55350 37728
rect 55310 37514 55338 37722
rect 55298 37508 55350 37514
rect 55298 37450 55350 37456
rect 55206 37440 55258 37446
rect 55206 37382 55258 37388
rect 55586 37378 55614 37910
rect 55022 37372 55074 37378
rect 55022 37314 55074 37320
rect 55482 37372 55534 37378
rect 55482 37314 55534 37320
rect 55574 37372 55626 37378
rect 55574 37314 55626 37320
rect 54930 36964 54982 36970
rect 54930 36906 54982 36912
rect 55494 36902 55522 37314
rect 55482 36896 55534 36902
rect 55482 36838 55534 36844
rect 52352 36799 52408 36808
rect 52446 36828 52498 36834
rect 52446 36770 52498 36776
rect 53456 36728 53512 36737
rect 52722 36692 52774 36698
rect 53456 36663 53512 36672
rect 52722 36634 52774 36640
rect 52734 36601 52762 36634
rect 53470 36630 53498 36663
rect 53366 36624 53418 36630
rect 52720 36592 52776 36601
rect 53366 36566 53418 36572
rect 53458 36624 53510 36630
rect 53458 36566 53510 36572
rect 52720 36527 52776 36536
rect 52262 36352 52314 36358
rect 52262 36294 52314 36300
rect 53378 36290 53406 36566
rect 54270 36524 54566 36544
rect 54326 36522 54350 36524
rect 54406 36522 54430 36524
rect 54486 36522 54510 36524
rect 54348 36470 54350 36522
rect 54412 36470 54424 36522
rect 54486 36470 54488 36522
rect 54326 36468 54350 36470
rect 54406 36468 54430 36470
rect 54486 36468 54510 36470
rect 54270 36448 54566 36468
rect 52722 36284 52774 36290
rect 52722 36226 52774 36232
rect 53366 36284 53418 36290
rect 53366 36226 53418 36232
rect 51894 36216 51946 36222
rect 51894 36158 51946 36164
rect 52078 36216 52130 36222
rect 52078 36158 52130 36164
rect 51526 36148 51578 36154
rect 51526 36090 51578 36096
rect 51618 36148 51670 36154
rect 51618 36090 51670 36096
rect 51538 35785 51566 36090
rect 51606 35980 51902 36000
rect 51662 35978 51686 35980
rect 51742 35978 51766 35980
rect 51822 35978 51846 35980
rect 51684 35926 51686 35978
rect 51748 35926 51760 35978
rect 51822 35926 51824 35978
rect 51662 35924 51686 35926
rect 51742 35924 51766 35926
rect 51822 35924 51846 35926
rect 51606 35904 51902 35924
rect 51524 35776 51580 35785
rect 51524 35711 51580 35720
rect 49410 35604 49462 35610
rect 49410 35546 49462 35552
rect 51986 35604 52038 35610
rect 51986 35546 52038 35552
rect 49422 35338 49450 35546
rect 51894 35536 51946 35542
rect 51894 35478 51946 35484
rect 48214 35332 48266 35338
rect 48214 35274 48266 35280
rect 49318 35332 49370 35338
rect 49318 35274 49370 35280
rect 49410 35332 49462 35338
rect 49410 35274 49462 35280
rect 47478 35264 47530 35270
rect 47478 35206 47530 35212
rect 47570 35196 47622 35202
rect 47570 35138 47622 35144
rect 47582 34522 47610 35138
rect 48226 34726 48254 35274
rect 49330 35202 49358 35274
rect 51906 35202 51934 35478
rect 49318 35196 49370 35202
rect 49318 35138 49370 35144
rect 51894 35196 51946 35202
rect 51894 35138 51946 35144
rect 51606 34892 51902 34912
rect 51662 34890 51686 34892
rect 51742 34890 51766 34892
rect 51822 34890 51846 34892
rect 51684 34838 51686 34890
rect 51748 34838 51760 34890
rect 51822 34838 51824 34890
rect 51662 34836 51686 34838
rect 51742 34836 51766 34838
rect 51822 34836 51846 34838
rect 51606 34816 51902 34836
rect 48214 34720 48266 34726
rect 48214 34662 48266 34668
rect 51894 34720 51946 34726
rect 51998 34674 52026 35546
rect 52090 35202 52118 36158
rect 52734 36086 52762 36226
rect 52354 36080 52406 36086
rect 52354 36022 52406 36028
rect 52722 36080 52774 36086
rect 52722 36022 52774 36028
rect 52366 35542 52394 36022
rect 52354 35536 52406 35542
rect 52354 35478 52406 35484
rect 52630 35536 52682 35542
rect 52630 35478 52682 35484
rect 52078 35196 52130 35202
rect 52078 35138 52130 35144
rect 52642 34998 52670 35478
rect 52734 35134 52762 36022
rect 53182 35672 53234 35678
rect 53182 35614 53234 35620
rect 52722 35128 52774 35134
rect 52722 35070 52774 35076
rect 52734 34998 52762 35070
rect 52630 34992 52682 34998
rect 52630 34934 52682 34940
rect 52722 34992 52774 34998
rect 52722 34934 52774 34940
rect 51946 34668 52026 34674
rect 51894 34662 52026 34668
rect 47662 34652 47714 34658
rect 51906 34646 52026 34662
rect 47662 34594 47714 34600
rect 47570 34516 47622 34522
rect 47570 34458 47622 34464
rect 47674 34182 47702 34594
rect 51526 34448 51578 34454
rect 51526 34390 51578 34396
rect 48942 34348 49238 34368
rect 48998 34346 49022 34348
rect 49078 34346 49102 34348
rect 49158 34346 49182 34348
rect 49020 34294 49022 34346
rect 49084 34294 49096 34346
rect 49158 34294 49160 34346
rect 48998 34292 49022 34294
rect 49078 34292 49102 34294
rect 49158 34292 49182 34294
rect 48942 34272 49238 34292
rect 51538 34250 51566 34390
rect 51526 34244 51578 34250
rect 51526 34186 51578 34192
rect 47662 34176 47714 34182
rect 47662 34118 47714 34124
rect 52446 34108 52498 34114
rect 52446 34050 52498 34056
rect 52458 33994 52486 34050
rect 52458 33966 52578 33994
rect 47202 33904 47254 33910
rect 47202 33846 47254 33852
rect 47110 33496 47162 33502
rect 47110 33438 47162 33444
rect 46926 33428 46978 33434
rect 46926 33370 46978 33376
rect 46742 32816 46794 32822
rect 46740 32784 46742 32793
rect 46834 32816 46886 32822
rect 46794 32784 46796 32793
rect 46278 32716 46574 32736
rect 46834 32758 46886 32764
rect 46740 32719 46796 32728
rect 46334 32714 46358 32716
rect 46414 32714 46438 32716
rect 46494 32714 46518 32716
rect 46356 32662 46358 32714
rect 46420 32662 46432 32714
rect 46494 32662 46496 32714
rect 46334 32660 46358 32662
rect 46414 32660 46438 32662
rect 46494 32660 46518 32662
rect 46278 32640 46574 32660
rect 46742 32408 46794 32414
rect 46742 32350 46794 32356
rect 46466 32340 46518 32346
rect 46466 32282 46518 32288
rect 46478 32249 46506 32282
rect 46464 32240 46520 32249
rect 46464 32175 46520 32184
rect 46754 31938 46782 32350
rect 46938 32074 46966 33370
rect 47018 33360 47070 33366
rect 47122 33337 47150 33438
rect 47018 33302 47070 33308
rect 47108 33328 47164 33337
rect 47030 32414 47058 33302
rect 47108 33263 47164 33272
rect 47214 33026 47242 33846
rect 51606 33804 51902 33824
rect 51662 33802 51686 33804
rect 51742 33802 51766 33804
rect 51822 33802 51846 33804
rect 51684 33750 51686 33802
rect 51748 33750 51760 33802
rect 51822 33750 51824 33802
rect 51662 33748 51686 33750
rect 51742 33748 51766 33750
rect 51822 33748 51846 33750
rect 51606 33728 51902 33748
rect 49318 33700 49370 33706
rect 49318 33642 49370 33648
rect 48858 33496 48910 33502
rect 48858 33438 48910 33444
rect 47478 33428 47530 33434
rect 47478 33370 47530 33376
rect 47490 33094 47518 33370
rect 47478 33088 47530 33094
rect 47478 33030 47530 33036
rect 47202 33020 47254 33026
rect 47202 32962 47254 32968
rect 47294 32952 47346 32958
rect 47292 32920 47294 32929
rect 47346 32920 47348 32929
rect 47292 32855 47348 32864
rect 47570 32816 47622 32822
rect 47384 32784 47440 32793
rect 47384 32719 47440 32728
rect 47568 32784 47570 32793
rect 47662 32816 47714 32822
rect 47622 32784 47624 32793
rect 47662 32758 47714 32764
rect 48582 32816 48634 32822
rect 48582 32758 48634 32764
rect 47568 32719 47624 32728
rect 47018 32408 47070 32414
rect 47202 32408 47254 32414
rect 47018 32350 47070 32356
rect 47200 32376 47202 32385
rect 47254 32376 47256 32385
rect 46926 32068 46978 32074
rect 46926 32010 46978 32016
rect 44718 31932 44770 31938
rect 44718 31874 44770 31880
rect 45178 31932 45230 31938
rect 45178 31874 45230 31880
rect 46098 31932 46150 31938
rect 46098 31874 46150 31880
rect 46742 31932 46794 31938
rect 46742 31874 46794 31880
rect 44730 31462 44758 31874
rect 46110 31734 46138 31874
rect 46098 31728 46150 31734
rect 46098 31670 46150 31676
rect 44718 31456 44770 31462
rect 44718 31398 44770 31404
rect 43614 30844 43666 30850
rect 43614 30786 43666 30792
rect 44442 30844 44494 30850
rect 44442 30786 44494 30792
rect 44626 30844 44678 30850
rect 44626 30786 44678 30792
rect 43442 30158 43562 30186
rect 43442 29762 43470 30158
rect 43626 30084 43654 30786
rect 46110 30714 46138 31670
rect 46278 31628 46574 31648
rect 46334 31626 46358 31628
rect 46414 31626 46438 31628
rect 46494 31626 46518 31628
rect 46356 31574 46358 31626
rect 46420 31574 46432 31626
rect 46494 31574 46496 31626
rect 46334 31572 46358 31574
rect 46414 31572 46438 31574
rect 46494 31572 46518 31574
rect 46278 31552 46574 31572
rect 46464 31424 46520 31433
rect 46464 31359 46466 31368
rect 46518 31359 46520 31368
rect 46466 31330 46518 31336
rect 46938 31326 46966 32010
rect 47030 31530 47058 32350
rect 47200 32311 47256 32320
rect 47018 31524 47070 31530
rect 47018 31466 47070 31472
rect 46926 31320 46978 31326
rect 46926 31262 46978 31268
rect 47398 31190 47426 32719
rect 47478 32408 47530 32414
rect 47674 32396 47702 32758
rect 48594 32550 48622 32758
rect 48398 32544 48450 32550
rect 48396 32512 48398 32521
rect 48582 32544 48634 32550
rect 48450 32512 48452 32521
rect 48030 32476 48082 32482
rect 48582 32486 48634 32492
rect 48870 32482 48898 33438
rect 48942 33260 49238 33280
rect 48998 33258 49022 33260
rect 49078 33258 49102 33260
rect 49158 33258 49182 33260
rect 49020 33206 49022 33258
rect 49084 33206 49096 33258
rect 49158 33206 49160 33258
rect 48998 33204 49022 33206
rect 49078 33204 49102 33206
rect 49158 33204 49182 33206
rect 48942 33184 49238 33204
rect 49330 33162 49358 33642
rect 52550 33570 52578 33966
rect 52538 33564 52590 33570
rect 52538 33506 52590 33512
rect 52262 33496 52314 33502
rect 52262 33438 52314 33444
rect 49686 33428 49738 33434
rect 49686 33370 49738 33376
rect 49318 33156 49370 33162
rect 49318 33098 49370 33104
rect 49698 33026 49726 33370
rect 49686 33020 49738 33026
rect 49686 32962 49738 32968
rect 49698 32482 49726 32962
rect 51434 32952 51486 32958
rect 51434 32894 51486 32900
rect 50606 32884 50658 32890
rect 50606 32826 50658 32832
rect 50618 32550 50646 32826
rect 50606 32544 50658 32550
rect 50606 32486 50658 32492
rect 48396 32447 48452 32456
rect 48858 32476 48910 32482
rect 48030 32418 48082 32424
rect 48858 32418 48910 32424
rect 49686 32476 49738 32482
rect 49686 32418 49738 32424
rect 47530 32368 47702 32396
rect 47478 32350 47530 32356
rect 47490 32006 47518 32350
rect 47570 32272 47622 32278
rect 47568 32240 47570 32249
rect 47622 32240 47624 32249
rect 47674 32226 47702 32368
rect 47936 32376 47992 32385
rect 47936 32311 47992 32320
rect 47950 32278 47978 32311
rect 48042 32278 48070 32418
rect 51066 32408 51118 32414
rect 51066 32350 51118 32356
rect 48398 32340 48450 32346
rect 48398 32282 48450 32288
rect 47754 32272 47806 32278
rect 47674 32220 47754 32226
rect 47674 32214 47806 32220
rect 47938 32272 47990 32278
rect 47938 32214 47990 32220
rect 48030 32272 48082 32278
rect 48030 32214 48082 32220
rect 47674 32198 47794 32214
rect 47568 32175 47624 32184
rect 47478 32000 47530 32006
rect 47478 31942 47530 31948
rect 47662 31864 47714 31870
rect 47662 31806 47714 31812
rect 47386 31184 47438 31190
rect 47386 31126 47438 31132
rect 47674 30782 47702 31806
rect 47662 30776 47714 30782
rect 47662 30718 47714 30724
rect 46098 30708 46150 30714
rect 46098 30650 46150 30656
rect 45454 30640 45506 30646
rect 45454 30582 45506 30588
rect 43706 30368 43758 30374
rect 43706 30310 43758 30316
rect 43982 30368 44034 30374
rect 43982 30310 44034 30316
rect 43718 30238 43746 30310
rect 43706 30232 43758 30238
rect 43706 30174 43758 30180
rect 43534 30056 43654 30084
rect 43534 29762 43562 30056
rect 43614 29996 43910 30016
rect 43670 29994 43694 29996
rect 43750 29994 43774 29996
rect 43830 29994 43854 29996
rect 43692 29942 43694 29994
rect 43756 29942 43768 29994
rect 43830 29942 43832 29994
rect 43670 29940 43694 29942
rect 43750 29940 43774 29942
rect 43830 29940 43854 29942
rect 43614 29920 43910 29940
rect 43994 29898 44022 30310
rect 44074 30164 44126 30170
rect 44074 30106 44126 30112
rect 43982 29892 44034 29898
rect 43982 29834 44034 29840
rect 43430 29756 43482 29762
rect 43430 29698 43482 29704
rect 43522 29756 43574 29762
rect 43522 29698 43574 29704
rect 43430 29008 43482 29014
rect 43430 28950 43482 28956
rect 43442 28062 43470 28950
rect 43534 28674 43562 29698
rect 44086 29354 44114 30106
rect 44166 30096 44218 30102
rect 44166 30038 44218 30044
rect 45362 30096 45414 30102
rect 45362 30038 45414 30044
rect 44178 29898 44206 30038
rect 44166 29892 44218 29898
rect 44166 29834 44218 29840
rect 44074 29348 44126 29354
rect 44074 29290 44126 29296
rect 43614 28908 43910 28928
rect 43670 28906 43694 28908
rect 43750 28906 43774 28908
rect 43830 28906 43854 28908
rect 43692 28854 43694 28906
rect 43756 28854 43768 28906
rect 43830 28854 43832 28906
rect 43670 28852 43694 28854
rect 43750 28852 43774 28854
rect 43830 28852 43854 28854
rect 43614 28832 43910 28852
rect 43798 28736 43850 28742
rect 43798 28678 43850 28684
rect 43522 28668 43574 28674
rect 43522 28610 43574 28616
rect 43810 28062 43838 28678
rect 43430 28056 43482 28062
rect 43798 28056 43850 28062
rect 43482 28016 43562 28044
rect 43430 27998 43482 28004
rect 43534 27722 43562 28016
rect 43798 27998 43850 28004
rect 43614 27820 43910 27840
rect 43670 27818 43694 27820
rect 43750 27818 43774 27820
rect 43830 27818 43854 27820
rect 43692 27766 43694 27818
rect 43756 27766 43768 27818
rect 43830 27766 43832 27818
rect 43670 27764 43694 27766
rect 43750 27764 43774 27766
rect 43830 27764 43854 27766
rect 43614 27744 43910 27764
rect 43522 27716 43574 27722
rect 43522 27658 43574 27664
rect 43534 27586 43562 27658
rect 43522 27580 43574 27586
rect 43522 27522 43574 27528
rect 43706 27580 43758 27586
rect 43706 27522 43758 27528
rect 43718 27382 43746 27522
rect 43706 27376 43758 27382
rect 43706 27318 43758 27324
rect 44178 27042 44206 29834
rect 44994 29280 45046 29286
rect 44994 29222 45046 29228
rect 45006 28198 45034 29222
rect 45374 29082 45402 30038
rect 45466 29218 45494 30582
rect 46278 30540 46574 30560
rect 46334 30538 46358 30540
rect 46414 30538 46438 30540
rect 46494 30538 46518 30540
rect 46356 30486 46358 30538
rect 46420 30486 46432 30538
rect 46494 30486 46496 30538
rect 46334 30484 46358 30486
rect 46414 30484 46438 30486
rect 46494 30484 46518 30486
rect 46278 30464 46574 30484
rect 47846 30232 47898 30238
rect 47846 30174 47898 30180
rect 47858 29558 47886 30174
rect 46834 29552 46886 29558
rect 46834 29494 46886 29500
rect 47846 29552 47898 29558
rect 47846 29494 47898 29500
rect 46278 29452 46574 29472
rect 46334 29450 46358 29452
rect 46414 29450 46438 29452
rect 46494 29450 46518 29452
rect 46356 29398 46358 29450
rect 46420 29398 46432 29450
rect 46494 29398 46496 29450
rect 46334 29396 46358 29398
rect 46414 29396 46438 29398
rect 46494 29396 46518 29398
rect 46278 29376 46574 29396
rect 45822 29280 45874 29286
rect 45822 29222 45874 29228
rect 46006 29280 46058 29286
rect 46006 29222 46058 29228
rect 45454 29212 45506 29218
rect 45454 29154 45506 29160
rect 45362 29076 45414 29082
rect 45362 29018 45414 29024
rect 45546 29076 45598 29082
rect 45546 29018 45598 29024
rect 45558 28810 45586 29018
rect 45546 28804 45598 28810
rect 45546 28746 45598 28752
rect 45270 28464 45322 28470
rect 45270 28406 45322 28412
rect 44994 28192 45046 28198
rect 44994 28134 45046 28140
rect 44442 28056 44494 28062
rect 44362 28016 44442 28044
rect 44362 27722 44390 28016
rect 44442 27998 44494 28004
rect 44350 27716 44402 27722
rect 44350 27658 44402 27664
rect 44362 27450 44390 27658
rect 45282 27450 45310 28406
rect 45834 28130 45862 29222
rect 46018 29121 46046 29222
rect 46846 29218 46874 29494
rect 47294 29348 47346 29354
rect 47294 29290 47346 29296
rect 46834 29212 46886 29218
rect 46834 29154 46886 29160
rect 47306 29150 47334 29290
rect 47294 29144 47346 29150
rect 46004 29112 46060 29121
rect 47294 29086 47346 29092
rect 46004 29047 46060 29056
rect 47754 28464 47806 28470
rect 47754 28406 47806 28412
rect 46278 28364 46574 28384
rect 46334 28362 46358 28364
rect 46414 28362 46438 28364
rect 46494 28362 46518 28364
rect 46356 28310 46358 28362
rect 46420 28310 46432 28362
rect 46494 28310 46496 28362
rect 46334 28308 46358 28310
rect 46414 28308 46438 28310
rect 46494 28308 46518 28310
rect 46278 28288 46574 28308
rect 46098 28260 46150 28266
rect 46098 28202 46150 28208
rect 45822 28124 45874 28130
rect 45822 28066 45874 28072
rect 45546 27580 45598 27586
rect 45546 27522 45598 27528
rect 45362 27512 45414 27518
rect 45362 27454 45414 27460
rect 44350 27444 44402 27450
rect 44350 27386 44402 27392
rect 45270 27444 45322 27450
rect 45270 27386 45322 27392
rect 44362 27042 44390 27386
rect 45374 27178 45402 27454
rect 45558 27382 45586 27522
rect 45546 27376 45598 27382
rect 45546 27318 45598 27324
rect 45362 27172 45414 27178
rect 45362 27114 45414 27120
rect 44166 27036 44218 27042
rect 44166 26978 44218 26984
rect 44350 27036 44402 27042
rect 44350 26978 44402 26984
rect 43614 26732 43910 26752
rect 43670 26730 43694 26732
rect 43750 26730 43774 26732
rect 43830 26730 43854 26732
rect 43692 26678 43694 26730
rect 43756 26678 43768 26730
rect 43830 26678 43832 26730
rect 43670 26676 43694 26678
rect 43750 26676 43774 26678
rect 43830 26676 43854 26678
rect 43614 26656 43910 26676
rect 46110 23613 46138 28202
rect 46282 27988 46334 27994
rect 46282 27930 46334 27936
rect 46294 27654 46322 27930
rect 46282 27648 46334 27654
rect 46282 27590 46334 27596
rect 47766 27586 47794 28406
rect 47858 28062 47886 29494
rect 47950 28606 47978 32214
rect 48410 31938 48438 32282
rect 48942 32172 49238 32192
rect 48998 32170 49022 32172
rect 49078 32170 49102 32172
rect 49158 32170 49182 32172
rect 49020 32118 49022 32170
rect 49084 32118 49096 32170
rect 49158 32118 49160 32170
rect 48998 32116 49022 32118
rect 49078 32116 49102 32118
rect 49158 32116 49182 32118
rect 48942 32096 49238 32116
rect 48398 31932 48450 31938
rect 48398 31874 48450 31880
rect 50790 31932 50842 31938
rect 50790 31874 50842 31880
rect 50802 31716 50830 31874
rect 51078 31870 51106 32350
rect 51066 31864 51118 31870
rect 51066 31806 51118 31812
rect 50974 31728 51026 31734
rect 50802 31688 50974 31716
rect 50974 31670 51026 31676
rect 50882 31456 50934 31462
rect 50882 31398 50934 31404
rect 48858 31388 48910 31394
rect 48858 31330 48910 31336
rect 48870 30782 48898 31330
rect 50894 31190 50922 31398
rect 51078 31258 51106 31806
rect 51446 31326 51474 32894
rect 51606 32716 51902 32736
rect 51662 32714 51686 32716
rect 51742 32714 51766 32716
rect 51822 32714 51846 32716
rect 51684 32662 51686 32714
rect 51748 32662 51760 32714
rect 51822 32662 51824 32714
rect 51662 32660 51686 32662
rect 51742 32660 51766 32662
rect 51822 32660 51846 32662
rect 51606 32640 51902 32660
rect 52274 32550 52302 33438
rect 52262 32544 52314 32550
rect 52262 32486 52314 32492
rect 51526 32408 51578 32414
rect 51526 32350 51578 32356
rect 51986 32408 52038 32414
rect 51986 32350 52038 32356
rect 51538 31530 51566 32350
rect 51998 31734 52026 32350
rect 52642 32278 52670 34934
rect 52630 32272 52682 32278
rect 52630 32214 52682 32220
rect 52734 31734 52762 34934
rect 53194 34726 53222 35614
rect 53274 35536 53326 35542
rect 53274 35478 53326 35484
rect 52814 34720 52866 34726
rect 52814 34662 52866 34668
rect 53182 34720 53234 34726
rect 53182 34662 53234 34668
rect 52826 34250 52854 34662
rect 52814 34244 52866 34250
rect 52814 34186 52866 34192
rect 52814 34108 52866 34114
rect 52814 34050 52866 34056
rect 52826 33910 52854 34050
rect 52814 33904 52866 33910
rect 52814 33846 52866 33852
rect 52906 33904 52958 33910
rect 52906 33846 52958 33852
rect 52918 33502 52946 33846
rect 52906 33496 52958 33502
rect 52906 33438 52958 33444
rect 52906 32816 52958 32822
rect 52906 32758 52958 32764
rect 52812 32512 52868 32521
rect 52812 32447 52868 32456
rect 51986 31728 52038 31734
rect 51986 31670 52038 31676
rect 52722 31728 52774 31734
rect 52722 31670 52774 31676
rect 51606 31628 51902 31648
rect 51662 31626 51686 31628
rect 51742 31626 51766 31628
rect 51822 31626 51846 31628
rect 51684 31574 51686 31626
rect 51748 31574 51760 31626
rect 51822 31574 51824 31626
rect 51662 31572 51686 31574
rect 51742 31572 51766 31574
rect 51822 31572 51846 31574
rect 51606 31552 51902 31572
rect 51526 31524 51578 31530
rect 51526 31466 51578 31472
rect 51434 31320 51486 31326
rect 51434 31262 51486 31268
rect 51066 31252 51118 31258
rect 51066 31194 51118 31200
rect 49778 31184 49830 31190
rect 49778 31126 49830 31132
rect 50882 31184 50934 31190
rect 50882 31126 50934 31132
rect 48942 31084 49238 31104
rect 48998 31082 49022 31084
rect 49078 31082 49102 31084
rect 49158 31082 49182 31084
rect 49020 31030 49022 31082
rect 49084 31030 49096 31082
rect 49158 31030 49160 31082
rect 48998 31028 49022 31030
rect 49078 31028 49102 31030
rect 49158 31028 49182 31030
rect 48942 31008 49238 31028
rect 48858 30776 48910 30782
rect 48858 30718 48910 30724
rect 48306 30640 48358 30646
rect 48306 30582 48358 30588
rect 48674 30640 48726 30646
rect 48674 30582 48726 30588
rect 49410 30640 49462 30646
rect 49410 30582 49462 30588
rect 48318 29354 48346 30582
rect 48686 30442 48714 30582
rect 48674 30436 48726 30442
rect 48674 30378 48726 30384
rect 48858 30164 48910 30170
rect 48858 30106 48910 30112
rect 48398 29552 48450 29558
rect 48398 29494 48450 29500
rect 48410 29354 48438 29494
rect 48122 29348 48174 29354
rect 48122 29290 48174 29296
rect 48306 29348 48358 29354
rect 48306 29290 48358 29296
rect 48398 29348 48450 29354
rect 48398 29290 48450 29296
rect 48582 29348 48634 29354
rect 48582 29290 48634 29296
rect 48134 29234 48162 29290
rect 48134 29218 48346 29234
rect 48134 29212 48358 29218
rect 48134 29206 48306 29212
rect 48306 29154 48358 29160
rect 48490 29212 48542 29218
rect 48490 29154 48542 29160
rect 47938 28600 47990 28606
rect 47938 28542 47990 28548
rect 48306 28124 48358 28130
rect 48306 28066 48358 28072
rect 47846 28056 47898 28062
rect 47846 27998 47898 28004
rect 48212 28024 48268 28033
rect 48212 27959 48268 27968
rect 48226 27926 48254 27959
rect 48214 27920 48266 27926
rect 48214 27862 48266 27868
rect 48214 27716 48266 27722
rect 48318 27704 48346 28066
rect 48398 27920 48450 27926
rect 48398 27862 48450 27868
rect 48266 27676 48346 27704
rect 48214 27658 48266 27664
rect 48410 27586 48438 27862
rect 48502 27654 48530 29154
rect 48490 27648 48542 27654
rect 48490 27590 48542 27596
rect 47754 27580 47806 27586
rect 47754 27522 47806 27528
rect 48398 27580 48450 27586
rect 48398 27522 48450 27528
rect 48396 27480 48452 27489
rect 48396 27415 48452 27424
rect 46278 27276 46574 27296
rect 46334 27274 46358 27276
rect 46414 27274 46438 27276
rect 46494 27274 46518 27276
rect 46356 27222 46358 27274
rect 46420 27222 46432 27274
rect 46494 27222 46496 27274
rect 46334 27220 46358 27222
rect 46414 27220 46438 27222
rect 46494 27220 46518 27222
rect 46278 27200 46574 27220
rect 48410 27042 48438 27415
rect 48398 27036 48450 27042
rect 48398 26978 48450 26984
rect 48594 26974 48622 29290
rect 48674 29144 48726 29150
rect 48674 29086 48726 29092
rect 48686 29014 48714 29086
rect 48674 29008 48726 29014
rect 48674 28950 48726 28956
rect 48686 27382 48714 28950
rect 48870 28470 48898 30106
rect 48942 29996 49238 30016
rect 48998 29994 49022 29996
rect 49078 29994 49102 29996
rect 49158 29994 49182 29996
rect 49020 29942 49022 29994
rect 49084 29942 49096 29994
rect 49158 29942 49160 29994
rect 48998 29940 49022 29942
rect 49078 29940 49102 29942
rect 49158 29940 49182 29942
rect 48942 29920 49238 29940
rect 49422 29898 49450 30582
rect 49410 29892 49462 29898
rect 49410 29834 49462 29840
rect 49686 29008 49738 29014
rect 49686 28950 49738 28956
rect 48942 28908 49238 28928
rect 48998 28906 49022 28908
rect 49078 28906 49102 28908
rect 49158 28906 49182 28908
rect 49020 28854 49022 28906
rect 49084 28854 49096 28906
rect 49158 28854 49160 28906
rect 48998 28852 49022 28854
rect 49078 28852 49102 28854
rect 49158 28852 49182 28854
rect 48942 28832 49238 28852
rect 49698 28674 49726 28950
rect 49318 28668 49370 28674
rect 49318 28610 49370 28616
rect 49686 28668 49738 28674
rect 49686 28610 49738 28616
rect 48858 28464 48910 28470
rect 48858 28406 48910 28412
rect 49330 28266 49358 28610
rect 49318 28260 49370 28266
rect 49318 28202 49370 28208
rect 48942 27820 49238 27840
rect 48998 27818 49022 27820
rect 49078 27818 49102 27820
rect 49158 27818 49182 27820
rect 49020 27766 49022 27818
rect 49084 27766 49096 27818
rect 49158 27766 49160 27818
rect 48998 27764 49022 27766
rect 49078 27764 49102 27766
rect 49158 27764 49182 27766
rect 48942 27744 49238 27764
rect 48674 27376 48726 27382
rect 48674 27318 48726 27324
rect 48686 27178 48714 27318
rect 48674 27172 48726 27178
rect 48674 27114 48726 27120
rect 48582 26968 48634 26974
rect 48582 26910 48634 26916
rect 49330 26906 49358 28202
rect 49790 27586 49818 31126
rect 50698 30776 50750 30782
rect 50698 30718 50750 30724
rect 50710 29762 50738 30718
rect 50790 29824 50842 29830
rect 50790 29766 50842 29772
rect 50698 29756 50750 29762
rect 50698 29698 50750 29704
rect 50802 29506 50830 29766
rect 50894 29762 50922 31126
rect 51606 30540 51902 30560
rect 51662 30538 51686 30540
rect 51742 30538 51766 30540
rect 51822 30538 51846 30540
rect 51684 30486 51686 30538
rect 51748 30486 51760 30538
rect 51822 30486 51824 30538
rect 51662 30484 51686 30486
rect 51742 30484 51766 30486
rect 51822 30484 51846 30486
rect 51606 30464 51902 30484
rect 51998 30238 52026 31670
rect 52170 30912 52222 30918
rect 52168 30880 52170 30889
rect 52222 30880 52224 30889
rect 52168 30815 52224 30824
rect 52826 30782 52854 32447
rect 52918 30782 52946 32758
rect 53194 32550 53222 34662
rect 53286 34658 53314 35478
rect 53378 35202 53406 36226
rect 54194 35876 54246 35882
rect 54194 35818 54246 35824
rect 53458 35672 53510 35678
rect 53510 35620 54050 35626
rect 53458 35614 54050 35620
rect 53470 35598 54050 35614
rect 54022 35542 54050 35598
rect 54206 35542 54234 35818
rect 55586 35814 55614 37314
rect 55574 35808 55626 35814
rect 55574 35750 55626 35756
rect 54654 35604 54706 35610
rect 54654 35546 54706 35552
rect 54010 35536 54062 35542
rect 54010 35478 54062 35484
rect 54194 35536 54246 35542
rect 54194 35478 54246 35484
rect 53366 35196 53418 35202
rect 53366 35138 53418 35144
rect 54022 34726 54050 35478
rect 54270 35436 54566 35456
rect 54326 35434 54350 35436
rect 54406 35434 54430 35436
rect 54486 35434 54510 35436
rect 54348 35382 54350 35434
rect 54412 35382 54424 35434
rect 54486 35382 54488 35434
rect 54326 35380 54350 35382
rect 54406 35380 54430 35382
rect 54486 35380 54510 35382
rect 54270 35360 54566 35380
rect 54102 35264 54154 35270
rect 54102 35206 54154 35212
rect 54114 34998 54142 35206
rect 54666 35134 54694 35546
rect 55862 35134 55890 39082
rect 56126 37712 56178 37718
rect 56126 37654 56178 37660
rect 56138 36834 56166 37654
rect 56126 36828 56178 36834
rect 56126 36770 56178 36776
rect 56138 36222 56166 36770
rect 56126 36216 56178 36222
rect 56126 36158 56178 36164
rect 54654 35128 54706 35134
rect 54654 35070 54706 35076
rect 55850 35128 55902 35134
rect 55850 35070 55902 35076
rect 54102 34992 54154 34998
rect 54102 34934 54154 34940
rect 54286 34992 54338 34998
rect 54286 34934 54338 34940
rect 55298 34992 55350 34998
rect 55298 34934 55350 34940
rect 54010 34720 54062 34726
rect 54010 34662 54062 34668
rect 53274 34652 53326 34658
rect 53274 34594 53326 34600
rect 54022 34590 54050 34662
rect 54010 34584 54062 34590
rect 54010 34526 54062 34532
rect 54298 34522 54326 34934
rect 55310 34794 55338 34934
rect 55298 34788 55350 34794
rect 55298 34730 55350 34736
rect 55390 34788 55442 34794
rect 55390 34730 55442 34736
rect 54286 34516 54338 34522
rect 54286 34458 54338 34464
rect 54194 34448 54246 34454
rect 54194 34390 54246 34396
rect 54654 34448 54706 34454
rect 54654 34390 54706 34396
rect 54206 34250 54234 34390
rect 54270 34348 54566 34368
rect 54326 34346 54350 34348
rect 54406 34346 54430 34348
rect 54486 34346 54510 34348
rect 54348 34294 54350 34346
rect 54412 34294 54424 34346
rect 54486 34294 54488 34346
rect 54326 34292 54350 34294
rect 54406 34292 54430 34294
rect 54486 34292 54510 34294
rect 54270 34272 54566 34292
rect 54194 34244 54246 34250
rect 54194 34186 54246 34192
rect 54666 34046 54694 34390
rect 55402 34114 55430 34730
rect 55390 34108 55442 34114
rect 55390 34050 55442 34056
rect 54654 34040 54706 34046
rect 54654 33982 54706 33988
rect 53458 33904 53510 33910
rect 53458 33846 53510 33852
rect 54654 33904 54706 33910
rect 54654 33846 54706 33852
rect 53470 33502 53498 33846
rect 54666 33706 54694 33846
rect 54654 33700 54706 33706
rect 54654 33642 54706 33648
rect 53642 33632 53694 33638
rect 54010 33632 54062 33638
rect 53694 33580 54010 33586
rect 53642 33574 54062 33580
rect 53654 33558 54050 33574
rect 53458 33496 53510 33502
rect 53458 33438 53510 33444
rect 54270 33260 54566 33280
rect 54326 33258 54350 33260
rect 54406 33258 54430 33260
rect 54486 33258 54510 33260
rect 54348 33206 54350 33258
rect 54412 33206 54424 33258
rect 54486 33206 54488 33258
rect 54326 33204 54350 33206
rect 54406 33204 54430 33206
rect 54486 33204 54510 33206
rect 54270 33184 54566 33204
rect 56598 32958 56626 39354
rect 56874 37854 56902 39490
rect 56934 39244 57230 39264
rect 56990 39242 57014 39244
rect 57070 39242 57094 39244
rect 57150 39242 57174 39244
rect 57012 39190 57014 39242
rect 57076 39190 57088 39242
rect 57150 39190 57152 39242
rect 56990 39188 57014 39190
rect 57070 39188 57094 39190
rect 57150 39188 57174 39190
rect 56934 39168 57230 39188
rect 56934 38156 57230 38176
rect 56990 38154 57014 38156
rect 57070 38154 57094 38156
rect 57150 38154 57174 38156
rect 57012 38102 57014 38154
rect 57076 38102 57088 38154
rect 57150 38102 57152 38154
rect 56990 38100 57014 38102
rect 57070 38100 57094 38102
rect 57150 38100 57174 38102
rect 56934 38080 57230 38100
rect 57138 37916 57190 37922
rect 57138 37858 57190 37864
rect 56862 37848 56914 37854
rect 56862 37790 56914 37796
rect 57150 37310 57178 37858
rect 56770 37304 56822 37310
rect 56770 37246 56822 37252
rect 57138 37304 57190 37310
rect 57138 37246 57190 37252
rect 56782 36290 56810 37246
rect 56934 37068 57230 37088
rect 56990 37066 57014 37068
rect 57070 37066 57094 37068
rect 57150 37066 57174 37068
rect 57012 37014 57014 37066
rect 57076 37014 57088 37066
rect 57150 37014 57152 37066
rect 56990 37012 57014 37014
rect 57070 37012 57094 37014
rect 57150 37012 57174 37014
rect 56934 36992 57230 37012
rect 57138 36760 57190 36766
rect 57138 36702 57190 36708
rect 56770 36284 56822 36290
rect 56770 36226 56822 36232
rect 57150 36222 57178 36702
rect 57138 36216 57190 36222
rect 57138 36158 57190 36164
rect 56934 35980 57230 36000
rect 56990 35978 57014 35980
rect 57070 35978 57094 35980
rect 57150 35978 57174 35980
rect 57012 35926 57014 35978
rect 57076 35926 57088 35978
rect 57150 35926 57152 35978
rect 56990 35924 57014 35926
rect 57070 35924 57094 35926
rect 57150 35924 57174 35926
rect 56934 35904 57230 35924
rect 56676 35776 56732 35785
rect 56676 35711 56732 35720
rect 56690 35678 56718 35711
rect 56678 35672 56730 35678
rect 56678 35614 56730 35620
rect 56934 34892 57230 34912
rect 56990 34890 57014 34892
rect 57070 34890 57094 34892
rect 57150 34890 57174 34892
rect 57012 34838 57014 34890
rect 57076 34838 57088 34890
rect 57150 34838 57152 34890
rect 56990 34836 57014 34838
rect 57070 34836 57094 34838
rect 57150 34836 57174 34838
rect 56934 34816 57230 34836
rect 56934 33804 57230 33824
rect 56990 33802 57014 33804
rect 57070 33802 57094 33804
rect 57150 33802 57174 33804
rect 57012 33750 57014 33802
rect 57076 33750 57088 33802
rect 57150 33750 57152 33802
rect 56990 33748 57014 33750
rect 57070 33748 57094 33750
rect 57150 33748 57174 33750
rect 56934 33728 57230 33748
rect 57334 32958 57362 39626
rect 57702 37922 57730 39950
rect 58622 39690 58650 43312
rect 59818 42154 59846 43312
rect 59542 42126 59846 42154
rect 58702 40976 58754 40982
rect 58702 40918 58754 40924
rect 58714 40642 58742 40918
rect 58702 40636 58754 40642
rect 58702 40578 58754 40584
rect 59542 40506 59570 42126
rect 59598 41964 59894 41984
rect 59654 41962 59678 41964
rect 59734 41962 59758 41964
rect 59814 41962 59838 41964
rect 59676 41910 59678 41962
rect 59740 41910 59752 41962
rect 59814 41910 59816 41962
rect 59654 41908 59678 41910
rect 59734 41908 59758 41910
rect 59814 41908 59838 41910
rect 59598 41888 59894 41908
rect 61106 41322 61134 43312
rect 62302 41610 62330 43312
rect 62302 41582 62698 41610
rect 62262 41420 62558 41440
rect 62318 41418 62342 41420
rect 62398 41418 62422 41420
rect 62478 41418 62502 41420
rect 62340 41366 62342 41418
rect 62404 41366 62416 41418
rect 62478 41366 62480 41418
rect 62318 41364 62342 41366
rect 62398 41364 62422 41366
rect 62478 41364 62502 41366
rect 62262 41344 62558 41364
rect 61094 41316 61146 41322
rect 61094 41258 61146 41264
rect 60266 41112 60318 41118
rect 61738 41112 61790 41118
rect 60266 41054 60318 41060
rect 61658 41060 61738 41066
rect 61658 41054 61790 41060
rect 59598 40876 59894 40896
rect 59654 40874 59678 40876
rect 59734 40874 59758 40876
rect 59814 40874 59838 40876
rect 59676 40822 59678 40874
rect 59740 40822 59752 40874
rect 59814 40822 59816 40874
rect 59654 40820 59678 40822
rect 59734 40820 59758 40822
rect 59814 40820 59838 40822
rect 59598 40800 59894 40820
rect 59530 40500 59582 40506
rect 59530 40442 59582 40448
rect 60278 40030 60306 41054
rect 61658 41038 61778 41054
rect 61658 40642 61686 41038
rect 61738 40976 61790 40982
rect 61738 40918 61790 40924
rect 61646 40636 61698 40642
rect 61646 40578 61698 40584
rect 61370 40568 61422 40574
rect 61370 40510 61422 40516
rect 61382 40234 61410 40510
rect 61370 40228 61422 40234
rect 61370 40170 61422 40176
rect 60266 40024 60318 40030
rect 60266 39966 60318 39972
rect 59990 39956 60042 39962
rect 59990 39898 60042 39904
rect 59598 39788 59894 39808
rect 59654 39786 59678 39788
rect 59734 39786 59758 39788
rect 59814 39786 59838 39788
rect 59676 39734 59678 39786
rect 59740 39734 59752 39786
rect 59814 39734 59816 39786
rect 59654 39732 59678 39734
rect 59734 39732 59758 39734
rect 59814 39732 59838 39734
rect 59598 39712 59894 39732
rect 58610 39684 58662 39690
rect 58610 39626 58662 39632
rect 60002 39010 60030 39898
rect 59990 39004 60042 39010
rect 59990 38946 60042 38952
rect 60278 38806 60306 39966
rect 60358 38936 60410 38942
rect 60358 38878 60410 38884
rect 61370 38936 61422 38942
rect 61370 38878 61422 38884
rect 60266 38800 60318 38806
rect 60186 38748 60266 38754
rect 60186 38742 60318 38748
rect 60186 38726 60306 38742
rect 59598 38700 59894 38720
rect 59654 38698 59678 38700
rect 59734 38698 59758 38700
rect 59814 38698 59838 38700
rect 59676 38646 59678 38698
rect 59740 38646 59752 38698
rect 59814 38646 59816 38698
rect 59654 38644 59678 38646
rect 59734 38644 59758 38646
rect 59814 38644 59838 38646
rect 59598 38624 59894 38644
rect 59070 38460 59122 38466
rect 59070 38402 59122 38408
rect 57966 38256 58018 38262
rect 57966 38198 58018 38204
rect 57690 37916 57742 37922
rect 57690 37858 57742 37864
rect 57872 37816 57928 37825
rect 57872 37751 57928 37760
rect 57780 37136 57836 37145
rect 57780 37071 57836 37080
rect 57794 36766 57822 37071
rect 57782 36760 57834 36766
rect 57688 36728 57744 36737
rect 57782 36702 57834 36708
rect 57688 36663 57690 36672
rect 57742 36663 57744 36672
rect 57690 36634 57742 36640
rect 57782 36624 57834 36630
rect 57782 36566 57834 36572
rect 57794 34658 57822 36566
rect 57886 35785 57914 37751
rect 57978 37378 58006 38198
rect 59082 37854 59110 38402
rect 58058 37848 58110 37854
rect 58058 37790 58110 37796
rect 58150 37848 58202 37854
rect 58150 37790 58202 37796
rect 58886 37848 58938 37854
rect 58886 37790 58938 37796
rect 59070 37848 59122 37854
rect 59070 37790 59122 37796
rect 59438 37848 59490 37854
rect 59438 37790 59490 37796
rect 58070 37718 58098 37790
rect 58058 37712 58110 37718
rect 58058 37654 58110 37660
rect 57966 37372 58018 37378
rect 57966 37314 58018 37320
rect 57964 37272 58020 37281
rect 57964 37207 57966 37216
rect 58018 37207 58020 37216
rect 57966 37178 58018 37184
rect 58070 36970 58098 37654
rect 57966 36964 58018 36970
rect 57966 36906 58018 36912
rect 58058 36964 58110 36970
rect 58058 36906 58110 36912
rect 57978 36850 58006 36906
rect 58162 36850 58190 37790
rect 58242 37440 58294 37446
rect 58242 37382 58294 37388
rect 58254 37174 58282 37382
rect 58898 37378 58926 37790
rect 59082 37718 59110 37790
rect 59070 37712 59122 37718
rect 59070 37654 59122 37660
rect 58610 37372 58662 37378
rect 58610 37314 58662 37320
rect 58886 37372 58938 37378
rect 58886 37314 58938 37320
rect 58242 37168 58294 37174
rect 58242 37110 58294 37116
rect 57978 36822 58190 36850
rect 58058 36760 58110 36766
rect 58058 36702 58110 36708
rect 58424 36728 58480 36737
rect 58070 36154 58098 36702
rect 58424 36663 58426 36672
rect 58478 36663 58480 36672
rect 58426 36634 58478 36640
rect 58622 36630 58650 37314
rect 59450 37242 59478 37790
rect 59598 37612 59894 37632
rect 59654 37610 59678 37612
rect 59734 37610 59758 37612
rect 59814 37610 59838 37612
rect 59676 37558 59678 37610
rect 59740 37558 59752 37610
rect 59814 37558 59816 37610
rect 59654 37556 59678 37558
rect 59734 37556 59758 37558
rect 59814 37556 59838 37558
rect 59598 37536 59894 37556
rect 60186 37378 60214 38726
rect 60370 37514 60398 38878
rect 61382 38534 61410 38878
rect 61658 38602 61686 40578
rect 61750 40574 61778 40918
rect 62670 40642 62698 41582
rect 62658 40636 62710 40642
rect 62658 40578 62710 40584
rect 62934 40636 62986 40642
rect 62934 40578 62986 40584
rect 61738 40568 61790 40574
rect 61738 40510 61790 40516
rect 62750 40568 62802 40574
rect 62750 40510 62802 40516
rect 62658 40432 62710 40438
rect 62658 40374 62710 40380
rect 62262 40332 62558 40352
rect 62318 40330 62342 40332
rect 62398 40330 62422 40332
rect 62478 40330 62502 40332
rect 62340 40278 62342 40330
rect 62404 40278 62416 40330
rect 62478 40278 62480 40330
rect 62318 40276 62342 40278
rect 62398 40276 62422 40278
rect 62478 40276 62502 40278
rect 62262 40256 62558 40276
rect 62106 40092 62158 40098
rect 62106 40034 62158 40040
rect 62118 39690 62146 40034
rect 62670 40030 62698 40374
rect 62658 40024 62710 40030
rect 62658 39966 62710 39972
rect 62106 39684 62158 39690
rect 62106 39626 62158 39632
rect 62762 39350 62790 40510
rect 62750 39344 62802 39350
rect 62750 39286 62802 39292
rect 62262 39244 62558 39264
rect 62318 39242 62342 39244
rect 62398 39242 62422 39244
rect 62478 39242 62502 39244
rect 62340 39190 62342 39242
rect 62404 39190 62416 39242
rect 62478 39190 62480 39242
rect 62318 39188 62342 39190
rect 62398 39188 62422 39190
rect 62478 39188 62502 39190
rect 62262 39168 62558 39188
rect 61646 38596 61698 38602
rect 61646 38538 61698 38544
rect 61370 38528 61422 38534
rect 61370 38470 61422 38476
rect 60634 38392 60686 38398
rect 60634 38334 60686 38340
rect 60542 37984 60594 37990
rect 60542 37926 60594 37932
rect 60358 37508 60410 37514
rect 60358 37450 60410 37456
rect 60554 37378 60582 37926
rect 60646 37922 60674 38334
rect 61738 38256 61790 38262
rect 61738 38198 61790 38204
rect 60634 37916 60686 37922
rect 60634 37858 60686 37864
rect 61750 37854 61778 38198
rect 62262 38156 62558 38176
rect 62318 38154 62342 38156
rect 62398 38154 62422 38156
rect 62478 38154 62502 38156
rect 62340 38102 62342 38154
rect 62404 38102 62416 38154
rect 62478 38102 62480 38154
rect 62318 38100 62342 38102
rect 62398 38100 62422 38102
rect 62478 38100 62502 38102
rect 62262 38080 62558 38100
rect 61738 37848 61790 37854
rect 61738 37790 61790 37796
rect 62106 37848 62158 37854
rect 62106 37790 62158 37796
rect 62474 37848 62526 37854
rect 62474 37790 62526 37796
rect 62118 37718 62146 37790
rect 61370 37712 61422 37718
rect 61370 37654 61422 37660
rect 62106 37712 62158 37718
rect 62106 37654 62158 37660
rect 61382 37514 61410 37654
rect 61370 37508 61422 37514
rect 61370 37450 61422 37456
rect 60174 37372 60226 37378
rect 60174 37314 60226 37320
rect 60358 37372 60410 37378
rect 60358 37314 60410 37320
rect 60542 37372 60594 37378
rect 60542 37314 60594 37320
rect 59622 37304 59674 37310
rect 59620 37272 59622 37281
rect 59674 37272 59676 37281
rect 59438 37236 59490 37242
rect 60370 37242 60398 37314
rect 59620 37207 59676 37216
rect 60358 37236 60410 37242
rect 59438 37178 59490 37184
rect 60358 37178 60410 37184
rect 60554 37174 60582 37314
rect 62118 37310 62146 37654
rect 62486 37446 62514 37790
rect 62474 37440 62526 37446
rect 62474 37382 62526 37388
rect 62106 37304 62158 37310
rect 62106 37246 62158 37252
rect 62118 37174 62146 37246
rect 60542 37168 60594 37174
rect 60542 37110 60594 37116
rect 61186 37168 61238 37174
rect 62106 37168 62158 37174
rect 61186 37110 61238 37116
rect 62104 37136 62106 37145
rect 62158 37136 62160 37145
rect 61198 36902 61226 37110
rect 62104 37071 62160 37080
rect 62262 37068 62558 37088
rect 62318 37066 62342 37068
rect 62398 37066 62422 37068
rect 62478 37066 62502 37068
rect 62340 37014 62342 37066
rect 62404 37014 62416 37066
rect 62478 37014 62480 37066
rect 62318 37012 62342 37014
rect 62398 37012 62422 37014
rect 62478 37012 62502 37014
rect 62262 36992 62558 37012
rect 62014 36964 62066 36970
rect 62014 36906 62066 36912
rect 61186 36896 61238 36902
rect 61186 36838 61238 36844
rect 58610 36624 58662 36630
rect 58610 36566 58662 36572
rect 62026 36578 62054 36906
rect 62474 36624 62526 36630
rect 62026 36572 62474 36578
rect 62026 36566 62526 36572
rect 62026 36550 62514 36566
rect 59598 36524 59894 36544
rect 59654 36522 59678 36524
rect 59734 36522 59758 36524
rect 59814 36522 59838 36524
rect 59676 36470 59678 36522
rect 59740 36470 59752 36522
rect 59814 36470 59816 36522
rect 59654 36468 59678 36470
rect 59734 36468 59758 36470
rect 59814 36468 59838 36470
rect 59598 36448 59894 36468
rect 61462 36352 61514 36358
rect 61462 36294 61514 36300
rect 61474 36154 61502 36294
rect 61830 36284 61882 36290
rect 61830 36226 61882 36232
rect 61554 36216 61606 36222
rect 61738 36216 61790 36222
rect 61606 36164 61738 36170
rect 61554 36158 61790 36164
rect 58058 36148 58110 36154
rect 58058 36090 58110 36096
rect 61462 36148 61514 36154
rect 61566 36142 61778 36158
rect 61462 36090 61514 36096
rect 59070 36080 59122 36086
rect 59070 36022 59122 36028
rect 57872 35776 57928 35785
rect 57872 35711 57874 35720
rect 57926 35711 57928 35720
rect 57874 35682 57926 35688
rect 57886 35651 57914 35682
rect 59082 35678 59110 36022
rect 61842 35746 61870 36226
rect 62564 36184 62620 36193
rect 62564 36119 62566 36128
rect 62618 36119 62620 36128
rect 62566 36090 62618 36096
rect 62262 35980 62558 36000
rect 62318 35978 62342 35980
rect 62398 35978 62422 35980
rect 62478 35978 62502 35980
rect 62340 35926 62342 35978
rect 62404 35926 62416 35978
rect 62478 35926 62480 35978
rect 62318 35924 62342 35926
rect 62398 35924 62422 35926
rect 62478 35924 62502 35926
rect 62262 35904 62558 35924
rect 62762 35898 62790 39286
rect 62946 38942 62974 40578
rect 63498 40234 63526 43312
rect 63578 40976 63630 40982
rect 63578 40918 63630 40924
rect 63590 40642 63618 40918
rect 63578 40636 63630 40642
rect 63578 40578 63630 40584
rect 64038 40432 64090 40438
rect 64038 40374 64090 40380
rect 63486 40228 63538 40234
rect 63486 40170 63538 40176
rect 64050 40166 64078 40374
rect 64038 40160 64090 40166
rect 64038 40102 64090 40108
rect 63118 39956 63170 39962
rect 63118 39898 63170 39904
rect 63026 39004 63078 39010
rect 63026 38946 63078 38952
rect 62934 38936 62986 38942
rect 62934 38878 62986 38884
rect 62934 36760 62986 36766
rect 62934 36702 62986 36708
rect 62762 35870 62882 35898
rect 59990 35740 60042 35746
rect 59990 35682 60042 35688
rect 61830 35740 61882 35746
rect 61830 35682 61882 35688
rect 58334 35672 58386 35678
rect 58334 35614 58386 35620
rect 58886 35672 58938 35678
rect 58886 35614 58938 35620
rect 59070 35672 59122 35678
rect 59070 35614 59122 35620
rect 57782 34652 57834 34658
rect 57782 34594 57834 34600
rect 58346 34590 58374 35614
rect 58898 34590 58926 35614
rect 59598 35436 59894 35456
rect 59654 35434 59678 35436
rect 59734 35434 59758 35436
rect 59814 35434 59838 35436
rect 59676 35382 59678 35434
rect 59740 35382 59752 35434
rect 59814 35382 59816 35434
rect 59654 35380 59678 35382
rect 59734 35380 59758 35382
rect 59814 35380 59838 35382
rect 59598 35360 59894 35380
rect 60002 34658 60030 35682
rect 60174 35672 60226 35678
rect 60174 35614 60226 35620
rect 62382 35672 62434 35678
rect 62382 35614 62434 35620
rect 62566 35672 62618 35678
rect 62566 35614 62618 35620
rect 59438 34652 59490 34658
rect 59438 34594 59490 34600
rect 59990 34652 60042 34658
rect 59990 34594 60042 34600
rect 57414 34584 57466 34590
rect 57414 34526 57466 34532
rect 58334 34584 58386 34590
rect 58426 34584 58478 34590
rect 58334 34526 58386 34532
rect 58424 34552 58426 34561
rect 58886 34584 58938 34590
rect 58478 34552 58480 34561
rect 57426 33026 57454 34526
rect 58886 34526 58938 34532
rect 58424 34487 58480 34496
rect 59450 33978 59478 34594
rect 60186 34590 60214 35614
rect 60266 35604 60318 35610
rect 60266 35546 60318 35552
rect 60174 34584 60226 34590
rect 60174 34526 60226 34532
rect 59598 34348 59894 34368
rect 59654 34346 59678 34348
rect 59734 34346 59758 34348
rect 59814 34346 59838 34348
rect 59676 34294 59678 34346
rect 59740 34294 59752 34346
rect 59814 34294 59816 34346
rect 59654 34292 59678 34294
rect 59734 34292 59758 34294
rect 59814 34292 59838 34294
rect 59598 34272 59894 34292
rect 59806 34040 59858 34046
rect 59858 34000 59938 34028
rect 59806 33982 59858 33988
rect 59910 33994 59938 34000
rect 59910 33978 60122 33994
rect 59438 33972 59490 33978
rect 59910 33972 60134 33978
rect 59910 33966 60082 33972
rect 59438 33914 59490 33920
rect 60082 33914 60134 33920
rect 59530 33904 59582 33910
rect 59530 33846 59582 33852
rect 59990 33904 60042 33910
rect 59990 33846 60042 33852
rect 58886 33700 58938 33706
rect 58938 33660 59202 33688
rect 58886 33642 58938 33648
rect 57874 33496 57926 33502
rect 57874 33438 57926 33444
rect 58426 33496 58478 33502
rect 58426 33438 58478 33444
rect 58518 33496 58570 33502
rect 58518 33438 58570 33444
rect 57598 33360 57650 33366
rect 57598 33302 57650 33308
rect 57610 33162 57638 33302
rect 57598 33156 57650 33162
rect 57598 33098 57650 33104
rect 57414 33020 57466 33026
rect 57414 32962 57466 32968
rect 56586 32952 56638 32958
rect 56586 32894 56638 32900
rect 57322 32952 57374 32958
rect 57322 32894 57374 32900
rect 54194 32884 54246 32890
rect 54194 32826 54246 32832
rect 53182 32544 53234 32550
rect 53182 32486 53234 32492
rect 53838 31938 54142 31954
rect 53642 31932 53694 31938
rect 53642 31874 53694 31880
rect 53838 31932 54154 31938
rect 53838 31926 54102 31932
rect 53654 31326 53682 31874
rect 53838 31734 53866 31926
rect 54102 31874 54154 31880
rect 54206 31818 54234 32826
rect 56934 32716 57230 32736
rect 56990 32714 57014 32716
rect 57070 32714 57094 32716
rect 57150 32714 57174 32716
rect 57012 32662 57014 32714
rect 57076 32662 57088 32714
rect 57150 32662 57152 32714
rect 56990 32660 57014 32662
rect 57070 32660 57094 32662
rect 57150 32660 57174 32662
rect 56934 32640 57230 32660
rect 57334 32482 57362 32894
rect 57886 32657 57914 33438
rect 57966 33360 58018 33366
rect 57966 33302 58018 33308
rect 57978 33026 58006 33302
rect 58438 33162 58466 33438
rect 58426 33156 58478 33162
rect 58426 33098 58478 33104
rect 57966 33020 58018 33026
rect 57966 32962 58018 32968
rect 58058 33020 58110 33026
rect 58058 32962 58110 32968
rect 58242 33020 58294 33026
rect 58242 32962 58294 32968
rect 57872 32648 57928 32657
rect 57872 32583 57928 32592
rect 57322 32476 57374 32482
rect 57322 32418 57374 32424
rect 58070 32414 58098 32962
rect 58254 32822 58282 32962
rect 58242 32816 58294 32822
rect 58242 32758 58294 32764
rect 58334 32816 58386 32822
rect 58334 32758 58386 32764
rect 58346 32482 58374 32758
rect 58438 32550 58466 33098
rect 58426 32544 58478 32550
rect 58426 32486 58478 32492
rect 58334 32476 58386 32482
rect 58334 32418 58386 32424
rect 58530 32414 58558 33438
rect 59174 33434 59202 33660
rect 59346 33496 59398 33502
rect 59346 33438 59398 33444
rect 59162 33428 59214 33434
rect 59162 33370 59214 33376
rect 59358 33162 59386 33438
rect 59438 33360 59490 33366
rect 59438 33302 59490 33308
rect 59346 33156 59398 33162
rect 59346 33098 59398 33104
rect 59450 33026 59478 33302
rect 59438 33020 59490 33026
rect 59438 32962 59490 32968
rect 58792 32920 58848 32929
rect 58792 32855 58848 32864
rect 58806 32822 58834 32855
rect 58794 32816 58846 32822
rect 58794 32758 58846 32764
rect 59346 32816 59398 32822
rect 59346 32758 59398 32764
rect 59358 32414 59386 32758
rect 59542 32550 59570 33846
rect 60002 33706 60030 33846
rect 60278 33706 60306 35546
rect 61922 35536 61974 35542
rect 61922 35478 61974 35484
rect 62106 35536 62158 35542
rect 62394 35513 62422 35614
rect 62578 35542 62606 35614
rect 62566 35536 62618 35542
rect 62106 35478 62158 35484
rect 62380 35504 62436 35513
rect 60816 35368 60872 35377
rect 60816 35303 60872 35312
rect 60830 35270 60858 35303
rect 60818 35264 60870 35270
rect 60818 35206 60870 35212
rect 61002 34788 61054 34794
rect 61002 34730 61054 34736
rect 61014 34250 61042 34730
rect 60450 34244 60502 34250
rect 60450 34186 60502 34192
rect 61002 34244 61054 34250
rect 61002 34186 61054 34192
rect 60462 33706 60490 34186
rect 59990 33700 60042 33706
rect 59990 33642 60042 33648
rect 60082 33700 60134 33706
rect 60082 33642 60134 33648
rect 60266 33700 60318 33706
rect 60266 33642 60318 33648
rect 60450 33700 60502 33706
rect 60450 33642 60502 33648
rect 59598 33260 59894 33280
rect 59654 33258 59678 33260
rect 59734 33258 59758 33260
rect 59814 33258 59838 33260
rect 59676 33206 59678 33258
rect 59740 33206 59752 33258
rect 59814 33206 59816 33258
rect 59654 33204 59678 33206
rect 59734 33204 59758 33206
rect 59814 33204 59838 33206
rect 59598 33184 59894 33204
rect 60094 33162 60122 33642
rect 60908 33600 60964 33609
rect 60908 33535 60964 33544
rect 60922 33502 60950 33535
rect 60910 33496 60962 33502
rect 60910 33438 60962 33444
rect 61934 33366 61962 35478
rect 62118 35338 62146 35478
rect 62566 35478 62618 35484
rect 62380 35439 62436 35448
rect 62106 35332 62158 35338
rect 62106 35274 62158 35280
rect 62566 35196 62618 35202
rect 62618 35156 62698 35184
rect 62566 35138 62618 35144
rect 62106 35128 62158 35134
rect 62106 35070 62158 35076
rect 62118 34658 62146 35070
rect 62262 34892 62558 34912
rect 62318 34890 62342 34892
rect 62398 34890 62422 34892
rect 62478 34890 62502 34892
rect 62340 34838 62342 34890
rect 62404 34838 62416 34890
rect 62478 34838 62480 34890
rect 62318 34836 62342 34838
rect 62398 34836 62422 34838
rect 62478 34836 62502 34838
rect 62262 34816 62558 34836
rect 62106 34652 62158 34658
rect 62106 34594 62158 34600
rect 62566 34584 62618 34590
rect 62670 34572 62698 35156
rect 62618 34544 62698 34572
rect 62566 34526 62618 34532
rect 62578 34454 62606 34526
rect 62566 34448 62618 34454
rect 62566 34390 62618 34396
rect 62262 33804 62558 33824
rect 62318 33802 62342 33804
rect 62398 33802 62422 33804
rect 62478 33802 62502 33804
rect 62340 33750 62342 33802
rect 62404 33750 62416 33802
rect 62478 33750 62480 33802
rect 62318 33748 62342 33750
rect 62398 33748 62422 33750
rect 62478 33748 62502 33750
rect 62262 33728 62558 33748
rect 62656 33736 62712 33745
rect 62656 33671 62712 33680
rect 62670 33638 62698 33671
rect 62658 33632 62710 33638
rect 62658 33574 62710 33580
rect 62854 33570 62882 35870
rect 62842 33564 62894 33570
rect 62842 33506 62894 33512
rect 61922 33360 61974 33366
rect 61922 33302 61974 33308
rect 60082 33156 60134 33162
rect 60082 33098 60134 33104
rect 60910 33156 60962 33162
rect 60910 33098 60962 33104
rect 60922 33026 60950 33098
rect 61094 33088 61146 33094
rect 61278 33088 61330 33094
rect 61146 33036 61278 33042
rect 61094 33030 61330 33036
rect 60174 33020 60226 33026
rect 60174 32962 60226 32968
rect 60358 33020 60410 33026
rect 60358 32962 60410 32968
rect 60910 33020 60962 33026
rect 61106 33014 61318 33030
rect 62750 33020 62802 33026
rect 60910 32962 60962 32968
rect 62750 32962 62802 32968
rect 59806 32884 59858 32890
rect 59806 32826 59858 32832
rect 59530 32544 59582 32550
rect 59818 32521 59846 32826
rect 60082 32612 60134 32618
rect 60082 32554 60134 32560
rect 59530 32486 59582 32492
rect 59804 32512 59860 32521
rect 59804 32447 59860 32456
rect 58058 32408 58110 32414
rect 58058 32350 58110 32356
rect 58518 32408 58570 32414
rect 58518 32350 58570 32356
rect 59346 32408 59398 32414
rect 59346 32350 59398 32356
rect 58426 32272 58478 32278
rect 58424 32240 58426 32249
rect 58478 32240 58480 32249
rect 54270 32172 54566 32192
rect 58424 32175 58480 32184
rect 54326 32170 54350 32172
rect 54406 32170 54430 32172
rect 54486 32170 54510 32172
rect 54348 32118 54350 32170
rect 54412 32118 54424 32170
rect 54486 32118 54488 32170
rect 54326 32116 54350 32118
rect 54406 32116 54430 32118
rect 54486 32116 54510 32118
rect 54270 32096 54566 32116
rect 57598 31932 57650 31938
rect 57598 31874 57650 31880
rect 57702 31926 58374 31954
rect 57610 31841 57638 31874
rect 57702 31870 57730 31926
rect 58346 31870 58374 31926
rect 58530 31870 58558 32350
rect 60094 32249 60122 32554
rect 58700 32240 58756 32249
rect 60080 32240 60136 32249
rect 58700 32175 58756 32184
rect 58714 32006 58742 32175
rect 59598 32172 59894 32192
rect 60080 32175 60136 32184
rect 59654 32170 59678 32172
rect 59734 32170 59758 32172
rect 59814 32170 59838 32172
rect 59676 32118 59678 32170
rect 59740 32118 59752 32170
rect 59814 32118 59816 32170
rect 59654 32116 59678 32118
rect 59734 32116 59758 32118
rect 59814 32116 59838 32118
rect 59598 32096 59894 32116
rect 58610 32000 58662 32006
rect 58608 31968 58610 31977
rect 58702 32000 58754 32006
rect 58662 31968 58664 31977
rect 58702 31942 58754 31948
rect 60186 31938 60214 32962
rect 60370 32822 60398 32962
rect 60358 32816 60410 32822
rect 60358 32758 60410 32764
rect 61370 32816 61422 32822
rect 61370 32758 61422 32764
rect 60370 32414 60398 32758
rect 61382 32414 61410 32758
rect 62262 32716 62558 32736
rect 62318 32714 62342 32716
rect 62398 32714 62422 32716
rect 62478 32714 62502 32716
rect 62340 32662 62342 32714
rect 62404 32662 62416 32714
rect 62478 32662 62480 32714
rect 62318 32660 62342 32662
rect 62398 32660 62422 32662
rect 62478 32660 62502 32662
rect 62012 32648 62068 32657
rect 62262 32640 62558 32660
rect 62012 32583 62068 32592
rect 60358 32408 60410 32414
rect 60358 32350 60410 32356
rect 61370 32408 61422 32414
rect 61370 32350 61422 32356
rect 58608 31903 58664 31912
rect 60174 31932 60226 31938
rect 60174 31874 60226 31880
rect 57690 31864 57742 31870
rect 57596 31832 57652 31841
rect 53930 31802 54326 31818
rect 53918 31796 54326 31802
rect 53970 31790 54326 31796
rect 53918 31738 53970 31744
rect 53826 31728 53878 31734
rect 53826 31670 53878 31676
rect 54010 31728 54062 31734
rect 54010 31670 54062 31676
rect 54194 31728 54246 31734
rect 54194 31670 54246 31676
rect 54022 31326 54050 31670
rect 54206 31546 54234 31670
rect 54114 31530 54234 31546
rect 54102 31524 54234 31530
rect 54154 31518 54234 31524
rect 54102 31466 54154 31472
rect 54298 31462 54326 31790
rect 57690 31806 57742 31812
rect 58334 31864 58386 31870
rect 58334 31806 58386 31812
rect 58518 31864 58570 31870
rect 58518 31806 58570 31812
rect 58884 31832 58940 31841
rect 57596 31767 57652 31776
rect 58150 31796 58202 31802
rect 58150 31738 58202 31744
rect 56934 31628 57230 31648
rect 56990 31626 57014 31628
rect 57070 31626 57094 31628
rect 57150 31626 57174 31628
rect 57012 31574 57014 31626
rect 57076 31574 57088 31626
rect 57150 31574 57152 31626
rect 56990 31572 57014 31574
rect 57070 31572 57094 31574
rect 57150 31572 57174 31574
rect 56934 31552 57230 31572
rect 54286 31456 54338 31462
rect 54286 31398 54338 31404
rect 54654 31456 54706 31462
rect 54654 31398 54706 31404
rect 54744 31424 54800 31433
rect 53642 31320 53694 31326
rect 53642 31262 53694 31268
rect 54010 31320 54062 31326
rect 54010 31262 54062 31268
rect 52814 30776 52866 30782
rect 52814 30718 52866 30724
rect 52906 30776 52958 30782
rect 52906 30718 52958 30724
rect 53654 30374 53682 31262
rect 53826 30912 53878 30918
rect 53826 30854 53878 30860
rect 53916 30880 53972 30889
rect 53642 30368 53694 30374
rect 53642 30310 53694 30316
rect 51066 30232 51118 30238
rect 51066 30174 51118 30180
rect 51986 30232 52038 30238
rect 51986 30174 52038 30180
rect 52630 30232 52682 30238
rect 52630 30174 52682 30180
rect 50882 29756 50934 29762
rect 50882 29698 50934 29704
rect 50802 29478 51014 29506
rect 50986 29354 51014 29478
rect 50882 29348 50934 29354
rect 50882 29290 50934 29296
rect 50974 29348 51026 29354
rect 50974 29290 51026 29296
rect 49962 29008 50014 29014
rect 49962 28950 50014 28956
rect 49974 28266 50002 28950
rect 50330 28736 50382 28742
rect 50330 28678 50382 28684
rect 50054 28668 50106 28674
rect 50054 28610 50106 28616
rect 49962 28260 50014 28266
rect 49962 28202 50014 28208
rect 50066 28062 50094 28610
rect 50342 28266 50370 28678
rect 50894 28538 50922 29290
rect 50422 28532 50474 28538
rect 50422 28474 50474 28480
rect 50882 28532 50934 28538
rect 50882 28474 50934 28480
rect 50434 28266 50462 28474
rect 50330 28260 50382 28266
rect 50330 28202 50382 28208
rect 50422 28260 50474 28266
rect 50422 28202 50474 28208
rect 50054 28056 50106 28062
rect 50054 27998 50106 28004
rect 50790 28056 50842 28062
rect 50790 27998 50842 28004
rect 50422 27988 50474 27994
rect 50422 27930 50474 27936
rect 50434 27897 50462 27930
rect 50420 27888 50476 27897
rect 50420 27823 50476 27832
rect 50146 27648 50198 27654
rect 50146 27590 50198 27596
rect 49778 27580 49830 27586
rect 49778 27522 49830 27528
rect 49790 27382 49818 27522
rect 49778 27376 49830 27382
rect 49778 27318 49830 27324
rect 50158 27042 50186 27590
rect 50238 27580 50290 27586
rect 50238 27522 50290 27528
rect 50146 27036 50198 27042
rect 50146 26978 50198 26984
rect 50250 26974 50278 27522
rect 50434 26974 50462 27823
rect 50802 27382 50830 27998
rect 51078 27926 51106 30174
rect 52446 29824 52498 29830
rect 52498 29784 52578 29812
rect 52446 29766 52498 29772
rect 52260 29656 52316 29665
rect 52260 29591 52262 29600
rect 52314 29591 52316 29600
rect 52262 29562 52314 29568
rect 52446 29552 52498 29558
rect 52446 29494 52498 29500
rect 51606 29452 51902 29472
rect 51662 29450 51686 29452
rect 51742 29450 51766 29452
rect 51822 29450 51846 29452
rect 51684 29398 51686 29450
rect 51748 29398 51760 29450
rect 51822 29398 51824 29450
rect 51662 29396 51686 29398
rect 51742 29396 51766 29398
rect 51822 29396 51846 29398
rect 51606 29376 51902 29396
rect 52354 29212 52406 29218
rect 52354 29154 52406 29160
rect 51158 29144 51210 29150
rect 51158 29086 51210 29092
rect 51802 29144 51854 29150
rect 51802 29086 51854 29092
rect 51066 27920 51118 27926
rect 51170 27897 51198 29086
rect 51814 28606 51842 29086
rect 52076 28704 52132 28713
rect 51894 28668 51946 28674
rect 51946 28628 52026 28656
rect 52076 28639 52078 28648
rect 51894 28610 51946 28616
rect 51802 28600 51854 28606
rect 51802 28542 51854 28548
rect 51606 28364 51902 28384
rect 51662 28362 51686 28364
rect 51742 28362 51766 28364
rect 51822 28362 51846 28364
rect 51684 28310 51686 28362
rect 51748 28310 51760 28362
rect 51822 28310 51824 28362
rect 51662 28308 51686 28310
rect 51742 28308 51766 28310
rect 51822 28308 51846 28310
rect 51606 28288 51902 28308
rect 51526 28192 51578 28198
rect 51526 28134 51578 28140
rect 51538 28033 51566 28134
rect 51524 28024 51580 28033
rect 51524 27959 51580 27968
rect 51250 27920 51302 27926
rect 51066 27862 51118 27868
rect 51156 27888 51212 27897
rect 50790 27376 50842 27382
rect 50790 27318 50842 27324
rect 51078 27081 51106 27862
rect 51250 27862 51302 27868
rect 51156 27823 51212 27832
rect 51262 27586 51290 27862
rect 51250 27580 51302 27586
rect 51618 27580 51670 27586
rect 51250 27522 51302 27528
rect 51538 27540 51618 27568
rect 51434 27512 51486 27518
rect 51434 27454 51486 27460
rect 51158 27376 51210 27382
rect 51158 27318 51210 27324
rect 51170 27110 51198 27318
rect 51158 27104 51210 27110
rect 51064 27072 51120 27081
rect 51158 27046 51210 27052
rect 51446 27042 51474 27454
rect 51538 27382 51566 27540
rect 51618 27522 51670 27528
rect 51526 27376 51578 27382
rect 51526 27318 51578 27324
rect 51606 27276 51902 27296
rect 51662 27274 51686 27276
rect 51742 27274 51766 27276
rect 51822 27274 51846 27276
rect 51684 27222 51686 27274
rect 51748 27222 51760 27274
rect 51822 27222 51824 27274
rect 51662 27220 51686 27222
rect 51742 27220 51766 27222
rect 51822 27220 51846 27222
rect 51606 27200 51902 27220
rect 51998 27194 52026 28628
rect 52130 28639 52132 28648
rect 52078 28610 52130 28616
rect 52090 28266 52118 28610
rect 52366 28606 52394 29154
rect 52458 28656 52486 29494
rect 52550 29150 52578 29784
rect 52642 29558 52670 30174
rect 53838 29762 53866 30854
rect 53916 30815 53972 30824
rect 53930 30306 53958 30815
rect 54022 30714 54050 31262
rect 54666 31258 54694 31398
rect 54744 31359 54746 31368
rect 54798 31359 54800 31368
rect 54746 31330 54798 31336
rect 57506 31320 57558 31326
rect 57504 31288 57506 31297
rect 57874 31320 57926 31326
rect 57558 31288 57560 31297
rect 54654 31252 54706 31258
rect 57874 31262 57926 31268
rect 57504 31223 57560 31232
rect 54654 31194 54706 31200
rect 54102 31184 54154 31190
rect 54102 31126 54154 31132
rect 54114 30850 54142 31126
rect 54270 31084 54566 31104
rect 54326 31082 54350 31084
rect 54406 31082 54430 31084
rect 54486 31082 54510 31084
rect 54348 31030 54350 31082
rect 54412 31030 54424 31082
rect 54486 31030 54488 31082
rect 54326 31028 54350 31030
rect 54406 31028 54430 31030
rect 54486 31028 54510 31030
rect 54270 31008 54566 31028
rect 54102 30844 54154 30850
rect 54102 30786 54154 30792
rect 54010 30708 54062 30714
rect 54010 30650 54062 30656
rect 53918 30300 53970 30306
rect 53918 30242 53970 30248
rect 54022 30238 54050 30650
rect 54010 30232 54062 30238
rect 54010 30174 54062 30180
rect 54194 30164 54246 30170
rect 54194 30106 54246 30112
rect 54010 30096 54062 30102
rect 54010 30038 54062 30044
rect 54102 30096 54154 30102
rect 54102 30038 54154 30044
rect 52814 29756 52866 29762
rect 52814 29698 52866 29704
rect 53826 29756 53878 29762
rect 53826 29698 53878 29704
rect 52630 29552 52682 29558
rect 52630 29494 52682 29500
rect 52538 29144 52590 29150
rect 52538 29086 52590 29092
rect 52628 29112 52684 29121
rect 52628 29047 52630 29056
rect 52682 29047 52684 29056
rect 52630 29018 52682 29024
rect 52826 28674 52854 29698
rect 53918 29620 53970 29626
rect 53918 29562 53970 29568
rect 53642 29144 53694 29150
rect 53642 29086 53694 29092
rect 52996 28704 53052 28713
rect 52814 28668 52866 28674
rect 52458 28628 52578 28656
rect 52354 28600 52406 28606
rect 52354 28542 52406 28548
rect 52078 28260 52130 28266
rect 52078 28202 52130 28208
rect 52550 28130 52578 28628
rect 52996 28639 53052 28648
rect 52814 28610 52866 28616
rect 53010 28606 53038 28639
rect 52998 28600 53050 28606
rect 52998 28542 53050 28548
rect 53654 28470 53682 29086
rect 53826 29008 53878 29014
rect 53826 28950 53878 28956
rect 53838 28674 53866 28950
rect 53826 28668 53878 28674
rect 53826 28610 53878 28616
rect 53826 28532 53878 28538
rect 53826 28474 53878 28480
rect 53642 28464 53694 28470
rect 53642 28406 53694 28412
rect 53838 28266 53866 28474
rect 53930 28266 53958 29562
rect 54022 29558 54050 30038
rect 54114 29898 54142 30038
rect 54206 29898 54234 30106
rect 54270 29996 54566 30016
rect 54326 29994 54350 29996
rect 54406 29994 54430 29996
rect 54486 29994 54510 29996
rect 54348 29942 54350 29994
rect 54412 29942 54424 29994
rect 54486 29942 54488 29994
rect 54326 29940 54350 29942
rect 54406 29940 54430 29942
rect 54486 29940 54510 29942
rect 54270 29920 54566 29940
rect 54666 29898 54694 31194
rect 54838 31184 54890 31190
rect 54838 31126 54890 31132
rect 54850 30850 54878 31126
rect 57886 30918 57914 31262
rect 57874 30912 57926 30918
rect 57874 30854 57926 30860
rect 58162 30850 58190 31738
rect 58346 30850 58374 31806
rect 58530 30850 58558 31806
rect 58884 31767 58940 31776
rect 58898 31734 58926 31767
rect 58610 31728 58662 31734
rect 58610 31670 58662 31676
rect 58794 31728 58846 31734
rect 58794 31670 58846 31676
rect 58886 31728 58938 31734
rect 58886 31670 58938 31676
rect 58622 31394 58650 31670
rect 58610 31388 58662 31394
rect 58610 31330 58662 31336
rect 54838 30844 54890 30850
rect 54838 30786 54890 30792
rect 58150 30844 58202 30850
rect 58150 30786 58202 30792
rect 58334 30844 58386 30850
rect 58334 30786 58386 30792
rect 58518 30844 58570 30850
rect 58518 30786 58570 30792
rect 56934 30540 57230 30560
rect 56990 30538 57014 30540
rect 57070 30538 57094 30540
rect 57150 30538 57174 30540
rect 57012 30486 57014 30538
rect 57076 30486 57088 30538
rect 57150 30486 57152 30538
rect 56990 30484 57014 30486
rect 57070 30484 57094 30486
rect 57150 30484 57174 30486
rect 56934 30464 57230 30484
rect 58610 30232 58662 30238
rect 58610 30174 58662 30180
rect 55022 30096 55074 30102
rect 55022 30038 55074 30044
rect 54102 29892 54154 29898
rect 54102 29834 54154 29840
rect 54194 29892 54246 29898
rect 54194 29834 54246 29840
rect 54654 29892 54706 29898
rect 54654 29834 54706 29840
rect 54102 29756 54154 29762
rect 54102 29698 54154 29704
rect 54010 29552 54062 29558
rect 54010 29494 54062 29500
rect 54022 28554 54050 29494
rect 54114 29354 54142 29698
rect 54102 29348 54154 29354
rect 54102 29290 54154 29296
rect 54114 29150 54142 29290
rect 54102 29144 54154 29150
rect 54102 29086 54154 29092
rect 54206 28674 54234 29834
rect 55034 29830 55062 30038
rect 58622 29898 58650 30174
rect 58610 29892 58662 29898
rect 58610 29834 58662 29840
rect 55022 29824 55074 29830
rect 55022 29766 55074 29772
rect 56402 29756 56454 29762
rect 56402 29698 56454 29704
rect 54468 29656 54524 29665
rect 54378 29620 54430 29626
rect 54468 29591 54470 29600
rect 54378 29562 54430 29568
rect 54522 29591 54524 29600
rect 54470 29562 54522 29568
rect 54286 29348 54338 29354
rect 54286 29290 54338 29296
rect 54298 29218 54326 29290
rect 54286 29212 54338 29218
rect 54286 29154 54338 29160
rect 54390 29150 54418 29562
rect 54930 29280 54982 29286
rect 54930 29222 54982 29228
rect 54378 29144 54430 29150
rect 54378 29086 54430 29092
rect 54270 28908 54566 28928
rect 54326 28906 54350 28908
rect 54406 28906 54430 28908
rect 54486 28906 54510 28908
rect 54348 28854 54350 28906
rect 54412 28854 54424 28906
rect 54486 28854 54488 28906
rect 54326 28852 54350 28854
rect 54406 28852 54430 28854
rect 54486 28852 54510 28854
rect 54270 28832 54566 28852
rect 54942 28810 54970 29222
rect 55298 29144 55350 29150
rect 55298 29086 55350 29092
rect 54930 28804 54982 28810
rect 54930 28746 54982 28752
rect 55310 28674 55338 29086
rect 56414 28810 56442 29698
rect 56934 29452 57230 29472
rect 56990 29450 57014 29452
rect 57070 29450 57094 29452
rect 57150 29450 57174 29452
rect 57012 29398 57014 29450
rect 57076 29398 57088 29450
rect 57150 29398 57152 29450
rect 56990 29396 57014 29398
rect 57070 29396 57094 29398
rect 57150 29396 57174 29398
rect 56934 29376 57230 29396
rect 58622 29218 58650 29834
rect 58610 29212 58662 29218
rect 58610 29154 58662 29160
rect 56584 29112 56640 29121
rect 56584 29047 56640 29056
rect 57506 29076 57558 29082
rect 56402 28804 56454 28810
rect 56402 28746 56454 28752
rect 56598 28742 56626 29047
rect 57506 29018 57558 29024
rect 56586 28736 56638 28742
rect 56586 28678 56638 28684
rect 57518 28674 57546 29018
rect 54194 28668 54246 28674
rect 54194 28610 54246 28616
rect 55298 28668 55350 28674
rect 55298 28610 55350 28616
rect 57506 28668 57558 28674
rect 57506 28610 57558 28616
rect 54286 28600 54338 28606
rect 54022 28548 54286 28554
rect 54022 28542 54338 28548
rect 56494 28600 56546 28606
rect 56494 28542 56546 28548
rect 54022 28526 54326 28542
rect 53826 28260 53878 28266
rect 53826 28202 53878 28208
rect 53918 28260 53970 28266
rect 53918 28202 53970 28208
rect 52538 28124 52590 28130
rect 52538 28066 52590 28072
rect 52906 28124 52958 28130
rect 52906 28066 52958 28072
rect 52078 28056 52130 28062
rect 52078 27998 52130 28004
rect 52354 28056 52406 28062
rect 52354 27998 52406 28004
rect 52090 27704 52118 27998
rect 52170 27716 52222 27722
rect 52090 27676 52170 27704
rect 52170 27658 52222 27664
rect 52366 27518 52394 27998
rect 52354 27512 52406 27518
rect 52918 27489 52946 28066
rect 53458 28056 53510 28062
rect 53458 27998 53510 28004
rect 53366 27920 53418 27926
rect 53366 27862 53418 27868
rect 53378 27586 53406 27862
rect 53366 27580 53418 27586
rect 53366 27522 53418 27528
rect 52354 27454 52406 27460
rect 52904 27480 52960 27489
rect 52904 27415 52960 27424
rect 51998 27166 52118 27194
rect 51064 27007 51120 27016
rect 51434 27036 51486 27042
rect 51078 26974 51106 27007
rect 52090 27024 52118 27166
rect 52906 27104 52958 27110
rect 52904 27072 52906 27081
rect 52958 27072 52960 27081
rect 52170 27036 52222 27042
rect 52090 26996 52170 27024
rect 51434 26978 51486 26984
rect 52904 27007 52960 27016
rect 52170 26978 52222 26984
rect 50238 26968 50290 26974
rect 50238 26910 50290 26916
rect 50422 26968 50474 26974
rect 50422 26910 50474 26916
rect 51066 26968 51118 26974
rect 51066 26910 51118 26916
rect 53470 26906 53498 27998
rect 53838 27654 53866 28202
rect 54008 27888 54064 27897
rect 54008 27823 54064 27832
rect 53734 27648 53786 27654
rect 53734 27590 53786 27596
rect 53826 27648 53878 27654
rect 53826 27590 53878 27596
rect 53746 27110 53774 27590
rect 54022 27586 54050 27823
rect 54270 27820 54566 27840
rect 54326 27818 54350 27820
rect 54406 27818 54430 27820
rect 54486 27818 54510 27820
rect 54348 27766 54350 27818
rect 54412 27766 54424 27818
rect 54486 27766 54488 27818
rect 54326 27764 54350 27766
rect 54406 27764 54430 27766
rect 54486 27764 54510 27766
rect 54270 27744 54566 27764
rect 54010 27580 54062 27586
rect 54010 27522 54062 27528
rect 55298 27512 55350 27518
rect 55298 27454 55350 27460
rect 55310 27178 55338 27454
rect 56506 27178 56534 28542
rect 56934 28364 57230 28384
rect 56990 28362 57014 28364
rect 57070 28362 57094 28364
rect 57150 28362 57174 28364
rect 57012 28310 57014 28362
rect 57076 28310 57088 28362
rect 57150 28310 57152 28362
rect 56990 28308 57014 28310
rect 57070 28308 57094 28310
rect 57150 28308 57174 28310
rect 56934 28288 57230 28308
rect 57518 28198 57546 28610
rect 57598 28464 57650 28470
rect 57598 28406 57650 28412
rect 57506 28192 57558 28198
rect 57506 28134 57558 28140
rect 57610 28130 57638 28406
rect 57598 28124 57650 28130
rect 57598 28066 57650 28072
rect 58426 28124 58478 28130
rect 58426 28066 58478 28072
rect 57414 28056 57466 28062
rect 57414 27998 57466 28004
rect 56862 27988 56914 27994
rect 56862 27930 56914 27936
rect 56954 27988 57006 27994
rect 56954 27930 57006 27936
rect 55298 27172 55350 27178
rect 55298 27114 55350 27120
rect 56494 27172 56546 27178
rect 56494 27114 56546 27120
rect 53734 27104 53786 27110
rect 53734 27046 53786 27052
rect 56506 27042 56534 27114
rect 56494 27036 56546 27042
rect 56494 26978 56546 26984
rect 56874 26974 56902 27930
rect 56966 27722 56994 27930
rect 57426 27722 57454 27998
rect 56954 27716 57006 27722
rect 56954 27658 57006 27664
rect 57414 27716 57466 27722
rect 57414 27658 57466 27664
rect 56966 27450 56994 27658
rect 57610 27568 57638 28066
rect 58334 28056 58386 28062
rect 58334 27998 58386 28004
rect 57690 27580 57742 27586
rect 57610 27540 57690 27568
rect 57690 27522 57742 27528
rect 56954 27444 57006 27450
rect 56954 27386 57006 27392
rect 56934 27276 57230 27296
rect 56990 27274 57014 27276
rect 57070 27274 57094 27276
rect 57150 27274 57174 27276
rect 57012 27222 57014 27274
rect 57076 27222 57088 27274
rect 57150 27222 57152 27274
rect 56990 27220 57014 27222
rect 57070 27220 57094 27222
rect 57150 27220 57174 27222
rect 56934 27200 57230 27220
rect 58346 27178 58374 27998
rect 58438 27518 58466 28066
rect 58806 27926 58834 31670
rect 60186 31326 60214 31874
rect 62026 31462 62054 32583
rect 62762 32550 62790 32962
rect 62854 32906 62882 33506
rect 62946 33026 62974 36702
rect 63038 36193 63066 38946
rect 63024 36184 63080 36193
rect 63024 36119 63080 36128
rect 63026 36080 63078 36086
rect 63026 36022 63078 36028
rect 63038 33502 63066 36022
rect 63130 35202 63158 39898
rect 64694 39554 64722 43312
rect 64926 41964 65222 41984
rect 64982 41962 65006 41964
rect 65062 41962 65086 41964
rect 65142 41962 65166 41964
rect 65004 41910 65006 41962
rect 65068 41910 65080 41962
rect 65142 41910 65144 41962
rect 64982 41908 65006 41910
rect 65062 41908 65086 41910
rect 65142 41908 65166 41910
rect 64926 41888 65222 41908
rect 65326 41656 65378 41662
rect 65326 41598 65378 41604
rect 65338 41118 65366 41598
rect 65326 41112 65378 41118
rect 65326 41054 65378 41060
rect 64926 40876 65222 40896
rect 64982 40874 65006 40876
rect 65062 40874 65086 40876
rect 65142 40874 65166 40876
rect 65004 40822 65006 40874
rect 65068 40822 65080 40874
rect 65142 40822 65144 40874
rect 64982 40820 65006 40822
rect 65062 40820 65086 40822
rect 65142 40820 65166 40822
rect 64926 40800 65222 40820
rect 64926 39788 65222 39808
rect 64982 39786 65006 39788
rect 65062 39786 65086 39788
rect 65142 39786 65166 39788
rect 65004 39734 65006 39786
rect 65068 39734 65080 39786
rect 65142 39734 65144 39786
rect 64982 39732 65006 39734
rect 65062 39732 65086 39734
rect 65142 39732 65166 39734
rect 64926 39712 65222 39732
rect 65338 39570 65366 41054
rect 65982 40098 66010 43312
rect 65970 40092 66022 40098
rect 65970 40034 66022 40040
rect 67178 39894 67206 43312
rect 67442 41520 67494 41526
rect 67442 41462 67494 41468
rect 67454 40234 67482 41462
rect 67590 41420 67886 41440
rect 67646 41418 67670 41420
rect 67726 41418 67750 41420
rect 67806 41418 67830 41420
rect 67668 41366 67670 41418
rect 67732 41366 67744 41418
rect 67806 41366 67808 41418
rect 67646 41364 67670 41366
rect 67726 41364 67750 41366
rect 67806 41364 67830 41366
rect 67590 41344 67886 41364
rect 68374 40642 68402 43312
rect 68546 41656 68598 41662
rect 68546 41598 68598 41604
rect 68362 40636 68414 40642
rect 68362 40578 68414 40584
rect 68178 40568 68230 40574
rect 68178 40510 68230 40516
rect 67590 40332 67886 40352
rect 67646 40330 67670 40332
rect 67726 40330 67750 40332
rect 67806 40330 67830 40332
rect 67668 40278 67670 40330
rect 67732 40278 67744 40330
rect 67806 40278 67808 40330
rect 67646 40276 67670 40278
rect 67726 40276 67750 40278
rect 67806 40276 67830 40278
rect 67590 40256 67886 40276
rect 67442 40228 67494 40234
rect 67442 40170 67494 40176
rect 67994 39956 68046 39962
rect 67994 39898 68046 39904
rect 67166 39888 67218 39894
rect 67166 39830 67218 39836
rect 64682 39548 64734 39554
rect 64682 39490 64734 39496
rect 65246 39542 65366 39570
rect 67808 39584 67864 39593
rect 68006 39554 68034 39898
rect 65246 39486 65274 39542
rect 67808 39519 67810 39528
rect 67862 39519 67864 39528
rect 67994 39548 68046 39554
rect 67810 39490 67862 39496
rect 67994 39490 68046 39496
rect 68190 39486 68218 40510
rect 68558 40098 68586 41598
rect 68546 40092 68598 40098
rect 68546 40034 68598 40040
rect 68454 40024 68506 40030
rect 68454 39966 68506 39972
rect 68270 39548 68322 39554
rect 68270 39490 68322 39496
rect 65234 39480 65286 39486
rect 65234 39422 65286 39428
rect 65510 39480 65562 39486
rect 65510 39422 65562 39428
rect 68178 39480 68230 39486
rect 68178 39422 68230 39428
rect 65522 39146 65550 39422
rect 66798 39344 66850 39350
rect 66798 39286 66850 39292
rect 67994 39344 68046 39350
rect 67994 39286 68046 39292
rect 65510 39140 65562 39146
rect 65510 39082 65562 39088
rect 66810 38942 66838 39286
rect 67590 39244 67886 39264
rect 67646 39242 67670 39244
rect 67726 39242 67750 39244
rect 67806 39242 67830 39244
rect 67668 39190 67670 39242
rect 67732 39190 67744 39242
rect 67806 39190 67808 39242
rect 67646 39188 67670 39190
rect 67726 39188 67750 39190
rect 67806 39188 67830 39190
rect 67590 39168 67886 39188
rect 64130 38936 64182 38942
rect 64130 38878 64182 38884
rect 64774 38936 64826 38942
rect 64774 38878 64826 38884
rect 66798 38936 66850 38942
rect 66798 38878 66850 38884
rect 63670 38868 63722 38874
rect 63670 38810 63722 38816
rect 63682 38602 63710 38810
rect 63670 38596 63722 38602
rect 63670 38538 63722 38544
rect 64142 38466 64170 38878
rect 64786 38806 64814 38878
rect 64774 38800 64826 38806
rect 64774 38742 64826 38748
rect 64926 38700 65222 38720
rect 64982 38698 65006 38700
rect 65062 38698 65086 38700
rect 65142 38698 65166 38700
rect 65004 38646 65006 38698
rect 65068 38646 65080 38698
rect 65142 38646 65144 38698
rect 64982 38644 65006 38646
rect 65062 38644 65086 38646
rect 65142 38644 65166 38646
rect 64926 38624 65222 38644
rect 64130 38460 64182 38466
rect 64130 38402 64182 38408
rect 67810 38460 67862 38466
rect 67810 38402 67862 38408
rect 67822 38346 67850 38402
rect 67822 38318 67942 38346
rect 63210 38256 63262 38262
rect 63210 38198 63262 38204
rect 63222 37174 63250 38198
rect 67590 38156 67886 38176
rect 67646 38154 67670 38156
rect 67726 38154 67750 38156
rect 67806 38154 67830 38156
rect 67668 38102 67670 38154
rect 67732 38102 67744 38154
rect 67806 38102 67808 38154
rect 67646 38100 67670 38102
rect 67726 38100 67750 38102
rect 67806 38100 67830 38102
rect 67590 38080 67886 38100
rect 63762 37712 63814 37718
rect 63762 37654 63814 37660
rect 63210 37168 63262 37174
rect 63210 37110 63262 37116
rect 63774 36766 63802 37654
rect 64926 37612 65222 37632
rect 64982 37610 65006 37612
rect 65062 37610 65086 37612
rect 65142 37610 65166 37612
rect 65004 37558 65006 37610
rect 65068 37558 65080 37610
rect 65142 37558 65144 37610
rect 64982 37556 65006 37558
rect 65062 37556 65086 37558
rect 65142 37556 65166 37558
rect 64926 37536 65222 37556
rect 67074 37372 67126 37378
rect 67074 37314 67126 37320
rect 67086 37174 67114 37314
rect 64038 37168 64090 37174
rect 64038 37110 64090 37116
rect 67074 37168 67126 37174
rect 67074 37110 67126 37116
rect 64050 36766 64078 37110
rect 67590 37068 67886 37088
rect 67646 37066 67670 37068
rect 67726 37066 67750 37068
rect 67806 37066 67830 37068
rect 67668 37014 67670 37066
rect 67732 37014 67744 37066
rect 67806 37014 67808 37066
rect 67646 37012 67670 37014
rect 67726 37012 67750 37014
rect 67806 37012 67830 37014
rect 67590 36992 67886 37012
rect 65602 36828 65654 36834
rect 65602 36770 65654 36776
rect 63762 36760 63814 36766
rect 63762 36702 63814 36708
rect 64038 36760 64090 36766
rect 64038 36702 64090 36708
rect 64926 36524 65222 36544
rect 64982 36522 65006 36524
rect 65062 36522 65086 36524
rect 65142 36522 65166 36524
rect 65004 36470 65006 36522
rect 65068 36470 65080 36522
rect 65142 36470 65144 36522
rect 64982 36468 65006 36470
rect 65062 36468 65086 36470
rect 65142 36468 65166 36470
rect 64926 36448 65222 36468
rect 65614 36426 65642 36770
rect 65970 36624 66022 36630
rect 65970 36566 66022 36572
rect 65602 36420 65654 36426
rect 65602 36362 65654 36368
rect 63302 36284 63354 36290
rect 63302 36226 63354 36232
rect 63210 36080 63262 36086
rect 63210 36022 63262 36028
rect 63222 35542 63250 36022
rect 63314 35678 63342 36226
rect 64130 36080 64182 36086
rect 64130 36022 64182 36028
rect 63946 35740 63998 35746
rect 63946 35682 63998 35688
rect 63302 35672 63354 35678
rect 63302 35614 63354 35620
rect 63210 35536 63262 35542
rect 63210 35478 63262 35484
rect 63578 35536 63630 35542
rect 63958 35513 63986 35682
rect 64142 35542 64170 36022
rect 64130 35536 64182 35542
rect 63578 35478 63630 35484
rect 63944 35504 64000 35513
rect 63300 35368 63356 35377
rect 63300 35303 63356 35312
rect 63314 35270 63342 35303
rect 63302 35264 63354 35270
rect 63302 35206 63354 35212
rect 63118 35196 63170 35202
rect 63118 35138 63170 35144
rect 63210 35196 63262 35202
rect 63210 35138 63262 35144
rect 63222 34590 63250 35138
rect 63394 35060 63446 35066
rect 63394 35002 63446 35008
rect 63406 34794 63434 35002
rect 63394 34788 63446 34794
rect 63394 34730 63446 34736
rect 63210 34584 63262 34590
rect 63210 34526 63262 34532
rect 63222 34454 63250 34526
rect 63210 34448 63262 34454
rect 63210 34390 63262 34396
rect 63486 34448 63538 34454
rect 63486 34390 63538 34396
rect 63498 33706 63526 34390
rect 63590 34182 63618 35478
rect 64130 35478 64182 35484
rect 63944 35439 64000 35448
rect 64142 35338 64170 35478
rect 64926 35436 65222 35456
rect 64982 35434 65006 35436
rect 65062 35434 65086 35436
rect 65142 35434 65166 35436
rect 65004 35382 65006 35434
rect 65068 35382 65080 35434
rect 65142 35382 65144 35434
rect 64982 35380 65006 35382
rect 65062 35380 65086 35382
rect 65142 35380 65166 35382
rect 64926 35360 65222 35380
rect 64038 35332 64090 35338
rect 64038 35274 64090 35280
rect 64130 35332 64182 35338
rect 64130 35274 64182 35280
rect 63854 34992 63906 34998
rect 63854 34934 63906 34940
rect 63670 34448 63722 34454
rect 63670 34390 63722 34396
rect 63578 34176 63630 34182
rect 63578 34118 63630 34124
rect 63682 34114 63710 34390
rect 63762 34244 63814 34250
rect 63762 34186 63814 34192
rect 63670 34108 63722 34114
rect 63670 34050 63722 34056
rect 63486 33700 63538 33706
rect 63486 33642 63538 33648
rect 63774 33638 63802 34186
rect 63866 34114 63894 34934
rect 63854 34108 63906 34114
rect 63854 34050 63906 34056
rect 63762 33632 63814 33638
rect 63762 33574 63814 33580
rect 63026 33496 63078 33502
rect 63026 33438 63078 33444
rect 63946 33496 63998 33502
rect 63946 33438 63998 33444
rect 62934 33020 62986 33026
rect 62934 32962 62986 32968
rect 63210 33020 63262 33026
rect 63210 32962 63262 32968
rect 63222 32906 63250 32962
rect 62854 32878 63250 32906
rect 63222 32793 63250 32878
rect 63854 32884 63906 32890
rect 63854 32826 63906 32832
rect 63208 32784 63264 32793
rect 63208 32719 63264 32728
rect 63392 32648 63448 32657
rect 63392 32583 63448 32592
rect 62750 32544 62802 32550
rect 62750 32486 62802 32492
rect 63406 32414 63434 32583
rect 63866 32414 63894 32826
rect 63302 32408 63354 32414
rect 63302 32350 63354 32356
rect 63394 32408 63446 32414
rect 63394 32350 63446 32356
rect 63854 32408 63906 32414
rect 63854 32350 63906 32356
rect 62106 32272 62158 32278
rect 62106 32214 62158 32220
rect 62014 31456 62066 31462
rect 62014 31398 62066 31404
rect 60174 31320 60226 31326
rect 60172 31288 60174 31297
rect 60226 31288 60228 31297
rect 60172 31223 60228 31232
rect 61830 31252 61882 31258
rect 61830 31194 61882 31200
rect 60358 31184 60410 31190
rect 60358 31126 60410 31132
rect 59598 31084 59894 31104
rect 59654 31082 59678 31084
rect 59734 31082 59758 31084
rect 59814 31082 59838 31084
rect 59676 31030 59678 31082
rect 59740 31030 59752 31082
rect 59814 31030 59816 31082
rect 59654 31028 59678 31030
rect 59734 31028 59758 31030
rect 59814 31028 59838 31030
rect 59598 31008 59894 31028
rect 59622 30640 59674 30646
rect 59622 30582 59674 30588
rect 59634 30306 59662 30582
rect 60174 30368 60226 30374
rect 60174 30310 60226 30316
rect 59622 30300 59674 30306
rect 59622 30242 59674 30248
rect 59162 30232 59214 30238
rect 59990 30232 60042 30238
rect 59162 30174 59214 30180
rect 59988 30200 59990 30209
rect 60042 30200 60044 30209
rect 59174 29150 59202 30174
rect 59530 30164 59582 30170
rect 59988 30135 60044 30144
rect 59530 30106 59582 30112
rect 59438 29212 59490 29218
rect 59438 29154 59490 29160
rect 58886 29144 58938 29150
rect 58886 29086 58938 29092
rect 59162 29144 59214 29150
rect 59162 29086 59214 29092
rect 58898 29014 58926 29086
rect 59450 29082 59478 29154
rect 59438 29076 59490 29082
rect 59438 29018 59490 29024
rect 58886 29008 58938 29014
rect 58886 28950 58938 28956
rect 59542 28674 59570 30106
rect 59598 29996 59894 30016
rect 59654 29994 59678 29996
rect 59734 29994 59758 29996
rect 59814 29994 59838 29996
rect 59676 29942 59678 29994
rect 59740 29942 59752 29994
rect 59814 29942 59816 29994
rect 59654 29940 59678 29942
rect 59734 29940 59758 29942
rect 59814 29940 59838 29942
rect 59598 29920 59894 29940
rect 60186 29898 60214 30310
rect 60370 29898 60398 31126
rect 61278 30708 61330 30714
rect 61278 30650 61330 30656
rect 60174 29892 60226 29898
rect 60174 29834 60226 29840
rect 60358 29892 60410 29898
rect 60358 29834 60410 29840
rect 61186 29892 61238 29898
rect 61186 29834 61238 29840
rect 60186 29286 60214 29834
rect 61198 29626 61226 29834
rect 61290 29694 61318 30650
rect 61278 29688 61330 29694
rect 61278 29630 61330 29636
rect 60450 29620 60502 29626
rect 60450 29562 60502 29568
rect 61186 29620 61238 29626
rect 61186 29562 61238 29568
rect 60358 29348 60410 29354
rect 60358 29290 60410 29296
rect 60174 29280 60226 29286
rect 60370 29257 60398 29290
rect 60174 29222 60226 29228
rect 60356 29248 60412 29257
rect 60356 29183 60412 29192
rect 60462 29150 60490 29562
rect 60726 29348 60778 29354
rect 60726 29290 60778 29296
rect 60450 29144 60502 29150
rect 60450 29086 60502 29092
rect 60738 29082 60766 29290
rect 60726 29076 60778 29082
rect 60726 29018 60778 29024
rect 59598 28908 59894 28928
rect 59654 28906 59678 28908
rect 59734 28906 59758 28908
rect 59814 28906 59838 28908
rect 59676 28854 59678 28906
rect 59740 28854 59752 28906
rect 59814 28854 59816 28906
rect 59654 28852 59678 28854
rect 59734 28852 59758 28854
rect 59814 28852 59838 28854
rect 59598 28832 59894 28852
rect 59530 28668 59582 28674
rect 59530 28610 59582 28616
rect 61198 28606 61226 29562
rect 61842 29218 61870 31194
rect 62026 30850 62054 31398
rect 62118 30918 62146 32214
rect 63314 32113 63342 32350
rect 63300 32104 63356 32113
rect 63300 32039 63356 32048
rect 63958 31870 63986 33438
rect 64050 32634 64078 35274
rect 65878 35196 65930 35202
rect 65878 35138 65930 35144
rect 64774 34720 64826 34726
rect 64774 34662 64826 34668
rect 64128 34552 64184 34561
rect 64128 34487 64184 34496
rect 64142 34182 64170 34487
rect 64786 34250 64814 34662
rect 64926 34348 65222 34368
rect 64982 34346 65006 34348
rect 65062 34346 65086 34348
rect 65142 34346 65166 34348
rect 65004 34294 65006 34346
rect 65068 34294 65080 34346
rect 65142 34294 65144 34346
rect 64982 34292 65006 34294
rect 65062 34292 65086 34294
rect 65142 34292 65166 34294
rect 64926 34272 65222 34292
rect 64774 34244 64826 34250
rect 64774 34186 64826 34192
rect 64130 34176 64182 34182
rect 64130 34118 64182 34124
rect 65602 34040 65654 34046
rect 65602 33982 65654 33988
rect 64130 33972 64182 33978
rect 64130 33914 64182 33920
rect 64142 33706 64170 33914
rect 64130 33700 64182 33706
rect 64130 33642 64182 33648
rect 65510 33428 65562 33434
rect 65510 33370 65562 33376
rect 64926 33260 65222 33280
rect 64982 33258 65006 33260
rect 65062 33258 65086 33260
rect 65142 33258 65166 33260
rect 65004 33206 65006 33258
rect 65068 33206 65080 33258
rect 65142 33206 65144 33258
rect 64982 33204 65006 33206
rect 65062 33204 65086 33206
rect 65142 33204 65166 33206
rect 64926 33184 65222 33204
rect 65522 33162 65550 33370
rect 65418 33156 65470 33162
rect 65418 33098 65470 33104
rect 65510 33156 65562 33162
rect 65510 33098 65562 33104
rect 65050 33020 65102 33026
rect 65102 32980 65182 33008
rect 65050 32962 65102 32968
rect 64680 32920 64736 32929
rect 64130 32884 64182 32890
rect 64130 32826 64182 32832
rect 64602 32864 64680 32872
rect 64602 32844 64682 32864
rect 64142 32793 64170 32826
rect 64128 32784 64184 32793
rect 64128 32719 64184 32728
rect 64050 32606 64170 32634
rect 64142 31870 64170 32606
rect 64498 32544 64550 32550
rect 64498 32486 64550 32492
rect 64510 32249 64538 32486
rect 64602 32346 64630 32844
rect 64734 32855 64736 32864
rect 65050 32884 65102 32890
rect 64682 32826 64734 32832
rect 65050 32826 65102 32832
rect 64680 32648 64736 32657
rect 64680 32583 64736 32592
rect 64694 32482 64722 32583
rect 64682 32476 64734 32482
rect 64682 32418 64734 32424
rect 64590 32340 64642 32346
rect 64590 32282 64642 32288
rect 64682 32272 64734 32278
rect 64496 32240 64552 32249
rect 65062 32260 65090 32826
rect 65154 32346 65182 32980
rect 65234 32816 65286 32822
rect 65234 32758 65286 32764
rect 65246 32414 65274 32758
rect 65234 32408 65286 32414
rect 65234 32350 65286 32356
rect 65430 32346 65458 33098
rect 65614 32958 65642 33982
rect 65786 33020 65838 33026
rect 65786 32962 65838 32968
rect 65602 32952 65654 32958
rect 65602 32894 65654 32900
rect 65798 32618 65826 32962
rect 65786 32612 65838 32618
rect 65786 32554 65838 32560
rect 65142 32340 65194 32346
rect 65142 32282 65194 32288
rect 65418 32340 65470 32346
rect 65418 32282 65470 32288
rect 64682 32214 64734 32220
rect 64786 32232 65090 32260
rect 65510 32272 65562 32278
rect 64496 32175 64552 32184
rect 64694 32113 64722 32214
rect 64680 32104 64736 32113
rect 64680 32039 64736 32048
rect 64694 31870 64722 32039
rect 63946 31864 63998 31870
rect 63946 31806 63998 31812
rect 64130 31864 64182 31870
rect 64130 31806 64182 31812
rect 64682 31864 64734 31870
rect 64682 31806 64734 31812
rect 63210 31728 63262 31734
rect 63210 31670 63262 31676
rect 63394 31728 63446 31734
rect 63394 31670 63446 31676
rect 62262 31628 62558 31648
rect 62318 31626 62342 31628
rect 62398 31626 62422 31628
rect 62478 31626 62502 31628
rect 62340 31574 62342 31626
rect 62404 31574 62416 31626
rect 62478 31574 62480 31626
rect 62318 31572 62342 31574
rect 62398 31572 62422 31574
rect 62478 31572 62502 31574
rect 62262 31552 62558 31572
rect 63222 31394 63250 31670
rect 63406 31530 63434 31670
rect 63394 31524 63446 31530
rect 63394 31466 63446 31472
rect 63210 31388 63262 31394
rect 63210 31330 63262 31336
rect 62750 31320 62802 31326
rect 62750 31262 62802 31268
rect 62106 30912 62158 30918
rect 62106 30854 62158 30860
rect 62014 30844 62066 30850
rect 62014 30786 62066 30792
rect 62658 30844 62710 30850
rect 62658 30786 62710 30792
rect 62262 30540 62558 30560
rect 62318 30538 62342 30540
rect 62398 30538 62422 30540
rect 62478 30538 62502 30540
rect 62340 30486 62342 30538
rect 62404 30486 62416 30538
rect 62478 30486 62480 30538
rect 62318 30484 62342 30486
rect 62398 30484 62422 30486
rect 62478 30484 62502 30486
rect 62262 30464 62558 30484
rect 62106 30436 62158 30442
rect 62106 30378 62158 30384
rect 62118 30345 62146 30378
rect 62104 30336 62160 30345
rect 62104 30271 62160 30280
rect 62290 30300 62342 30306
rect 62290 30242 62342 30248
rect 62302 29626 62330 30242
rect 62670 30238 62698 30786
rect 62658 30232 62710 30238
rect 62658 30174 62710 30180
rect 62566 30164 62618 30170
rect 62566 30106 62618 30112
rect 62290 29620 62342 29626
rect 62290 29562 62342 29568
rect 62578 29540 62606 30106
rect 62762 29694 62790 31262
rect 63394 30912 63446 30918
rect 63394 30854 63446 30860
rect 63026 30844 63078 30850
rect 63026 30786 63078 30792
rect 63038 30374 63066 30786
rect 63026 30368 63078 30374
rect 63026 30310 63078 30316
rect 63118 30164 63170 30170
rect 63118 30106 63170 30112
rect 63130 29762 63158 30106
rect 63406 30102 63434 30854
rect 63946 30164 63998 30170
rect 63946 30106 63998 30112
rect 63394 30096 63446 30102
rect 63394 30038 63446 30044
rect 63118 29756 63170 29762
rect 63118 29698 63170 29704
rect 62750 29688 62802 29694
rect 62750 29630 62802 29636
rect 63958 29558 63986 30106
rect 62842 29552 62894 29558
rect 62578 29512 62790 29540
rect 62262 29452 62558 29472
rect 62318 29450 62342 29452
rect 62398 29450 62422 29452
rect 62478 29450 62502 29452
rect 62340 29398 62342 29450
rect 62404 29398 62416 29450
rect 62478 29398 62480 29450
rect 62318 29396 62342 29398
rect 62398 29396 62422 29398
rect 62478 29396 62502 29398
rect 62262 29376 62558 29396
rect 61830 29212 61882 29218
rect 61830 29154 61882 29160
rect 62106 29076 62158 29082
rect 62106 29018 62158 29024
rect 61186 28600 61238 28606
rect 61186 28542 61238 28548
rect 59806 28464 59858 28470
rect 59806 28406 59858 28412
rect 59818 28266 59846 28406
rect 59806 28260 59858 28266
rect 59806 28202 59858 28208
rect 58794 27920 58846 27926
rect 58794 27862 58846 27868
rect 58806 27654 58834 27862
rect 59598 27820 59894 27840
rect 59654 27818 59678 27820
rect 59734 27818 59758 27820
rect 59814 27818 59838 27820
rect 59676 27766 59678 27818
rect 59740 27766 59752 27818
rect 59814 27766 59816 27818
rect 59654 27764 59678 27766
rect 59734 27764 59758 27766
rect 59814 27764 59838 27766
rect 59598 27744 59894 27764
rect 58794 27648 58846 27654
rect 58794 27590 58846 27596
rect 58426 27512 58478 27518
rect 58426 27454 58478 27460
rect 58334 27172 58386 27178
rect 58334 27114 58386 27120
rect 61198 27042 61226 28542
rect 62118 27654 62146 29018
rect 62658 29008 62710 29014
rect 62658 28950 62710 28956
rect 62670 28538 62698 28950
rect 62762 28742 62790 29512
rect 62842 29494 62894 29500
rect 63946 29552 63998 29558
rect 63946 29494 63998 29500
rect 62854 29150 62882 29494
rect 62934 29348 62986 29354
rect 62934 29290 62986 29296
rect 62842 29144 62894 29150
rect 62842 29086 62894 29092
rect 62750 28736 62802 28742
rect 62750 28678 62802 28684
rect 62658 28532 62710 28538
rect 62658 28474 62710 28480
rect 62262 28364 62558 28384
rect 62318 28362 62342 28364
rect 62398 28362 62422 28364
rect 62478 28362 62502 28364
rect 62340 28310 62342 28362
rect 62404 28310 62416 28362
rect 62478 28310 62480 28362
rect 62318 28308 62342 28310
rect 62398 28308 62422 28310
rect 62478 28308 62502 28310
rect 62262 28288 62558 28308
rect 62658 28056 62710 28062
rect 62762 28044 62790 28678
rect 62946 28554 62974 29290
rect 63210 29008 63262 29014
rect 63210 28950 63262 28956
rect 63222 28674 63250 28950
rect 63210 28668 63262 28674
rect 63210 28610 63262 28616
rect 63302 28668 63354 28674
rect 63302 28610 63354 28616
rect 63314 28554 63342 28610
rect 62946 28526 63342 28554
rect 62946 28062 62974 28526
rect 63958 28266 63986 29494
rect 64496 29248 64552 29257
rect 64496 29183 64552 29192
rect 64510 29082 64538 29183
rect 64498 29076 64550 29082
rect 64498 29018 64550 29024
rect 64406 29008 64458 29014
rect 64406 28950 64458 28956
rect 64418 28742 64446 28950
rect 64406 28736 64458 28742
rect 64406 28678 64458 28684
rect 64222 28600 64274 28606
rect 64222 28542 64274 28548
rect 64130 28464 64182 28470
rect 64130 28406 64182 28412
rect 63946 28260 63998 28266
rect 63946 28202 63998 28208
rect 62710 28016 62790 28044
rect 62934 28056 62986 28062
rect 62658 27998 62710 28004
rect 62934 27998 62986 28004
rect 64142 27994 64170 28406
rect 64234 28266 64262 28542
rect 64786 28538 64814 32232
rect 65510 32214 65562 32220
rect 64926 32172 65222 32192
rect 64982 32170 65006 32172
rect 65062 32170 65086 32172
rect 65142 32170 65166 32172
rect 65004 32118 65006 32170
rect 65068 32118 65080 32170
rect 65142 32118 65144 32170
rect 64982 32116 65006 32118
rect 65062 32116 65086 32118
rect 65142 32116 65166 32118
rect 64926 32096 65222 32116
rect 65522 31977 65550 32214
rect 65508 31968 65564 31977
rect 65508 31903 65564 31912
rect 65890 31190 65918 35138
rect 65982 34998 66010 36566
rect 66522 36148 66574 36154
rect 66522 36090 66574 36096
rect 65970 34992 66022 34998
rect 65970 34934 66022 34940
rect 66062 33972 66114 33978
rect 66062 33914 66114 33920
rect 65968 33736 66024 33745
rect 65968 33671 65970 33680
rect 66022 33671 66024 33680
rect 65970 33642 66022 33648
rect 66074 33638 66102 33914
rect 66062 33632 66114 33638
rect 66062 33574 66114 33580
rect 65970 33564 66022 33570
rect 65970 33506 66022 33512
rect 65982 33366 66010 33506
rect 65970 33360 66022 33366
rect 65970 33302 66022 33308
rect 65970 33156 66022 33162
rect 65970 33098 66022 33104
rect 65982 32822 66010 33098
rect 66534 33026 66562 36090
rect 67590 35980 67886 36000
rect 67646 35978 67670 35980
rect 67726 35978 67750 35980
rect 67806 35978 67830 35980
rect 67668 35926 67670 35978
rect 67732 35926 67744 35978
rect 67806 35926 67808 35978
rect 67646 35924 67670 35926
rect 67726 35924 67750 35926
rect 67806 35924 67830 35926
rect 67590 35904 67886 35924
rect 67442 35808 67494 35814
rect 67442 35750 67494 35756
rect 66890 35604 66942 35610
rect 66942 35564 67022 35592
rect 66890 35546 66942 35552
rect 66522 33020 66574 33026
rect 66522 32962 66574 32968
rect 66890 32952 66942 32958
rect 66890 32894 66942 32900
rect 65970 32816 66022 32822
rect 66706 32816 66758 32822
rect 65970 32758 66022 32764
rect 66704 32784 66706 32793
rect 66758 32784 66760 32793
rect 66704 32719 66760 32728
rect 65970 32544 66022 32550
rect 65970 32486 66022 32492
rect 65982 32414 66010 32486
rect 65970 32408 66022 32414
rect 65970 32350 66022 32356
rect 66902 32346 66930 32894
rect 66890 32340 66942 32346
rect 66890 32282 66942 32288
rect 66902 31734 66930 32282
rect 66890 31728 66942 31734
rect 66890 31670 66942 31676
rect 65878 31184 65930 31190
rect 65878 31126 65930 31132
rect 66062 31184 66114 31190
rect 66062 31126 66114 31132
rect 64926 31084 65222 31104
rect 64982 31082 65006 31084
rect 65062 31082 65086 31084
rect 65142 31082 65166 31084
rect 65004 31030 65006 31082
rect 65068 31030 65080 31082
rect 65142 31030 65144 31082
rect 64982 31028 65006 31030
rect 65062 31028 65086 31030
rect 65142 31028 65166 31030
rect 64926 31008 65222 31028
rect 65416 30336 65472 30345
rect 65416 30271 65472 30280
rect 65430 30170 65458 30271
rect 65786 30232 65838 30238
rect 65786 30174 65838 30180
rect 65418 30164 65470 30170
rect 65418 30106 65470 30112
rect 64926 29996 65222 30016
rect 64982 29994 65006 29996
rect 65062 29994 65086 29996
rect 65142 29994 65166 29996
rect 65004 29942 65006 29994
rect 65068 29942 65080 29994
rect 65142 29942 65144 29994
rect 64982 29940 65006 29942
rect 65062 29940 65086 29942
rect 65142 29940 65166 29942
rect 64926 29920 65222 29940
rect 65798 29830 65826 30174
rect 65786 29824 65838 29830
rect 65786 29766 65838 29772
rect 65326 29756 65378 29762
rect 65326 29698 65378 29704
rect 65338 29150 65366 29698
rect 65326 29144 65378 29150
rect 65326 29086 65378 29092
rect 64926 28908 65222 28928
rect 64982 28906 65006 28908
rect 65062 28906 65086 28908
rect 65142 28906 65166 28908
rect 65004 28854 65006 28906
rect 65068 28854 65080 28906
rect 65142 28854 65144 28906
rect 64982 28852 65006 28854
rect 65062 28852 65086 28854
rect 65142 28852 65166 28854
rect 64926 28832 65222 28852
rect 64774 28532 64826 28538
rect 64774 28474 64826 28480
rect 64222 28260 64274 28266
rect 64222 28202 64274 28208
rect 65890 28198 65918 31126
rect 66074 30714 66102 31126
rect 66994 30782 67022 35564
rect 67454 34130 67482 35750
rect 67914 35746 67942 38318
rect 68006 37922 68034 39286
rect 68282 39146 68310 39490
rect 68270 39140 68322 39146
rect 68270 39082 68322 39088
rect 68362 38800 68414 38806
rect 68362 38742 68414 38748
rect 68374 38466 68402 38742
rect 68362 38460 68414 38466
rect 68362 38402 68414 38408
rect 68270 38256 68322 38262
rect 68270 38198 68322 38204
rect 68282 37922 68310 38198
rect 67994 37916 68046 37922
rect 67994 37858 68046 37864
rect 68270 37916 68322 37922
rect 68270 37858 68322 37864
rect 68176 37408 68232 37417
rect 68176 37343 68232 37352
rect 68362 37372 68414 37378
rect 68190 37310 68218 37343
rect 68362 37314 68414 37320
rect 68178 37304 68230 37310
rect 68178 37246 68230 37252
rect 68270 37304 68322 37310
rect 68270 37246 68322 37252
rect 68282 37156 68310 37246
rect 68098 37128 68310 37156
rect 68098 36902 68126 37128
rect 68086 36896 68138 36902
rect 68086 36838 68138 36844
rect 68178 36896 68230 36902
rect 68178 36838 68230 36844
rect 68190 36426 68218 36838
rect 68374 36766 68402 37314
rect 68466 37242 68494 39966
rect 68638 38936 68690 38942
rect 68638 38878 68690 38884
rect 69006 38936 69058 38942
rect 69006 38878 69058 38884
rect 68650 38602 68678 38878
rect 68638 38596 68690 38602
rect 68638 38538 68690 38544
rect 68546 38256 68598 38262
rect 68546 38198 68598 38204
rect 68558 37310 68586 38198
rect 68546 37304 68598 37310
rect 68546 37246 68598 37252
rect 68454 37236 68506 37242
rect 68454 37178 68506 37184
rect 68650 37174 68678 38538
rect 69018 37990 69046 38878
rect 69098 38460 69150 38466
rect 69098 38402 69150 38408
rect 69110 38058 69138 38402
rect 69662 38262 69690 43312
rect 70254 41964 70550 41984
rect 70310 41962 70334 41964
rect 70390 41962 70414 41964
rect 70470 41962 70494 41964
rect 70332 41910 70334 41962
rect 70396 41910 70408 41962
rect 70470 41910 70472 41962
rect 70310 41908 70334 41910
rect 70390 41908 70414 41910
rect 70470 41908 70494 41910
rect 70254 41888 70550 41908
rect 70858 40930 70886 43312
rect 70858 40902 71254 40930
rect 70254 40876 70550 40896
rect 70310 40874 70334 40876
rect 70390 40874 70414 40876
rect 70470 40874 70494 40876
rect 70332 40822 70334 40874
rect 70396 40822 70408 40874
rect 70470 40822 70472 40874
rect 70310 40820 70334 40822
rect 70390 40820 70414 40822
rect 70470 40820 70494 40822
rect 70254 40800 70550 40820
rect 71122 40772 71174 40778
rect 71122 40714 71174 40720
rect 70754 40636 70806 40642
rect 70754 40578 70806 40584
rect 69926 40568 69978 40574
rect 69926 40510 69978 40516
rect 69938 39350 69966 40510
rect 70254 39788 70550 39808
rect 70310 39786 70334 39788
rect 70390 39786 70414 39788
rect 70470 39786 70494 39788
rect 70332 39734 70334 39786
rect 70396 39734 70408 39786
rect 70470 39734 70472 39786
rect 70310 39732 70334 39734
rect 70390 39732 70414 39734
rect 70470 39732 70494 39734
rect 70254 39712 70550 39732
rect 70766 39622 70794 40578
rect 71134 39894 71162 40714
rect 71226 40642 71254 40902
rect 71214 40636 71266 40642
rect 71214 40578 71266 40584
rect 72054 40098 72082 43312
rect 73250 41526 73278 43312
rect 73238 41520 73290 41526
rect 73238 41462 73290 41468
rect 72918 41420 73214 41440
rect 72974 41418 72998 41420
rect 73054 41418 73078 41420
rect 73134 41418 73158 41420
rect 72996 41366 72998 41418
rect 73060 41366 73072 41418
rect 73134 41366 73136 41418
rect 72974 41364 72998 41366
rect 73054 41364 73078 41366
rect 73134 41364 73158 41366
rect 72918 41344 73214 41364
rect 73698 41112 73750 41118
rect 73698 41054 73750 41060
rect 73882 41112 73934 41118
rect 73882 41054 73934 41060
rect 73710 40574 73738 41054
rect 73606 40568 73658 40574
rect 73606 40510 73658 40516
rect 73698 40568 73750 40574
rect 73698 40510 73750 40516
rect 72226 40432 72278 40438
rect 72226 40374 72278 40380
rect 72238 40234 72266 40374
rect 72918 40332 73214 40352
rect 72974 40330 72998 40332
rect 73054 40330 73078 40332
rect 73134 40330 73158 40332
rect 72996 40278 72998 40330
rect 73060 40278 73072 40330
rect 73134 40278 73136 40330
rect 72974 40276 72998 40278
rect 73054 40276 73078 40278
rect 73134 40276 73158 40278
rect 72918 40256 73214 40276
rect 72226 40228 72278 40234
rect 72226 40170 72278 40176
rect 72042 40092 72094 40098
rect 72042 40034 72094 40040
rect 73330 40092 73382 40098
rect 73330 40034 73382 40040
rect 71214 40024 71266 40030
rect 71214 39966 71266 39972
rect 71582 40024 71634 40030
rect 71582 39966 71634 39972
rect 72870 40024 72922 40030
rect 72870 39966 72922 39972
rect 71122 39888 71174 39894
rect 71122 39830 71174 39836
rect 70754 39616 70806 39622
rect 70754 39558 70806 39564
rect 70846 39548 70898 39554
rect 70846 39490 70898 39496
rect 69926 39344 69978 39350
rect 69926 39286 69978 39292
rect 70858 39332 70886 39490
rect 71226 39486 71254 39966
rect 71214 39480 71266 39486
rect 71214 39422 71266 39428
rect 71306 39344 71358 39350
rect 70858 39304 71306 39332
rect 69650 38256 69702 38262
rect 69650 38198 69702 38204
rect 69098 38052 69150 38058
rect 69098 37994 69150 38000
rect 69006 37984 69058 37990
rect 69006 37926 69058 37932
rect 69018 37446 69046 37926
rect 69938 37922 69966 39286
rect 70858 39078 70886 39304
rect 71306 39286 71358 39292
rect 70846 39072 70898 39078
rect 70846 39014 70898 39020
rect 70254 38700 70550 38720
rect 70310 38698 70334 38700
rect 70390 38698 70414 38700
rect 70470 38698 70494 38700
rect 70332 38646 70334 38698
rect 70396 38646 70408 38698
rect 70470 38646 70472 38698
rect 70310 38644 70334 38646
rect 70390 38644 70414 38646
rect 70470 38644 70494 38646
rect 70254 38624 70550 38644
rect 69926 37916 69978 37922
rect 69926 37858 69978 37864
rect 70254 37612 70550 37632
rect 70310 37610 70334 37612
rect 70390 37610 70414 37612
rect 70470 37610 70494 37612
rect 70332 37558 70334 37610
rect 70396 37558 70408 37610
rect 70470 37558 70472 37610
rect 70310 37556 70334 37558
rect 70390 37556 70414 37558
rect 70470 37556 70494 37558
rect 70254 37536 70550 37556
rect 71594 37446 71622 39966
rect 72778 39956 72830 39962
rect 72778 39898 72830 39904
rect 72410 38596 72462 38602
rect 72410 38538 72462 38544
rect 72422 38482 72450 38538
rect 72422 38466 72634 38482
rect 72422 38460 72646 38466
rect 72422 38454 72594 38460
rect 72594 38402 72646 38408
rect 72226 38256 72278 38262
rect 72226 38198 72278 38204
rect 72238 38058 72266 38198
rect 72226 38052 72278 38058
rect 72226 37994 72278 38000
rect 72226 37712 72278 37718
rect 72226 37654 72278 37660
rect 69006 37440 69058 37446
rect 71582 37440 71634 37446
rect 69006 37382 69058 37388
rect 69280 37408 69336 37417
rect 69190 37372 69242 37378
rect 71582 37382 71634 37388
rect 69280 37343 69282 37352
rect 69190 37314 69242 37320
rect 69334 37343 69336 37352
rect 69650 37372 69702 37378
rect 69282 37314 69334 37320
rect 69650 37314 69702 37320
rect 69202 37281 69230 37314
rect 69188 37272 69244 37281
rect 69188 37207 69244 37216
rect 69282 37236 69334 37242
rect 69282 37178 69334 37184
rect 68638 37168 68690 37174
rect 68638 37110 68690 37116
rect 68730 36896 68782 36902
rect 68730 36838 68782 36844
rect 68742 36766 68770 36838
rect 69190 36828 69242 36834
rect 69190 36770 69242 36776
rect 68362 36760 68414 36766
rect 68362 36702 68414 36708
rect 68730 36760 68782 36766
rect 68730 36702 68782 36708
rect 68912 36728 68968 36737
rect 68178 36420 68230 36426
rect 68178 36362 68230 36368
rect 68374 35814 68402 36702
rect 68912 36663 68914 36672
rect 68966 36663 68968 36672
rect 68914 36634 68966 36640
rect 69202 36290 69230 36770
rect 69190 36284 69242 36290
rect 69190 36226 69242 36232
rect 69006 36080 69058 36086
rect 69006 36022 69058 36028
rect 68362 35808 68414 35814
rect 67992 35776 68048 35785
rect 67902 35740 67954 35746
rect 68362 35750 68414 35756
rect 67992 35711 68048 35720
rect 67902 35682 67954 35688
rect 67902 35128 67954 35134
rect 67902 35070 67954 35076
rect 67590 34892 67886 34912
rect 67646 34890 67670 34892
rect 67726 34890 67750 34892
rect 67806 34890 67830 34892
rect 67668 34838 67670 34890
rect 67732 34838 67744 34890
rect 67806 34838 67808 34890
rect 67646 34836 67670 34838
rect 67726 34836 67750 34838
rect 67806 34836 67830 34838
rect 67590 34816 67886 34836
rect 67810 34584 67862 34590
rect 67810 34526 67862 34532
rect 67914 34538 67942 35070
rect 68006 34726 68034 35711
rect 68914 35672 68966 35678
rect 69018 35626 69046 36022
rect 69294 35746 69322 37178
rect 69662 36306 69690 37314
rect 70018 37168 70070 37174
rect 70018 37110 70070 37116
rect 69662 36278 69782 36306
rect 69650 36216 69702 36222
rect 69650 36158 69702 36164
rect 69374 36148 69426 36154
rect 69374 36090 69426 36096
rect 69282 35740 69334 35746
rect 69282 35682 69334 35688
rect 68966 35620 69046 35626
rect 68914 35614 69046 35620
rect 68926 35598 69046 35614
rect 68362 35196 68414 35202
rect 68362 35138 68414 35144
rect 68178 35128 68230 35134
rect 68178 35070 68230 35076
rect 67994 34720 68046 34726
rect 67994 34662 68046 34668
rect 68190 34590 68218 35070
rect 68374 34998 68402 35138
rect 68362 34992 68414 34998
rect 68362 34934 68414 34940
rect 68178 34584 68230 34590
rect 67822 34436 67850 34526
rect 67914 34510 68034 34538
rect 68178 34526 68230 34532
rect 68270 34584 68322 34590
rect 68270 34526 68322 34532
rect 67822 34408 67942 34436
rect 67454 34114 67666 34130
rect 67454 34108 67678 34114
rect 67454 34102 67626 34108
rect 67626 34050 67678 34056
rect 67914 33978 67942 34408
rect 67902 33972 67954 33978
rect 67902 33914 67954 33920
rect 67590 33804 67886 33824
rect 67646 33802 67670 33804
rect 67726 33802 67750 33804
rect 67806 33802 67830 33804
rect 67668 33750 67670 33802
rect 67732 33750 67744 33802
rect 67806 33750 67808 33802
rect 67646 33748 67670 33750
rect 67726 33748 67750 33750
rect 67806 33748 67830 33750
rect 67590 33728 67886 33748
rect 67534 33360 67586 33366
rect 67534 33302 67586 33308
rect 67074 33020 67126 33026
rect 67074 32962 67126 32968
rect 67442 33020 67494 33026
rect 67442 32962 67494 32968
rect 67086 32929 67114 32962
rect 67454 32929 67482 32962
rect 67072 32920 67128 32929
rect 67072 32855 67128 32864
rect 67440 32920 67496 32929
rect 67440 32855 67496 32864
rect 67546 32804 67574 33302
rect 67270 32776 67574 32804
rect 67270 32634 67298 32776
rect 67590 32716 67886 32736
rect 67646 32714 67670 32716
rect 67726 32714 67750 32716
rect 67806 32714 67830 32716
rect 67668 32662 67670 32714
rect 67732 32662 67744 32714
rect 67806 32662 67808 32714
rect 67646 32660 67670 32662
rect 67726 32660 67750 32662
rect 67806 32660 67830 32662
rect 67590 32640 67886 32660
rect 67086 32606 67298 32634
rect 66522 30776 66574 30782
rect 66522 30718 66574 30724
rect 66798 30776 66850 30782
rect 66982 30776 67034 30782
rect 66798 30718 66850 30724
rect 66902 30736 66982 30764
rect 66062 30708 66114 30714
rect 66062 30650 66114 30656
rect 66074 30374 66102 30650
rect 66062 30368 66114 30374
rect 66062 30310 66114 30316
rect 66534 30306 66562 30718
rect 66522 30300 66574 30306
rect 66522 30242 66574 30248
rect 66614 30300 66666 30306
rect 66614 30242 66666 30248
rect 66626 30209 66654 30242
rect 66612 30200 66668 30209
rect 66612 30135 66668 30144
rect 66810 29898 66838 30718
rect 66902 30238 66930 30736
rect 66982 30718 67034 30724
rect 66890 30232 66942 30238
rect 66890 30174 66942 30180
rect 66798 29892 66850 29898
rect 66798 29834 66850 29840
rect 65878 28192 65930 28198
rect 65878 28134 65930 28140
rect 64130 27988 64182 27994
rect 64130 27930 64182 27936
rect 62106 27648 62158 27654
rect 62106 27590 62158 27596
rect 64142 27586 64170 27930
rect 64926 27820 65222 27840
rect 64982 27818 65006 27820
rect 65062 27818 65086 27820
rect 65142 27818 65166 27820
rect 65004 27766 65006 27818
rect 65068 27766 65080 27818
rect 65142 27766 65144 27818
rect 64982 27764 65006 27766
rect 65062 27764 65086 27766
rect 65142 27764 65166 27766
rect 64926 27744 65222 27764
rect 63302 27580 63354 27586
rect 63302 27522 63354 27528
rect 64130 27580 64182 27586
rect 64130 27522 64182 27528
rect 62658 27512 62710 27518
rect 62658 27454 62710 27460
rect 62262 27276 62558 27296
rect 62318 27274 62342 27276
rect 62398 27274 62422 27276
rect 62478 27274 62502 27276
rect 62340 27222 62342 27274
rect 62404 27222 62416 27274
rect 62478 27222 62480 27274
rect 62318 27220 62342 27222
rect 62398 27220 62422 27222
rect 62478 27220 62502 27222
rect 62262 27200 62558 27220
rect 62670 27042 62698 27454
rect 63314 27042 63342 27522
rect 63394 27512 63446 27518
rect 63394 27454 63446 27460
rect 63406 27110 63434 27454
rect 63394 27104 63446 27110
rect 63394 27046 63446 27052
rect 64142 27042 64170 27522
rect 67086 27518 67114 32606
rect 67914 32521 67942 33914
rect 67900 32512 67956 32521
rect 67900 32447 67956 32456
rect 67164 32376 67220 32385
rect 67164 32311 67220 32320
rect 67178 30170 67206 32311
rect 67590 31628 67886 31648
rect 67646 31626 67670 31628
rect 67726 31626 67750 31628
rect 67806 31626 67830 31628
rect 67668 31574 67670 31626
rect 67732 31574 67744 31626
rect 67806 31574 67808 31626
rect 67646 31572 67670 31574
rect 67726 31572 67750 31574
rect 67806 31572 67830 31574
rect 67590 31552 67886 31572
rect 67902 31456 67954 31462
rect 67902 31398 67954 31404
rect 67258 30640 67310 30646
rect 67258 30582 67310 30588
rect 67270 30170 67298 30582
rect 67590 30540 67886 30560
rect 67646 30538 67670 30540
rect 67726 30538 67750 30540
rect 67806 30538 67830 30540
rect 67668 30486 67670 30538
rect 67732 30486 67744 30538
rect 67806 30486 67808 30538
rect 67646 30484 67670 30486
rect 67726 30484 67750 30486
rect 67806 30484 67830 30486
rect 67590 30464 67886 30484
rect 67350 30436 67402 30442
rect 67350 30378 67402 30384
rect 67166 30164 67218 30170
rect 67166 30106 67218 30112
rect 67258 30164 67310 30170
rect 67258 30106 67310 30112
rect 67166 29552 67218 29558
rect 67166 29494 67218 29500
rect 67178 28674 67206 29494
rect 67270 29354 67298 30106
rect 67362 29558 67390 30378
rect 67718 30096 67770 30102
rect 67718 30038 67770 30044
rect 67730 29762 67758 30038
rect 67442 29756 67494 29762
rect 67442 29698 67494 29704
rect 67718 29756 67770 29762
rect 67718 29698 67770 29704
rect 67350 29552 67402 29558
rect 67350 29494 67402 29500
rect 67258 29348 67310 29354
rect 67258 29290 67310 29296
rect 67454 29218 67482 29698
rect 67590 29452 67886 29472
rect 67646 29450 67670 29452
rect 67726 29450 67750 29452
rect 67806 29450 67830 29452
rect 67668 29398 67670 29450
rect 67732 29398 67744 29450
rect 67806 29398 67808 29450
rect 67646 29396 67670 29398
rect 67726 29396 67750 29398
rect 67806 29396 67830 29398
rect 67590 29376 67886 29396
rect 67442 29212 67494 29218
rect 67442 29154 67494 29160
rect 67914 29150 67942 31398
rect 67902 29144 67954 29150
rect 67902 29086 67954 29092
rect 67914 28810 67942 29086
rect 68006 28810 68034 34510
rect 68282 34182 68310 34526
rect 68270 34176 68322 34182
rect 68270 34118 68322 34124
rect 68086 32816 68138 32822
rect 68086 32758 68138 32764
rect 68098 31326 68126 32758
rect 68374 32385 68402 34934
rect 68914 34584 68966 34590
rect 68914 34526 68966 34532
rect 68638 34108 68690 34114
rect 68926 34096 68954 34526
rect 68690 34068 68954 34096
rect 68638 34050 68690 34056
rect 68650 33978 68678 34050
rect 68638 33972 68690 33978
rect 68638 33914 68690 33920
rect 68730 33972 68782 33978
rect 68730 33914 68782 33920
rect 68742 33570 68770 33914
rect 68730 33564 68782 33570
rect 68730 33506 68782 33512
rect 69018 33502 69046 35598
rect 69282 35128 69334 35134
rect 69282 35070 69334 35076
rect 69294 34726 69322 35070
rect 69282 34720 69334 34726
rect 69282 34662 69334 34668
rect 68638 33496 68690 33502
rect 68638 33438 68690 33444
rect 69006 33496 69058 33502
rect 69006 33438 69058 33444
rect 68650 33366 68678 33438
rect 69098 33428 69150 33434
rect 69098 33370 69150 33376
rect 68638 33360 68690 33366
rect 68638 33302 68690 33308
rect 69110 33026 69138 33370
rect 68546 33020 68598 33026
rect 68546 32962 68598 32968
rect 69098 33020 69150 33026
rect 69098 32962 69150 32968
rect 68558 32890 68586 32962
rect 69386 32890 69414 36090
rect 69558 35672 69610 35678
rect 69558 35614 69610 35620
rect 69570 35338 69598 35614
rect 69662 35338 69690 36158
rect 69558 35332 69610 35338
rect 69558 35274 69610 35280
rect 69650 35332 69702 35338
rect 69650 35274 69702 35280
rect 69754 35066 69782 36278
rect 69926 35128 69978 35134
rect 69926 35070 69978 35076
rect 69742 35060 69794 35066
rect 69742 35002 69794 35008
rect 69466 34788 69518 34794
rect 69466 34730 69518 34736
rect 69478 34454 69506 34730
rect 69650 34584 69702 34590
rect 69650 34526 69702 34532
rect 69662 34454 69690 34526
rect 69466 34448 69518 34454
rect 69466 34390 69518 34396
rect 69650 34448 69702 34454
rect 69650 34390 69702 34396
rect 69662 34182 69690 34390
rect 69650 34176 69702 34182
rect 69650 34118 69702 34124
rect 69938 33366 69966 35070
rect 69926 33360 69978 33366
rect 69926 33302 69978 33308
rect 69740 33056 69796 33065
rect 69740 32991 69796 33000
rect 69754 32906 69782 32991
rect 68546 32884 68598 32890
rect 68546 32826 68598 32832
rect 69282 32884 69334 32890
rect 69282 32826 69334 32832
rect 69374 32884 69426 32890
rect 69754 32878 69874 32906
rect 69374 32826 69426 32832
rect 68558 32550 68586 32826
rect 68730 32816 68782 32822
rect 68730 32758 68782 32764
rect 68546 32544 68598 32550
rect 68546 32486 68598 32492
rect 68360 32376 68416 32385
rect 68360 32311 68416 32320
rect 68362 31932 68414 31938
rect 68362 31874 68414 31880
rect 68374 31462 68402 31874
rect 68638 31796 68690 31802
rect 68638 31738 68690 31744
rect 68650 31530 68678 31738
rect 68638 31524 68690 31530
rect 68638 31466 68690 31472
rect 68362 31456 68414 31462
rect 68362 31398 68414 31404
rect 68086 31320 68138 31326
rect 68086 31262 68138 31268
rect 68178 31184 68230 31190
rect 68178 31126 68230 31132
rect 68190 30986 68218 31126
rect 68178 30980 68230 30986
rect 68178 30922 68230 30928
rect 68638 30164 68690 30170
rect 68638 30106 68690 30112
rect 68650 29830 68678 30106
rect 68638 29824 68690 29830
rect 68638 29766 68690 29772
rect 68650 29694 68678 29766
rect 68638 29688 68690 29694
rect 68638 29630 68690 29636
rect 68086 29620 68138 29626
rect 68086 29562 68138 29568
rect 68178 29620 68230 29626
rect 68178 29562 68230 29568
rect 68098 29354 68126 29562
rect 68086 29348 68138 29354
rect 68086 29290 68138 29296
rect 68190 29150 68218 29562
rect 68178 29144 68230 29150
rect 68178 29086 68230 29092
rect 68638 29144 68690 29150
rect 68638 29086 68690 29092
rect 67902 28804 67954 28810
rect 67902 28746 67954 28752
rect 67994 28804 68046 28810
rect 67994 28746 68046 28752
rect 67166 28668 67218 28674
rect 67166 28610 67218 28616
rect 67590 28364 67886 28384
rect 67646 28362 67670 28364
rect 67726 28362 67750 28364
rect 67806 28362 67830 28364
rect 67668 28310 67670 28362
rect 67732 28310 67744 28362
rect 67806 28310 67808 28362
rect 67646 28308 67670 28310
rect 67726 28308 67750 28310
rect 67806 28308 67830 28310
rect 67590 28288 67886 28308
rect 67914 27722 67942 28746
rect 68006 28130 68034 28746
rect 68176 28160 68232 28169
rect 67994 28124 68046 28130
rect 68176 28095 68232 28104
rect 67994 28066 68046 28072
rect 67902 27716 67954 27722
rect 67902 27658 67954 27664
rect 65418 27512 65470 27518
rect 65418 27454 65470 27460
rect 67074 27512 67126 27518
rect 67074 27454 67126 27460
rect 67994 27512 68046 27518
rect 67994 27454 68046 27460
rect 68190 27466 68218 28095
rect 68650 27994 68678 29086
rect 68638 27988 68690 27994
rect 68638 27930 68690 27936
rect 68270 27920 68322 27926
rect 68270 27862 68322 27868
rect 68282 27586 68310 27862
rect 68270 27580 68322 27586
rect 68270 27522 68322 27528
rect 61186 27036 61238 27042
rect 61186 26978 61238 26984
rect 62658 27036 62710 27042
rect 62658 26978 62710 26984
rect 63302 27036 63354 27042
rect 63302 26978 63354 26984
rect 64130 27036 64182 27042
rect 64130 26978 64182 26984
rect 65430 26974 65458 27454
rect 66154 27444 66206 27450
rect 66154 27386 66206 27392
rect 66166 27110 66194 27386
rect 67590 27276 67886 27296
rect 67646 27274 67670 27276
rect 67726 27274 67750 27276
rect 67806 27274 67830 27276
rect 67668 27222 67670 27274
rect 67732 27222 67744 27274
rect 67806 27222 67808 27274
rect 67646 27220 67670 27222
rect 67726 27220 67750 27222
rect 67806 27220 67830 27222
rect 67590 27200 67886 27220
rect 66154 27104 66206 27110
rect 66154 27046 66206 27052
rect 68006 27042 68034 27454
rect 68190 27438 68494 27466
rect 67994 27036 68046 27042
rect 67994 26978 68046 26984
rect 56862 26968 56914 26974
rect 56862 26910 56914 26916
rect 65418 26968 65470 26974
rect 65418 26910 65470 26916
rect 49318 26900 49370 26906
rect 49318 26842 49370 26848
rect 53458 26900 53510 26906
rect 53458 26842 53510 26848
rect 50330 26832 50382 26838
rect 50422 26832 50474 26838
rect 50382 26780 50422 26786
rect 50330 26774 50474 26780
rect 50342 26758 50462 26774
rect 48942 26732 49238 26752
rect 48998 26730 49022 26732
rect 49078 26730 49102 26732
rect 49158 26730 49182 26732
rect 49020 26678 49022 26730
rect 49084 26678 49096 26730
rect 49158 26678 49160 26730
rect 48998 26676 49022 26678
rect 49078 26676 49102 26678
rect 49158 26676 49182 26678
rect 48942 26656 49238 26676
rect 54270 26732 54566 26752
rect 54326 26730 54350 26732
rect 54406 26730 54430 26732
rect 54486 26730 54510 26732
rect 54348 26678 54350 26730
rect 54412 26678 54424 26730
rect 54486 26678 54488 26730
rect 54326 26676 54350 26678
rect 54406 26676 54430 26678
rect 54486 26676 54510 26678
rect 54270 26656 54566 26676
rect 59598 26732 59894 26752
rect 59654 26730 59678 26732
rect 59734 26730 59758 26732
rect 59814 26730 59838 26732
rect 59676 26678 59678 26730
rect 59740 26678 59752 26730
rect 59814 26678 59816 26730
rect 59654 26676 59678 26678
rect 59734 26676 59758 26678
rect 59814 26676 59838 26678
rect 59598 26656 59894 26676
rect 64926 26732 65222 26752
rect 64982 26730 65006 26732
rect 65062 26730 65086 26732
rect 65142 26730 65166 26732
rect 65004 26678 65006 26730
rect 65068 26678 65080 26730
rect 65142 26678 65144 26730
rect 64982 26676 65006 26678
rect 65062 26676 65086 26678
rect 65142 26676 65166 26678
rect 64926 26656 65222 26676
rect 67074 26288 67126 26294
rect 67074 26230 67126 26236
rect 46096 23604 46152 23613
rect 43522 23568 43574 23574
rect 46096 23539 46152 23548
rect 43522 23510 43574 23516
rect 43534 23001 43562 23510
rect 43520 22992 43576 23001
rect 43520 22927 43576 22936
rect 67086 21890 67114 26230
rect 67086 21862 67206 21890
rect 67074 21800 67126 21806
rect 67074 21742 67126 21748
rect 67086 20689 67114 21742
rect 67178 21369 67206 21862
rect 67164 21360 67220 21369
rect 67164 21295 67220 21304
rect 67072 20680 67128 20689
rect 67072 20615 67128 20624
rect 43258 18734 43378 18762
rect 40950 18572 41246 18592
rect 41006 18570 41030 18572
rect 41086 18570 41110 18572
rect 41166 18570 41190 18572
rect 41028 18518 41030 18570
rect 41092 18518 41104 18570
rect 41166 18518 41168 18570
rect 41006 18516 41030 18518
rect 41086 18516 41110 18518
rect 41166 18516 41190 18518
rect 40950 18496 41246 18516
rect 40762 18264 40814 18270
rect 40762 18206 40814 18212
rect 39198 17788 39250 17794
rect 39198 17730 39250 17736
rect 40670 17788 40722 17794
rect 40670 17730 40722 17736
rect 39210 17250 39238 17730
rect 40774 17726 40802 18206
rect 42050 18128 42102 18134
rect 42050 18070 42102 18076
rect 42062 17969 42090 18070
rect 42048 17960 42104 17969
rect 42048 17895 42050 17904
rect 42102 17895 42104 17904
rect 42050 17866 42102 17872
rect 42062 17835 42090 17866
rect 40762 17720 40814 17726
rect 40762 17662 40814 17668
rect 40950 17484 41246 17504
rect 41006 17482 41030 17484
rect 41086 17482 41110 17484
rect 41166 17482 41190 17484
rect 41028 17430 41030 17482
rect 41092 17430 41104 17482
rect 41166 17430 41168 17482
rect 41006 17428 41030 17430
rect 41086 17428 41110 17430
rect 41166 17428 41190 17430
rect 40950 17408 41246 17428
rect 39750 17312 39802 17318
rect 39750 17254 39802 17260
rect 39198 17244 39250 17250
rect 39198 17186 39250 17192
rect 38738 17176 38790 17182
rect 38738 17118 38790 17124
rect 38828 17144 38884 17153
rect 38286 16940 38582 16960
rect 38342 16938 38366 16940
rect 38422 16938 38446 16940
rect 38502 16938 38526 16940
rect 38364 16886 38366 16938
rect 38428 16886 38440 16938
rect 38502 16886 38504 16938
rect 38342 16884 38366 16886
rect 38422 16884 38446 16886
rect 38502 16884 38526 16886
rect 38286 16864 38582 16884
rect 38750 16706 38778 17118
rect 38828 17079 38830 17088
rect 38882 17079 38884 17088
rect 38830 17050 38882 17056
rect 39762 16842 39790 17254
rect 39842 17176 39894 17182
rect 40762 17176 40814 17182
rect 39842 17118 39894 17124
rect 40760 17144 40762 17153
rect 40814 17144 40816 17153
rect 39854 17046 39882 17118
rect 40760 17079 40816 17088
rect 39842 17040 39894 17046
rect 39842 16982 39894 16988
rect 41038 17040 41090 17046
rect 41038 16982 41090 16988
rect 39750 16836 39802 16842
rect 39750 16778 39802 16784
rect 38646 16700 38698 16706
rect 38646 16642 38698 16648
rect 38738 16700 38790 16706
rect 38738 16642 38790 16648
rect 38002 16292 38054 16298
rect 38002 16234 38054 16240
rect 37726 15952 37778 15958
rect 37726 15894 37778 15900
rect 37082 15612 37134 15618
rect 37082 15554 37134 15560
rect 37358 15612 37410 15618
rect 37358 15554 37410 15560
rect 35622 15308 35918 15328
rect 35678 15306 35702 15308
rect 35758 15306 35782 15308
rect 35838 15306 35862 15308
rect 35700 15254 35702 15306
rect 35764 15254 35776 15306
rect 35838 15254 35840 15306
rect 35678 15252 35702 15254
rect 35758 15252 35782 15254
rect 35838 15252 35862 15254
rect 35622 15232 35918 15252
rect 37094 15210 37122 15554
rect 37082 15204 37134 15210
rect 37082 15146 37134 15152
rect 37738 15074 37766 15894
rect 38286 15852 38582 15872
rect 38342 15850 38366 15852
rect 38422 15850 38446 15852
rect 38502 15850 38526 15852
rect 38364 15798 38366 15850
rect 38428 15798 38440 15850
rect 38502 15798 38504 15850
rect 38342 15796 38366 15798
rect 38422 15796 38446 15798
rect 38502 15796 38526 15798
rect 38286 15776 38582 15796
rect 38658 15414 38686 16642
rect 39762 16638 39790 16778
rect 41050 16706 41078 16982
rect 41038 16700 41090 16706
rect 41038 16642 41090 16648
rect 39750 16632 39802 16638
rect 41682 16632 41734 16638
rect 39750 16574 39802 16580
rect 41680 16600 41682 16609
rect 41734 16600 41736 16609
rect 41680 16535 41736 16544
rect 40950 16396 41246 16416
rect 41006 16394 41030 16396
rect 41086 16394 41110 16396
rect 41166 16394 41190 16396
rect 41028 16342 41030 16394
rect 41092 16342 41104 16394
rect 41166 16342 41168 16394
rect 41006 16340 41030 16342
rect 41086 16340 41110 16342
rect 41166 16340 41190 16342
rect 40950 16320 41246 16340
rect 38922 16088 38974 16094
rect 38922 16030 38974 16036
rect 38646 15408 38698 15414
rect 38646 15350 38698 15356
rect 37726 15068 37778 15074
rect 37726 15010 37778 15016
rect 38934 14938 38962 16030
rect 40950 15308 41246 15328
rect 41006 15306 41030 15308
rect 41086 15306 41110 15308
rect 41166 15306 41190 15308
rect 41028 15254 41030 15306
rect 41092 15254 41104 15306
rect 41166 15254 41168 15306
rect 41006 15252 41030 15254
rect 41086 15252 41110 15254
rect 41166 15252 41190 15254
rect 40950 15232 41246 15252
rect 38922 14932 38974 14938
rect 38922 14874 38974 14880
rect 34414 14864 34466 14870
rect 34412 14832 34414 14841
rect 34466 14832 34468 14841
rect 34412 14767 34468 14776
rect 38286 14764 38582 14784
rect 38342 14762 38366 14764
rect 38422 14762 38446 14764
rect 38502 14762 38526 14764
rect 38364 14710 38366 14762
rect 38428 14710 38440 14762
rect 38502 14710 38504 14762
rect 38342 14708 38366 14710
rect 38422 14708 38446 14710
rect 38502 14708 38526 14710
rect 38286 14688 38582 14708
rect 35622 14220 35918 14240
rect 35678 14218 35702 14220
rect 35758 14218 35782 14220
rect 35838 14218 35862 14220
rect 35700 14166 35702 14218
rect 35764 14166 35776 14218
rect 35838 14166 35840 14218
rect 35678 14164 35702 14166
rect 35758 14164 35782 14166
rect 35838 14164 35862 14166
rect 35622 14144 35918 14164
rect 38286 13676 38582 13696
rect 38342 13674 38366 13676
rect 38422 13674 38446 13676
rect 38502 13674 38526 13676
rect 38364 13622 38366 13674
rect 38428 13622 38440 13674
rect 38502 13622 38504 13674
rect 38342 13620 38366 13622
rect 38422 13620 38446 13622
rect 38502 13620 38526 13622
rect 38286 13600 38582 13620
rect 35622 13132 35918 13152
rect 35678 13130 35702 13132
rect 35758 13130 35782 13132
rect 35838 13130 35862 13132
rect 35700 13078 35702 13130
rect 35764 13078 35776 13130
rect 35838 13078 35840 13130
rect 35678 13076 35702 13078
rect 35758 13076 35782 13078
rect 35838 13076 35862 13078
rect 35622 13056 35918 13076
rect 38286 12588 38582 12608
rect 38342 12586 38366 12588
rect 38422 12586 38446 12588
rect 38502 12586 38526 12588
rect 38364 12534 38366 12586
rect 38428 12534 38440 12586
rect 38502 12534 38504 12586
rect 38342 12532 38366 12534
rect 38422 12532 38446 12534
rect 38502 12532 38526 12534
rect 38286 12512 38582 12532
rect 35622 12044 35918 12064
rect 35678 12042 35702 12044
rect 35758 12042 35782 12044
rect 35838 12042 35862 12044
rect 35700 11990 35702 12042
rect 35764 11990 35776 12042
rect 35838 11990 35840 12042
rect 35678 11988 35702 11990
rect 35758 11988 35782 11990
rect 35838 11988 35862 11990
rect 35622 11968 35918 11988
rect 38934 11674 38962 14874
rect 40950 14220 41246 14240
rect 41006 14218 41030 14220
rect 41086 14218 41110 14220
rect 41166 14218 41190 14220
rect 41028 14166 41030 14218
rect 41092 14166 41104 14218
rect 41166 14166 41168 14218
rect 41006 14164 41030 14166
rect 41086 14164 41110 14166
rect 41166 14164 41190 14166
rect 40950 14144 41246 14164
rect 40950 13132 41246 13152
rect 41006 13130 41030 13132
rect 41086 13130 41110 13132
rect 41166 13130 41190 13132
rect 41028 13078 41030 13130
rect 41092 13078 41104 13130
rect 41166 13078 41168 13130
rect 41006 13076 41030 13078
rect 41086 13076 41110 13078
rect 41166 13076 41190 13078
rect 40950 13056 41246 13076
rect 40950 12044 41246 12064
rect 41006 12042 41030 12044
rect 41086 12042 41110 12044
rect 41166 12042 41190 12044
rect 41028 11990 41030 12042
rect 41092 11990 41104 12042
rect 41166 11990 41168 12042
rect 41006 11988 41030 11990
rect 41086 11988 41110 11990
rect 41166 11988 41190 11990
rect 40950 11968 41246 11988
rect 38922 11668 38974 11674
rect 38922 11610 38974 11616
rect 38286 11500 38582 11520
rect 38342 11498 38366 11500
rect 38422 11498 38446 11500
rect 38502 11498 38526 11500
rect 38364 11446 38366 11498
rect 38428 11446 38440 11498
rect 38502 11446 38504 11498
rect 38342 11444 38366 11446
rect 38422 11444 38446 11446
rect 38502 11444 38526 11446
rect 38286 11424 38582 11444
rect 35622 10956 35918 10976
rect 35678 10954 35702 10956
rect 35758 10954 35782 10956
rect 35838 10954 35862 10956
rect 35700 10902 35702 10954
rect 35764 10902 35776 10954
rect 35838 10902 35840 10954
rect 35678 10900 35702 10902
rect 35758 10900 35782 10902
rect 35838 10900 35862 10902
rect 35622 10880 35918 10900
rect 40950 10956 41246 10976
rect 41006 10954 41030 10956
rect 41086 10954 41110 10956
rect 41166 10954 41190 10956
rect 41028 10902 41030 10954
rect 41092 10902 41104 10954
rect 41166 10902 41168 10954
rect 41006 10900 41030 10902
rect 41086 10900 41110 10902
rect 41166 10900 41190 10902
rect 40950 10880 41246 10900
rect 34414 10512 34466 10518
rect 34412 10480 34414 10489
rect 34466 10480 34468 10489
rect 34412 10415 34468 10424
rect 38286 10412 38582 10432
rect 38342 10410 38366 10412
rect 38422 10410 38446 10412
rect 38502 10410 38526 10412
rect 38364 10358 38366 10410
rect 38428 10358 38440 10410
rect 38502 10358 38504 10410
rect 38342 10356 38366 10358
rect 38422 10356 38446 10358
rect 38502 10356 38526 10358
rect 38286 10336 38582 10356
rect 11190 10188 11270 10194
rect 11138 10182 11270 10188
rect 6078 10172 6130 10178
rect 11150 10166 11270 10182
rect 6078 10114 6130 10120
rect 7090 9968 7142 9974
rect 7090 9910 7142 9916
rect 3654 9868 3950 9888
rect 3710 9866 3734 9868
rect 3790 9866 3814 9868
rect 3870 9866 3894 9868
rect 3732 9814 3734 9866
rect 3796 9814 3808 9866
rect 3870 9814 3872 9866
rect 3710 9812 3734 9814
rect 3790 9812 3814 9814
rect 3870 9812 3894 9814
rect 3654 9792 3950 9812
rect 6318 9324 6614 9344
rect 6374 9322 6398 9324
rect 6454 9322 6478 9324
rect 6534 9322 6558 9324
rect 6396 9270 6398 9322
rect 6460 9270 6472 9322
rect 6534 9270 6536 9322
rect 6374 9268 6398 9270
rect 6454 9268 6478 9270
rect 6534 9268 6558 9270
rect 6318 9248 6614 9268
rect 3654 8780 3950 8800
rect 3710 8778 3734 8780
rect 3790 8778 3814 8780
rect 3870 8778 3894 8780
rect 3732 8726 3734 8778
rect 3796 8726 3808 8778
rect 3870 8726 3872 8778
rect 3710 8724 3734 8726
rect 3790 8724 3814 8726
rect 3870 8724 3894 8726
rect 3654 8704 3950 8724
rect 6318 8236 6614 8256
rect 6374 8234 6398 8236
rect 6454 8234 6478 8236
rect 6534 8234 6558 8236
rect 6396 8182 6398 8234
rect 6460 8182 6472 8234
rect 6534 8182 6536 8234
rect 6374 8180 6398 8182
rect 6454 8180 6478 8182
rect 6534 8180 6558 8182
rect 6318 8160 6614 8180
rect 3654 7692 3950 7712
rect 3710 7690 3734 7692
rect 3790 7690 3814 7692
rect 3870 7690 3894 7692
rect 3732 7638 3734 7690
rect 3796 7638 3808 7690
rect 3870 7638 3872 7690
rect 3710 7636 3734 7638
rect 3790 7636 3814 7638
rect 3870 7636 3894 7638
rect 3654 7616 3950 7636
rect 6318 7148 6614 7168
rect 6374 7146 6398 7148
rect 6454 7146 6478 7148
rect 6534 7146 6558 7148
rect 6396 7094 6398 7146
rect 6460 7094 6472 7146
rect 6534 7094 6536 7146
rect 6374 7092 6398 7094
rect 6454 7092 6478 7094
rect 6534 7092 6558 7094
rect 6318 7072 6614 7092
rect 3654 6604 3950 6624
rect 3710 6602 3734 6604
rect 3790 6602 3814 6604
rect 3870 6602 3894 6604
rect 3732 6550 3734 6602
rect 3796 6550 3808 6602
rect 3870 6550 3872 6602
rect 3710 6548 3734 6550
rect 3790 6548 3814 6550
rect 3870 6548 3894 6550
rect 3654 6528 3950 6548
rect 6318 6060 6614 6080
rect 6374 6058 6398 6060
rect 6454 6058 6478 6060
rect 6534 6058 6558 6060
rect 6396 6006 6398 6058
rect 6460 6006 6472 6058
rect 6534 6006 6536 6058
rect 6374 6004 6398 6006
rect 6454 6004 6478 6006
rect 6534 6004 6558 6006
rect 6318 5984 6614 6004
rect 3654 5516 3950 5536
rect 3710 5514 3734 5516
rect 3790 5514 3814 5516
rect 3870 5514 3894 5516
rect 3732 5462 3734 5514
rect 3796 5462 3808 5514
rect 3870 5462 3872 5514
rect 3710 5460 3734 5462
rect 3790 5460 3814 5462
rect 3870 5460 3894 5462
rect 3654 5440 3950 5460
rect 6318 4972 6614 4992
rect 6374 4970 6398 4972
rect 6454 4970 6478 4972
rect 6534 4970 6558 4972
rect 6396 4918 6398 4970
rect 6460 4918 6472 4970
rect 6534 4918 6536 4970
rect 6374 4916 6398 4918
rect 6454 4916 6478 4918
rect 6534 4916 6558 4918
rect 6318 4896 6614 4916
rect 3654 4428 3950 4448
rect 3710 4426 3734 4428
rect 3790 4426 3814 4428
rect 3870 4426 3894 4428
rect 3732 4374 3734 4426
rect 3796 4374 3808 4426
rect 3870 4374 3872 4426
rect 3710 4372 3734 4374
rect 3790 4372 3814 4374
rect 3870 4372 3894 4374
rect 3654 4352 3950 4372
rect 6318 3884 6614 3904
rect 6374 3882 6398 3884
rect 6454 3882 6478 3884
rect 6534 3882 6558 3884
rect 6396 3830 6398 3882
rect 6460 3830 6472 3882
rect 6534 3830 6536 3882
rect 6374 3828 6398 3830
rect 6454 3828 6478 3830
rect 6534 3828 6558 3830
rect 6318 3808 6614 3828
rect 3654 3340 3950 3360
rect 3710 3338 3734 3340
rect 3790 3338 3814 3340
rect 3870 3338 3894 3340
rect 3732 3286 3734 3338
rect 3796 3286 3808 3338
rect 3870 3286 3872 3338
rect 3710 3284 3734 3286
rect 3790 3284 3814 3286
rect 3870 3284 3894 3286
rect 3654 3264 3950 3284
rect 6318 2796 6614 2816
rect 6374 2794 6398 2796
rect 6454 2794 6478 2796
rect 6534 2794 6558 2796
rect 6396 2742 6398 2794
rect 6460 2742 6472 2794
rect 6534 2742 6536 2794
rect 6374 2740 6398 2742
rect 6454 2740 6478 2742
rect 6534 2740 6558 2742
rect 6318 2720 6614 2740
rect 3654 2252 3950 2272
rect 3710 2250 3734 2252
rect 3790 2250 3814 2252
rect 3870 2250 3894 2252
rect 3732 2198 3734 2250
rect 3796 2198 3808 2250
rect 3870 2198 3872 2250
rect 3710 2196 3734 2198
rect 3790 2196 3814 2198
rect 3870 2196 3894 2198
rect 3654 2176 3950 2196
rect 7102 2154 7130 9910
rect 35622 9868 35918 9888
rect 35678 9866 35702 9868
rect 35758 9866 35782 9868
rect 35838 9866 35862 9868
rect 35700 9814 35702 9866
rect 35764 9814 35776 9866
rect 35838 9814 35840 9866
rect 35678 9812 35702 9814
rect 35758 9812 35782 9814
rect 35838 9812 35862 9814
rect 35622 9792 35918 9812
rect 40950 9868 41246 9888
rect 41006 9866 41030 9868
rect 41086 9866 41110 9868
rect 41166 9866 41190 9868
rect 41028 9814 41030 9866
rect 41092 9814 41104 9866
rect 41166 9814 41168 9866
rect 41006 9812 41030 9814
rect 41086 9812 41110 9814
rect 41166 9812 41190 9814
rect 40950 9792 41246 9812
rect 38286 9324 38582 9344
rect 38342 9322 38366 9324
rect 38422 9322 38446 9324
rect 38502 9322 38526 9324
rect 38364 9270 38366 9322
rect 38428 9270 38440 9322
rect 38502 9270 38504 9322
rect 38342 9268 38366 9270
rect 38422 9268 38446 9270
rect 38502 9268 38526 9270
rect 38286 9248 38582 9268
rect 35622 8780 35918 8800
rect 35678 8778 35702 8780
rect 35758 8778 35782 8780
rect 35838 8778 35862 8780
rect 35700 8726 35702 8778
rect 35764 8726 35776 8778
rect 35838 8726 35840 8778
rect 35678 8724 35702 8726
rect 35758 8724 35782 8726
rect 35838 8724 35862 8726
rect 35622 8704 35918 8724
rect 40950 8780 41246 8800
rect 41006 8778 41030 8780
rect 41086 8778 41110 8780
rect 41166 8778 41190 8780
rect 41028 8726 41030 8778
rect 41092 8726 41104 8778
rect 41166 8726 41168 8778
rect 41006 8724 41030 8726
rect 41086 8724 41110 8726
rect 41166 8724 41190 8726
rect 40950 8704 41246 8724
rect 38286 8236 38582 8256
rect 38342 8234 38366 8236
rect 38422 8234 38446 8236
rect 38502 8234 38526 8236
rect 38364 8182 38366 8234
rect 38428 8182 38440 8234
rect 38502 8182 38504 8234
rect 38342 8180 38366 8182
rect 38422 8180 38446 8182
rect 38502 8180 38526 8182
rect 38286 8160 38582 8180
rect 35622 7692 35918 7712
rect 35678 7690 35702 7692
rect 35758 7690 35782 7692
rect 35838 7690 35862 7692
rect 35700 7638 35702 7690
rect 35764 7638 35776 7690
rect 35838 7638 35840 7690
rect 35678 7636 35702 7638
rect 35758 7636 35782 7638
rect 35838 7636 35862 7638
rect 35622 7616 35918 7636
rect 40950 7692 41246 7712
rect 41006 7690 41030 7692
rect 41086 7690 41110 7692
rect 41166 7690 41190 7692
rect 41028 7638 41030 7690
rect 41092 7638 41104 7690
rect 41166 7638 41168 7690
rect 41006 7636 41030 7638
rect 41086 7636 41110 7638
rect 41166 7636 41190 7638
rect 40950 7616 41246 7636
rect 38286 7148 38582 7168
rect 38342 7146 38366 7148
rect 38422 7146 38446 7148
rect 38502 7146 38526 7148
rect 38364 7094 38366 7146
rect 38428 7094 38440 7146
rect 38502 7094 38504 7146
rect 38342 7092 38366 7094
rect 38422 7092 38446 7094
rect 38502 7092 38526 7094
rect 38286 7072 38582 7092
rect 35622 6604 35918 6624
rect 35678 6602 35702 6604
rect 35758 6602 35782 6604
rect 35838 6602 35862 6604
rect 35700 6550 35702 6602
rect 35764 6550 35776 6602
rect 35838 6550 35840 6602
rect 35678 6548 35702 6550
rect 35758 6548 35782 6550
rect 35838 6548 35862 6550
rect 35622 6528 35918 6548
rect 40950 6604 41246 6624
rect 41006 6602 41030 6604
rect 41086 6602 41110 6604
rect 41166 6602 41190 6604
rect 41028 6550 41030 6602
rect 41092 6550 41104 6602
rect 41166 6550 41168 6602
rect 41006 6548 41030 6550
rect 41086 6548 41110 6550
rect 41166 6548 41190 6550
rect 40950 6528 41246 6548
rect 38286 6060 38582 6080
rect 38342 6058 38366 6060
rect 38422 6058 38446 6060
rect 38502 6058 38526 6060
rect 38364 6006 38366 6058
rect 38428 6006 38440 6058
rect 38502 6006 38504 6058
rect 38342 6004 38366 6006
rect 38422 6004 38446 6006
rect 38502 6004 38526 6006
rect 38286 5984 38582 6004
rect 35622 5516 35918 5536
rect 35678 5514 35702 5516
rect 35758 5514 35782 5516
rect 35838 5514 35862 5516
rect 35700 5462 35702 5514
rect 35764 5462 35776 5514
rect 35838 5462 35840 5514
rect 35678 5460 35702 5462
rect 35758 5460 35782 5462
rect 35838 5460 35862 5462
rect 35622 5440 35918 5460
rect 40950 5516 41246 5536
rect 41006 5514 41030 5516
rect 41086 5514 41110 5516
rect 41166 5514 41190 5516
rect 41028 5462 41030 5514
rect 41092 5462 41104 5514
rect 41166 5462 41168 5514
rect 41006 5460 41030 5462
rect 41086 5460 41110 5462
rect 41166 5460 41190 5462
rect 40950 5440 41246 5460
rect 38286 4972 38582 4992
rect 38342 4970 38366 4972
rect 38422 4970 38446 4972
rect 38502 4970 38526 4972
rect 38364 4918 38366 4970
rect 38428 4918 38440 4970
rect 38502 4918 38504 4970
rect 38342 4916 38366 4918
rect 38422 4916 38446 4918
rect 38502 4916 38526 4918
rect 38286 4896 38582 4916
rect 35622 4428 35918 4448
rect 35678 4426 35702 4428
rect 35758 4426 35782 4428
rect 35838 4426 35862 4428
rect 35700 4374 35702 4426
rect 35764 4374 35776 4426
rect 35838 4374 35840 4426
rect 35678 4372 35702 4374
rect 35758 4372 35782 4374
rect 35838 4372 35862 4374
rect 35622 4352 35918 4372
rect 40950 4428 41246 4448
rect 41006 4426 41030 4428
rect 41086 4426 41110 4428
rect 41166 4426 41190 4428
rect 41028 4374 41030 4426
rect 41092 4374 41104 4426
rect 41166 4374 41168 4426
rect 41006 4372 41030 4374
rect 41086 4372 41110 4374
rect 41166 4372 41190 4374
rect 40950 4352 41246 4372
rect 38286 3884 38582 3904
rect 38342 3882 38366 3884
rect 38422 3882 38446 3884
rect 38502 3882 38526 3884
rect 38364 3830 38366 3882
rect 38428 3830 38440 3882
rect 38502 3830 38504 3882
rect 38342 3828 38366 3830
rect 38422 3828 38446 3830
rect 38502 3828 38526 3830
rect 38286 3808 38582 3828
rect 35622 3340 35918 3360
rect 35678 3338 35702 3340
rect 35758 3338 35782 3340
rect 35838 3338 35862 3340
rect 35700 3286 35702 3338
rect 35764 3286 35776 3338
rect 35838 3286 35840 3338
rect 35678 3284 35702 3286
rect 35758 3284 35782 3286
rect 35838 3284 35862 3286
rect 35622 3264 35918 3284
rect 40950 3340 41246 3360
rect 41006 3338 41030 3340
rect 41086 3338 41110 3340
rect 41166 3338 41190 3340
rect 41028 3286 41030 3338
rect 41092 3286 41104 3338
rect 41166 3286 41168 3338
rect 41006 3284 41030 3286
rect 41086 3284 41110 3286
rect 41166 3284 41190 3286
rect 40950 3264 41246 3284
rect 38286 2796 38582 2816
rect 38342 2794 38366 2796
rect 38422 2794 38446 2796
rect 38502 2794 38526 2796
rect 38364 2742 38366 2794
rect 38428 2742 38440 2794
rect 38502 2742 38504 2794
rect 38342 2740 38366 2742
rect 38422 2740 38446 2742
rect 38502 2740 38526 2742
rect 38286 2720 38582 2740
rect 43258 2698 43286 18734
rect 43338 18672 43390 18678
rect 43338 18614 43390 18620
rect 43350 17017 43378 18614
rect 43522 18332 43574 18338
rect 43522 18274 43574 18280
rect 43534 18105 43562 18274
rect 67086 18105 67114 20615
rect 68190 20281 68218 27438
rect 68270 27376 68322 27382
rect 68270 27318 68322 27324
rect 68282 27042 68310 27318
rect 68466 27042 68494 27438
rect 68742 27382 68770 32758
rect 68822 32408 68874 32414
rect 68822 32350 68874 32356
rect 68834 31870 68862 32350
rect 69190 32340 69242 32346
rect 69190 32282 69242 32288
rect 69202 32090 69230 32282
rect 69294 32260 69322 32826
rect 69386 32414 69414 32826
rect 69742 32816 69794 32822
rect 69742 32758 69794 32764
rect 69754 32414 69782 32758
rect 69846 32414 69874 32878
rect 69374 32408 69426 32414
rect 69374 32350 69426 32356
rect 69742 32408 69794 32414
rect 69742 32350 69794 32356
rect 69834 32408 69886 32414
rect 69834 32350 69886 32356
rect 69846 32260 69874 32350
rect 69294 32232 69506 32260
rect 69202 32062 69414 32090
rect 69004 31968 69060 31977
rect 69386 31938 69414 32062
rect 69004 31903 69006 31912
rect 69058 31903 69060 31912
rect 69190 31932 69242 31938
rect 69006 31874 69058 31880
rect 69190 31874 69242 31880
rect 69374 31932 69426 31938
rect 69374 31874 69426 31880
rect 68822 31864 68874 31870
rect 68874 31824 68954 31852
rect 68822 31806 68874 31812
rect 68926 31734 68954 31824
rect 68822 31728 68874 31734
rect 68822 31670 68874 31676
rect 68914 31728 68966 31734
rect 68914 31670 68966 31676
rect 68834 31462 68862 31670
rect 69202 31530 69230 31874
rect 69190 31524 69242 31530
rect 69190 31466 69242 31472
rect 68822 31456 68874 31462
rect 68822 31398 68874 31404
rect 69190 30640 69242 30646
rect 69190 30582 69242 30588
rect 69006 29756 69058 29762
rect 69006 29698 69058 29704
rect 69098 29756 69150 29762
rect 69098 29698 69150 29704
rect 69018 29150 69046 29698
rect 69110 29218 69138 29698
rect 69098 29212 69150 29218
rect 69098 29154 69150 29160
rect 69006 29144 69058 29150
rect 69006 29086 69058 29092
rect 69018 28810 69046 29086
rect 69202 29014 69230 30582
rect 69478 29286 69506 32232
rect 69570 32232 69874 32260
rect 69570 29558 69598 32232
rect 69650 32000 69702 32006
rect 69648 31968 69650 31977
rect 69702 31968 69704 31977
rect 70030 31938 70058 37110
rect 72238 36834 72266 37654
rect 72502 37440 72554 37446
rect 72502 37382 72554 37388
rect 72514 36970 72542 37382
rect 72606 37378 72634 38402
rect 72790 37786 72818 39898
rect 72882 39554 72910 39966
rect 72870 39548 72922 39554
rect 72870 39490 72922 39496
rect 72918 39244 73214 39264
rect 72974 39242 72998 39244
rect 73054 39242 73078 39244
rect 73134 39242 73158 39244
rect 72996 39190 72998 39242
rect 73060 39190 73072 39242
rect 73134 39190 73136 39242
rect 72974 39188 72998 39190
rect 73054 39188 73078 39190
rect 73134 39188 73158 39190
rect 72918 39168 73214 39188
rect 72918 38156 73214 38176
rect 72974 38154 72998 38156
rect 73054 38154 73078 38156
rect 73134 38154 73158 38156
rect 72996 38102 72998 38154
rect 73060 38102 73072 38154
rect 73134 38102 73136 38154
rect 72974 38100 72998 38102
rect 73054 38100 73078 38102
rect 73134 38100 73158 38102
rect 72918 38080 73214 38100
rect 73054 37984 73106 37990
rect 73054 37926 73106 37932
rect 72778 37780 72830 37786
rect 72778 37722 72830 37728
rect 73066 37378 73094 37926
rect 72594 37372 72646 37378
rect 72594 37314 72646 37320
rect 73054 37372 73106 37378
rect 73054 37314 73106 37320
rect 72606 36970 72634 37314
rect 72918 37068 73214 37088
rect 72974 37066 72998 37068
rect 73054 37066 73078 37068
rect 73134 37066 73158 37068
rect 72996 37014 72998 37066
rect 73060 37014 73072 37066
rect 73134 37014 73136 37066
rect 72974 37012 72998 37014
rect 73054 37012 73078 37014
rect 73134 37012 73158 37014
rect 72918 36992 73214 37012
rect 72502 36964 72554 36970
rect 72502 36906 72554 36912
rect 72594 36964 72646 36970
rect 72594 36906 72646 36912
rect 72226 36828 72278 36834
rect 72226 36770 72278 36776
rect 70254 36524 70550 36544
rect 70310 36522 70334 36524
rect 70390 36522 70414 36524
rect 70470 36522 70494 36524
rect 70332 36470 70334 36522
rect 70396 36470 70408 36522
rect 70470 36470 70472 36522
rect 70310 36468 70334 36470
rect 70390 36468 70414 36470
rect 70470 36468 70494 36470
rect 70254 36448 70550 36468
rect 73342 36290 73370 40034
rect 73618 39894 73646 40510
rect 73710 40438 73738 40510
rect 73698 40432 73750 40438
rect 73698 40374 73750 40380
rect 73606 39888 73658 39894
rect 73606 39830 73658 39836
rect 73894 39622 73922 41054
rect 74066 40024 74118 40030
rect 74066 39966 74118 39972
rect 73882 39616 73934 39622
rect 73882 39558 73934 39564
rect 73422 39548 73474 39554
rect 73422 39490 73474 39496
rect 73434 38534 73462 39490
rect 74078 39146 74106 39966
rect 74538 39962 74566 43312
rect 75734 42154 75762 43312
rect 75734 42126 75946 42154
rect 75582 41964 75878 41984
rect 75638 41962 75662 41964
rect 75718 41962 75742 41964
rect 75798 41962 75822 41964
rect 75660 41910 75662 41962
rect 75724 41910 75736 41962
rect 75798 41910 75800 41962
rect 75638 41908 75662 41910
rect 75718 41908 75742 41910
rect 75798 41908 75822 41910
rect 75582 41888 75878 41908
rect 75582 40876 75878 40896
rect 75638 40874 75662 40876
rect 75718 40874 75742 40876
rect 75798 40874 75822 40876
rect 75660 40822 75662 40874
rect 75724 40822 75736 40874
rect 75798 40822 75800 40874
rect 75638 40820 75662 40822
rect 75718 40820 75742 40822
rect 75798 40820 75822 40822
rect 75582 40800 75878 40820
rect 74710 40432 74762 40438
rect 74710 40374 74762 40380
rect 74722 40166 74750 40374
rect 75918 40234 75946 42126
rect 76930 41202 76958 43312
rect 78218 41610 78246 43312
rect 78218 41582 78614 41610
rect 78246 41420 78542 41440
rect 78302 41418 78326 41420
rect 78382 41418 78406 41420
rect 78462 41418 78486 41420
rect 78324 41366 78326 41418
rect 78388 41366 78400 41418
rect 78462 41366 78464 41418
rect 78302 41364 78326 41366
rect 78382 41364 78406 41366
rect 78462 41364 78486 41366
rect 78246 41344 78542 41364
rect 76930 41174 77142 41202
rect 75998 40976 76050 40982
rect 75998 40918 76050 40924
rect 76010 40574 76038 40918
rect 75998 40568 76050 40574
rect 75998 40510 76050 40516
rect 76366 40568 76418 40574
rect 76366 40510 76418 40516
rect 76010 40438 76038 40510
rect 75998 40432 76050 40438
rect 75998 40374 76050 40380
rect 75906 40228 75958 40234
rect 75906 40170 75958 40176
rect 74710 40160 74762 40166
rect 74710 40102 74762 40108
rect 75446 40092 75498 40098
rect 75446 40034 75498 40040
rect 75262 40024 75314 40030
rect 75262 39966 75314 39972
rect 74526 39956 74578 39962
rect 74526 39898 74578 39904
rect 75274 39894 75302 39966
rect 75458 39894 75486 40034
rect 76274 39956 76326 39962
rect 76274 39898 76326 39904
rect 74158 39888 74210 39894
rect 74158 39830 74210 39836
rect 75262 39888 75314 39894
rect 75262 39830 75314 39836
rect 75446 39888 75498 39894
rect 75446 39830 75498 39836
rect 74066 39140 74118 39146
rect 74066 39082 74118 39088
rect 74170 39010 74198 39830
rect 75458 39593 75486 39830
rect 75582 39788 75878 39808
rect 75638 39786 75662 39788
rect 75718 39786 75742 39788
rect 75798 39786 75822 39788
rect 75660 39734 75662 39786
rect 75724 39734 75736 39786
rect 75798 39734 75800 39786
rect 75638 39732 75662 39734
rect 75718 39732 75742 39734
rect 75798 39732 75822 39734
rect 75582 39712 75878 39732
rect 75444 39584 75500 39593
rect 75444 39519 75500 39528
rect 75458 39146 75486 39519
rect 75446 39140 75498 39146
rect 75446 39082 75498 39088
rect 73974 39004 74026 39010
rect 73974 38946 74026 38952
rect 74158 39004 74210 39010
rect 74158 38946 74210 38952
rect 73698 38936 73750 38942
rect 73698 38878 73750 38884
rect 73422 38528 73474 38534
rect 73422 38470 73474 38476
rect 73710 38466 73738 38878
rect 73790 38868 73842 38874
rect 73790 38810 73842 38816
rect 73802 38534 73830 38810
rect 73790 38528 73842 38534
rect 73790 38470 73842 38476
rect 73698 38460 73750 38466
rect 73698 38402 73750 38408
rect 73802 37990 73830 38470
rect 73790 37984 73842 37990
rect 73790 37926 73842 37932
rect 73986 37854 74014 38946
rect 76286 38942 76314 39898
rect 76274 38936 76326 38942
rect 76274 38878 76326 38884
rect 75582 38700 75878 38720
rect 75638 38698 75662 38700
rect 75718 38698 75742 38700
rect 75798 38698 75822 38700
rect 75660 38646 75662 38698
rect 75724 38646 75736 38698
rect 75798 38646 75800 38698
rect 75638 38644 75662 38646
rect 75718 38644 75742 38646
rect 75798 38644 75822 38646
rect 75582 38624 75878 38644
rect 74250 38596 74302 38602
rect 74250 38538 74302 38544
rect 73974 37848 74026 37854
rect 74158 37848 74210 37854
rect 74026 37796 74158 37802
rect 73974 37790 74210 37796
rect 73882 37780 73934 37786
rect 73986 37774 74198 37790
rect 73882 37722 73934 37728
rect 73894 37378 73922 37722
rect 74066 37712 74118 37718
rect 74066 37654 74118 37660
rect 74158 37712 74210 37718
rect 74158 37654 74210 37660
rect 73698 37372 73750 37378
rect 73698 37314 73750 37320
rect 73882 37372 73934 37378
rect 73882 37314 73934 37320
rect 73606 37304 73658 37310
rect 73606 37246 73658 37252
rect 73618 36290 73646 37246
rect 73330 36284 73382 36290
rect 73330 36226 73382 36232
rect 73606 36284 73658 36290
rect 73606 36226 73658 36232
rect 70110 36148 70162 36154
rect 70110 36090 70162 36096
rect 70122 35542 70150 36090
rect 72918 35980 73214 36000
rect 72974 35978 72998 35980
rect 73054 35978 73078 35980
rect 73134 35978 73158 35980
rect 72996 35926 72998 35978
rect 73060 35926 73072 35978
rect 73134 35926 73136 35978
rect 72974 35924 72998 35926
rect 73054 35924 73078 35926
rect 73134 35924 73158 35926
rect 72918 35904 73214 35924
rect 73342 35746 73370 36226
rect 73238 35740 73290 35746
rect 73238 35682 73290 35688
rect 73330 35740 73382 35746
rect 73330 35682 73382 35688
rect 70662 35604 70714 35610
rect 70662 35546 70714 35552
rect 70110 35536 70162 35542
rect 70110 35478 70162 35484
rect 70254 35436 70550 35456
rect 70310 35434 70334 35436
rect 70390 35434 70414 35436
rect 70470 35434 70494 35436
rect 70332 35382 70334 35434
rect 70396 35382 70408 35434
rect 70470 35382 70472 35434
rect 70310 35380 70334 35382
rect 70390 35380 70414 35382
rect 70470 35380 70494 35382
rect 70254 35360 70550 35380
rect 70674 35202 70702 35546
rect 73250 35202 73278 35682
rect 70662 35196 70714 35202
rect 70662 35138 70714 35144
rect 73238 35196 73290 35202
rect 73238 35138 73290 35144
rect 72918 34892 73214 34912
rect 72974 34890 72998 34892
rect 73054 34890 73078 34892
rect 73134 34890 73158 34892
rect 72996 34838 72998 34890
rect 73060 34838 73072 34890
rect 73134 34838 73136 34890
rect 72974 34836 72998 34838
rect 73054 34836 73078 34838
rect 73134 34836 73158 34838
rect 72918 34816 73214 34836
rect 70254 34348 70550 34368
rect 70310 34346 70334 34348
rect 70390 34346 70414 34348
rect 70470 34346 70494 34348
rect 70332 34294 70334 34346
rect 70396 34294 70408 34346
rect 70470 34294 70472 34346
rect 70310 34292 70334 34294
rect 70390 34292 70414 34294
rect 70470 34292 70494 34294
rect 70254 34272 70550 34292
rect 72918 33804 73214 33824
rect 72974 33802 72998 33804
rect 73054 33802 73078 33804
rect 73134 33802 73158 33804
rect 72996 33750 72998 33802
rect 73060 33750 73072 33802
rect 73134 33750 73136 33802
rect 72974 33748 72998 33750
rect 73054 33748 73078 33750
rect 73134 33748 73158 33750
rect 72918 33728 73214 33748
rect 73618 33706 73646 36226
rect 73710 35746 73738 37314
rect 73974 37304 74026 37310
rect 73974 37246 74026 37252
rect 73986 36902 74014 37246
rect 74078 36902 74106 37654
rect 74170 37281 74198 37654
rect 74262 37378 74290 38538
rect 74986 38460 75038 38466
rect 74986 38402 75038 38408
rect 75446 38460 75498 38466
rect 75446 38402 75498 38408
rect 74710 38392 74762 38398
rect 74710 38334 74762 38340
rect 74722 37854 74750 38334
rect 74998 37854 75026 38402
rect 74710 37848 74762 37854
rect 74710 37790 74762 37796
rect 74986 37848 75038 37854
rect 74986 37790 75038 37796
rect 74434 37440 74486 37446
rect 74434 37382 74486 37388
rect 74250 37372 74302 37378
rect 74250 37314 74302 37320
rect 74156 37272 74212 37281
rect 74156 37207 74212 37216
rect 74250 37236 74302 37242
rect 73974 36896 74026 36902
rect 73974 36838 74026 36844
rect 74066 36896 74118 36902
rect 74066 36838 74118 36844
rect 73986 35762 74014 36838
rect 74170 36290 74198 37207
rect 74250 37178 74302 37184
rect 74262 36737 74290 37178
rect 74248 36728 74304 36737
rect 74248 36663 74304 36672
rect 74158 36284 74210 36290
rect 74158 36226 74210 36232
rect 73698 35740 73750 35746
rect 73698 35682 73750 35688
rect 73802 35734 74382 35762
rect 73710 34182 73738 35682
rect 73802 35678 73830 35734
rect 74354 35678 74382 35734
rect 73790 35672 73842 35678
rect 73790 35614 73842 35620
rect 74342 35672 74394 35678
rect 74342 35614 74394 35620
rect 74066 35536 74118 35542
rect 74066 35478 74118 35484
rect 74158 35536 74210 35542
rect 74158 35478 74210 35484
rect 73974 35196 74026 35202
rect 73974 35138 74026 35144
rect 73986 34658 74014 35138
rect 74078 34810 74106 35478
rect 74170 35202 74198 35478
rect 74158 35196 74210 35202
rect 74158 35138 74210 35144
rect 74078 34782 74290 34810
rect 74158 34720 74210 34726
rect 74158 34662 74210 34668
rect 73974 34652 74026 34658
rect 73974 34594 74026 34600
rect 73698 34176 73750 34182
rect 73698 34118 73750 34124
rect 73710 34046 73738 34118
rect 73882 34108 73934 34114
rect 73882 34050 73934 34056
rect 73698 34040 73750 34046
rect 73698 33982 73750 33988
rect 73894 33910 73922 34050
rect 74066 34040 74118 34046
rect 74064 34008 74066 34017
rect 74118 34008 74120 34017
rect 74064 33943 74120 33952
rect 73882 33904 73934 33910
rect 73882 33846 73934 33852
rect 73606 33700 73658 33706
rect 73606 33642 73658 33648
rect 73618 33570 73646 33642
rect 73606 33564 73658 33570
rect 73606 33506 73658 33512
rect 73894 33502 73922 33846
rect 74170 33570 74198 34662
rect 74158 33564 74210 33570
rect 74158 33506 74210 33512
rect 73882 33496 73934 33502
rect 73882 33438 73934 33444
rect 73894 33366 73922 33438
rect 72134 33360 72186 33366
rect 72134 33302 72186 33308
rect 73882 33360 73934 33366
rect 73882 33302 73934 33308
rect 70254 33260 70550 33280
rect 70310 33258 70334 33260
rect 70390 33258 70414 33260
rect 70470 33258 70494 33260
rect 70332 33206 70334 33258
rect 70396 33206 70408 33258
rect 70470 33206 70472 33258
rect 70310 33204 70334 33206
rect 70390 33204 70414 33206
rect 70470 33204 70494 33206
rect 70254 33184 70550 33204
rect 71214 32884 71266 32890
rect 71214 32826 71266 32832
rect 71226 32550 71254 32826
rect 71214 32544 71266 32550
rect 71214 32486 71266 32492
rect 71226 32414 71254 32486
rect 71214 32408 71266 32414
rect 71214 32350 71266 32356
rect 70254 32172 70550 32192
rect 70310 32170 70334 32172
rect 70390 32170 70414 32172
rect 70470 32170 70494 32172
rect 70332 32118 70334 32170
rect 70396 32118 70408 32170
rect 70470 32118 70472 32170
rect 70310 32116 70334 32118
rect 70390 32116 70414 32118
rect 70470 32116 70494 32118
rect 70254 32096 70550 32116
rect 69648 31903 69704 31912
rect 69834 31932 69886 31938
rect 69834 31874 69886 31880
rect 70018 31932 70070 31938
rect 70018 31874 70070 31880
rect 69846 31734 69874 31874
rect 69834 31728 69886 31734
rect 69834 31670 69886 31676
rect 70254 31084 70550 31104
rect 70310 31082 70334 31084
rect 70390 31082 70414 31084
rect 70470 31082 70494 31084
rect 70332 31030 70334 31082
rect 70396 31030 70408 31082
rect 70470 31030 70472 31082
rect 70310 31028 70334 31030
rect 70390 31028 70414 31030
rect 70470 31028 70494 31030
rect 70254 31008 70550 31028
rect 71226 30850 71254 32350
rect 72146 31938 72174 33302
rect 72918 32716 73214 32736
rect 72974 32714 72998 32716
rect 73054 32714 73078 32716
rect 73134 32714 73158 32716
rect 72996 32662 72998 32714
rect 73060 32662 73072 32714
rect 73134 32662 73136 32714
rect 72974 32660 72998 32662
rect 73054 32660 73078 32662
rect 73134 32660 73158 32662
rect 72918 32640 73214 32660
rect 73802 32470 74198 32498
rect 73698 32408 73750 32414
rect 73696 32376 73698 32385
rect 73750 32376 73752 32385
rect 73696 32311 73752 32320
rect 71766 31932 71818 31938
rect 71766 31874 71818 31880
rect 72134 31932 72186 31938
rect 72134 31874 72186 31880
rect 71674 31524 71726 31530
rect 71674 31466 71726 31472
rect 69926 30844 69978 30850
rect 69926 30786 69978 30792
rect 71214 30844 71266 30850
rect 71214 30786 71266 30792
rect 69832 30336 69888 30345
rect 69832 30271 69834 30280
rect 69886 30271 69888 30280
rect 69834 30242 69886 30248
rect 69938 30238 69966 30786
rect 71398 30776 71450 30782
rect 71398 30718 71450 30724
rect 70754 30436 70806 30442
rect 70754 30378 70806 30384
rect 71030 30436 71082 30442
rect 71030 30378 71082 30384
rect 69926 30232 69978 30238
rect 69926 30174 69978 30180
rect 70766 30102 70794 30378
rect 70846 30300 70898 30306
rect 70846 30242 70898 30248
rect 70018 30096 70070 30102
rect 70018 30038 70070 30044
rect 70754 30096 70806 30102
rect 70754 30038 70806 30044
rect 70030 29694 70058 30038
rect 70254 29996 70550 30016
rect 70310 29994 70334 29996
rect 70390 29994 70414 29996
rect 70470 29994 70494 29996
rect 70332 29942 70334 29994
rect 70396 29942 70408 29994
rect 70470 29942 70472 29994
rect 70310 29940 70334 29942
rect 70390 29940 70414 29942
rect 70470 29940 70494 29942
rect 70254 29920 70550 29940
rect 70858 29762 70886 30242
rect 71042 30238 71070 30378
rect 71030 30232 71082 30238
rect 71030 30174 71082 30180
rect 71410 29830 71438 30718
rect 71398 29824 71450 29830
rect 71398 29766 71450 29772
rect 70846 29756 70898 29762
rect 70846 29698 70898 29704
rect 69650 29688 69702 29694
rect 69650 29630 69702 29636
rect 70018 29688 70070 29694
rect 70018 29630 70070 29636
rect 69558 29552 69610 29558
rect 69558 29494 69610 29500
rect 69466 29280 69518 29286
rect 69662 29234 69690 29630
rect 69742 29552 69794 29558
rect 69742 29494 69794 29500
rect 69466 29222 69518 29228
rect 69570 29206 69690 29234
rect 69570 29150 69598 29206
rect 69558 29144 69610 29150
rect 69754 29098 69782 29494
rect 69558 29086 69610 29092
rect 69466 29076 69518 29082
rect 69466 29018 69518 29024
rect 69190 29008 69242 29014
rect 69190 28950 69242 28956
rect 69006 28804 69058 28810
rect 69006 28746 69058 28752
rect 69478 28742 69506 29018
rect 69466 28736 69518 28742
rect 69466 28678 69518 28684
rect 69374 28668 69426 28674
rect 69374 28610 69426 28616
rect 68730 27376 68782 27382
rect 68730 27318 68782 27324
rect 69386 27110 69414 28610
rect 69570 28062 69598 29086
rect 69662 29070 69782 29098
rect 69558 28056 69610 28062
rect 69558 27998 69610 28004
rect 69662 27874 69690 29070
rect 69742 28532 69794 28538
rect 69742 28474 69794 28480
rect 69754 28062 69782 28474
rect 69742 28056 69794 28062
rect 69742 27998 69794 28004
rect 69662 27846 69782 27874
rect 69754 27722 69782 27846
rect 69742 27716 69794 27722
rect 69742 27658 69794 27664
rect 69374 27104 69426 27110
rect 69374 27046 69426 27052
rect 68270 27036 68322 27042
rect 68270 26978 68322 26984
rect 68454 27036 68506 27042
rect 68454 26978 68506 26984
rect 68362 26968 68414 26974
rect 68362 26910 68414 26916
rect 68270 23772 68322 23778
rect 68270 23714 68322 23720
rect 68176 20272 68232 20281
rect 68176 20207 68232 20216
rect 67166 20032 67218 20038
rect 67164 20000 67166 20009
rect 67218 20000 67220 20009
rect 67164 19935 67220 19944
rect 68282 19193 68310 23714
rect 68374 23545 68402 26910
rect 68360 23536 68416 23545
rect 68360 23471 68416 23480
rect 68268 19184 68324 19193
rect 68268 19119 68324 19128
rect 68268 18504 68324 18513
rect 68268 18439 68324 18448
rect 43520 18096 43576 18105
rect 43520 18031 43576 18040
rect 67072 18096 67128 18105
rect 67072 18031 67128 18040
rect 68282 17969 68310 18439
rect 68268 17960 68324 17969
rect 68268 17895 68324 17904
rect 43336 17008 43392 17017
rect 43336 16943 43392 16952
rect 43522 15408 43574 15414
rect 43522 15350 43574 15356
rect 43534 14841 43562 15350
rect 43520 14832 43576 14841
rect 43520 14767 43576 14776
rect 43522 11668 43574 11674
rect 43522 11610 43574 11616
rect 43534 10489 43562 11610
rect 68282 10489 68310 17895
rect 68360 16600 68416 16609
rect 68360 16535 68416 16544
rect 68374 15890 68402 16535
rect 68362 15884 68414 15890
rect 68362 15826 68414 15832
rect 43520 10480 43576 10489
rect 43520 10415 43576 10424
rect 68268 10480 68324 10489
rect 68268 10415 68324 10424
rect 43246 2692 43298 2698
rect 43246 2634 43298 2640
rect 31390 2358 31418 2389
rect 31378 2352 31430 2358
rect 31376 2320 31378 2329
rect 43258 2329 43286 2634
rect 69754 2329 69782 27658
rect 70030 27450 70058 29630
rect 71030 29552 71082 29558
rect 71030 29494 71082 29500
rect 70254 28908 70550 28928
rect 70310 28906 70334 28908
rect 70390 28906 70414 28908
rect 70470 28906 70494 28908
rect 70332 28854 70334 28906
rect 70396 28854 70408 28906
rect 70470 28854 70472 28906
rect 70310 28852 70334 28854
rect 70390 28852 70414 28854
rect 70470 28852 70494 28854
rect 70254 28832 70550 28852
rect 71042 28198 71070 29494
rect 71122 29144 71174 29150
rect 71122 29086 71174 29092
rect 71030 28192 71082 28198
rect 71030 28134 71082 28140
rect 70110 27988 70162 27994
rect 70110 27930 70162 27936
rect 70122 27654 70150 27930
rect 70254 27820 70550 27840
rect 70310 27818 70334 27820
rect 70390 27818 70414 27820
rect 70470 27818 70494 27820
rect 70332 27766 70334 27818
rect 70396 27766 70408 27818
rect 70470 27766 70472 27818
rect 70310 27764 70334 27766
rect 70390 27764 70414 27766
rect 70470 27764 70494 27766
rect 70254 27744 70550 27764
rect 70110 27648 70162 27654
rect 70110 27590 70162 27596
rect 70018 27444 70070 27450
rect 70018 27386 70070 27392
rect 71134 27110 71162 29086
rect 71686 28674 71714 31466
rect 71778 31326 71806 31874
rect 72918 31628 73214 31648
rect 72974 31626 72998 31628
rect 73054 31626 73078 31628
rect 73134 31626 73158 31628
rect 72996 31574 72998 31626
rect 73060 31574 73072 31626
rect 73134 31574 73136 31626
rect 72974 31572 72998 31574
rect 73054 31572 73078 31574
rect 73134 31572 73158 31574
rect 72918 31552 73214 31572
rect 73802 31394 73830 32470
rect 74170 32414 74198 32470
rect 73974 32408 74026 32414
rect 73974 32350 74026 32356
rect 74158 32408 74210 32414
rect 74158 32350 74210 32356
rect 73882 31728 73934 31734
rect 73882 31670 73934 31676
rect 73790 31388 73842 31394
rect 73790 31330 73842 31336
rect 71766 31320 71818 31326
rect 71766 31262 71818 31268
rect 71778 30782 71806 31262
rect 73238 31184 73290 31190
rect 73238 31126 73290 31132
rect 71766 30776 71818 30782
rect 71766 30718 71818 30724
rect 72318 30776 72370 30782
rect 72318 30718 72370 30724
rect 72330 30238 72358 30718
rect 72918 30540 73214 30560
rect 72974 30538 72998 30540
rect 73054 30538 73078 30540
rect 73134 30538 73158 30540
rect 72996 30486 72998 30538
rect 73060 30486 73072 30538
rect 73134 30486 73136 30538
rect 72974 30484 72998 30486
rect 73054 30484 73078 30486
rect 73134 30484 73158 30486
rect 72918 30464 73214 30484
rect 72318 30232 72370 30238
rect 72318 30174 72370 30180
rect 72778 30232 72830 30238
rect 72778 30174 72830 30180
rect 72790 29762 72818 30174
rect 72778 29756 72830 29762
rect 72778 29698 72830 29704
rect 73250 29558 73278 31126
rect 73894 30238 73922 31670
rect 73986 31530 74014 32350
rect 74262 31938 74290 34782
rect 74342 34516 74394 34522
rect 74342 34458 74394 34464
rect 74354 33910 74382 34458
rect 74342 33904 74394 33910
rect 74342 33846 74394 33852
rect 74446 33586 74474 37382
rect 74722 36834 74750 37790
rect 74998 37378 75026 37790
rect 75354 37780 75406 37786
rect 75354 37722 75406 37728
rect 75366 37378 75394 37722
rect 75458 37514 75486 38402
rect 76378 37718 76406 40510
rect 77114 40030 77142 41174
rect 78586 40642 78614 41582
rect 78114 40636 78166 40642
rect 78114 40578 78166 40584
rect 78574 40636 78626 40642
rect 78574 40578 78626 40584
rect 78126 40438 78154 40578
rect 78114 40432 78166 40438
rect 78114 40374 78166 40380
rect 79218 40432 79270 40438
rect 79218 40374 79270 40380
rect 77102 40024 77154 40030
rect 77102 39966 77154 39972
rect 77654 39956 77706 39962
rect 77654 39898 77706 39904
rect 77206 39678 77602 39706
rect 77206 39554 77234 39678
rect 77470 39616 77522 39622
rect 77470 39558 77522 39564
rect 77194 39548 77246 39554
rect 77194 39490 77246 39496
rect 76458 38936 76510 38942
rect 76458 38878 76510 38884
rect 77102 38936 77154 38942
rect 77102 38878 77154 38884
rect 76470 38602 76498 38878
rect 77114 38602 77142 38878
rect 77482 38806 77510 39558
rect 77574 39486 77602 39678
rect 77666 39554 77694 39898
rect 77654 39548 77706 39554
rect 77654 39490 77706 39496
rect 77562 39480 77614 39486
rect 77562 39422 77614 39428
rect 77470 38800 77522 38806
rect 77470 38742 77522 38748
rect 76458 38596 76510 38602
rect 76458 38538 76510 38544
rect 77102 38596 77154 38602
rect 77102 38538 77154 38544
rect 77482 38262 77510 38742
rect 77470 38256 77522 38262
rect 77470 38198 77522 38204
rect 76642 37916 76694 37922
rect 76826 37916 76878 37922
rect 76694 37876 76826 37904
rect 76642 37858 76694 37864
rect 76826 37858 76878 37864
rect 76458 37848 76510 37854
rect 76458 37790 76510 37796
rect 76366 37712 76418 37718
rect 76366 37654 76418 37660
rect 75582 37612 75878 37632
rect 75638 37610 75662 37612
rect 75718 37610 75742 37612
rect 75798 37610 75822 37612
rect 75660 37558 75662 37610
rect 75724 37558 75736 37610
rect 75798 37558 75800 37610
rect 75638 37556 75662 37558
rect 75718 37556 75742 37558
rect 75798 37556 75822 37558
rect 75582 37536 75878 37556
rect 75446 37508 75498 37514
rect 75446 37450 75498 37456
rect 75906 37440 75958 37446
rect 75906 37382 75958 37388
rect 74986 37372 75038 37378
rect 74986 37314 75038 37320
rect 75354 37372 75406 37378
rect 75354 37314 75406 37320
rect 74710 36828 74762 36834
rect 74710 36770 74762 36776
rect 75582 36524 75878 36544
rect 75638 36522 75662 36524
rect 75718 36522 75742 36524
rect 75798 36522 75822 36524
rect 75660 36470 75662 36522
rect 75724 36470 75736 36522
rect 75798 36470 75800 36522
rect 75638 36468 75662 36470
rect 75718 36468 75742 36470
rect 75798 36468 75822 36470
rect 75582 36448 75878 36468
rect 75262 36284 75314 36290
rect 75262 36226 75314 36232
rect 74526 36080 74578 36086
rect 74526 36022 74578 36028
rect 74538 34658 74566 36022
rect 75274 35814 75302 36226
rect 75262 35808 75314 35814
rect 75262 35750 75314 35756
rect 75446 35536 75498 35542
rect 75446 35478 75498 35484
rect 75458 35338 75486 35478
rect 75582 35436 75878 35456
rect 75638 35434 75662 35436
rect 75718 35434 75742 35436
rect 75798 35434 75822 35436
rect 75660 35382 75662 35434
rect 75724 35382 75736 35434
rect 75798 35382 75800 35434
rect 75638 35380 75662 35382
rect 75718 35380 75742 35382
rect 75798 35380 75822 35382
rect 75582 35360 75878 35380
rect 75446 35332 75498 35338
rect 75446 35274 75498 35280
rect 75446 34992 75498 34998
rect 75446 34934 75498 34940
rect 74526 34652 74578 34658
rect 74526 34594 74578 34600
rect 75354 34448 75406 34454
rect 75354 34390 75406 34396
rect 74354 33558 74750 33586
rect 74354 32890 74382 33558
rect 74434 33496 74486 33502
rect 74434 33438 74486 33444
rect 74446 33026 74474 33438
rect 74722 33026 74750 33558
rect 75366 33502 75394 34390
rect 75458 34114 75486 34934
rect 75582 34348 75878 34368
rect 75638 34346 75662 34348
rect 75718 34346 75742 34348
rect 75798 34346 75822 34348
rect 75660 34294 75662 34346
rect 75724 34294 75736 34346
rect 75798 34294 75800 34346
rect 75638 34292 75662 34294
rect 75718 34292 75742 34294
rect 75798 34292 75822 34294
rect 75582 34272 75878 34292
rect 75446 34108 75498 34114
rect 75446 34050 75498 34056
rect 75354 33496 75406 33502
rect 75354 33438 75406 33444
rect 75582 33260 75878 33280
rect 75638 33258 75662 33260
rect 75718 33258 75742 33260
rect 75798 33258 75822 33260
rect 75660 33206 75662 33258
rect 75724 33206 75736 33258
rect 75798 33206 75800 33258
rect 75638 33204 75662 33206
rect 75718 33204 75742 33206
rect 75798 33204 75822 33206
rect 75582 33184 75878 33204
rect 74434 33020 74486 33026
rect 74434 32962 74486 32968
rect 74710 33020 74762 33026
rect 74710 32962 74762 32968
rect 74342 32884 74394 32890
rect 74342 32826 74394 32832
rect 74526 32884 74578 32890
rect 74526 32826 74578 32832
rect 74538 32618 74566 32826
rect 74526 32612 74578 32618
rect 74526 32554 74578 32560
rect 74618 32476 74670 32482
rect 74618 32418 74670 32424
rect 74630 32385 74658 32418
rect 74616 32376 74672 32385
rect 74616 32311 74672 32320
rect 74722 32006 74750 32962
rect 75354 32952 75406 32958
rect 75354 32894 75406 32900
rect 75366 32414 75394 32894
rect 75918 32822 75946 37382
rect 76470 36766 76498 37790
rect 76734 37712 76786 37718
rect 76654 37672 76734 37700
rect 76654 37174 76682 37672
rect 76734 37654 76786 37660
rect 77482 37310 77510 38198
rect 77930 37916 77982 37922
rect 77930 37858 77982 37864
rect 77470 37304 77522 37310
rect 77470 37246 77522 37252
rect 77482 37174 77510 37246
rect 76642 37168 76694 37174
rect 76642 37110 76694 37116
rect 76734 37168 76786 37174
rect 76734 37110 76786 37116
rect 77470 37168 77522 37174
rect 77470 37110 77522 37116
rect 76458 36760 76510 36766
rect 76458 36702 76510 36708
rect 76746 36630 76774 37110
rect 76734 36624 76786 36630
rect 76734 36566 76786 36572
rect 76746 35134 76774 36566
rect 76734 35128 76786 35134
rect 76734 35070 76786 35076
rect 77942 34114 77970 37858
rect 78126 37174 78154 40374
rect 78246 40332 78542 40352
rect 78302 40330 78326 40332
rect 78382 40330 78406 40332
rect 78462 40330 78486 40332
rect 78324 40278 78326 40330
rect 78388 40278 78400 40330
rect 78462 40278 78464 40330
rect 78302 40276 78326 40278
rect 78382 40276 78406 40278
rect 78462 40276 78486 40278
rect 78246 40256 78542 40276
rect 79230 39418 79258 40374
rect 79414 39690 79442 43312
rect 79494 41112 79546 41118
rect 79494 41054 79546 41060
rect 79506 40710 79534 41054
rect 79494 40704 79546 40710
rect 79494 40646 79546 40652
rect 80610 40642 80638 43312
rect 80910 41964 81206 41984
rect 80966 41962 80990 41964
rect 81046 41962 81070 41964
rect 81126 41962 81150 41964
rect 80988 41910 80990 41962
rect 81052 41910 81064 41962
rect 81126 41910 81128 41962
rect 80966 41908 80990 41910
rect 81046 41908 81070 41910
rect 81126 41908 81150 41910
rect 80910 41888 81206 41908
rect 81150 41112 81202 41118
rect 81426 41112 81478 41118
rect 81202 41060 81282 41066
rect 81150 41054 81282 41060
rect 81426 41054 81478 41060
rect 81162 41038 81282 41054
rect 80910 40876 81206 40896
rect 80966 40874 80990 40876
rect 81046 40874 81070 40876
rect 81126 40874 81150 40876
rect 80988 40822 80990 40874
rect 81052 40822 81064 40874
rect 81126 40822 81128 40874
rect 80966 40820 80990 40822
rect 81046 40820 81070 40822
rect 81126 40820 81150 40822
rect 80910 40800 81206 40820
rect 81150 40704 81202 40710
rect 81254 40658 81282 41038
rect 81202 40652 81282 40658
rect 81150 40646 81282 40652
rect 80598 40636 80650 40642
rect 80598 40578 80650 40584
rect 80874 40636 80926 40642
rect 80874 40578 80926 40584
rect 81162 40630 81282 40646
rect 80886 40438 80914 40578
rect 80874 40432 80926 40438
rect 80874 40374 80926 40380
rect 81162 40030 81190 40630
rect 79862 40024 79914 40030
rect 79862 39966 79914 39972
rect 81150 40024 81202 40030
rect 81150 39966 81202 39972
rect 79402 39684 79454 39690
rect 79402 39626 79454 39632
rect 79218 39412 79270 39418
rect 79218 39354 79270 39360
rect 79874 39350 79902 39966
rect 80910 39788 81206 39808
rect 80966 39786 80990 39788
rect 81046 39786 81070 39788
rect 81126 39786 81150 39788
rect 80988 39734 80990 39786
rect 81052 39734 81064 39786
rect 81126 39734 81128 39786
rect 80966 39732 80990 39734
rect 81046 39732 81070 39734
rect 81126 39732 81150 39734
rect 80910 39712 81206 39732
rect 79862 39344 79914 39350
rect 79862 39286 79914 39292
rect 78246 39244 78542 39264
rect 78302 39242 78326 39244
rect 78382 39242 78406 39244
rect 78462 39242 78486 39244
rect 78324 39190 78326 39242
rect 78388 39190 78400 39242
rect 78462 39190 78464 39242
rect 78302 39188 78326 39190
rect 78382 39188 78406 39190
rect 78462 39188 78486 39190
rect 78246 39168 78542 39188
rect 79218 38256 79270 38262
rect 79218 38198 79270 38204
rect 78246 38156 78542 38176
rect 78302 38154 78326 38156
rect 78382 38154 78406 38156
rect 78462 38154 78486 38156
rect 78324 38102 78326 38154
rect 78388 38102 78400 38154
rect 78462 38102 78464 38154
rect 78302 38100 78326 38102
rect 78382 38100 78406 38102
rect 78462 38100 78486 38102
rect 78246 38080 78542 38100
rect 79230 37854 79258 38198
rect 79218 37848 79270 37854
rect 79218 37790 79270 37796
rect 78114 37168 78166 37174
rect 78114 37110 78166 37116
rect 79218 37168 79270 37174
rect 79218 37110 79270 37116
rect 78246 37068 78542 37088
rect 78302 37066 78326 37068
rect 78382 37066 78406 37068
rect 78462 37066 78486 37068
rect 78324 37014 78326 37066
rect 78388 37014 78400 37066
rect 78462 37014 78464 37066
rect 78302 37012 78326 37014
rect 78382 37012 78406 37014
rect 78462 37012 78486 37014
rect 78246 36992 78542 37012
rect 79230 36766 79258 37110
rect 79310 36828 79362 36834
rect 79310 36770 79362 36776
rect 79218 36760 79270 36766
rect 79218 36702 79270 36708
rect 78246 35980 78542 36000
rect 78302 35978 78326 35980
rect 78382 35978 78406 35980
rect 78462 35978 78486 35980
rect 78324 35926 78326 35978
rect 78388 35926 78400 35978
rect 78462 35926 78464 35978
rect 78302 35924 78326 35926
rect 78382 35924 78406 35926
rect 78462 35924 78486 35926
rect 78246 35904 78542 35924
rect 78246 34892 78542 34912
rect 78302 34890 78326 34892
rect 78382 34890 78406 34892
rect 78462 34890 78486 34892
rect 78324 34838 78326 34890
rect 78388 34838 78400 34890
rect 78462 34838 78464 34890
rect 78302 34836 78326 34838
rect 78382 34836 78406 34838
rect 78462 34836 78486 34838
rect 78246 34816 78542 34836
rect 76090 34108 76142 34114
rect 76090 34050 76142 34056
rect 77930 34108 77982 34114
rect 77930 34050 77982 34056
rect 78574 34108 78626 34114
rect 78574 34050 78626 34056
rect 75630 32816 75682 32822
rect 75630 32758 75682 32764
rect 75906 32816 75958 32822
rect 75906 32758 75958 32764
rect 75642 32414 75670 32758
rect 75918 32482 75946 32758
rect 76102 32482 76130 34050
rect 77838 33088 77890 33094
rect 77838 33030 77890 33036
rect 76826 33020 76878 33026
rect 76826 32962 76878 32968
rect 76642 32816 76694 32822
rect 76642 32758 76694 32764
rect 76274 32612 76326 32618
rect 76274 32554 76326 32560
rect 75906 32476 75958 32482
rect 75906 32418 75958 32424
rect 76090 32476 76142 32482
rect 76090 32418 76142 32424
rect 76286 32414 76314 32554
rect 76654 32414 76682 32758
rect 76838 32414 76866 32962
rect 77850 32906 77878 33030
rect 77942 33026 77970 34050
rect 78246 33804 78542 33824
rect 78302 33802 78326 33804
rect 78382 33802 78406 33804
rect 78462 33802 78486 33804
rect 78324 33750 78326 33802
rect 78388 33750 78400 33802
rect 78462 33750 78464 33802
rect 78302 33748 78326 33750
rect 78382 33748 78406 33750
rect 78462 33748 78486 33750
rect 78246 33728 78542 33748
rect 78586 33570 78614 34050
rect 78942 33904 78994 33910
rect 78942 33846 78994 33852
rect 78574 33564 78626 33570
rect 78574 33506 78626 33512
rect 78586 33094 78614 33506
rect 78574 33088 78626 33094
rect 78574 33030 78626 33036
rect 77930 33020 77982 33026
rect 77930 32962 77982 32968
rect 78206 33020 78258 33026
rect 78206 32962 78258 32968
rect 78218 32906 78246 32962
rect 77850 32878 78246 32906
rect 78246 32716 78542 32736
rect 78302 32714 78326 32716
rect 78382 32714 78406 32716
rect 78462 32714 78486 32716
rect 78324 32662 78326 32714
rect 78388 32662 78400 32714
rect 78462 32662 78464 32714
rect 78302 32660 78326 32662
rect 78382 32660 78406 32662
rect 78462 32660 78486 32662
rect 78246 32640 78542 32660
rect 75354 32408 75406 32414
rect 75354 32350 75406 32356
rect 75630 32408 75682 32414
rect 75630 32350 75682 32356
rect 76274 32408 76326 32414
rect 76274 32350 76326 32356
rect 76642 32408 76694 32414
rect 76642 32350 76694 32356
rect 76826 32408 76878 32414
rect 76826 32350 76878 32356
rect 74986 32272 75038 32278
rect 74986 32214 75038 32220
rect 74710 32000 74762 32006
rect 74710 31942 74762 31948
rect 74998 31938 75026 32214
rect 75582 32172 75878 32192
rect 75638 32170 75662 32172
rect 75718 32170 75742 32172
rect 75798 32170 75822 32172
rect 75660 32118 75662 32170
rect 75724 32118 75736 32170
rect 75798 32118 75800 32170
rect 75638 32116 75662 32118
rect 75718 32116 75742 32118
rect 75798 32116 75822 32118
rect 75582 32096 75878 32116
rect 76838 32006 76866 32350
rect 76918 32272 76970 32278
rect 76918 32214 76970 32220
rect 76826 32000 76878 32006
rect 76826 31942 76878 31948
rect 74250 31932 74302 31938
rect 74250 31874 74302 31880
rect 74986 31932 75038 31938
rect 74986 31874 75038 31880
rect 75446 31864 75498 31870
rect 75446 31806 75498 31812
rect 75354 31728 75406 31734
rect 75354 31670 75406 31676
rect 73974 31524 74026 31530
rect 73974 31466 74026 31472
rect 75366 31326 75394 31670
rect 74158 31320 74210 31326
rect 74158 31262 74210 31268
rect 75354 31320 75406 31326
rect 75354 31262 75406 31268
rect 74170 30850 74198 31262
rect 74342 31252 74394 31258
rect 74342 31194 74394 31200
rect 74158 30844 74210 30850
rect 74158 30786 74210 30792
rect 74354 30714 74382 31194
rect 75366 31002 75394 31262
rect 75274 30974 75394 31002
rect 75274 30918 75302 30974
rect 75262 30912 75314 30918
rect 75262 30854 75314 30860
rect 75078 30844 75130 30850
rect 75078 30786 75130 30792
rect 74342 30708 74394 30714
rect 74342 30650 74394 30656
rect 74434 30708 74486 30714
rect 74434 30650 74486 30656
rect 73882 30232 73934 30238
rect 73882 30174 73934 30180
rect 74354 30102 74382 30650
rect 74446 30442 74474 30650
rect 74434 30436 74486 30442
rect 74434 30378 74486 30384
rect 74526 30436 74578 30442
rect 74526 30378 74578 30384
rect 74538 30345 74566 30378
rect 74524 30336 74580 30345
rect 74524 30271 74580 30280
rect 75090 30170 75118 30786
rect 75458 30714 75486 31806
rect 76550 31320 76602 31326
rect 76550 31262 76602 31268
rect 75582 31084 75878 31104
rect 75638 31082 75662 31084
rect 75718 31082 75742 31084
rect 75798 31082 75822 31084
rect 75660 31030 75662 31082
rect 75724 31030 75736 31082
rect 75798 31030 75800 31082
rect 75638 31028 75662 31030
rect 75718 31028 75742 31030
rect 75798 31028 75822 31030
rect 75582 31008 75878 31028
rect 75538 30844 75590 30850
rect 75538 30786 75590 30792
rect 75446 30708 75498 30714
rect 75446 30650 75498 30656
rect 75550 30306 75578 30786
rect 75538 30300 75590 30306
rect 75538 30242 75590 30248
rect 75998 30232 76050 30238
rect 75998 30174 76050 30180
rect 76182 30232 76234 30238
rect 76182 30174 76234 30180
rect 75078 30164 75130 30170
rect 75078 30106 75130 30112
rect 74158 30096 74210 30102
rect 74158 30038 74210 30044
rect 74342 30096 74394 30102
rect 74342 30038 74394 30044
rect 74710 30096 74762 30102
rect 74710 30038 74762 30044
rect 74170 29830 74198 30038
rect 74158 29824 74210 29830
rect 74158 29766 74210 29772
rect 74354 29762 74382 30038
rect 74342 29756 74394 29762
rect 74342 29698 74394 29704
rect 74722 29694 74750 30038
rect 74984 29792 75040 29801
rect 74984 29727 74986 29736
rect 75038 29727 75040 29736
rect 74986 29698 75038 29704
rect 74710 29688 74762 29694
rect 74710 29630 74762 29636
rect 73238 29552 73290 29558
rect 73238 29494 73290 29500
rect 72918 29452 73214 29472
rect 72974 29450 72998 29452
rect 73054 29450 73078 29452
rect 73134 29450 73158 29452
rect 72996 29398 72998 29450
rect 73060 29398 73072 29450
rect 73134 29398 73136 29450
rect 72974 29396 72998 29398
rect 73054 29396 73078 29398
rect 73134 29396 73158 29398
rect 72918 29376 73214 29396
rect 73250 28742 73278 29494
rect 74998 29218 75026 29698
rect 75090 29694 75118 30106
rect 75354 30096 75406 30102
rect 75906 30096 75958 30102
rect 75406 30056 75486 30084
rect 75354 30038 75406 30044
rect 75170 29756 75222 29762
rect 75170 29698 75222 29704
rect 75078 29688 75130 29694
rect 75078 29630 75130 29636
rect 75182 29626 75210 29698
rect 75458 29676 75486 30056
rect 75906 30038 75958 30044
rect 75582 29996 75878 30016
rect 75638 29994 75662 29996
rect 75718 29994 75742 29996
rect 75798 29994 75822 29996
rect 75660 29942 75662 29994
rect 75724 29942 75736 29994
rect 75798 29942 75800 29994
rect 75638 29940 75662 29942
rect 75718 29940 75742 29942
rect 75798 29940 75822 29942
rect 75582 29920 75878 29940
rect 75918 29830 75946 30038
rect 76010 29830 76038 30174
rect 75906 29824 75958 29830
rect 75906 29766 75958 29772
rect 75998 29824 76050 29830
rect 75998 29766 76050 29772
rect 75538 29688 75590 29694
rect 75458 29648 75538 29676
rect 75538 29630 75590 29636
rect 75998 29688 76050 29694
rect 76194 29676 76222 30174
rect 76274 29824 76326 29830
rect 76274 29766 76326 29772
rect 76050 29648 76222 29676
rect 75998 29630 76050 29636
rect 75170 29620 75222 29626
rect 75170 29562 75222 29568
rect 74986 29212 75038 29218
rect 74986 29154 75038 29160
rect 74250 29144 74302 29150
rect 74250 29086 74302 29092
rect 73698 29008 73750 29014
rect 73698 28950 73750 28956
rect 73238 28736 73290 28742
rect 73238 28678 73290 28684
rect 71674 28668 71726 28674
rect 71674 28610 71726 28616
rect 73606 28668 73658 28674
rect 73606 28610 73658 28616
rect 71686 27586 71714 28610
rect 72686 28464 72738 28470
rect 72686 28406 72738 28412
rect 72698 28062 72726 28406
rect 72918 28364 73214 28384
rect 72974 28362 72998 28364
rect 73054 28362 73078 28364
rect 73134 28362 73158 28364
rect 72996 28310 72998 28362
rect 73060 28310 73072 28362
rect 73134 28310 73136 28362
rect 72974 28308 72998 28310
rect 73054 28308 73078 28310
rect 73134 28308 73158 28310
rect 72918 28288 73214 28308
rect 73330 28192 73382 28198
rect 73330 28134 73382 28140
rect 72686 28056 72738 28062
rect 72686 27998 72738 28004
rect 73054 27988 73106 27994
rect 73054 27930 73106 27936
rect 73066 27654 73094 27930
rect 73054 27648 73106 27654
rect 73054 27590 73106 27596
rect 71674 27580 71726 27586
rect 71674 27522 71726 27528
rect 72318 27512 72370 27518
rect 72318 27454 72370 27460
rect 71950 27376 72002 27382
rect 71950 27318 72002 27324
rect 71122 27104 71174 27110
rect 71122 27046 71174 27052
rect 70110 27036 70162 27042
rect 70110 26978 70162 26984
rect 70018 26900 70070 26906
rect 70018 26842 70070 26848
rect 69926 26832 69978 26838
rect 69926 26774 69978 26780
rect 69938 26294 69966 26774
rect 69926 26288 69978 26294
rect 69926 26230 69978 26236
rect 70030 24186 70058 26842
rect 70122 25562 70150 26978
rect 71962 26906 71990 27318
rect 72330 27042 72358 27454
rect 72918 27276 73214 27296
rect 72974 27274 72998 27276
rect 73054 27274 73078 27276
rect 73134 27274 73158 27276
rect 72996 27222 72998 27274
rect 73060 27222 73072 27274
rect 73134 27222 73136 27274
rect 72974 27220 72998 27222
rect 73054 27220 73078 27222
rect 73134 27220 73158 27222
rect 72918 27200 73214 27220
rect 72318 27036 72370 27042
rect 72318 26978 72370 26984
rect 73342 26974 73370 28134
rect 73618 28130 73646 28610
rect 73606 28124 73658 28130
rect 73606 28066 73658 28072
rect 73710 28062 73738 28950
rect 73882 28736 73934 28742
rect 73882 28678 73934 28684
rect 73698 28056 73750 28062
rect 73698 27998 73750 28004
rect 73790 28056 73842 28062
rect 73790 27998 73842 28004
rect 73710 27586 73738 27998
rect 73698 27580 73750 27586
rect 73698 27522 73750 27528
rect 73802 27382 73830 27998
rect 73894 27382 73922 28678
rect 74066 28600 74118 28606
rect 74066 28542 74118 28548
rect 74078 28130 74106 28542
rect 74262 28266 74290 29086
rect 74618 29076 74670 29082
rect 74618 29018 74670 29024
rect 74630 28810 74658 29018
rect 75582 28908 75878 28928
rect 75638 28906 75662 28908
rect 75718 28906 75742 28908
rect 75798 28906 75822 28908
rect 75660 28854 75662 28906
rect 75724 28854 75736 28906
rect 75798 28854 75800 28906
rect 75638 28852 75662 28854
rect 75718 28852 75742 28854
rect 75798 28852 75822 28854
rect 75582 28832 75878 28852
rect 74618 28804 74670 28810
rect 74618 28746 74670 28752
rect 74250 28260 74302 28266
rect 74250 28202 74302 28208
rect 74066 28124 74118 28130
rect 74066 28066 74118 28072
rect 75582 27820 75878 27840
rect 75638 27818 75662 27820
rect 75718 27818 75742 27820
rect 75798 27818 75822 27820
rect 75660 27766 75662 27818
rect 75724 27766 75736 27818
rect 75798 27766 75800 27818
rect 75638 27764 75662 27766
rect 75718 27764 75742 27766
rect 75798 27764 75822 27766
rect 75582 27744 75878 27764
rect 76194 27722 76222 29648
rect 76286 29558 76314 29766
rect 76562 29626 76590 31262
rect 76930 30442 76958 32214
rect 78586 32006 78614 33030
rect 77470 32000 77522 32006
rect 77470 31942 77522 31948
rect 78574 32000 78626 32006
rect 78574 31942 78626 31948
rect 77378 31932 77430 31938
rect 77378 31874 77430 31880
rect 77102 31728 77154 31734
rect 77102 31670 77154 31676
rect 77114 30782 77142 31670
rect 77102 30776 77154 30782
rect 77102 30718 77154 30724
rect 77010 30708 77062 30714
rect 77010 30650 77062 30656
rect 76918 30436 76970 30442
rect 76918 30378 76970 30384
rect 76918 30300 76970 30306
rect 76918 30242 76970 30248
rect 76642 30232 76694 30238
rect 76642 30174 76694 30180
rect 76654 29801 76682 30174
rect 76640 29792 76696 29801
rect 76640 29727 76696 29736
rect 76930 29694 76958 30242
rect 77022 29694 77050 30650
rect 77114 30442 77142 30718
rect 77102 30436 77154 30442
rect 77102 30378 77154 30384
rect 77390 29898 77418 31874
rect 77482 30850 77510 31942
rect 78246 31628 78542 31648
rect 78302 31626 78326 31628
rect 78382 31626 78406 31628
rect 78462 31626 78486 31628
rect 78324 31574 78326 31626
rect 78388 31574 78400 31626
rect 78462 31574 78464 31626
rect 78302 31572 78326 31574
rect 78382 31572 78406 31574
rect 78462 31572 78486 31574
rect 78246 31552 78542 31572
rect 77470 30844 77522 30850
rect 77470 30786 77522 30792
rect 77482 30238 77510 30786
rect 78114 30776 78166 30782
rect 78114 30718 78166 30724
rect 77746 30640 77798 30646
rect 77746 30582 77798 30588
rect 78022 30640 78074 30646
rect 78022 30582 78074 30588
rect 77758 30306 77786 30582
rect 78034 30442 78062 30582
rect 78022 30436 78074 30442
rect 78022 30378 78074 30384
rect 77746 30300 77798 30306
rect 77746 30242 77798 30248
rect 77470 30232 77522 30238
rect 77470 30174 77522 30180
rect 78022 30164 78074 30170
rect 78022 30106 78074 30112
rect 77378 29892 77430 29898
rect 77378 29834 77430 29840
rect 77746 29892 77798 29898
rect 77746 29834 77798 29840
rect 76918 29688 76970 29694
rect 76918 29630 76970 29636
rect 77010 29688 77062 29694
rect 77010 29630 77062 29636
rect 76550 29620 76602 29626
rect 76550 29562 76602 29568
rect 76274 29552 76326 29558
rect 76274 29494 76326 29500
rect 76918 29552 76970 29558
rect 76918 29494 76970 29500
rect 76930 29286 76958 29494
rect 76918 29280 76970 29286
rect 76918 29222 76970 29228
rect 77758 29150 77786 29834
rect 78034 29762 78062 30106
rect 78126 29898 78154 30718
rect 78246 30540 78542 30560
rect 78302 30538 78326 30540
rect 78382 30538 78406 30540
rect 78462 30538 78486 30540
rect 78324 30486 78326 30538
rect 78388 30486 78400 30538
rect 78462 30486 78464 30538
rect 78302 30484 78326 30486
rect 78382 30484 78406 30486
rect 78462 30484 78486 30486
rect 78246 30464 78542 30484
rect 78114 29892 78166 29898
rect 78114 29834 78166 29840
rect 78022 29756 78074 29762
rect 78022 29698 78074 29704
rect 78246 29452 78542 29472
rect 78302 29450 78326 29452
rect 78382 29450 78406 29452
rect 78462 29450 78486 29452
rect 78324 29398 78326 29450
rect 78388 29398 78400 29450
rect 78462 29398 78464 29450
rect 78302 29396 78326 29398
rect 78382 29396 78406 29398
rect 78462 29396 78486 29398
rect 78246 29376 78542 29396
rect 77746 29144 77798 29150
rect 77746 29086 77798 29092
rect 77562 29008 77614 29014
rect 77562 28950 77614 28956
rect 77574 28062 77602 28950
rect 78246 28364 78542 28384
rect 78302 28362 78326 28364
rect 78382 28362 78406 28364
rect 78462 28362 78486 28364
rect 78324 28310 78326 28362
rect 78388 28310 78400 28362
rect 78462 28310 78464 28362
rect 78302 28308 78326 28310
rect 78382 28308 78406 28310
rect 78462 28308 78486 28310
rect 78246 28288 78542 28308
rect 77562 28056 77614 28062
rect 77562 27998 77614 28004
rect 76182 27716 76234 27722
rect 76182 27658 76234 27664
rect 78586 27568 78614 31942
rect 78850 31864 78902 31870
rect 78850 31806 78902 31812
rect 78666 31728 78718 31734
rect 78666 31670 78718 31676
rect 78678 31530 78706 31670
rect 78666 31524 78718 31530
rect 78666 31466 78718 31472
rect 78862 30646 78890 31806
rect 78850 30640 78902 30646
rect 78850 30582 78902 30588
rect 78954 29762 78982 33846
rect 79322 33502 79350 36770
rect 79874 33502 79902 39286
rect 80414 38800 80466 38806
rect 80414 38742 80466 38748
rect 80426 38466 80454 38742
rect 80910 38700 81206 38720
rect 80966 38698 80990 38700
rect 81046 38698 81070 38700
rect 81126 38698 81150 38700
rect 80988 38646 80990 38698
rect 81052 38646 81064 38698
rect 81126 38646 81128 38698
rect 80966 38644 80990 38646
rect 81046 38644 81070 38646
rect 81126 38644 81150 38646
rect 80910 38624 81206 38644
rect 80414 38460 80466 38466
rect 80414 38402 80466 38408
rect 80322 37168 80374 37174
rect 80322 37110 80374 37116
rect 80334 36970 80362 37110
rect 80322 36964 80374 36970
rect 80322 36906 80374 36912
rect 80230 35536 80282 35542
rect 80230 35478 80282 35484
rect 80242 34590 80270 35478
rect 80230 34584 80282 34590
rect 80230 34526 80282 34532
rect 79954 34176 80006 34182
rect 79954 34118 80006 34124
rect 79966 33502 79994 34118
rect 80426 34114 80454 38402
rect 80910 37612 81206 37632
rect 80966 37610 80990 37612
rect 81046 37610 81070 37612
rect 81126 37610 81150 37612
rect 80988 37558 80990 37610
rect 81052 37558 81064 37610
rect 81126 37558 81128 37610
rect 80966 37556 80990 37558
rect 81046 37556 81070 37558
rect 81126 37556 81150 37558
rect 80910 37536 81206 37556
rect 80910 36524 81206 36544
rect 80966 36522 80990 36524
rect 81046 36522 81070 36524
rect 81126 36522 81150 36524
rect 80988 36470 80990 36522
rect 81052 36470 81064 36522
rect 81126 36470 81128 36522
rect 80966 36468 80990 36470
rect 81046 36468 81070 36470
rect 81126 36468 81150 36470
rect 80910 36448 81206 36468
rect 80690 35876 80742 35882
rect 80690 35818 80742 35824
rect 80702 35338 80730 35818
rect 80910 35436 81206 35456
rect 80966 35434 80990 35436
rect 81046 35434 81070 35436
rect 81126 35434 81150 35436
rect 80988 35382 80990 35434
rect 81052 35382 81064 35434
rect 81126 35382 81128 35434
rect 80966 35380 80990 35382
rect 81046 35380 81070 35382
rect 81126 35380 81150 35382
rect 80910 35360 81206 35380
rect 80690 35332 80742 35338
rect 80690 35274 80742 35280
rect 80702 34250 80730 35274
rect 80874 35264 80926 35270
rect 80874 35206 80926 35212
rect 80886 34726 80914 35206
rect 81150 35196 81202 35202
rect 81150 35138 81202 35144
rect 81162 34726 81190 35138
rect 80874 34720 80926 34726
rect 80874 34662 80926 34668
rect 81150 34720 81202 34726
rect 81150 34662 81202 34668
rect 81334 34652 81386 34658
rect 81334 34594 81386 34600
rect 80782 34584 80834 34590
rect 80782 34526 80834 34532
rect 81242 34584 81294 34590
rect 81242 34526 81294 34532
rect 80794 34454 80822 34526
rect 80782 34448 80834 34454
rect 80782 34390 80834 34396
rect 80910 34348 81206 34368
rect 80966 34346 80990 34348
rect 81046 34346 81070 34348
rect 81126 34346 81150 34348
rect 80988 34294 80990 34346
rect 81052 34294 81064 34346
rect 81126 34294 81128 34346
rect 80966 34292 80990 34294
rect 81046 34292 81070 34294
rect 81126 34292 81150 34294
rect 80910 34272 81206 34292
rect 80690 34244 80742 34250
rect 80690 34186 80742 34192
rect 81254 34182 81282 34526
rect 81346 34454 81374 34594
rect 81334 34448 81386 34454
rect 81334 34390 81386 34396
rect 81242 34176 81294 34182
rect 81242 34118 81294 34124
rect 80414 34108 80466 34114
rect 80414 34050 80466 34056
rect 80426 33570 80454 34050
rect 80414 33564 80466 33570
rect 80414 33506 80466 33512
rect 79310 33496 79362 33502
rect 79310 33438 79362 33444
rect 79862 33496 79914 33502
rect 79862 33438 79914 33444
rect 79954 33496 80006 33502
rect 79954 33438 80006 33444
rect 80598 33496 80650 33502
rect 80598 33438 80650 33444
rect 79322 31938 79350 33438
rect 79874 32482 79902 33438
rect 79862 32476 79914 32482
rect 79862 32418 79914 32424
rect 80414 32408 80466 32414
rect 80414 32350 80466 32356
rect 80426 31938 80454 32350
rect 79310 31932 79362 31938
rect 79310 31874 79362 31880
rect 79678 31932 79730 31938
rect 79678 31874 79730 31880
rect 80414 31932 80466 31938
rect 80414 31874 80466 31880
rect 79690 30986 79718 31874
rect 80610 31734 80638 33438
rect 80910 33260 81206 33280
rect 80966 33258 80990 33260
rect 81046 33258 81070 33260
rect 81126 33258 81150 33260
rect 80988 33206 80990 33258
rect 81052 33206 81064 33258
rect 81126 33206 81128 33258
rect 80966 33204 80990 33206
rect 81046 33204 81070 33206
rect 81126 33204 81150 33206
rect 80910 33184 81206 33204
rect 81438 32906 81466 41054
rect 81806 35678 81834 43312
rect 83094 41322 83122 43312
rect 84290 43242 84318 43312
rect 84290 43214 84410 43242
rect 83574 41420 83870 41440
rect 83630 41418 83654 41420
rect 83710 41418 83734 41420
rect 83790 41418 83814 41420
rect 83652 41366 83654 41418
rect 83716 41366 83728 41418
rect 83790 41366 83792 41418
rect 83630 41364 83654 41366
rect 83710 41364 83734 41366
rect 83790 41364 83814 41366
rect 83574 41344 83870 41364
rect 83082 41316 83134 41322
rect 83082 41258 83134 41264
rect 83634 41180 83686 41186
rect 83634 41122 83686 41128
rect 82346 40772 82398 40778
rect 82346 40714 82398 40720
rect 82070 40636 82122 40642
rect 82070 40578 82122 40584
rect 82082 39554 82110 40578
rect 82358 40098 82386 40714
rect 82530 40636 82582 40642
rect 82530 40578 82582 40584
rect 82346 40092 82398 40098
rect 82346 40034 82398 40040
rect 82070 39548 82122 39554
rect 82070 39490 82122 39496
rect 82070 38052 82122 38058
rect 82070 37994 82122 38000
rect 82082 37378 82110 37994
rect 82162 37848 82214 37854
rect 82162 37790 82214 37796
rect 82070 37372 82122 37378
rect 82070 37314 82122 37320
rect 82174 36970 82202 37790
rect 82162 36964 82214 36970
rect 82162 36906 82214 36912
rect 82174 36426 82202 36906
rect 82542 36426 82570 40578
rect 83646 40574 83674 41122
rect 83634 40568 83686 40574
rect 83634 40510 83686 40516
rect 84186 40568 84238 40574
rect 84186 40510 84238 40516
rect 83574 40332 83870 40352
rect 83630 40330 83654 40332
rect 83710 40330 83734 40332
rect 83790 40330 83814 40332
rect 83652 40278 83654 40330
rect 83716 40278 83728 40330
rect 83790 40278 83792 40330
rect 83630 40276 83654 40278
rect 83710 40276 83734 40278
rect 83790 40276 83814 40278
rect 83574 40256 83870 40276
rect 83726 40160 83778 40166
rect 83726 40102 83778 40108
rect 82806 39888 82858 39894
rect 82806 39830 82858 39836
rect 82818 38466 82846 39830
rect 83738 39622 83766 40102
rect 83910 40024 83962 40030
rect 83910 39966 83962 39972
rect 83726 39616 83778 39622
rect 83726 39558 83778 39564
rect 83922 39554 83950 39966
rect 84198 39690 84226 40510
rect 84186 39684 84238 39690
rect 84186 39626 84238 39632
rect 83910 39548 83962 39554
rect 83910 39490 83962 39496
rect 83574 39244 83870 39264
rect 83630 39242 83654 39244
rect 83710 39242 83734 39244
rect 83790 39242 83814 39244
rect 83652 39190 83654 39242
rect 83716 39190 83728 39242
rect 83790 39190 83792 39242
rect 83630 39188 83654 39190
rect 83710 39188 83734 39190
rect 83790 39188 83814 39190
rect 83574 39168 83870 39188
rect 82806 38460 82858 38466
rect 82806 38402 82858 38408
rect 83266 38460 83318 38466
rect 83266 38402 83318 38408
rect 82818 37990 82846 38402
rect 82806 37984 82858 37990
rect 82806 37926 82858 37932
rect 83278 37514 83306 38402
rect 83574 38156 83870 38176
rect 83630 38154 83654 38156
rect 83710 38154 83734 38156
rect 83790 38154 83814 38156
rect 83652 38102 83654 38154
rect 83716 38102 83728 38154
rect 83790 38102 83792 38154
rect 83630 38100 83654 38102
rect 83710 38100 83734 38102
rect 83790 38100 83814 38102
rect 83574 38080 83870 38100
rect 84278 37780 84330 37786
rect 84278 37722 84330 37728
rect 84002 37712 84054 37718
rect 84002 37654 84054 37660
rect 83266 37508 83318 37514
rect 83266 37450 83318 37456
rect 82714 37168 82766 37174
rect 82714 37110 82766 37116
rect 83910 37168 83962 37174
rect 83910 37110 83962 37116
rect 82726 36766 82754 37110
rect 83574 37068 83870 37088
rect 83630 37066 83654 37068
rect 83710 37066 83734 37068
rect 83790 37066 83814 37068
rect 83652 37014 83654 37066
rect 83716 37014 83728 37066
rect 83790 37014 83792 37066
rect 83630 37012 83654 37014
rect 83710 37012 83734 37014
rect 83790 37012 83814 37014
rect 83574 36992 83870 37012
rect 82714 36760 82766 36766
rect 82714 36702 82766 36708
rect 82162 36420 82214 36426
rect 82162 36362 82214 36368
rect 82530 36420 82582 36426
rect 82530 36362 82582 36368
rect 82726 36290 82754 36702
rect 83082 36624 83134 36630
rect 83082 36566 83134 36572
rect 83094 36290 83122 36566
rect 82714 36284 82766 36290
rect 82714 36226 82766 36232
rect 83082 36284 83134 36290
rect 83082 36226 83134 36232
rect 82530 36216 82582 36222
rect 82530 36158 82582 36164
rect 81794 35672 81846 35678
rect 81794 35614 81846 35620
rect 82070 35672 82122 35678
rect 82070 35614 82122 35620
rect 81702 35536 81754 35542
rect 81702 35478 81754 35484
rect 81518 33700 81570 33706
rect 81518 33642 81570 33648
rect 81346 32878 81466 32906
rect 81530 32890 81558 33642
rect 81714 33638 81742 35478
rect 82082 35270 82110 35614
rect 82070 35264 82122 35270
rect 82070 35206 82122 35212
rect 82542 34590 82570 36158
rect 82714 36148 82766 36154
rect 82714 36090 82766 36096
rect 82726 35678 82754 36090
rect 83574 35980 83870 36000
rect 83630 35978 83654 35980
rect 83710 35978 83734 35980
rect 83790 35978 83814 35980
rect 83652 35926 83654 35978
rect 83716 35926 83728 35978
rect 83790 35926 83792 35978
rect 83630 35924 83654 35926
rect 83710 35924 83734 35926
rect 83790 35924 83814 35926
rect 83574 35904 83870 35924
rect 82714 35672 82766 35678
rect 82714 35614 82766 35620
rect 82530 34584 82582 34590
rect 82530 34526 82582 34532
rect 82346 34448 82398 34454
rect 82346 34390 82398 34396
rect 81702 33632 81754 33638
rect 81702 33574 81754 33580
rect 82358 33502 82386 34390
rect 82346 33496 82398 33502
rect 82346 33438 82398 33444
rect 82254 33428 82306 33434
rect 82254 33370 82306 33376
rect 81518 32884 81570 32890
rect 81346 32346 81374 32878
rect 81518 32826 81570 32832
rect 81426 32816 81478 32822
rect 81426 32758 81478 32764
rect 81438 32550 81466 32758
rect 81426 32544 81478 32550
rect 81426 32486 81478 32492
rect 82266 32346 82294 33370
rect 82542 32414 82570 34526
rect 82726 34454 82754 35614
rect 83542 35604 83594 35610
rect 83542 35546 83594 35552
rect 83554 35202 83582 35546
rect 83922 35338 83950 37110
rect 84014 36902 84042 37654
rect 84290 37378 84318 37722
rect 84278 37372 84330 37378
rect 84278 37314 84330 37320
rect 84002 36896 84054 36902
rect 84002 36838 84054 36844
rect 83910 35332 83962 35338
rect 83910 35274 83962 35280
rect 83542 35196 83594 35202
rect 83542 35138 83594 35144
rect 84278 35060 84330 35066
rect 84278 35002 84330 35008
rect 82898 34992 82950 34998
rect 82898 34934 82950 34940
rect 82714 34448 82766 34454
rect 82714 34390 82766 34396
rect 82714 33428 82766 33434
rect 82714 33370 82766 33376
rect 82622 32476 82674 32482
rect 82622 32418 82674 32424
rect 82530 32408 82582 32414
rect 82530 32350 82582 32356
rect 81334 32340 81386 32346
rect 81334 32282 81386 32288
rect 82254 32340 82306 32346
rect 82254 32282 82306 32288
rect 80910 32172 81206 32192
rect 80966 32170 80990 32172
rect 81046 32170 81070 32172
rect 81126 32170 81150 32172
rect 80988 32118 80990 32170
rect 81052 32118 81064 32170
rect 81126 32118 81128 32170
rect 80966 32116 80990 32118
rect 81046 32116 81070 32118
rect 81126 32116 81150 32118
rect 80910 32096 81206 32116
rect 80598 31728 80650 31734
rect 80598 31670 80650 31676
rect 80610 31258 80638 31670
rect 82634 31326 82662 32418
rect 82726 32414 82754 33370
rect 82910 33162 82938 34934
rect 83574 34892 83870 34912
rect 83630 34890 83654 34892
rect 83710 34890 83734 34892
rect 83790 34890 83814 34892
rect 83652 34838 83654 34890
rect 83716 34838 83728 34890
rect 83790 34838 83792 34890
rect 83630 34836 83654 34838
rect 83710 34836 83734 34838
rect 83790 34836 83814 34838
rect 83574 34816 83870 34836
rect 84290 34794 84318 35002
rect 84278 34788 84330 34794
rect 84278 34730 84330 34736
rect 83574 33804 83870 33824
rect 83630 33802 83654 33804
rect 83710 33802 83734 33804
rect 83790 33802 83814 33804
rect 83652 33750 83654 33802
rect 83716 33750 83728 33802
rect 83790 33750 83792 33802
rect 83630 33748 83654 33750
rect 83710 33748 83734 33750
rect 83790 33748 83814 33750
rect 83574 33728 83870 33748
rect 84382 33473 84410 43214
rect 85014 40976 85066 40982
rect 85014 40918 85066 40924
rect 85026 40642 85054 40918
rect 85486 40642 85514 43312
rect 91650 42154 91678 43312
rect 91282 42126 91678 42154
rect 86238 41964 86534 41984
rect 86294 41962 86318 41964
rect 86374 41962 86398 41964
rect 86454 41962 86478 41964
rect 86316 41910 86318 41962
rect 86380 41910 86392 41962
rect 86454 41910 86456 41962
rect 86294 41908 86318 41910
rect 86374 41908 86398 41910
rect 86454 41908 86478 41910
rect 86238 41888 86534 41908
rect 88142 41656 88194 41662
rect 88142 41598 88194 41604
rect 89338 41656 89390 41662
rect 89338 41598 89390 41604
rect 85658 41112 85710 41118
rect 85658 41054 85710 41060
rect 85014 40636 85066 40642
rect 85014 40578 85066 40584
rect 85474 40636 85526 40642
rect 85474 40578 85526 40584
rect 84462 39548 84514 39554
rect 84462 39490 84514 39496
rect 84474 36834 84502 39490
rect 84922 37848 84974 37854
rect 85026 37836 85054 40578
rect 85670 39894 85698 41054
rect 88154 40982 88182 41598
rect 88902 41420 89198 41440
rect 88958 41418 88982 41420
rect 89038 41418 89062 41420
rect 89118 41418 89142 41420
rect 88980 41366 88982 41418
rect 89044 41366 89056 41418
rect 89118 41366 89120 41418
rect 88958 41364 88982 41366
rect 89038 41364 89062 41366
rect 89118 41364 89142 41366
rect 88902 41344 89198 41364
rect 88142 40976 88194 40982
rect 88142 40918 88194 40924
rect 86238 40876 86534 40896
rect 86294 40874 86318 40876
rect 86374 40874 86398 40876
rect 86454 40874 86478 40876
rect 86316 40822 86318 40874
rect 86380 40822 86392 40874
rect 86454 40822 86456 40874
rect 86294 40820 86318 40822
rect 86374 40820 86398 40822
rect 86454 40820 86478 40822
rect 86238 40800 86534 40820
rect 88154 40778 88182 40918
rect 88142 40772 88194 40778
rect 88142 40714 88194 40720
rect 88154 40574 88182 40714
rect 88142 40568 88194 40574
rect 88510 40568 88562 40574
rect 88194 40516 88366 40522
rect 88142 40510 88366 40516
rect 88510 40510 88562 40516
rect 88154 40494 88366 40510
rect 88142 40432 88194 40438
rect 88142 40374 88194 40380
rect 85842 40024 85894 40030
rect 85842 39966 85894 39972
rect 85658 39888 85710 39894
rect 85658 39830 85710 39836
rect 85106 38392 85158 38398
rect 85106 38334 85158 38340
rect 85118 37922 85146 38334
rect 85290 38256 85342 38262
rect 85290 38198 85342 38204
rect 85106 37916 85158 37922
rect 85106 37858 85158 37864
rect 84974 37808 85054 37836
rect 84922 37790 84974 37796
rect 84462 36828 84514 36834
rect 84462 36770 84514 36776
rect 85302 36630 85330 38198
rect 85474 36896 85526 36902
rect 85474 36838 85526 36844
rect 85486 36766 85514 36838
rect 85474 36760 85526 36766
rect 85474 36702 85526 36708
rect 85290 36624 85342 36630
rect 85290 36566 85342 36572
rect 84646 34992 84698 34998
rect 84646 34934 84698 34940
rect 84658 34590 84686 34934
rect 84646 34584 84698 34590
rect 84646 34526 84698 34532
rect 85302 33706 85330 36566
rect 85486 35746 85514 36702
rect 85658 36080 85710 36086
rect 85658 36022 85710 36028
rect 85474 35740 85526 35746
rect 85474 35682 85526 35688
rect 85670 35678 85698 36022
rect 85854 35882 85882 39966
rect 86238 39788 86534 39808
rect 86294 39786 86318 39788
rect 86374 39786 86398 39788
rect 86454 39786 86478 39788
rect 86316 39734 86318 39786
rect 86380 39734 86392 39786
rect 86454 39734 86456 39786
rect 86294 39732 86318 39734
rect 86374 39732 86398 39734
rect 86454 39732 86478 39734
rect 86238 39712 86534 39732
rect 88154 39486 88182 40374
rect 88338 39622 88366 40494
rect 88418 40092 88470 40098
rect 88418 40034 88470 40040
rect 88234 39616 88286 39622
rect 88234 39558 88286 39564
rect 88326 39616 88378 39622
rect 88326 39558 88378 39564
rect 88142 39480 88194 39486
rect 88142 39422 88194 39428
rect 86238 38700 86534 38720
rect 86294 38698 86318 38700
rect 86374 38698 86398 38700
rect 86454 38698 86478 38700
rect 86316 38646 86318 38698
rect 86380 38646 86392 38698
rect 86454 38646 86456 38698
rect 86294 38644 86318 38646
rect 86374 38644 86398 38646
rect 86454 38644 86478 38646
rect 86238 38624 86534 38644
rect 86394 38460 86446 38466
rect 86394 38402 86446 38408
rect 86406 38058 86434 38402
rect 86394 38052 86446 38058
rect 86394 37994 86446 38000
rect 86578 37780 86630 37786
rect 86578 37722 86630 37728
rect 86238 37612 86534 37632
rect 86294 37610 86318 37612
rect 86374 37610 86398 37612
rect 86454 37610 86478 37612
rect 86316 37558 86318 37610
rect 86380 37558 86392 37610
rect 86454 37558 86456 37610
rect 86294 37556 86318 37558
rect 86374 37556 86398 37558
rect 86454 37556 86478 37558
rect 86238 37536 86534 37556
rect 86590 37394 86618 37722
rect 86406 37366 86618 37394
rect 85934 36760 85986 36766
rect 85934 36702 85986 36708
rect 85946 36630 85974 36702
rect 86406 36698 86434 37366
rect 86578 37168 86630 37174
rect 86578 37110 86630 37116
rect 86590 36834 86618 37110
rect 86578 36828 86630 36834
rect 86578 36770 86630 36776
rect 86026 36692 86078 36698
rect 86026 36634 86078 36640
rect 86394 36692 86446 36698
rect 86394 36634 86446 36640
rect 85934 36624 85986 36630
rect 85934 36566 85986 36572
rect 86038 36290 86066 36634
rect 86238 36524 86534 36544
rect 86294 36522 86318 36524
rect 86374 36522 86398 36524
rect 86454 36522 86478 36524
rect 86316 36470 86318 36522
rect 86380 36470 86392 36522
rect 86454 36470 86456 36522
rect 86294 36468 86318 36470
rect 86374 36468 86398 36470
rect 86454 36468 86478 36470
rect 86238 36448 86534 36468
rect 88246 36426 88274 39558
rect 88430 38602 88458 40034
rect 88522 39690 88550 40510
rect 88902 40332 89198 40352
rect 88958 40330 88982 40332
rect 89038 40330 89062 40332
rect 89118 40330 89142 40332
rect 88980 40278 88982 40330
rect 89044 40278 89056 40330
rect 89118 40278 89120 40330
rect 88958 40276 88982 40278
rect 89038 40276 89062 40278
rect 89118 40276 89142 40278
rect 88902 40256 89198 40276
rect 89350 40098 89378 41598
rect 90994 40568 91046 40574
rect 90994 40510 91046 40516
rect 91006 40438 91034 40510
rect 90166 40432 90218 40438
rect 90166 40374 90218 40380
rect 90534 40432 90586 40438
rect 90534 40374 90586 40380
rect 90994 40432 91046 40438
rect 90994 40374 91046 40380
rect 89338 40092 89390 40098
rect 89338 40034 89390 40040
rect 88786 40024 88838 40030
rect 88786 39966 88838 39972
rect 88694 39956 88746 39962
rect 88694 39898 88746 39904
rect 88510 39684 88562 39690
rect 88510 39626 88562 39632
rect 88706 39554 88734 39898
rect 88694 39548 88746 39554
rect 88694 39490 88746 39496
rect 88602 39480 88654 39486
rect 88602 39422 88654 39428
rect 88418 38596 88470 38602
rect 88418 38538 88470 38544
rect 88430 37514 88458 38538
rect 88614 37922 88642 39422
rect 88694 38392 88746 38398
rect 88694 38334 88746 38340
rect 88602 37916 88654 37922
rect 88602 37858 88654 37864
rect 88510 37848 88562 37854
rect 88510 37790 88562 37796
rect 88418 37508 88470 37514
rect 88418 37450 88470 37456
rect 88326 37304 88378 37310
rect 88326 37246 88378 37252
rect 88338 36970 88366 37246
rect 88326 36964 88378 36970
rect 88326 36906 88378 36912
rect 88234 36420 88286 36426
rect 88234 36362 88286 36368
rect 86026 36284 86078 36290
rect 86026 36226 86078 36232
rect 85842 35876 85894 35882
rect 85842 35818 85894 35824
rect 86038 35678 86066 36226
rect 88246 35746 88274 36362
rect 86578 35740 86630 35746
rect 86578 35682 86630 35688
rect 88234 35740 88286 35746
rect 88234 35682 88286 35688
rect 85658 35672 85710 35678
rect 85658 35614 85710 35620
rect 86026 35672 86078 35678
rect 86026 35614 86078 35620
rect 85670 33706 85698 35614
rect 86590 35610 86618 35682
rect 88338 35678 88366 36906
rect 88522 36902 88550 37790
rect 88510 36896 88562 36902
rect 88510 36838 88562 36844
rect 88706 36290 88734 38334
rect 88798 36970 88826 39966
rect 90178 39622 90206 40374
rect 90546 40166 90574 40374
rect 90534 40160 90586 40166
rect 90534 40102 90586 40108
rect 90166 39616 90218 39622
rect 90166 39558 90218 39564
rect 88902 39244 89198 39264
rect 88958 39242 88982 39244
rect 89038 39242 89062 39244
rect 89118 39242 89142 39244
rect 88980 39190 88982 39242
rect 89044 39190 89056 39242
rect 89118 39190 89120 39242
rect 88958 39188 88982 39190
rect 89038 39188 89062 39190
rect 89118 39188 89142 39190
rect 88902 39168 89198 39188
rect 90178 39146 90206 39558
rect 90166 39140 90218 39146
rect 90166 39082 90218 39088
rect 90178 39010 90206 39082
rect 90166 39004 90218 39010
rect 90166 38946 90218 38952
rect 89890 38460 89942 38466
rect 89890 38402 89942 38408
rect 88902 38156 89198 38176
rect 88958 38154 88982 38156
rect 89038 38154 89062 38156
rect 89118 38154 89142 38156
rect 88980 38102 88982 38154
rect 89044 38102 89056 38154
rect 89118 38102 89120 38154
rect 88958 38100 88982 38102
rect 89038 38100 89062 38102
rect 89118 38100 89142 38102
rect 88902 38080 89198 38100
rect 89522 37916 89574 37922
rect 89522 37858 89574 37864
rect 89246 37780 89298 37786
rect 89246 37722 89298 37728
rect 88902 37068 89198 37088
rect 88958 37066 88982 37068
rect 89038 37066 89062 37068
rect 89118 37066 89142 37068
rect 88980 37014 88982 37066
rect 89044 37014 89056 37066
rect 89118 37014 89120 37066
rect 88958 37012 88982 37014
rect 89038 37012 89062 37014
rect 89118 37012 89142 37014
rect 88902 36992 89198 37012
rect 88786 36964 88838 36970
rect 88786 36906 88838 36912
rect 89258 36766 89286 37722
rect 89534 37378 89562 37858
rect 89902 37854 89930 38402
rect 90178 38058 90206 38946
rect 90718 38936 90770 38942
rect 90718 38878 90770 38884
rect 90730 38602 90758 38878
rect 90718 38596 90770 38602
rect 90718 38538 90770 38544
rect 90166 38052 90218 38058
rect 90166 37994 90218 38000
rect 89890 37848 89942 37854
rect 89890 37790 89942 37796
rect 90350 37848 90402 37854
rect 90350 37790 90402 37796
rect 90718 37848 90770 37854
rect 90718 37790 90770 37796
rect 89522 37372 89574 37378
rect 89522 37314 89574 37320
rect 89534 37242 89562 37314
rect 89522 37236 89574 37242
rect 89522 37178 89574 37184
rect 90258 37236 90310 37242
rect 90258 37178 90310 37184
rect 88786 36760 88838 36766
rect 88786 36702 88838 36708
rect 89246 36760 89298 36766
rect 89246 36702 89298 36708
rect 89522 36760 89574 36766
rect 89522 36702 89574 36708
rect 88694 36284 88746 36290
rect 88694 36226 88746 36232
rect 88798 35678 88826 36702
rect 89534 36290 89562 36702
rect 89522 36284 89574 36290
rect 89522 36226 89574 36232
rect 88902 35980 89198 36000
rect 88958 35978 88982 35980
rect 89038 35978 89062 35980
rect 89118 35978 89142 35980
rect 88980 35926 88982 35978
rect 89044 35926 89056 35978
rect 89118 35926 89120 35978
rect 88958 35924 88982 35926
rect 89038 35924 89062 35926
rect 89118 35924 89142 35926
rect 88902 35904 89198 35924
rect 88326 35672 88378 35678
rect 88326 35614 88378 35620
rect 88786 35672 88838 35678
rect 88786 35614 88838 35620
rect 86578 35604 86630 35610
rect 86578 35546 86630 35552
rect 87774 35604 87826 35610
rect 87774 35546 87826 35552
rect 86238 35436 86534 35456
rect 86294 35434 86318 35436
rect 86374 35434 86398 35436
rect 86454 35434 86478 35436
rect 86316 35382 86318 35434
rect 86380 35382 86392 35434
rect 86454 35382 86456 35434
rect 86294 35380 86318 35382
rect 86374 35380 86398 35382
rect 86454 35380 86478 35382
rect 86238 35360 86534 35380
rect 86590 34590 86618 35546
rect 86670 35536 86722 35542
rect 86670 35478 86722 35484
rect 86578 34584 86630 34590
rect 86578 34526 86630 34532
rect 86590 34454 86618 34526
rect 86026 34448 86078 34454
rect 86026 34390 86078 34396
rect 86578 34448 86630 34454
rect 86578 34390 86630 34396
rect 85290 33700 85342 33706
rect 85290 33642 85342 33648
rect 85658 33700 85710 33706
rect 85658 33642 85710 33648
rect 86038 33502 86066 34390
rect 86238 34348 86534 34368
rect 86294 34346 86318 34348
rect 86374 34346 86398 34348
rect 86454 34346 86478 34348
rect 86316 34294 86318 34346
rect 86380 34294 86392 34346
rect 86454 34294 86456 34346
rect 86294 34292 86318 34294
rect 86374 34292 86398 34294
rect 86454 34292 86478 34294
rect 86238 34272 86534 34292
rect 86026 33496 86078 33502
rect 84368 33464 84424 33473
rect 84368 33399 84424 33408
rect 86024 33464 86026 33473
rect 86078 33464 86080 33473
rect 86024 33399 86080 33408
rect 84186 33360 84238 33366
rect 84186 33302 84238 33308
rect 82898 33156 82950 33162
rect 82898 33098 82950 33104
rect 82806 33020 82858 33026
rect 82806 32962 82858 32968
rect 83266 33020 83318 33026
rect 83266 32962 83318 32968
rect 83634 33020 83686 33026
rect 83634 32962 83686 32968
rect 83910 33020 83962 33026
rect 83910 32962 83962 32968
rect 82714 32408 82766 32414
rect 82714 32350 82766 32356
rect 82818 32006 82846 32962
rect 83082 32816 83134 32822
rect 83082 32758 83134 32764
rect 83094 32618 83122 32758
rect 83082 32612 83134 32618
rect 83082 32554 83134 32560
rect 82990 32340 83042 32346
rect 82990 32282 83042 32288
rect 82806 32000 82858 32006
rect 82806 31942 82858 31948
rect 83002 31530 83030 32282
rect 83278 32074 83306 32962
rect 83646 32890 83674 32962
rect 83450 32884 83502 32890
rect 83450 32826 83502 32832
rect 83634 32884 83686 32890
rect 83634 32826 83686 32832
rect 83462 32532 83490 32826
rect 83574 32716 83870 32736
rect 83630 32714 83654 32716
rect 83710 32714 83734 32716
rect 83790 32714 83814 32716
rect 83652 32662 83654 32714
rect 83716 32662 83728 32714
rect 83790 32662 83792 32714
rect 83630 32660 83654 32662
rect 83710 32660 83734 32662
rect 83790 32660 83814 32662
rect 83574 32640 83870 32660
rect 83542 32544 83594 32550
rect 83462 32504 83542 32532
rect 83542 32486 83594 32492
rect 83634 32408 83686 32414
rect 83634 32350 83686 32356
rect 83450 32340 83502 32346
rect 83450 32282 83502 32288
rect 83266 32068 83318 32074
rect 83266 32010 83318 32016
rect 83278 31938 83306 32010
rect 83266 31932 83318 31938
rect 83266 31874 83318 31880
rect 83462 31870 83490 32282
rect 83646 31938 83674 32350
rect 83922 31938 83950 32962
rect 84094 32816 84146 32822
rect 84094 32758 84146 32764
rect 83634 31932 83686 31938
rect 83634 31874 83686 31880
rect 83910 31932 83962 31938
rect 83910 31874 83962 31880
rect 83450 31864 83502 31870
rect 83450 31806 83502 31812
rect 83574 31628 83870 31648
rect 83630 31626 83654 31628
rect 83710 31626 83734 31628
rect 83790 31626 83814 31628
rect 83652 31574 83654 31626
rect 83716 31574 83728 31626
rect 83790 31574 83792 31626
rect 83630 31572 83654 31574
rect 83710 31572 83734 31574
rect 83790 31572 83814 31574
rect 83574 31552 83870 31572
rect 82990 31524 83042 31530
rect 82990 31466 83042 31472
rect 81518 31320 81570 31326
rect 81518 31262 81570 31268
rect 82622 31320 82674 31326
rect 82622 31262 82674 31268
rect 80598 31252 80650 31258
rect 80598 31194 80650 31200
rect 80322 31184 80374 31190
rect 80322 31126 80374 31132
rect 80506 31184 80558 31190
rect 80506 31126 80558 31132
rect 79678 30980 79730 30986
rect 79678 30922 79730 30928
rect 79494 30096 79546 30102
rect 79494 30038 79546 30044
rect 79126 29892 79178 29898
rect 79126 29834 79178 29840
rect 78942 29756 78994 29762
rect 78942 29698 78994 29704
rect 78954 29218 78982 29698
rect 79138 29694 79166 29834
rect 79126 29688 79178 29694
rect 79126 29630 79178 29636
rect 78942 29212 78994 29218
rect 78942 29154 78994 29160
rect 79138 28198 79166 29630
rect 79506 29014 79534 30038
rect 79690 29830 79718 30922
rect 80334 30889 80362 31126
rect 80320 30880 80376 30889
rect 80320 30815 80376 30824
rect 79770 30164 79822 30170
rect 79770 30106 79822 30112
rect 79678 29824 79730 29830
rect 79678 29766 79730 29772
rect 79494 29008 79546 29014
rect 79494 28950 79546 28956
rect 79506 28674 79534 28950
rect 79218 28668 79270 28674
rect 79218 28610 79270 28616
rect 79494 28668 79546 28674
rect 79494 28610 79546 28616
rect 79126 28192 79178 28198
rect 79126 28134 79178 28140
rect 78666 27580 78718 27586
rect 78586 27540 78666 27568
rect 78666 27522 78718 27528
rect 75630 27512 75682 27518
rect 75630 27454 75682 27460
rect 75538 27444 75590 27450
rect 75538 27386 75590 27392
rect 73790 27376 73842 27382
rect 73790 27318 73842 27324
rect 73882 27376 73934 27382
rect 73882 27318 73934 27324
rect 73894 27058 73922 27318
rect 73618 27042 73922 27058
rect 73606 27036 73922 27042
rect 73658 27030 73922 27036
rect 73606 26978 73658 26984
rect 73894 26974 73922 27030
rect 75550 26974 75578 27386
rect 75642 27110 75670 27454
rect 78246 27276 78542 27296
rect 78302 27274 78326 27276
rect 78382 27274 78406 27276
rect 78462 27274 78486 27276
rect 78324 27222 78326 27274
rect 78388 27222 78400 27274
rect 78462 27222 78464 27274
rect 78302 27220 78326 27222
rect 78382 27220 78406 27222
rect 78462 27220 78486 27222
rect 78246 27200 78542 27220
rect 75630 27104 75682 27110
rect 75630 27046 75682 27052
rect 73330 26968 73382 26974
rect 73330 26910 73382 26916
rect 73882 26968 73934 26974
rect 73882 26910 73934 26916
rect 75538 26968 75590 26974
rect 75538 26910 75590 26916
rect 78678 26906 78706 27522
rect 79034 27376 79086 27382
rect 79034 27318 79086 27324
rect 79046 26974 79074 27318
rect 79230 27110 79258 28610
rect 79782 28130 79810 30106
rect 80322 29824 80374 29830
rect 80322 29766 80374 29772
rect 79862 29144 79914 29150
rect 79862 29086 79914 29092
rect 79770 28124 79822 28130
rect 79770 28066 79822 28072
rect 79874 27926 79902 29086
rect 80334 29082 80362 29766
rect 80138 29076 80190 29082
rect 80138 29018 80190 29024
rect 80322 29076 80374 29082
rect 80322 29018 80374 29024
rect 80150 28962 80178 29018
rect 80150 28934 80270 28962
rect 80138 27988 80190 27994
rect 80138 27930 80190 27936
rect 79862 27920 79914 27926
rect 79862 27862 79914 27868
rect 79874 27568 79902 27862
rect 80150 27722 80178 27930
rect 80138 27716 80190 27722
rect 80138 27658 80190 27664
rect 79954 27580 80006 27586
rect 79782 27540 79954 27568
rect 79782 27450 79810 27540
rect 79954 27522 80006 27528
rect 80242 27518 80270 28934
rect 80334 27586 80362 29018
rect 80414 28600 80466 28606
rect 80414 28542 80466 28548
rect 80426 28266 80454 28542
rect 80414 28260 80466 28266
rect 80414 28202 80466 28208
rect 80322 27580 80374 27586
rect 80322 27522 80374 27528
rect 80230 27512 80282 27518
rect 80230 27454 80282 27460
rect 80518 27450 80546 31126
rect 80610 30714 80638 31194
rect 80782 31184 80834 31190
rect 80782 31126 80834 31132
rect 80794 30850 80822 31126
rect 80910 31084 81206 31104
rect 80966 31082 80990 31084
rect 81046 31082 81070 31084
rect 81126 31082 81150 31084
rect 80988 31030 80990 31082
rect 81052 31030 81064 31082
rect 81126 31030 81128 31082
rect 80966 31028 80990 31030
rect 81046 31028 81070 31030
rect 81126 31028 81150 31030
rect 80910 31008 81206 31028
rect 80964 30880 81020 30889
rect 80782 30844 80834 30850
rect 81530 30850 81558 31262
rect 80964 30815 80966 30824
rect 80782 30786 80834 30792
rect 81018 30815 81020 30824
rect 81518 30844 81570 30850
rect 80966 30786 81018 30792
rect 81518 30786 81570 30792
rect 82070 30844 82122 30850
rect 82070 30786 82122 30792
rect 81058 30776 81110 30782
rect 81058 30718 81110 30724
rect 80598 30708 80650 30714
rect 80598 30650 80650 30656
rect 81070 30238 81098 30718
rect 82082 30442 82110 30786
rect 83574 30540 83870 30560
rect 83630 30538 83654 30540
rect 83710 30538 83734 30540
rect 83790 30538 83814 30540
rect 83652 30486 83654 30538
rect 83716 30486 83728 30538
rect 83790 30486 83792 30538
rect 83630 30484 83654 30486
rect 83710 30484 83734 30486
rect 83790 30484 83814 30486
rect 83574 30464 83870 30484
rect 82070 30436 82122 30442
rect 82070 30378 82122 30384
rect 81058 30232 81110 30238
rect 81058 30174 81110 30180
rect 80910 29996 81206 30016
rect 80966 29994 80990 29996
rect 81046 29994 81070 29996
rect 81126 29994 81150 29996
rect 80988 29942 80990 29994
rect 81052 29942 81064 29994
rect 81126 29942 81128 29994
rect 80966 29940 80990 29942
rect 81046 29940 81070 29942
rect 81126 29940 81150 29942
rect 80910 29920 81206 29940
rect 84106 29898 84134 32758
rect 84094 29892 84146 29898
rect 84094 29834 84146 29840
rect 84198 29762 84226 33302
rect 86238 33260 86534 33280
rect 86294 33258 86318 33260
rect 86374 33258 86398 33260
rect 86454 33258 86478 33260
rect 86316 33206 86318 33258
rect 86380 33206 86392 33258
rect 86454 33206 86456 33258
rect 86294 33204 86318 33206
rect 86374 33204 86398 33206
rect 86454 33204 86478 33206
rect 86238 33184 86534 33204
rect 86118 32884 86170 32890
rect 86118 32826 86170 32832
rect 84278 32816 84330 32822
rect 84278 32758 84330 32764
rect 84290 32618 84318 32758
rect 84278 32612 84330 32618
rect 84278 32554 84330 32560
rect 86130 32414 86158 32826
rect 86590 32550 86618 34390
rect 86682 33434 86710 35478
rect 87786 34590 87814 35546
rect 88798 34794 88826 35614
rect 89982 35604 90034 35610
rect 89982 35546 90034 35552
rect 89522 35536 89574 35542
rect 89522 35478 89574 35484
rect 89534 35338 89562 35478
rect 89522 35332 89574 35338
rect 89522 35274 89574 35280
rect 89994 35202 90022 35546
rect 89982 35196 90034 35202
rect 89982 35138 90034 35144
rect 88902 34892 89198 34912
rect 88958 34890 88982 34892
rect 89038 34890 89062 34892
rect 89118 34890 89142 34892
rect 88980 34838 88982 34890
rect 89044 34838 89056 34890
rect 89118 34838 89120 34890
rect 88958 34836 88982 34838
rect 89038 34836 89062 34838
rect 89118 34836 89142 34838
rect 88902 34816 89198 34836
rect 88786 34788 88838 34794
rect 88786 34730 88838 34736
rect 87774 34584 87826 34590
rect 87774 34526 87826 34532
rect 87958 34516 88010 34522
rect 87958 34458 88010 34464
rect 86670 33428 86722 33434
rect 86670 33370 86722 33376
rect 86682 32822 86710 33370
rect 87590 33360 87642 33366
rect 87590 33302 87642 33308
rect 87498 33020 87550 33026
rect 87498 32962 87550 32968
rect 87406 32952 87458 32958
rect 87406 32894 87458 32900
rect 87418 32822 87446 32894
rect 86670 32816 86722 32822
rect 86670 32758 86722 32764
rect 87406 32816 87458 32822
rect 87406 32758 87458 32764
rect 86578 32544 86630 32550
rect 86578 32486 86630 32492
rect 86118 32408 86170 32414
rect 86682 32362 86710 32758
rect 87418 32414 87446 32758
rect 86118 32350 86170 32356
rect 86590 32334 86710 32362
rect 87406 32408 87458 32414
rect 87406 32350 87458 32356
rect 86238 32172 86534 32192
rect 86294 32170 86318 32172
rect 86374 32170 86398 32172
rect 86454 32170 86478 32172
rect 86316 32118 86318 32170
rect 86380 32118 86392 32170
rect 86454 32118 86456 32170
rect 86294 32116 86318 32118
rect 86374 32116 86398 32118
rect 86454 32116 86478 32118
rect 86238 32096 86534 32116
rect 84830 32068 84882 32074
rect 84830 32010 84882 32016
rect 84370 31796 84422 31802
rect 84370 31738 84422 31744
rect 84278 31728 84330 31734
rect 84278 31670 84330 31676
rect 84290 31462 84318 31670
rect 84382 31462 84410 31738
rect 84278 31456 84330 31462
rect 84278 31398 84330 31404
rect 84370 31456 84422 31462
rect 84370 31398 84422 31404
rect 84842 30986 84870 32010
rect 86238 31084 86534 31104
rect 86294 31082 86318 31084
rect 86374 31082 86398 31084
rect 86454 31082 86478 31084
rect 86316 31030 86318 31082
rect 86380 31030 86392 31082
rect 86454 31030 86456 31082
rect 86294 31028 86318 31030
rect 86374 31028 86398 31030
rect 86454 31028 86478 31030
rect 86238 31008 86534 31028
rect 84830 30980 84882 30986
rect 84830 30922 84882 30928
rect 86118 30640 86170 30646
rect 86118 30582 86170 30588
rect 86026 30232 86078 30238
rect 86026 30174 86078 30180
rect 85198 30096 85250 30102
rect 85198 30038 85250 30044
rect 84554 29892 84606 29898
rect 84554 29834 84606 29840
rect 84186 29756 84238 29762
rect 84186 29698 84238 29704
rect 80598 29688 80650 29694
rect 80598 29630 80650 29636
rect 80610 27722 80638 29630
rect 83174 29620 83226 29626
rect 83174 29562 83226 29568
rect 81242 29144 81294 29150
rect 81242 29086 81294 29092
rect 80910 28908 81206 28928
rect 80966 28906 80990 28908
rect 81046 28906 81070 28908
rect 81126 28906 81150 28908
rect 80988 28854 80990 28906
rect 81052 28854 81064 28906
rect 81126 28854 81128 28906
rect 80966 28852 80990 28854
rect 81046 28852 81070 28854
rect 81126 28852 81150 28854
rect 80910 28832 81206 28852
rect 81254 28810 81282 29086
rect 81426 29076 81478 29082
rect 81426 29018 81478 29024
rect 81334 29008 81386 29014
rect 81334 28950 81386 28956
rect 81242 28804 81294 28810
rect 81242 28746 81294 28752
rect 81242 28192 81294 28198
rect 81242 28134 81294 28140
rect 81254 27994 81282 28134
rect 81346 28062 81374 28950
rect 81334 28056 81386 28062
rect 81334 27998 81386 28004
rect 81242 27988 81294 27994
rect 81242 27930 81294 27936
rect 80910 27820 81206 27840
rect 80966 27818 80990 27820
rect 81046 27818 81070 27820
rect 81126 27818 81150 27820
rect 80988 27766 80990 27818
rect 81052 27766 81064 27818
rect 81126 27766 81128 27818
rect 80966 27764 80990 27766
rect 81046 27764 81070 27766
rect 81126 27764 81150 27766
rect 80910 27744 81206 27764
rect 80598 27716 80650 27722
rect 80598 27658 80650 27664
rect 81438 27654 81466 29018
rect 83186 28198 83214 29562
rect 83574 29452 83870 29472
rect 83630 29450 83654 29452
rect 83710 29450 83734 29452
rect 83790 29450 83814 29452
rect 83652 29398 83654 29450
rect 83716 29398 83728 29450
rect 83790 29398 83792 29450
rect 83630 29396 83654 29398
rect 83710 29396 83734 29398
rect 83790 29396 83814 29398
rect 83574 29376 83870 29396
rect 84094 29076 84146 29082
rect 84094 29018 84146 29024
rect 83574 28364 83870 28384
rect 83630 28362 83654 28364
rect 83710 28362 83734 28364
rect 83790 28362 83814 28364
rect 83652 28310 83654 28362
rect 83716 28310 83728 28362
rect 83790 28310 83792 28362
rect 83630 28308 83654 28310
rect 83710 28308 83734 28310
rect 83790 28308 83814 28310
rect 83574 28288 83870 28308
rect 83174 28192 83226 28198
rect 83174 28134 83226 28140
rect 83266 27988 83318 27994
rect 83266 27930 83318 27936
rect 81426 27648 81478 27654
rect 81426 27590 81478 27596
rect 83278 27586 83306 27930
rect 83266 27580 83318 27586
rect 83266 27522 83318 27528
rect 84106 27518 84134 29018
rect 84198 28810 84226 29698
rect 84566 29082 84594 29834
rect 84922 29280 84974 29286
rect 84922 29222 84974 29228
rect 84830 29144 84882 29150
rect 84830 29086 84882 29092
rect 84554 29076 84606 29082
rect 84554 29018 84606 29024
rect 84186 28804 84238 28810
rect 84186 28746 84238 28752
rect 84554 28600 84606 28606
rect 84554 28542 84606 28548
rect 84566 28130 84594 28542
rect 84554 28124 84606 28130
rect 84554 28066 84606 28072
rect 84842 27654 84870 29086
rect 84934 28062 84962 29222
rect 85210 28470 85238 30038
rect 86038 29694 86066 30174
rect 86130 29762 86158 30582
rect 86238 29996 86534 30016
rect 86294 29994 86318 29996
rect 86374 29994 86398 29996
rect 86454 29994 86478 29996
rect 86316 29942 86318 29994
rect 86380 29942 86392 29994
rect 86454 29942 86456 29994
rect 86294 29940 86318 29942
rect 86374 29940 86398 29942
rect 86454 29940 86478 29942
rect 86238 29920 86534 29940
rect 86118 29756 86170 29762
rect 86118 29698 86170 29704
rect 85842 29688 85894 29694
rect 85842 29630 85894 29636
rect 86026 29688 86078 29694
rect 86026 29630 86078 29636
rect 85854 29286 85882 29630
rect 86394 29348 86446 29354
rect 86394 29290 86446 29296
rect 85842 29280 85894 29286
rect 85842 29222 85894 29228
rect 86406 29234 86434 29290
rect 86590 29234 86618 32334
rect 87418 32074 87446 32350
rect 87510 32278 87538 32962
rect 87602 32414 87630 33302
rect 87970 33026 87998 34458
rect 90270 34182 90298 37178
rect 90258 34176 90310 34182
rect 90258 34118 90310 34124
rect 89798 34108 89850 34114
rect 89798 34050 89850 34056
rect 88418 34040 88470 34046
rect 88418 33982 88470 33988
rect 87958 33020 88010 33026
rect 87958 32962 88010 32968
rect 87590 32408 87642 32414
rect 87590 32350 87642 32356
rect 87498 32272 87550 32278
rect 87498 32214 87550 32220
rect 87406 32068 87458 32074
rect 87406 32010 87458 32016
rect 88326 31728 88378 31734
rect 88326 31670 88378 31676
rect 88338 31530 88366 31670
rect 88430 31530 88458 33982
rect 88902 33804 89198 33824
rect 88958 33802 88982 33804
rect 89038 33802 89062 33804
rect 89118 33802 89142 33804
rect 88980 33750 88982 33802
rect 89044 33750 89056 33802
rect 89118 33750 89120 33802
rect 88958 33748 88982 33750
rect 89038 33748 89062 33750
rect 89118 33748 89142 33750
rect 88902 33728 89198 33748
rect 89810 33502 89838 34050
rect 90270 34046 90298 34118
rect 90258 34040 90310 34046
rect 90258 33982 90310 33988
rect 90362 33570 90390 37790
rect 90730 37514 90758 37790
rect 90718 37508 90770 37514
rect 90718 37450 90770 37456
rect 90442 36148 90494 36154
rect 90442 36090 90494 36096
rect 90350 33564 90402 33570
rect 90350 33506 90402 33512
rect 89798 33496 89850 33502
rect 89798 33438 89850 33444
rect 88902 32716 89198 32736
rect 88958 32714 88982 32716
rect 89038 32714 89062 32716
rect 89118 32714 89142 32716
rect 88980 32662 88982 32714
rect 89044 32662 89056 32714
rect 89118 32662 89120 32714
rect 88958 32660 88982 32662
rect 89038 32660 89062 32662
rect 89118 32660 89142 32662
rect 88902 32640 89198 32660
rect 89062 32476 89114 32482
rect 89062 32418 89114 32424
rect 89074 32074 89102 32418
rect 89062 32068 89114 32074
rect 89062 32010 89114 32016
rect 89706 31864 89758 31870
rect 89706 31806 89758 31812
rect 88902 31628 89198 31648
rect 88958 31626 88982 31628
rect 89038 31626 89062 31628
rect 89118 31626 89142 31628
rect 88980 31574 88982 31626
rect 89044 31574 89056 31626
rect 89118 31574 89120 31626
rect 88958 31572 88982 31574
rect 89038 31572 89062 31574
rect 89118 31572 89142 31574
rect 88902 31552 89198 31572
rect 88326 31524 88378 31530
rect 88326 31466 88378 31472
rect 88418 31524 88470 31530
rect 88418 31466 88470 31472
rect 88338 31326 88366 31466
rect 88326 31320 88378 31326
rect 88326 31262 88378 31268
rect 87682 30980 87734 30986
rect 87682 30922 87734 30928
rect 86762 30776 86814 30782
rect 86762 30718 86814 30724
rect 86774 30442 86802 30718
rect 86762 30436 86814 30442
rect 86762 30378 86814 30384
rect 86670 29824 86722 29830
rect 86670 29766 86722 29772
rect 86682 29354 86710 29766
rect 86774 29354 86802 30378
rect 87590 30096 87642 30102
rect 87590 30038 87642 30044
rect 86670 29348 86722 29354
rect 86670 29290 86722 29296
rect 86762 29348 86814 29354
rect 86762 29290 86814 29296
rect 86406 29206 86618 29234
rect 86774 29150 86802 29290
rect 86762 29144 86814 29150
rect 86762 29086 86814 29092
rect 86238 28908 86534 28928
rect 86294 28906 86318 28908
rect 86374 28906 86398 28908
rect 86454 28906 86478 28908
rect 86316 28854 86318 28906
rect 86380 28854 86392 28906
rect 86454 28854 86456 28906
rect 86294 28852 86318 28854
rect 86374 28852 86398 28854
rect 86454 28852 86478 28854
rect 86238 28832 86534 28852
rect 85198 28464 85250 28470
rect 85198 28406 85250 28412
rect 85566 28464 85618 28470
rect 85566 28406 85618 28412
rect 84922 28056 84974 28062
rect 84922 27998 84974 28004
rect 85014 28056 85066 28062
rect 85014 27998 85066 28004
rect 84830 27648 84882 27654
rect 84830 27590 84882 27596
rect 84094 27512 84146 27518
rect 84094 27454 84146 27460
rect 79770 27444 79822 27450
rect 79770 27386 79822 27392
rect 80506 27444 80558 27450
rect 80506 27386 80558 27392
rect 79218 27104 79270 27110
rect 79218 27046 79270 27052
rect 79230 26974 79258 27046
rect 79034 26968 79086 26974
rect 79034 26910 79086 26916
rect 79218 26968 79270 26974
rect 79218 26910 79270 26916
rect 80518 26906 80546 27386
rect 83574 27276 83870 27296
rect 83630 27274 83654 27276
rect 83710 27274 83734 27276
rect 83790 27274 83814 27276
rect 83652 27222 83654 27274
rect 83716 27222 83728 27274
rect 83790 27222 83792 27274
rect 83630 27220 83654 27222
rect 83710 27220 83734 27222
rect 83790 27220 83814 27222
rect 83574 27200 83870 27220
rect 84106 26974 84134 27454
rect 84094 26968 84146 26974
rect 84094 26910 84146 26916
rect 84842 26906 84870 27590
rect 85026 27450 85054 27998
rect 85014 27444 85066 27450
rect 85014 27386 85066 27392
rect 85578 26974 85606 28406
rect 87602 28130 87630 30038
rect 87694 29762 87722 30922
rect 88430 30850 88458 31466
rect 89338 31456 89390 31462
rect 89338 31398 89390 31404
rect 89246 30912 89298 30918
rect 89246 30854 89298 30860
rect 88418 30844 88470 30850
rect 88418 30786 88470 30792
rect 88786 30844 88838 30850
rect 88786 30786 88838 30792
rect 88798 30238 88826 30786
rect 88902 30540 89198 30560
rect 88958 30538 88982 30540
rect 89038 30538 89062 30540
rect 89118 30538 89142 30540
rect 88980 30486 88982 30538
rect 89044 30486 89056 30538
rect 89118 30486 89120 30538
rect 88958 30484 88982 30486
rect 89038 30484 89062 30486
rect 89118 30484 89142 30486
rect 88902 30464 89198 30484
rect 89258 30238 89286 30854
rect 88510 30232 88562 30238
rect 88510 30174 88562 30180
rect 88786 30232 88838 30238
rect 88786 30174 88838 30180
rect 89246 30232 89298 30238
rect 89246 30174 89298 30180
rect 88522 29898 88550 30174
rect 87774 29892 87826 29898
rect 87774 29834 87826 29840
rect 88510 29892 88562 29898
rect 88510 29834 88562 29840
rect 87682 29756 87734 29762
rect 87682 29698 87734 29704
rect 87786 29082 87814 29834
rect 88902 29452 89198 29472
rect 88958 29450 88982 29452
rect 89038 29450 89062 29452
rect 89118 29450 89142 29452
rect 88980 29398 88982 29450
rect 89044 29398 89056 29450
rect 89118 29398 89120 29450
rect 88958 29396 88982 29398
rect 89038 29396 89062 29398
rect 89118 29396 89142 29398
rect 88902 29376 89198 29396
rect 87774 29076 87826 29082
rect 87774 29018 87826 29024
rect 89258 28810 89286 30174
rect 89246 28804 89298 28810
rect 89246 28746 89298 28752
rect 88902 28364 89198 28384
rect 88958 28362 88982 28364
rect 89038 28362 89062 28364
rect 89118 28362 89142 28364
rect 88980 28310 88982 28362
rect 89044 28310 89056 28362
rect 89118 28310 89120 28362
rect 88958 28308 88982 28310
rect 89038 28308 89062 28310
rect 89118 28308 89142 28310
rect 88902 28288 89198 28308
rect 87590 28124 87642 28130
rect 87590 28066 87642 28072
rect 85750 28056 85802 28062
rect 85750 27998 85802 28004
rect 86118 28056 86170 28062
rect 86118 27998 86170 28004
rect 85762 27518 85790 27998
rect 86130 27586 86158 27998
rect 86578 27988 86630 27994
rect 86578 27930 86630 27936
rect 86238 27820 86534 27840
rect 86294 27818 86318 27820
rect 86374 27818 86398 27820
rect 86454 27818 86478 27820
rect 86316 27766 86318 27818
rect 86380 27766 86392 27818
rect 86454 27766 86456 27818
rect 86294 27764 86318 27766
rect 86374 27764 86398 27766
rect 86454 27764 86478 27766
rect 86238 27744 86534 27764
rect 86118 27580 86170 27586
rect 86118 27522 86170 27528
rect 85750 27512 85802 27518
rect 85750 27454 85802 27460
rect 85762 27042 85790 27454
rect 86590 27042 86618 27930
rect 87602 27382 87630 28066
rect 89350 28062 89378 31398
rect 89718 30986 89746 31806
rect 89706 30980 89758 30986
rect 89706 30922 89758 30928
rect 89614 30844 89666 30850
rect 89614 30786 89666 30792
rect 89626 30442 89654 30786
rect 89614 30436 89666 30442
rect 89614 30378 89666 30384
rect 89338 28056 89390 28062
rect 89338 27998 89390 28004
rect 89614 28056 89666 28062
rect 89614 27998 89666 28004
rect 89246 27988 89298 27994
rect 89246 27930 89298 27936
rect 89258 27586 89286 27930
rect 87682 27580 87734 27586
rect 87682 27522 87734 27528
rect 89246 27580 89298 27586
rect 89246 27522 89298 27528
rect 87590 27376 87642 27382
rect 87590 27318 87642 27324
rect 87694 27110 87722 27522
rect 89338 27376 89390 27382
rect 89338 27318 89390 27324
rect 88902 27276 89198 27296
rect 88958 27274 88982 27276
rect 89038 27274 89062 27276
rect 89118 27274 89142 27276
rect 88980 27222 88982 27274
rect 89044 27222 89056 27274
rect 89118 27222 89120 27274
rect 88958 27220 88982 27222
rect 89038 27220 89062 27222
rect 89118 27220 89142 27222
rect 88902 27200 89198 27220
rect 87682 27104 87734 27110
rect 87682 27046 87734 27052
rect 89350 27042 89378 27318
rect 85750 27036 85802 27042
rect 85750 26978 85802 26984
rect 86578 27036 86630 27042
rect 86578 26978 86630 26984
rect 89338 27036 89390 27042
rect 89338 26978 89390 26984
rect 85566 26968 85618 26974
rect 85566 26910 85618 26916
rect 89626 26906 89654 27998
rect 89810 27654 89838 33438
rect 90454 31938 90482 36090
rect 90718 36080 90770 36086
rect 90718 36022 90770 36028
rect 90730 35746 90758 36022
rect 90718 35740 90770 35746
rect 90718 35682 90770 35688
rect 91282 35241 91310 42126
rect 91566 41964 91862 41984
rect 91622 41962 91646 41964
rect 91702 41962 91726 41964
rect 91782 41962 91806 41964
rect 91644 41910 91646 41962
rect 91708 41910 91720 41962
rect 91782 41910 91784 41962
rect 91622 41908 91646 41910
rect 91702 41908 91726 41910
rect 91782 41908 91806 41910
rect 91566 41888 91862 41908
rect 91566 40876 91862 40896
rect 91622 40874 91646 40876
rect 91702 40874 91726 40876
rect 91782 40874 91806 40876
rect 91644 40822 91646 40874
rect 91708 40822 91720 40874
rect 91782 40822 91784 40874
rect 91622 40820 91646 40822
rect 91702 40820 91726 40822
rect 91782 40820 91806 40822
rect 91566 40800 91862 40820
rect 92846 40438 92874 43312
rect 94042 43242 94070 43312
rect 93306 43214 94070 43242
rect 92834 40432 92886 40438
rect 92834 40374 92886 40380
rect 91566 39788 91862 39808
rect 91622 39786 91646 39788
rect 91702 39786 91726 39788
rect 91782 39786 91806 39788
rect 91644 39734 91646 39786
rect 91708 39734 91720 39786
rect 91782 39734 91784 39786
rect 91622 39732 91646 39734
rect 91702 39732 91726 39734
rect 91782 39732 91806 39734
rect 91566 39712 91862 39732
rect 91454 38800 91506 38806
rect 91454 38742 91506 38748
rect 91466 38466 91494 38742
rect 91566 38700 91862 38720
rect 91622 38698 91646 38700
rect 91702 38698 91726 38700
rect 91782 38698 91806 38700
rect 91644 38646 91646 38698
rect 91708 38646 91720 38698
rect 91782 38646 91784 38698
rect 91622 38644 91646 38646
rect 91702 38644 91726 38646
rect 91782 38644 91806 38646
rect 91566 38624 91862 38644
rect 91454 38460 91506 38466
rect 91454 38402 91506 38408
rect 91362 37712 91414 37718
rect 91362 37654 91414 37660
rect 91374 37378 91402 37654
rect 91566 37612 91862 37632
rect 91622 37610 91646 37612
rect 91702 37610 91726 37612
rect 91782 37610 91806 37612
rect 91644 37558 91646 37610
rect 91708 37558 91720 37610
rect 91782 37558 91784 37610
rect 91622 37556 91646 37558
rect 91702 37556 91726 37558
rect 91782 37556 91806 37558
rect 91566 37536 91862 37556
rect 91362 37372 91414 37378
rect 91362 37314 91414 37320
rect 91566 36524 91862 36544
rect 91622 36522 91646 36524
rect 91702 36522 91726 36524
rect 91782 36522 91806 36524
rect 91644 36470 91646 36522
rect 91708 36470 91720 36522
rect 91782 36470 91784 36522
rect 91622 36468 91646 36470
rect 91702 36468 91726 36470
rect 91782 36468 91806 36470
rect 91566 36448 91862 36468
rect 91362 36284 91414 36290
rect 91362 36226 91414 36232
rect 91374 35882 91402 36226
rect 91362 35876 91414 35882
rect 91362 35818 91414 35824
rect 91566 35436 91862 35456
rect 91622 35434 91646 35436
rect 91702 35434 91726 35436
rect 91782 35434 91806 35436
rect 91644 35382 91646 35434
rect 91708 35382 91720 35434
rect 91782 35382 91784 35434
rect 91622 35380 91646 35382
rect 91702 35380 91726 35382
rect 91782 35380 91806 35382
rect 91566 35360 91862 35380
rect 91268 35232 91324 35241
rect 91268 35167 91324 35176
rect 90626 34992 90678 34998
rect 90626 34934 90678 34940
rect 91086 34992 91138 34998
rect 91086 34934 91138 34940
rect 90638 33638 90666 34934
rect 90718 34788 90770 34794
rect 90718 34730 90770 34736
rect 90626 33632 90678 33638
rect 90626 33574 90678 33580
rect 90442 31932 90494 31938
rect 90442 31874 90494 31880
rect 90730 31394 90758 34730
rect 91098 34590 91126 34934
rect 91086 34584 91138 34590
rect 91086 34526 91138 34532
rect 91566 34348 91862 34368
rect 91622 34346 91646 34348
rect 91702 34346 91726 34348
rect 91782 34346 91806 34348
rect 91644 34294 91646 34346
rect 91708 34294 91720 34346
rect 91782 34294 91784 34346
rect 91622 34292 91646 34294
rect 91702 34292 91726 34294
rect 91782 34292 91806 34294
rect 91566 34272 91862 34292
rect 91362 33972 91414 33978
rect 91362 33914 91414 33920
rect 91374 33609 91402 33914
rect 91360 33600 91416 33609
rect 91360 33535 91416 33544
rect 91566 33260 91862 33280
rect 91622 33258 91646 33260
rect 91702 33258 91726 33260
rect 91782 33258 91806 33260
rect 91644 33206 91646 33258
rect 91708 33206 91720 33258
rect 91782 33206 91784 33258
rect 91622 33204 91646 33206
rect 91702 33204 91726 33206
rect 91782 33204 91806 33206
rect 91566 33184 91862 33204
rect 91084 32648 91140 32657
rect 91084 32583 91140 32592
rect 90718 31388 90770 31394
rect 90718 31330 90770 31336
rect 90902 31320 90954 31326
rect 90902 31262 90954 31268
rect 90914 30850 90942 31262
rect 90902 30844 90954 30850
rect 90902 30786 90954 30792
rect 90442 30232 90494 30238
rect 90442 30174 90494 30180
rect 90994 30232 91046 30238
rect 90994 30174 91046 30180
rect 90074 28668 90126 28674
rect 90074 28610 90126 28616
rect 90350 28668 90402 28674
rect 90350 28610 90402 28616
rect 90086 28198 90114 28610
rect 90362 28266 90390 28610
rect 90350 28260 90402 28266
rect 90350 28202 90402 28208
rect 90074 28192 90126 28198
rect 90074 28134 90126 28140
rect 90086 27722 90114 28134
rect 90362 28130 90390 28202
rect 90350 28124 90402 28130
rect 90350 28066 90402 28072
rect 90074 27716 90126 27722
rect 90074 27658 90126 27664
rect 89798 27648 89850 27654
rect 89798 27590 89850 27596
rect 90362 27586 90390 28066
rect 90350 27580 90402 27586
rect 90350 27522 90402 27528
rect 90454 26974 90482 30174
rect 90534 29756 90586 29762
rect 90534 29698 90586 29704
rect 90626 29756 90678 29762
rect 90626 29698 90678 29704
rect 90546 27722 90574 29698
rect 90638 29014 90666 29698
rect 90810 29552 90862 29558
rect 90810 29494 90862 29500
rect 90822 29150 90850 29494
rect 91006 29354 91034 30174
rect 90994 29348 91046 29354
rect 90994 29290 91046 29296
rect 91098 29218 91126 32583
rect 91566 32172 91862 32192
rect 91622 32170 91646 32172
rect 91702 32170 91726 32172
rect 91782 32170 91806 32172
rect 91644 32118 91646 32170
rect 91708 32118 91720 32170
rect 91782 32118 91784 32170
rect 91622 32116 91646 32118
rect 91702 32116 91726 32118
rect 91782 32116 91806 32118
rect 91566 32096 91862 32116
rect 91362 31932 91414 31938
rect 91546 31932 91598 31938
rect 91414 31892 91546 31920
rect 91362 31874 91414 31880
rect 91466 31326 91494 31892
rect 91546 31874 91598 31880
rect 91454 31320 91506 31326
rect 91454 31262 91506 31268
rect 91362 30844 91414 30850
rect 91362 30786 91414 30792
rect 91374 30442 91402 30786
rect 91466 30646 91494 31262
rect 91566 31084 91862 31104
rect 91622 31082 91646 31084
rect 91702 31082 91726 31084
rect 91782 31082 91806 31084
rect 91644 31030 91646 31082
rect 91708 31030 91720 31082
rect 91782 31030 91784 31082
rect 91622 31028 91646 31030
rect 91702 31028 91726 31030
rect 91782 31028 91806 31030
rect 91566 31008 91862 31028
rect 91454 30640 91506 30646
rect 91454 30582 91506 30588
rect 91362 30436 91414 30442
rect 91362 30378 91414 30384
rect 91086 29212 91138 29218
rect 91086 29154 91138 29160
rect 91466 29150 91494 30582
rect 93306 30306 93334 43214
rect 93294 30300 93346 30306
rect 93294 30242 93346 30248
rect 91566 29996 91862 30016
rect 91622 29994 91646 29996
rect 91702 29994 91726 29996
rect 91782 29994 91806 29996
rect 91644 29942 91646 29994
rect 91708 29942 91720 29994
rect 91782 29942 91784 29994
rect 91622 29940 91646 29942
rect 91702 29940 91726 29942
rect 91782 29940 91806 29942
rect 91566 29920 91862 29940
rect 90810 29144 90862 29150
rect 90810 29086 90862 29092
rect 91454 29144 91506 29150
rect 91454 29086 91506 29092
rect 91914 29144 91966 29150
rect 91914 29086 91966 29092
rect 90718 29076 90770 29082
rect 90718 29018 90770 29024
rect 90626 29008 90678 29014
rect 90626 28950 90678 28956
rect 90638 28538 90666 28950
rect 90730 28810 90758 29018
rect 91566 28908 91862 28928
rect 91622 28906 91646 28908
rect 91702 28906 91726 28908
rect 91782 28906 91806 28908
rect 91644 28854 91646 28906
rect 91708 28854 91720 28906
rect 91782 28854 91784 28906
rect 91622 28852 91646 28854
rect 91702 28852 91726 28854
rect 91782 28852 91806 28854
rect 91566 28832 91862 28852
rect 90718 28804 90770 28810
rect 90718 28746 90770 28752
rect 91926 28690 91954 29086
rect 91834 28674 91954 28690
rect 91086 28668 91138 28674
rect 91086 28610 91138 28616
rect 91822 28668 91954 28674
rect 91874 28662 91954 28668
rect 91822 28610 91874 28616
rect 90626 28532 90678 28538
rect 90626 28474 90678 28480
rect 91098 28062 91126 28610
rect 91086 28056 91138 28062
rect 91086 27998 91138 28004
rect 91098 27722 91126 27998
rect 91566 27820 91862 27840
rect 91622 27818 91646 27820
rect 91702 27818 91726 27820
rect 91782 27818 91806 27820
rect 91644 27766 91646 27818
rect 91708 27766 91720 27818
rect 91782 27766 91784 27818
rect 91622 27764 91646 27766
rect 91702 27764 91726 27766
rect 91782 27764 91806 27766
rect 91566 27744 91862 27764
rect 90534 27716 90586 27722
rect 90534 27658 90586 27664
rect 91086 27716 91138 27722
rect 91086 27658 91138 27664
rect 91178 27172 91230 27178
rect 91178 27114 91230 27120
rect 90442 26968 90494 26974
rect 90442 26910 90494 26916
rect 70846 26900 70898 26906
rect 70846 26842 70898 26848
rect 70938 26900 70990 26906
rect 70938 26842 70990 26848
rect 71214 26900 71266 26906
rect 71214 26842 71266 26848
rect 71306 26900 71358 26906
rect 71306 26842 71358 26848
rect 71490 26900 71542 26906
rect 71490 26842 71542 26848
rect 71950 26900 72002 26906
rect 71950 26842 72002 26848
rect 78666 26900 78718 26906
rect 78666 26842 78718 26848
rect 80506 26900 80558 26906
rect 80506 26842 80558 26848
rect 84830 26900 84882 26906
rect 84830 26842 84882 26848
rect 89614 26900 89666 26906
rect 89614 26842 89666 26848
rect 70254 26732 70550 26752
rect 70310 26730 70334 26732
rect 70390 26730 70414 26732
rect 70470 26730 70494 26732
rect 70332 26678 70334 26730
rect 70396 26678 70408 26730
rect 70470 26678 70472 26730
rect 70310 26676 70334 26678
rect 70390 26676 70414 26678
rect 70470 26676 70494 26678
rect 70254 26656 70550 26676
rect 70122 25546 70242 25562
rect 70122 25540 70254 25546
rect 70122 25534 70202 25540
rect 70202 25482 70254 25488
rect 70018 24180 70070 24186
rect 70018 24122 70070 24128
rect 70030 23001 70058 24122
rect 70016 22992 70072 23001
rect 70016 22927 70072 22936
rect 70214 22525 70242 25482
rect 70200 22516 70256 22525
rect 70200 22451 70256 22460
rect 70478 20032 70530 20038
rect 70478 19974 70530 19980
rect 70386 18876 70438 18882
rect 70386 18818 70438 18824
rect 70398 18513 70426 18818
rect 70384 18504 70440 18513
rect 70384 18439 70440 18448
rect 70490 17085 70518 19974
rect 70858 18882 70886 26842
rect 70950 23778 70978 26842
rect 70938 23772 70990 23778
rect 70938 23714 70990 23720
rect 71226 21806 71254 26842
rect 71214 21800 71266 21806
rect 71214 21742 71266 21748
rect 71318 20038 71346 26842
rect 71306 20032 71358 20038
rect 71306 19974 71358 19980
rect 70846 18876 70898 18882
rect 70846 18818 70898 18824
rect 70476 17076 70532 17085
rect 70476 17011 70532 17020
rect 71502 15890 71530 26842
rect 75582 26732 75878 26752
rect 75638 26730 75662 26732
rect 75718 26730 75742 26732
rect 75798 26730 75822 26732
rect 75660 26678 75662 26730
rect 75724 26678 75736 26730
rect 75798 26678 75800 26730
rect 75638 26676 75662 26678
rect 75718 26676 75742 26678
rect 75798 26676 75822 26678
rect 75582 26656 75878 26676
rect 80910 26732 81206 26752
rect 80966 26730 80990 26732
rect 81046 26730 81070 26732
rect 81126 26730 81150 26732
rect 80988 26678 80990 26730
rect 81052 26678 81064 26730
rect 81126 26678 81128 26730
rect 80966 26676 80990 26678
rect 81046 26676 81070 26678
rect 81126 26676 81150 26678
rect 80910 26656 81206 26676
rect 86238 26732 86534 26752
rect 86294 26730 86318 26732
rect 86374 26730 86398 26732
rect 86454 26730 86478 26732
rect 86316 26678 86318 26730
rect 86380 26678 86392 26730
rect 86454 26678 86456 26730
rect 86294 26676 86318 26678
rect 86374 26676 86398 26678
rect 86454 26676 86478 26678
rect 86238 26656 86534 26676
rect 70478 15884 70530 15890
rect 70478 15826 70530 15832
rect 71490 15884 71542 15890
rect 71490 15826 71542 15832
rect 70490 14909 70518 15826
rect 70476 14900 70532 14909
rect 70476 14835 70532 14844
rect 91190 9537 91218 27114
rect 91566 26732 91862 26752
rect 91622 26730 91646 26732
rect 91702 26730 91726 26732
rect 91782 26730 91806 26732
rect 91644 26678 91646 26730
rect 91708 26678 91720 26730
rect 91782 26678 91784 26730
rect 91622 26676 91646 26678
rect 91702 26676 91726 26678
rect 91782 26676 91806 26678
rect 91566 26656 91862 26676
rect 91176 9528 91232 9537
rect 91176 9463 91232 9472
rect 31430 2320 31432 2329
rect 43244 2320 43300 2329
rect 31376 2255 31432 2264
rect 31390 2154 31418 2255
rect 35622 2252 35918 2272
rect 35678 2250 35702 2252
rect 35758 2250 35782 2252
rect 35838 2250 35862 2252
rect 35700 2198 35702 2250
rect 35764 2198 35776 2250
rect 35838 2198 35840 2250
rect 35678 2196 35702 2198
rect 35758 2196 35782 2198
rect 35838 2196 35862 2198
rect 35622 2176 35918 2196
rect 40950 2252 41246 2272
rect 43244 2255 43300 2264
rect 69740 2320 69796 2329
rect 69740 2255 69796 2264
rect 41006 2250 41030 2252
rect 41086 2250 41110 2252
rect 41166 2250 41190 2252
rect 41028 2198 41030 2250
rect 41092 2198 41104 2250
rect 41166 2198 41168 2250
rect 41006 2196 41030 2198
rect 41086 2196 41110 2198
rect 41166 2196 41190 2198
rect 40950 2176 41246 2196
rect 7090 2148 7142 2154
rect 7090 2090 7142 2096
rect 31378 2148 31430 2154
rect 31378 2090 31430 2096
rect 6318 1708 6614 1728
rect 6374 1706 6398 1708
rect 6454 1706 6478 1708
rect 6534 1706 6558 1708
rect 6396 1654 6398 1706
rect 6460 1654 6472 1706
rect 6534 1654 6536 1706
rect 6374 1652 6398 1654
rect 6454 1652 6478 1654
rect 6534 1652 6558 1654
rect 6318 1632 6614 1652
rect 38286 1708 38582 1728
rect 38342 1706 38366 1708
rect 38422 1706 38446 1708
rect 38502 1706 38526 1708
rect 38364 1654 38366 1706
rect 38428 1654 38440 1706
rect 38502 1654 38504 1706
rect 38342 1652 38366 1654
rect 38422 1652 38446 1654
rect 38502 1652 38526 1654
rect 38286 1632 38582 1652
rect 3654 1164 3950 1184
rect 3710 1162 3734 1164
rect 3790 1162 3814 1164
rect 3870 1162 3894 1164
rect 3732 1110 3734 1162
rect 3796 1110 3808 1162
rect 3870 1110 3872 1162
rect 3710 1108 3734 1110
rect 3790 1108 3814 1110
rect 3870 1108 3894 1110
rect 3654 1088 3950 1108
rect 35622 1164 35918 1184
rect 35678 1162 35702 1164
rect 35758 1162 35782 1164
rect 35838 1162 35862 1164
rect 35700 1110 35702 1162
rect 35764 1110 35776 1162
rect 35838 1110 35840 1162
rect 35678 1108 35702 1110
rect 35758 1108 35782 1110
rect 35838 1108 35862 1110
rect 35622 1088 35918 1108
rect 40950 1164 41246 1184
rect 41006 1162 41030 1164
rect 41086 1162 41110 1164
rect 41166 1162 41190 1164
rect 41028 1110 41030 1162
rect 41092 1110 41104 1162
rect 41166 1110 41168 1162
rect 41006 1108 41030 1110
rect 41086 1108 41110 1110
rect 41166 1108 41190 1110
rect 40950 1088 41246 1108
rect 6318 620 6614 640
rect 6374 618 6398 620
rect 6454 618 6478 620
rect 6534 618 6558 620
rect 6396 566 6398 618
rect 6460 566 6472 618
rect 6534 566 6536 618
rect 6374 564 6398 566
rect 6454 564 6478 566
rect 6534 564 6558 566
rect 6318 544 6614 564
rect 38286 620 38582 640
rect 38342 618 38366 620
rect 38422 618 38446 620
rect 38502 618 38526 620
rect 38364 566 38366 618
rect 38428 566 38440 618
rect 38502 566 38504 618
rect 38342 564 38366 566
rect 38422 564 38446 566
rect 38502 564 38526 566
rect 38286 544 38582 564
rect 3654 76 3950 96
rect 3710 74 3734 76
rect 3790 74 3814 76
rect 3870 74 3894 76
rect 3732 22 3734 74
rect 3796 22 3808 74
rect 3870 22 3872 74
rect 3710 20 3734 22
rect 3790 20 3814 22
rect 3870 20 3894 22
rect 3654 0 3950 20
rect 35622 76 35918 96
rect 35678 74 35702 76
rect 35758 74 35782 76
rect 35838 74 35862 76
rect 35700 22 35702 74
rect 35764 22 35776 74
rect 35838 22 35840 74
rect 35678 20 35702 22
rect 35758 20 35782 22
rect 35838 20 35862 22
rect 35622 0 35918 20
rect 40950 76 41246 96
rect 41006 74 41030 76
rect 41086 74 41110 76
rect 41166 74 41190 76
rect 41028 22 41030 74
rect 41092 22 41104 74
rect 41166 22 41168 74
rect 41006 20 41030 22
rect 41086 20 41110 22
rect 41166 20 41190 22
rect 40950 0 41246 20
<< via2 >>
rect 3654 41418 3710 41420
rect 3734 41418 3790 41420
rect 3814 41418 3870 41420
rect 3894 41418 3950 41420
rect 3654 41366 3680 41418
rect 3680 41366 3710 41418
rect 3734 41366 3744 41418
rect 3744 41366 3790 41418
rect 3814 41366 3860 41418
rect 3860 41366 3870 41418
rect 3894 41366 3924 41418
rect 3924 41366 3950 41418
rect 3654 41364 3710 41366
rect 3734 41364 3790 41366
rect 3814 41364 3870 41366
rect 3894 41364 3950 41366
rect 3654 40330 3710 40332
rect 3734 40330 3790 40332
rect 3814 40330 3870 40332
rect 3894 40330 3950 40332
rect 3654 40278 3680 40330
rect 3680 40278 3710 40330
rect 3734 40278 3744 40330
rect 3744 40278 3790 40330
rect 3814 40278 3860 40330
rect 3860 40278 3870 40330
rect 3894 40278 3924 40330
rect 3924 40278 3950 40330
rect 3654 40276 3710 40278
rect 3734 40276 3790 40278
rect 3814 40276 3870 40278
rect 3894 40276 3950 40278
rect 3654 39242 3710 39244
rect 3734 39242 3790 39244
rect 3814 39242 3870 39244
rect 3894 39242 3950 39244
rect 3654 39190 3680 39242
rect 3680 39190 3710 39242
rect 3734 39190 3744 39242
rect 3744 39190 3790 39242
rect 3814 39190 3860 39242
rect 3860 39190 3870 39242
rect 3894 39190 3924 39242
rect 3924 39190 3950 39242
rect 3654 39188 3710 39190
rect 3734 39188 3790 39190
rect 3814 39188 3870 39190
rect 3894 39188 3950 39190
rect 3654 38154 3710 38156
rect 3734 38154 3790 38156
rect 3814 38154 3870 38156
rect 3894 38154 3950 38156
rect 3654 38102 3680 38154
rect 3680 38102 3710 38154
rect 3734 38102 3744 38154
rect 3744 38102 3790 38154
rect 3814 38102 3860 38154
rect 3860 38102 3870 38154
rect 3894 38102 3924 38154
rect 3924 38102 3950 38154
rect 3654 38100 3710 38102
rect 3734 38100 3790 38102
rect 3814 38100 3870 38102
rect 3894 38100 3950 38102
rect 3654 37066 3710 37068
rect 3734 37066 3790 37068
rect 3814 37066 3870 37068
rect 3894 37066 3950 37068
rect 3654 37014 3680 37066
rect 3680 37014 3710 37066
rect 3734 37014 3744 37066
rect 3744 37014 3790 37066
rect 3814 37014 3860 37066
rect 3860 37014 3870 37066
rect 3894 37014 3924 37066
rect 3924 37014 3950 37066
rect 3654 37012 3710 37014
rect 3734 37012 3790 37014
rect 3814 37012 3870 37014
rect 3894 37012 3950 37014
rect 3654 35978 3710 35980
rect 3734 35978 3790 35980
rect 3814 35978 3870 35980
rect 3894 35978 3950 35980
rect 3654 35926 3680 35978
rect 3680 35926 3710 35978
rect 3734 35926 3744 35978
rect 3744 35926 3790 35978
rect 3814 35926 3860 35978
rect 3860 35926 3870 35978
rect 3894 35926 3924 35978
rect 3924 35926 3950 35978
rect 3654 35924 3710 35926
rect 3734 35924 3790 35926
rect 3814 35924 3870 35926
rect 3894 35924 3950 35926
rect 3654 34890 3710 34892
rect 3734 34890 3790 34892
rect 3814 34890 3870 34892
rect 3894 34890 3950 34892
rect 3654 34838 3680 34890
rect 3680 34838 3710 34890
rect 3734 34838 3744 34890
rect 3744 34838 3790 34890
rect 3814 34838 3860 34890
rect 3860 34838 3870 34890
rect 3894 34838 3924 34890
rect 3924 34838 3950 34890
rect 3654 34836 3710 34838
rect 3734 34836 3790 34838
rect 3814 34836 3870 34838
rect 3894 34836 3950 34838
rect 3654 33802 3710 33804
rect 3734 33802 3790 33804
rect 3814 33802 3870 33804
rect 3894 33802 3950 33804
rect 3654 33750 3680 33802
rect 3680 33750 3710 33802
rect 3734 33750 3744 33802
rect 3744 33750 3790 33802
rect 3814 33750 3860 33802
rect 3860 33750 3870 33802
rect 3894 33750 3924 33802
rect 3924 33750 3950 33802
rect 3654 33748 3710 33750
rect 3734 33748 3790 33750
rect 3814 33748 3870 33750
rect 3894 33748 3950 33750
rect 3654 32714 3710 32716
rect 3734 32714 3790 32716
rect 3814 32714 3870 32716
rect 3894 32714 3950 32716
rect 3654 32662 3680 32714
rect 3680 32662 3710 32714
rect 3734 32662 3744 32714
rect 3744 32662 3790 32714
rect 3814 32662 3860 32714
rect 3860 32662 3870 32714
rect 3894 32662 3924 32714
rect 3924 32662 3950 32714
rect 3654 32660 3710 32662
rect 3734 32660 3790 32662
rect 3814 32660 3870 32662
rect 3894 32660 3950 32662
rect 6318 41962 6374 41964
rect 6398 41962 6454 41964
rect 6478 41962 6534 41964
rect 6558 41962 6614 41964
rect 6318 41910 6344 41962
rect 6344 41910 6374 41962
rect 6398 41910 6408 41962
rect 6408 41910 6454 41962
rect 6478 41910 6524 41962
rect 6524 41910 6534 41962
rect 6558 41910 6588 41962
rect 6588 41910 6614 41962
rect 6318 41908 6374 41910
rect 6398 41908 6454 41910
rect 6478 41908 6534 41910
rect 6558 41908 6614 41910
rect 6318 40874 6374 40876
rect 6398 40874 6454 40876
rect 6478 40874 6534 40876
rect 6558 40874 6614 40876
rect 6318 40822 6344 40874
rect 6344 40822 6374 40874
rect 6398 40822 6408 40874
rect 6408 40822 6454 40874
rect 6478 40822 6524 40874
rect 6524 40822 6534 40874
rect 6558 40822 6588 40874
rect 6588 40822 6614 40874
rect 6318 40820 6374 40822
rect 6398 40820 6454 40822
rect 6478 40820 6534 40822
rect 6558 40820 6614 40822
rect 6318 39786 6374 39788
rect 6398 39786 6454 39788
rect 6478 39786 6534 39788
rect 6558 39786 6614 39788
rect 6318 39734 6344 39786
rect 6344 39734 6374 39786
rect 6398 39734 6408 39786
rect 6408 39734 6454 39786
rect 6478 39734 6524 39786
rect 6524 39734 6534 39786
rect 6558 39734 6588 39786
rect 6588 39734 6614 39786
rect 6318 39732 6374 39734
rect 6398 39732 6454 39734
rect 6478 39732 6534 39734
rect 6558 39732 6614 39734
rect 3654 31626 3710 31628
rect 3734 31626 3790 31628
rect 3814 31626 3870 31628
rect 3894 31626 3950 31628
rect 3654 31574 3680 31626
rect 3680 31574 3710 31626
rect 3734 31574 3744 31626
rect 3744 31574 3790 31626
rect 3814 31574 3860 31626
rect 3860 31574 3870 31626
rect 3894 31574 3924 31626
rect 3924 31574 3950 31626
rect 3654 31572 3710 31574
rect 3734 31572 3790 31574
rect 3814 31572 3870 31574
rect 3894 31572 3950 31574
rect 3654 30538 3710 30540
rect 3734 30538 3790 30540
rect 3814 30538 3870 30540
rect 3894 30538 3950 30540
rect 3654 30486 3680 30538
rect 3680 30486 3710 30538
rect 3734 30486 3744 30538
rect 3744 30486 3790 30538
rect 3814 30486 3860 30538
rect 3860 30486 3870 30538
rect 3894 30486 3924 30538
rect 3924 30486 3950 30538
rect 3654 30484 3710 30486
rect 3734 30484 3790 30486
rect 3814 30484 3870 30486
rect 3894 30484 3950 30486
rect 3654 29450 3710 29452
rect 3734 29450 3790 29452
rect 3814 29450 3870 29452
rect 3894 29450 3950 29452
rect 3654 29398 3680 29450
rect 3680 29398 3710 29450
rect 3734 29398 3744 29450
rect 3744 29398 3790 29450
rect 3814 29398 3860 29450
rect 3860 29398 3870 29450
rect 3894 29398 3924 29450
rect 3924 29398 3950 29450
rect 3654 29396 3710 29398
rect 3734 29396 3790 29398
rect 3814 29396 3870 29398
rect 3894 29396 3950 29398
rect 3654 28362 3710 28364
rect 3734 28362 3790 28364
rect 3814 28362 3870 28364
rect 3894 28362 3950 28364
rect 3654 28310 3680 28362
rect 3680 28310 3710 28362
rect 3734 28310 3744 28362
rect 3744 28310 3790 28362
rect 3814 28310 3860 28362
rect 3860 28310 3870 28362
rect 3894 28310 3924 28362
rect 3924 28310 3950 28362
rect 3654 28308 3710 28310
rect 3734 28308 3790 28310
rect 3814 28308 3870 28310
rect 3894 28308 3950 28310
rect 3654 27274 3710 27276
rect 3734 27274 3790 27276
rect 3814 27274 3870 27276
rect 3894 27274 3950 27276
rect 3654 27222 3680 27274
rect 3680 27222 3710 27274
rect 3734 27222 3744 27274
rect 3744 27222 3790 27274
rect 3814 27222 3860 27274
rect 3860 27222 3870 27274
rect 3894 27222 3924 27274
rect 3924 27222 3950 27274
rect 3654 27220 3710 27222
rect 3734 27220 3790 27222
rect 3814 27220 3870 27222
rect 3894 27220 3950 27222
rect 3654 26186 3710 26188
rect 3734 26186 3790 26188
rect 3814 26186 3870 26188
rect 3894 26186 3950 26188
rect 3654 26134 3680 26186
rect 3680 26134 3710 26186
rect 3734 26134 3744 26186
rect 3744 26134 3790 26186
rect 3814 26134 3860 26186
rect 3860 26134 3870 26186
rect 3894 26134 3924 26186
rect 3924 26134 3950 26186
rect 3654 26132 3710 26134
rect 3734 26132 3790 26134
rect 3814 26132 3870 26134
rect 3894 26132 3950 26134
rect 3654 25098 3710 25100
rect 3734 25098 3790 25100
rect 3814 25098 3870 25100
rect 3894 25098 3950 25100
rect 3654 25046 3680 25098
rect 3680 25046 3710 25098
rect 3734 25046 3744 25098
rect 3744 25046 3790 25098
rect 3814 25046 3860 25098
rect 3860 25046 3870 25098
rect 3894 25046 3924 25098
rect 3924 25046 3950 25098
rect 3654 25044 3710 25046
rect 3734 25044 3790 25046
rect 3814 25044 3870 25046
rect 3894 25044 3950 25046
rect 3654 24010 3710 24012
rect 3734 24010 3790 24012
rect 3814 24010 3870 24012
rect 3894 24010 3950 24012
rect 3654 23958 3680 24010
rect 3680 23958 3710 24010
rect 3734 23958 3744 24010
rect 3744 23958 3790 24010
rect 3814 23958 3860 24010
rect 3860 23958 3870 24010
rect 3894 23958 3924 24010
rect 3924 23958 3950 24010
rect 3654 23956 3710 23958
rect 3734 23956 3790 23958
rect 3814 23956 3870 23958
rect 3894 23956 3950 23958
rect 3654 22922 3710 22924
rect 3734 22922 3790 22924
rect 3814 22922 3870 22924
rect 3894 22922 3950 22924
rect 3654 22870 3680 22922
rect 3680 22870 3710 22922
rect 3734 22870 3744 22922
rect 3744 22870 3790 22922
rect 3814 22870 3860 22922
rect 3860 22870 3870 22922
rect 3894 22870 3924 22922
rect 3924 22870 3950 22922
rect 3654 22868 3710 22870
rect 3734 22868 3790 22870
rect 3814 22868 3870 22870
rect 3894 22868 3950 22870
rect 3500 22700 3502 22720
rect 3502 22700 3554 22720
rect 3554 22700 3556 22720
rect 3500 22664 3556 22700
rect 3654 21834 3710 21836
rect 3734 21834 3790 21836
rect 3814 21834 3870 21836
rect 3894 21834 3950 21836
rect 3654 21782 3680 21834
rect 3680 21782 3710 21834
rect 3734 21782 3744 21834
rect 3744 21782 3790 21834
rect 3814 21782 3860 21834
rect 3860 21782 3870 21834
rect 3894 21782 3924 21834
rect 3924 21782 3950 21834
rect 3654 21780 3710 21782
rect 3734 21780 3790 21782
rect 3814 21780 3870 21782
rect 3894 21780 3950 21782
rect 3654 20746 3710 20748
rect 3734 20746 3790 20748
rect 3814 20746 3870 20748
rect 3894 20746 3950 20748
rect 3654 20694 3680 20746
rect 3680 20694 3710 20746
rect 3734 20694 3744 20746
rect 3744 20694 3790 20746
rect 3814 20694 3860 20746
rect 3860 20694 3870 20746
rect 3894 20694 3924 20746
rect 3924 20694 3950 20746
rect 3654 20692 3710 20694
rect 3734 20692 3790 20694
rect 3814 20692 3870 20694
rect 3894 20692 3950 20694
rect 3654 19658 3710 19660
rect 3734 19658 3790 19660
rect 3814 19658 3870 19660
rect 3894 19658 3950 19660
rect 3654 19606 3680 19658
rect 3680 19606 3710 19658
rect 3734 19606 3744 19658
rect 3744 19606 3790 19658
rect 3814 19606 3860 19658
rect 3860 19606 3870 19658
rect 3894 19606 3924 19658
rect 3924 19606 3950 19658
rect 3654 19604 3710 19606
rect 3734 19604 3790 19606
rect 3814 19604 3870 19606
rect 3894 19604 3950 19606
rect 4144 19300 4146 19320
rect 4146 19300 4198 19320
rect 4198 19300 4200 19320
rect 4144 19264 4200 19300
rect 3654 18570 3710 18572
rect 3734 18570 3790 18572
rect 3814 18570 3870 18572
rect 3894 18570 3950 18572
rect 3654 18518 3680 18570
rect 3680 18518 3710 18570
rect 3734 18518 3744 18570
rect 3744 18518 3790 18570
rect 3814 18518 3860 18570
rect 3860 18518 3870 18570
rect 3894 18518 3924 18570
rect 3924 18518 3950 18570
rect 3654 18516 3710 18518
rect 3734 18516 3790 18518
rect 3814 18516 3870 18518
rect 3894 18516 3950 18518
rect 3654 17482 3710 17484
rect 3734 17482 3790 17484
rect 3814 17482 3870 17484
rect 3894 17482 3950 17484
rect 3654 17430 3680 17482
rect 3680 17430 3710 17482
rect 3734 17430 3744 17482
rect 3744 17430 3790 17482
rect 3814 17430 3860 17482
rect 3860 17430 3870 17482
rect 3894 17430 3924 17482
rect 3924 17430 3950 17482
rect 3654 17428 3710 17430
rect 3734 17428 3790 17430
rect 3814 17428 3870 17430
rect 3894 17428 3950 17430
rect 3654 16394 3710 16396
rect 3734 16394 3790 16396
rect 3814 16394 3870 16396
rect 3894 16394 3950 16396
rect 3654 16342 3680 16394
rect 3680 16342 3710 16394
rect 3734 16342 3744 16394
rect 3744 16342 3790 16394
rect 3814 16342 3860 16394
rect 3860 16342 3870 16394
rect 3894 16342 3924 16394
rect 3924 16342 3950 16394
rect 3654 16340 3710 16342
rect 3734 16340 3790 16342
rect 3814 16340 3870 16342
rect 3894 16340 3950 16342
rect 6318 38698 6374 38700
rect 6398 38698 6454 38700
rect 6478 38698 6534 38700
rect 6558 38698 6614 38700
rect 6318 38646 6344 38698
rect 6344 38646 6374 38698
rect 6398 38646 6408 38698
rect 6408 38646 6454 38698
rect 6478 38646 6524 38698
rect 6524 38646 6534 38698
rect 6558 38646 6588 38698
rect 6588 38646 6614 38698
rect 6318 38644 6374 38646
rect 6398 38644 6454 38646
rect 6478 38644 6534 38646
rect 6558 38644 6614 38646
rect 6318 37610 6374 37612
rect 6398 37610 6454 37612
rect 6478 37610 6534 37612
rect 6558 37610 6614 37612
rect 6318 37558 6344 37610
rect 6344 37558 6374 37610
rect 6398 37558 6408 37610
rect 6408 37558 6454 37610
rect 6478 37558 6524 37610
rect 6524 37558 6534 37610
rect 6558 37558 6588 37610
rect 6588 37558 6614 37610
rect 6318 37556 6374 37558
rect 6398 37556 6454 37558
rect 6478 37556 6534 37558
rect 6558 37556 6614 37558
rect 6318 36522 6374 36524
rect 6398 36522 6454 36524
rect 6478 36522 6534 36524
rect 6558 36522 6614 36524
rect 6318 36470 6344 36522
rect 6344 36470 6374 36522
rect 6398 36470 6408 36522
rect 6408 36470 6454 36522
rect 6478 36470 6524 36522
rect 6524 36470 6534 36522
rect 6558 36470 6588 36522
rect 6588 36470 6614 36522
rect 6318 36468 6374 36470
rect 6398 36468 6454 36470
rect 6478 36468 6534 36470
rect 6558 36468 6614 36470
rect 6318 35434 6374 35436
rect 6398 35434 6454 35436
rect 6478 35434 6534 35436
rect 6558 35434 6614 35436
rect 6318 35382 6344 35434
rect 6344 35382 6374 35434
rect 6398 35382 6408 35434
rect 6408 35382 6454 35434
rect 6478 35382 6524 35434
rect 6524 35382 6534 35434
rect 6558 35382 6588 35434
rect 6588 35382 6614 35434
rect 6318 35380 6374 35382
rect 6398 35380 6454 35382
rect 6478 35380 6534 35382
rect 6558 35380 6614 35382
rect 8982 41418 9038 41420
rect 9062 41418 9118 41420
rect 9142 41418 9198 41420
rect 9222 41418 9278 41420
rect 8982 41366 9008 41418
rect 9008 41366 9038 41418
rect 9062 41366 9072 41418
rect 9072 41366 9118 41418
rect 9142 41366 9188 41418
rect 9188 41366 9198 41418
rect 9222 41366 9252 41418
rect 9252 41366 9278 41418
rect 8982 41364 9038 41366
rect 9062 41364 9118 41366
rect 9142 41364 9198 41366
rect 9222 41364 9278 41366
rect 8982 40330 9038 40332
rect 9062 40330 9118 40332
rect 9142 40330 9198 40332
rect 9222 40330 9278 40332
rect 8982 40278 9008 40330
rect 9008 40278 9038 40330
rect 9062 40278 9072 40330
rect 9072 40278 9118 40330
rect 9142 40278 9188 40330
rect 9188 40278 9198 40330
rect 9222 40278 9252 40330
rect 9252 40278 9278 40330
rect 8982 40276 9038 40278
rect 9062 40276 9118 40278
rect 9142 40276 9198 40278
rect 9222 40276 9278 40278
rect 11646 41962 11702 41964
rect 11726 41962 11782 41964
rect 11806 41962 11862 41964
rect 11886 41962 11942 41964
rect 11646 41910 11672 41962
rect 11672 41910 11702 41962
rect 11726 41910 11736 41962
rect 11736 41910 11782 41962
rect 11806 41910 11852 41962
rect 11852 41910 11862 41962
rect 11886 41910 11916 41962
rect 11916 41910 11942 41962
rect 11646 41908 11702 41910
rect 11726 41908 11782 41910
rect 11806 41908 11862 41910
rect 11886 41908 11942 41910
rect 11646 40874 11702 40876
rect 11726 40874 11782 40876
rect 11806 40874 11862 40876
rect 11886 40874 11942 40876
rect 11646 40822 11672 40874
rect 11672 40822 11702 40874
rect 11726 40822 11736 40874
rect 11736 40822 11782 40874
rect 11806 40822 11852 40874
rect 11852 40822 11862 40874
rect 11886 40822 11916 40874
rect 11916 40822 11942 40874
rect 11646 40820 11702 40822
rect 11726 40820 11782 40822
rect 11806 40820 11862 40822
rect 11886 40820 11942 40822
rect 14310 41418 14366 41420
rect 14390 41418 14446 41420
rect 14470 41418 14526 41420
rect 14550 41418 14606 41420
rect 14310 41366 14336 41418
rect 14336 41366 14366 41418
rect 14390 41366 14400 41418
rect 14400 41366 14446 41418
rect 14470 41366 14516 41418
rect 14516 41366 14526 41418
rect 14550 41366 14580 41418
rect 14580 41366 14606 41418
rect 14310 41364 14366 41366
rect 14390 41364 14446 41366
rect 14470 41364 14526 41366
rect 14550 41364 14606 41366
rect 11646 39786 11702 39788
rect 11726 39786 11782 39788
rect 11806 39786 11862 39788
rect 11886 39786 11942 39788
rect 11646 39734 11672 39786
rect 11672 39734 11702 39786
rect 11726 39734 11736 39786
rect 11736 39734 11782 39786
rect 11806 39734 11852 39786
rect 11852 39734 11862 39786
rect 11886 39734 11916 39786
rect 11916 39734 11942 39786
rect 11646 39732 11702 39734
rect 11726 39732 11782 39734
rect 11806 39732 11862 39734
rect 11886 39732 11942 39734
rect 8982 39242 9038 39244
rect 9062 39242 9118 39244
rect 9142 39242 9198 39244
rect 9222 39242 9278 39244
rect 8982 39190 9008 39242
rect 9008 39190 9038 39242
rect 9062 39190 9072 39242
rect 9072 39190 9118 39242
rect 9142 39190 9188 39242
rect 9188 39190 9198 39242
rect 9222 39190 9252 39242
rect 9252 39190 9278 39242
rect 8982 39188 9038 39190
rect 9062 39188 9118 39190
rect 9142 39188 9198 39190
rect 9222 39188 9278 39190
rect 8982 38154 9038 38156
rect 9062 38154 9118 38156
rect 9142 38154 9198 38156
rect 9222 38154 9278 38156
rect 8982 38102 9008 38154
rect 9008 38102 9038 38154
rect 9062 38102 9072 38154
rect 9072 38102 9118 38154
rect 9142 38102 9188 38154
rect 9188 38102 9198 38154
rect 9222 38102 9252 38154
rect 9252 38102 9278 38154
rect 8982 38100 9038 38102
rect 9062 38100 9118 38102
rect 9142 38100 9198 38102
rect 9222 38100 9278 38102
rect 9112 37932 9114 37952
rect 9114 37932 9166 37952
rect 9166 37932 9168 37952
rect 9112 37896 9168 37932
rect 8982 37066 9038 37068
rect 9062 37066 9118 37068
rect 9142 37066 9198 37068
rect 9222 37066 9278 37068
rect 8982 37014 9008 37066
rect 9008 37014 9038 37066
rect 9062 37014 9072 37066
rect 9072 37014 9118 37066
rect 9142 37014 9188 37066
rect 9188 37014 9198 37066
rect 9222 37014 9252 37066
rect 9252 37014 9278 37066
rect 8982 37012 9038 37014
rect 9062 37012 9118 37014
rect 9142 37012 9198 37014
rect 9222 37012 9278 37014
rect 8982 35978 9038 35980
rect 9062 35978 9118 35980
rect 9142 35978 9198 35980
rect 9222 35978 9278 35980
rect 8982 35926 9008 35978
rect 9008 35926 9038 35978
rect 9062 35926 9072 35978
rect 9072 35926 9118 35978
rect 9142 35926 9188 35978
rect 9188 35926 9198 35978
rect 9222 35926 9252 35978
rect 9252 35926 9278 35978
rect 8982 35924 9038 35926
rect 9062 35924 9118 35926
rect 9142 35924 9198 35926
rect 9222 35924 9278 35926
rect 6318 34346 6374 34348
rect 6398 34346 6454 34348
rect 6478 34346 6534 34348
rect 6558 34346 6614 34348
rect 6318 34294 6344 34346
rect 6344 34294 6374 34346
rect 6398 34294 6408 34346
rect 6408 34294 6454 34346
rect 6478 34294 6524 34346
rect 6524 34294 6534 34346
rect 6558 34294 6588 34346
rect 6588 34294 6614 34346
rect 6318 34292 6374 34294
rect 6398 34292 6454 34294
rect 6478 34292 6534 34294
rect 6558 34292 6614 34294
rect 6318 33258 6374 33260
rect 6398 33258 6454 33260
rect 6478 33258 6534 33260
rect 6558 33258 6614 33260
rect 6318 33206 6344 33258
rect 6344 33206 6374 33258
rect 6398 33206 6408 33258
rect 6408 33206 6454 33258
rect 6478 33206 6524 33258
rect 6524 33206 6534 33258
rect 6558 33206 6588 33258
rect 6588 33206 6614 33258
rect 6318 33204 6374 33206
rect 6398 33204 6454 33206
rect 6478 33204 6534 33206
rect 6558 33204 6614 33206
rect 6318 32170 6374 32172
rect 6398 32170 6454 32172
rect 6478 32170 6534 32172
rect 6558 32170 6614 32172
rect 6318 32118 6344 32170
rect 6344 32118 6374 32170
rect 6398 32118 6408 32170
rect 6408 32118 6454 32170
rect 6478 32118 6524 32170
rect 6524 32118 6534 32170
rect 6558 32118 6588 32170
rect 6588 32118 6614 32170
rect 6318 32116 6374 32118
rect 6398 32116 6454 32118
rect 6478 32116 6534 32118
rect 6558 32116 6614 32118
rect 6318 31082 6374 31084
rect 6398 31082 6454 31084
rect 6478 31082 6534 31084
rect 6558 31082 6614 31084
rect 6318 31030 6344 31082
rect 6344 31030 6374 31082
rect 6398 31030 6408 31082
rect 6408 31030 6454 31082
rect 6478 31030 6524 31082
rect 6524 31030 6534 31082
rect 6558 31030 6588 31082
rect 6588 31030 6614 31082
rect 6318 31028 6374 31030
rect 6398 31028 6454 31030
rect 6478 31028 6534 31030
rect 6558 31028 6614 31030
rect 6318 29994 6374 29996
rect 6398 29994 6454 29996
rect 6478 29994 6534 29996
rect 6558 29994 6614 29996
rect 6318 29942 6344 29994
rect 6344 29942 6374 29994
rect 6398 29942 6408 29994
rect 6408 29942 6454 29994
rect 6478 29942 6524 29994
rect 6524 29942 6534 29994
rect 6558 29942 6588 29994
rect 6588 29942 6614 29994
rect 6318 29940 6374 29942
rect 6398 29940 6454 29942
rect 6478 29940 6534 29942
rect 6558 29940 6614 29942
rect 6318 28906 6374 28908
rect 6398 28906 6454 28908
rect 6478 28906 6534 28908
rect 6558 28906 6614 28908
rect 6318 28854 6344 28906
rect 6344 28854 6374 28906
rect 6398 28854 6408 28906
rect 6408 28854 6454 28906
rect 6478 28854 6524 28906
rect 6524 28854 6534 28906
rect 6558 28854 6588 28906
rect 6588 28854 6614 28906
rect 6318 28852 6374 28854
rect 6398 28852 6454 28854
rect 6478 28852 6534 28854
rect 6558 28852 6614 28854
rect 6318 27818 6374 27820
rect 6398 27818 6454 27820
rect 6478 27818 6534 27820
rect 6558 27818 6614 27820
rect 6318 27766 6344 27818
rect 6344 27766 6374 27818
rect 6398 27766 6408 27818
rect 6408 27766 6454 27818
rect 6478 27766 6524 27818
rect 6524 27766 6534 27818
rect 6558 27766 6588 27818
rect 6588 27766 6614 27818
rect 6318 27764 6374 27766
rect 6398 27764 6454 27766
rect 6478 27764 6534 27766
rect 6558 27764 6614 27766
rect 6318 26730 6374 26732
rect 6398 26730 6454 26732
rect 6478 26730 6534 26732
rect 6558 26730 6614 26732
rect 6318 26678 6344 26730
rect 6344 26678 6374 26730
rect 6398 26678 6408 26730
rect 6408 26678 6454 26730
rect 6478 26678 6524 26730
rect 6524 26678 6534 26730
rect 6558 26678 6588 26730
rect 6588 26678 6614 26730
rect 6318 26676 6374 26678
rect 6398 26676 6454 26678
rect 6478 26676 6534 26678
rect 6558 26676 6614 26678
rect 6318 25642 6374 25644
rect 6398 25642 6454 25644
rect 6478 25642 6534 25644
rect 6558 25642 6614 25644
rect 6318 25590 6344 25642
rect 6344 25590 6374 25642
rect 6398 25590 6408 25642
rect 6408 25590 6454 25642
rect 6478 25590 6524 25642
rect 6524 25590 6534 25642
rect 6558 25590 6588 25642
rect 6588 25590 6614 25642
rect 6318 25588 6374 25590
rect 6398 25588 6454 25590
rect 6478 25588 6534 25590
rect 6558 25588 6614 25590
rect 6318 24554 6374 24556
rect 6398 24554 6454 24556
rect 6478 24554 6534 24556
rect 6558 24554 6614 24556
rect 6318 24502 6344 24554
rect 6344 24502 6374 24554
rect 6398 24502 6408 24554
rect 6408 24502 6454 24554
rect 6478 24502 6524 24554
rect 6524 24502 6534 24554
rect 6558 24502 6588 24554
rect 6588 24502 6614 24554
rect 6318 24500 6374 24502
rect 6398 24500 6454 24502
rect 6478 24500 6534 24502
rect 6558 24500 6614 24502
rect 6318 23466 6374 23468
rect 6398 23466 6454 23468
rect 6478 23466 6534 23468
rect 6558 23466 6614 23468
rect 6318 23414 6344 23466
rect 6344 23414 6374 23466
rect 6398 23414 6408 23466
rect 6408 23414 6454 23466
rect 6478 23414 6524 23466
rect 6524 23414 6534 23466
rect 6558 23414 6588 23466
rect 6588 23414 6614 23466
rect 6318 23412 6374 23414
rect 6398 23412 6454 23414
rect 6478 23412 6534 23414
rect 6558 23412 6614 23414
rect 6318 22378 6374 22380
rect 6398 22378 6454 22380
rect 6478 22378 6534 22380
rect 6558 22378 6614 22380
rect 6318 22326 6344 22378
rect 6344 22326 6374 22378
rect 6398 22326 6408 22378
rect 6408 22326 6454 22378
rect 6478 22326 6524 22378
rect 6524 22326 6534 22378
rect 6558 22326 6588 22378
rect 6588 22326 6614 22378
rect 6318 22324 6374 22326
rect 6398 22324 6454 22326
rect 6478 22324 6534 22326
rect 6558 22324 6614 22326
rect 6318 21290 6374 21292
rect 6398 21290 6454 21292
rect 6478 21290 6534 21292
rect 6558 21290 6614 21292
rect 6318 21238 6344 21290
rect 6344 21238 6374 21290
rect 6398 21238 6408 21290
rect 6408 21238 6454 21290
rect 6478 21238 6524 21290
rect 6524 21238 6534 21290
rect 6558 21238 6588 21290
rect 6588 21238 6614 21290
rect 6318 21236 6374 21238
rect 6398 21236 6454 21238
rect 6478 21236 6534 21238
rect 6558 21236 6614 21238
rect 8982 34890 9038 34892
rect 9062 34890 9118 34892
rect 9142 34890 9198 34892
rect 9222 34890 9278 34892
rect 8982 34838 9008 34890
rect 9008 34838 9038 34890
rect 9062 34838 9072 34890
rect 9072 34838 9118 34890
rect 9142 34838 9188 34890
rect 9188 34838 9198 34890
rect 9222 34838 9252 34890
rect 9252 34838 9278 34890
rect 8982 34836 9038 34838
rect 9062 34836 9118 34838
rect 9142 34836 9198 34838
rect 9222 34836 9278 34838
rect 11646 38698 11702 38700
rect 11726 38698 11782 38700
rect 11806 38698 11862 38700
rect 11886 38698 11942 38700
rect 11646 38646 11672 38698
rect 11672 38646 11702 38698
rect 11726 38646 11736 38698
rect 11736 38646 11782 38698
rect 11806 38646 11852 38698
rect 11852 38646 11862 38698
rect 11886 38646 11916 38698
rect 11916 38646 11942 38698
rect 11646 38644 11702 38646
rect 11726 38644 11782 38646
rect 11806 38644 11862 38646
rect 11886 38644 11942 38646
rect 14310 40330 14366 40332
rect 14390 40330 14446 40332
rect 14470 40330 14526 40332
rect 14550 40330 14606 40332
rect 14310 40278 14336 40330
rect 14336 40278 14366 40330
rect 14390 40278 14400 40330
rect 14400 40278 14446 40330
rect 14470 40278 14516 40330
rect 14516 40278 14526 40330
rect 14550 40278 14580 40330
rect 14580 40278 14606 40330
rect 14310 40276 14366 40278
rect 14390 40276 14446 40278
rect 14470 40276 14526 40278
rect 14550 40276 14606 40278
rect 11646 37610 11702 37612
rect 11726 37610 11782 37612
rect 11806 37610 11862 37612
rect 11886 37610 11942 37612
rect 11646 37558 11672 37610
rect 11672 37558 11702 37610
rect 11726 37558 11736 37610
rect 11736 37558 11782 37610
rect 11806 37558 11852 37610
rect 11852 37558 11862 37610
rect 11886 37558 11916 37610
rect 11916 37558 11942 37610
rect 11646 37556 11702 37558
rect 11726 37556 11782 37558
rect 11806 37556 11862 37558
rect 11886 37556 11942 37558
rect 11646 36522 11702 36524
rect 11726 36522 11782 36524
rect 11806 36522 11862 36524
rect 11886 36522 11942 36524
rect 11646 36470 11672 36522
rect 11672 36470 11702 36522
rect 11726 36470 11736 36522
rect 11736 36470 11782 36522
rect 11806 36470 11852 36522
rect 11852 36470 11862 36522
rect 11886 36470 11916 36522
rect 11916 36470 11942 36522
rect 11646 36468 11702 36470
rect 11726 36468 11782 36470
rect 11806 36468 11862 36470
rect 11886 36468 11942 36470
rect 11646 35434 11702 35436
rect 11726 35434 11782 35436
rect 11806 35434 11862 35436
rect 11886 35434 11942 35436
rect 11646 35382 11672 35434
rect 11672 35382 11702 35434
rect 11726 35382 11736 35434
rect 11736 35382 11782 35434
rect 11806 35382 11852 35434
rect 11852 35382 11862 35434
rect 11886 35382 11916 35434
rect 11916 35382 11942 35434
rect 11646 35380 11702 35382
rect 11726 35380 11782 35382
rect 11806 35380 11862 35382
rect 11886 35380 11942 35382
rect 8982 33802 9038 33804
rect 9062 33802 9118 33804
rect 9142 33802 9198 33804
rect 9222 33802 9278 33804
rect 8982 33750 9008 33802
rect 9008 33750 9038 33802
rect 9062 33750 9072 33802
rect 9072 33750 9118 33802
rect 9142 33750 9188 33802
rect 9188 33750 9198 33802
rect 9222 33750 9252 33802
rect 9252 33750 9278 33802
rect 8982 33748 9038 33750
rect 9062 33748 9118 33750
rect 9142 33748 9198 33750
rect 9222 33748 9278 33750
rect 8982 32714 9038 32716
rect 9062 32714 9118 32716
rect 9142 32714 9198 32716
rect 9222 32714 9278 32716
rect 8982 32662 9008 32714
rect 9008 32662 9038 32714
rect 9062 32662 9072 32714
rect 9072 32662 9118 32714
rect 9142 32662 9188 32714
rect 9188 32662 9198 32714
rect 9222 32662 9252 32714
rect 9252 32662 9278 32714
rect 8982 32660 9038 32662
rect 9062 32660 9118 32662
rect 9142 32660 9198 32662
rect 9222 32660 9278 32662
rect 8982 31626 9038 31628
rect 9062 31626 9118 31628
rect 9142 31626 9198 31628
rect 9222 31626 9278 31628
rect 8982 31574 9008 31626
rect 9008 31574 9038 31626
rect 9062 31574 9072 31626
rect 9072 31574 9118 31626
rect 9142 31574 9188 31626
rect 9188 31574 9198 31626
rect 9222 31574 9252 31626
rect 9252 31574 9278 31626
rect 8982 31572 9038 31574
rect 9062 31572 9118 31574
rect 9142 31572 9198 31574
rect 9222 31572 9278 31574
rect 8982 30538 9038 30540
rect 9062 30538 9118 30540
rect 9142 30538 9198 30540
rect 9222 30538 9278 30540
rect 8982 30486 9008 30538
rect 9008 30486 9038 30538
rect 9062 30486 9072 30538
rect 9072 30486 9118 30538
rect 9142 30486 9188 30538
rect 9188 30486 9198 30538
rect 9222 30486 9252 30538
rect 9252 30486 9278 30538
rect 8982 30484 9038 30486
rect 9062 30484 9118 30486
rect 9142 30484 9198 30486
rect 9222 30484 9278 30486
rect 8982 29450 9038 29452
rect 9062 29450 9118 29452
rect 9142 29450 9198 29452
rect 9222 29450 9278 29452
rect 8982 29398 9008 29450
rect 9008 29398 9038 29450
rect 9062 29398 9072 29450
rect 9072 29398 9118 29450
rect 9142 29398 9188 29450
rect 9188 29398 9198 29450
rect 9222 29398 9252 29450
rect 9252 29398 9278 29450
rect 8982 29396 9038 29398
rect 9062 29396 9118 29398
rect 9142 29396 9198 29398
rect 9222 29396 9278 29398
rect 8982 28362 9038 28364
rect 9062 28362 9118 28364
rect 9142 28362 9198 28364
rect 9222 28362 9278 28364
rect 8982 28310 9008 28362
rect 9008 28310 9038 28362
rect 9062 28310 9072 28362
rect 9072 28310 9118 28362
rect 9142 28310 9188 28362
rect 9188 28310 9198 28362
rect 9222 28310 9252 28362
rect 9252 28310 9278 28362
rect 8982 28308 9038 28310
rect 9062 28308 9118 28310
rect 9142 28308 9198 28310
rect 9222 28308 9278 28310
rect 8982 27274 9038 27276
rect 9062 27274 9118 27276
rect 9142 27274 9198 27276
rect 9222 27274 9278 27276
rect 8982 27222 9008 27274
rect 9008 27222 9038 27274
rect 9062 27222 9072 27274
rect 9072 27222 9118 27274
rect 9142 27222 9188 27274
rect 9188 27222 9198 27274
rect 9222 27222 9252 27274
rect 9252 27222 9278 27274
rect 8982 27220 9038 27222
rect 9062 27220 9118 27222
rect 9142 27220 9198 27222
rect 9222 27220 9278 27222
rect 10124 27424 10180 27480
rect 6318 20202 6374 20204
rect 6398 20202 6454 20204
rect 6478 20202 6534 20204
rect 6558 20202 6614 20204
rect 6318 20150 6344 20202
rect 6344 20150 6374 20202
rect 6398 20150 6408 20202
rect 6408 20150 6454 20202
rect 6478 20150 6524 20202
rect 6524 20150 6534 20202
rect 6558 20150 6588 20202
rect 6588 20150 6614 20202
rect 6318 20148 6374 20150
rect 6398 20148 6454 20150
rect 6478 20148 6534 20150
rect 6558 20148 6614 20150
rect 6812 19980 6814 20000
rect 6814 19980 6866 20000
rect 6866 19980 6868 20000
rect 6812 19944 6868 19980
rect 6318 19114 6374 19116
rect 6398 19114 6454 19116
rect 6478 19114 6534 19116
rect 6558 19114 6614 19116
rect 6318 19062 6344 19114
rect 6344 19062 6374 19114
rect 6398 19062 6408 19114
rect 6408 19062 6454 19114
rect 6478 19062 6524 19114
rect 6524 19062 6534 19114
rect 6558 19062 6588 19114
rect 6588 19062 6614 19114
rect 6318 19060 6374 19062
rect 6398 19060 6454 19062
rect 6478 19060 6534 19062
rect 6558 19060 6614 19062
rect 6318 18026 6374 18028
rect 6398 18026 6454 18028
rect 6478 18026 6534 18028
rect 6558 18026 6614 18028
rect 6318 17974 6344 18026
rect 6344 17974 6374 18026
rect 6398 17974 6408 18026
rect 6408 17974 6454 18026
rect 6478 17974 6524 18026
rect 6524 17974 6534 18026
rect 6558 17974 6588 18026
rect 6588 17974 6614 18026
rect 6318 17972 6374 17974
rect 6398 17972 6454 17974
rect 6478 17972 6534 17974
rect 6558 17972 6614 17974
rect 5064 17224 5120 17280
rect 5708 16580 5710 16600
rect 5710 16580 5762 16600
rect 5762 16580 5764 16600
rect 5708 16544 5764 16580
rect 7272 17532 7274 17552
rect 7274 17532 7326 17552
rect 7326 17532 7328 17552
rect 7272 17496 7328 17532
rect 6318 16938 6374 16940
rect 6398 16938 6454 16940
rect 6478 16938 6534 16940
rect 6558 16938 6614 16940
rect 6318 16886 6344 16938
rect 6344 16886 6374 16938
rect 6398 16886 6408 16938
rect 6408 16886 6454 16938
rect 6478 16886 6524 16938
rect 6524 16886 6534 16938
rect 6558 16886 6588 16938
rect 6588 16886 6614 16938
rect 6318 16884 6374 16886
rect 6398 16884 6454 16886
rect 6478 16884 6534 16886
rect 6558 16884 6614 16886
rect 6318 15850 6374 15852
rect 6398 15850 6454 15852
rect 6478 15850 6534 15852
rect 6558 15850 6614 15852
rect 6318 15798 6344 15850
rect 6344 15798 6374 15850
rect 6398 15798 6408 15850
rect 6408 15798 6454 15850
rect 6478 15798 6524 15850
rect 6524 15798 6534 15850
rect 6558 15798 6588 15850
rect 6588 15798 6614 15850
rect 6318 15796 6374 15798
rect 6398 15796 6454 15798
rect 6478 15796 6534 15798
rect 6558 15796 6614 15798
rect 3654 15306 3710 15308
rect 3734 15306 3790 15308
rect 3814 15306 3870 15308
rect 3894 15306 3950 15308
rect 3654 15254 3680 15306
rect 3680 15254 3710 15306
rect 3734 15254 3744 15306
rect 3744 15254 3790 15306
rect 3814 15254 3860 15306
rect 3860 15254 3870 15306
rect 3894 15254 3924 15306
rect 3924 15254 3950 15306
rect 3654 15252 3710 15254
rect 3734 15252 3790 15254
rect 3814 15252 3870 15254
rect 3894 15252 3950 15254
rect 6318 14762 6374 14764
rect 6398 14762 6454 14764
rect 6478 14762 6534 14764
rect 6558 14762 6614 14764
rect 6318 14710 6344 14762
rect 6344 14710 6374 14762
rect 6398 14710 6408 14762
rect 6408 14710 6454 14762
rect 6478 14710 6524 14762
rect 6524 14710 6534 14762
rect 6558 14710 6588 14762
rect 6588 14710 6614 14762
rect 6318 14708 6374 14710
rect 6398 14708 6454 14710
rect 6478 14708 6534 14710
rect 6558 14708 6614 14710
rect 3654 14218 3710 14220
rect 3734 14218 3790 14220
rect 3814 14218 3870 14220
rect 3894 14218 3950 14220
rect 3654 14166 3680 14218
rect 3680 14166 3710 14218
rect 3734 14166 3744 14218
rect 3744 14166 3790 14218
rect 3814 14166 3860 14218
rect 3860 14166 3870 14218
rect 3894 14166 3924 14218
rect 3924 14166 3950 14218
rect 3654 14164 3710 14166
rect 3734 14164 3790 14166
rect 3814 14164 3870 14166
rect 3894 14164 3950 14166
rect 3654 13130 3710 13132
rect 3734 13130 3790 13132
rect 3814 13130 3870 13132
rect 3894 13130 3950 13132
rect 3654 13078 3680 13130
rect 3680 13078 3710 13130
rect 3734 13078 3744 13130
rect 3744 13078 3790 13130
rect 3814 13078 3860 13130
rect 3860 13078 3870 13130
rect 3894 13078 3924 13130
rect 3924 13078 3950 13130
rect 3654 13076 3710 13078
rect 3734 13076 3790 13078
rect 3814 13076 3870 13078
rect 3894 13076 3950 13078
rect 3654 12042 3710 12044
rect 3734 12042 3790 12044
rect 3814 12042 3870 12044
rect 3894 12042 3950 12044
rect 3654 11990 3680 12042
rect 3680 11990 3710 12042
rect 3734 11990 3744 12042
rect 3744 11990 3790 12042
rect 3814 11990 3860 12042
rect 3860 11990 3870 12042
rect 3894 11990 3924 12042
rect 3924 11990 3950 12042
rect 3654 11988 3710 11990
rect 3734 11988 3790 11990
rect 3814 11988 3870 11990
rect 3894 11988 3950 11990
rect 3654 10954 3710 10956
rect 3734 10954 3790 10956
rect 3814 10954 3870 10956
rect 3894 10954 3950 10956
rect 3654 10902 3680 10954
rect 3680 10902 3710 10954
rect 3734 10902 3744 10954
rect 3744 10902 3790 10954
rect 3814 10902 3860 10954
rect 3860 10902 3870 10954
rect 3894 10902 3924 10954
rect 3924 10902 3950 10954
rect 3654 10900 3710 10902
rect 3734 10900 3790 10902
rect 3814 10900 3870 10902
rect 3894 10900 3950 10902
rect 6996 15184 7052 15240
rect 7364 14524 7420 14560
rect 7364 14504 7366 14524
rect 7366 14504 7418 14524
rect 7418 14504 7420 14524
rect 6318 13674 6374 13676
rect 6398 13674 6454 13676
rect 6478 13674 6534 13676
rect 6558 13674 6614 13676
rect 6318 13622 6344 13674
rect 6344 13622 6374 13674
rect 6398 13622 6408 13674
rect 6408 13622 6454 13674
rect 6478 13622 6524 13674
rect 6524 13622 6534 13674
rect 6558 13622 6588 13674
rect 6588 13622 6614 13674
rect 6318 13620 6374 13622
rect 6398 13620 6454 13622
rect 6478 13620 6534 13622
rect 6558 13620 6614 13622
rect 6318 12586 6374 12588
rect 6398 12586 6454 12588
rect 6478 12586 6534 12588
rect 6558 12586 6614 12588
rect 6318 12534 6344 12586
rect 6344 12534 6374 12586
rect 6398 12534 6408 12586
rect 6408 12534 6454 12586
rect 6478 12534 6524 12586
rect 6524 12534 6534 12586
rect 6558 12534 6588 12586
rect 6588 12534 6614 12586
rect 6318 12532 6374 12534
rect 6398 12532 6454 12534
rect 6478 12532 6534 12534
rect 6558 12532 6614 12534
rect 6318 11498 6374 11500
rect 6398 11498 6454 11500
rect 6478 11498 6534 11500
rect 6558 11498 6614 11500
rect 6318 11446 6344 11498
rect 6344 11446 6374 11498
rect 6398 11446 6408 11498
rect 6408 11446 6454 11498
rect 6478 11446 6524 11498
rect 6524 11446 6534 11498
rect 6558 11446 6588 11498
rect 6588 11446 6614 11498
rect 6318 11444 6374 11446
rect 6398 11444 6454 11446
rect 6478 11444 6534 11446
rect 6558 11444 6614 11446
rect 6318 10410 6374 10412
rect 6398 10410 6454 10412
rect 6478 10410 6534 10412
rect 6558 10410 6614 10412
rect 6318 10358 6344 10410
rect 6344 10358 6374 10410
rect 6398 10358 6408 10410
rect 6408 10358 6454 10410
rect 6478 10358 6524 10410
rect 6524 10358 6534 10410
rect 6558 10358 6588 10410
rect 6588 10358 6614 10410
rect 6318 10356 6374 10358
rect 6398 10356 6454 10358
rect 6478 10356 6534 10358
rect 6558 10356 6614 10358
rect 11646 34346 11702 34348
rect 11726 34346 11782 34348
rect 11806 34346 11862 34348
rect 11886 34346 11942 34348
rect 11646 34294 11672 34346
rect 11672 34294 11702 34346
rect 11726 34294 11736 34346
rect 11736 34294 11782 34346
rect 11806 34294 11852 34346
rect 11852 34294 11862 34346
rect 11886 34294 11916 34346
rect 11916 34294 11942 34346
rect 11646 34292 11702 34294
rect 11726 34292 11782 34294
rect 11806 34292 11862 34294
rect 11886 34292 11942 34294
rect 11646 33258 11702 33260
rect 11726 33258 11782 33260
rect 11806 33258 11862 33260
rect 11886 33258 11942 33260
rect 11646 33206 11672 33258
rect 11672 33206 11702 33258
rect 11726 33206 11736 33258
rect 11736 33206 11782 33258
rect 11806 33206 11852 33258
rect 11852 33206 11862 33258
rect 11886 33206 11916 33258
rect 11916 33206 11942 33258
rect 11646 33204 11702 33206
rect 11726 33204 11782 33206
rect 11806 33204 11862 33206
rect 11886 33204 11942 33206
rect 11646 32170 11702 32172
rect 11726 32170 11782 32172
rect 11806 32170 11862 32172
rect 11886 32170 11942 32172
rect 11646 32118 11672 32170
rect 11672 32118 11702 32170
rect 11726 32118 11736 32170
rect 11736 32118 11782 32170
rect 11806 32118 11852 32170
rect 11852 32118 11862 32170
rect 11886 32118 11916 32170
rect 11916 32118 11942 32170
rect 11646 32116 11702 32118
rect 11726 32116 11782 32118
rect 11806 32116 11862 32118
rect 11886 32116 11942 32118
rect 11646 31082 11702 31084
rect 11726 31082 11782 31084
rect 11806 31082 11862 31084
rect 11886 31082 11942 31084
rect 11646 31030 11672 31082
rect 11672 31030 11702 31082
rect 11726 31030 11736 31082
rect 11736 31030 11782 31082
rect 11806 31030 11852 31082
rect 11852 31030 11862 31082
rect 11886 31030 11916 31082
rect 11916 31030 11942 31082
rect 11646 31028 11702 31030
rect 11726 31028 11782 31030
rect 11806 31028 11862 31030
rect 11886 31028 11942 31030
rect 11646 29994 11702 29996
rect 11726 29994 11782 29996
rect 11806 29994 11862 29996
rect 11886 29994 11942 29996
rect 11646 29942 11672 29994
rect 11672 29942 11702 29994
rect 11726 29942 11736 29994
rect 11736 29942 11782 29994
rect 11806 29942 11852 29994
rect 11852 29942 11862 29994
rect 11886 29942 11916 29994
rect 11916 29942 11942 29994
rect 11646 29940 11702 29942
rect 11726 29940 11782 29942
rect 11806 29940 11862 29942
rect 11886 29940 11942 29942
rect 11646 28906 11702 28908
rect 11726 28906 11782 28908
rect 11806 28906 11862 28908
rect 11886 28906 11942 28908
rect 11646 28854 11672 28906
rect 11672 28854 11702 28906
rect 11726 28854 11736 28906
rect 11736 28854 11782 28906
rect 11806 28854 11852 28906
rect 11852 28854 11862 28906
rect 11886 28854 11916 28906
rect 11916 28854 11942 28906
rect 11646 28852 11702 28854
rect 11726 28852 11782 28854
rect 11806 28852 11862 28854
rect 11886 28852 11942 28854
rect 11646 27818 11702 27820
rect 11726 27818 11782 27820
rect 11806 27818 11862 27820
rect 11886 27818 11942 27820
rect 11646 27766 11672 27818
rect 11672 27766 11702 27818
rect 11726 27766 11736 27818
rect 11736 27766 11782 27818
rect 11806 27766 11852 27818
rect 11852 27766 11862 27818
rect 11886 27766 11916 27818
rect 11916 27766 11942 27818
rect 11646 27764 11702 27766
rect 11726 27764 11782 27766
rect 11806 27764 11862 27766
rect 11886 27764 11942 27766
rect 12700 28104 12756 28160
rect 14310 39242 14366 39244
rect 14390 39242 14446 39244
rect 14470 39242 14526 39244
rect 14550 39242 14606 39244
rect 14310 39190 14336 39242
rect 14336 39190 14366 39242
rect 14390 39190 14400 39242
rect 14400 39190 14446 39242
rect 14470 39190 14516 39242
rect 14516 39190 14526 39242
rect 14550 39190 14580 39242
rect 14580 39190 14606 39242
rect 14310 39188 14366 39190
rect 14390 39188 14446 39190
rect 14470 39188 14526 39190
rect 14550 39188 14606 39190
rect 14310 38154 14366 38156
rect 14390 38154 14446 38156
rect 14470 38154 14526 38156
rect 14550 38154 14606 38156
rect 14310 38102 14336 38154
rect 14336 38102 14366 38154
rect 14390 38102 14400 38154
rect 14400 38102 14446 38154
rect 14470 38102 14516 38154
rect 14516 38102 14526 38154
rect 14550 38102 14580 38154
rect 14580 38102 14606 38154
rect 14310 38100 14366 38102
rect 14390 38100 14446 38102
rect 14470 38100 14526 38102
rect 14550 38100 14606 38102
rect 14310 37066 14366 37068
rect 14390 37066 14446 37068
rect 14470 37066 14526 37068
rect 14550 37066 14606 37068
rect 14310 37014 14336 37066
rect 14336 37014 14366 37066
rect 14390 37014 14400 37066
rect 14400 37014 14446 37066
rect 14470 37014 14516 37066
rect 14516 37014 14526 37066
rect 14550 37014 14580 37066
rect 14580 37014 14606 37066
rect 14310 37012 14366 37014
rect 14390 37012 14446 37014
rect 14470 37012 14526 37014
rect 14550 37012 14606 37014
rect 14310 35978 14366 35980
rect 14390 35978 14446 35980
rect 14470 35978 14526 35980
rect 14550 35978 14606 35980
rect 14310 35926 14336 35978
rect 14336 35926 14366 35978
rect 14390 35926 14400 35978
rect 14400 35926 14446 35978
rect 14470 35926 14516 35978
rect 14516 35926 14526 35978
rect 14550 35926 14580 35978
rect 14580 35926 14606 35978
rect 14310 35924 14366 35926
rect 14390 35924 14446 35926
rect 14470 35924 14526 35926
rect 14550 35924 14606 35926
rect 14724 35196 14780 35232
rect 14724 35176 14726 35196
rect 14726 35176 14778 35196
rect 14778 35176 14780 35196
rect 15092 35212 15094 35232
rect 15094 35212 15146 35232
rect 15146 35212 15148 35232
rect 15092 35176 15148 35212
rect 14310 34890 14366 34892
rect 14390 34890 14446 34892
rect 14470 34890 14526 34892
rect 14550 34890 14606 34892
rect 14310 34838 14336 34890
rect 14336 34838 14366 34890
rect 14390 34838 14400 34890
rect 14400 34838 14446 34890
rect 14470 34838 14516 34890
rect 14516 34838 14526 34890
rect 14550 34838 14580 34890
rect 14580 34838 14606 34890
rect 14310 34836 14366 34838
rect 14390 34836 14446 34838
rect 14470 34836 14526 34838
rect 14550 34836 14606 34838
rect 14310 33802 14366 33804
rect 14390 33802 14446 33804
rect 14470 33802 14526 33804
rect 14550 33802 14606 33804
rect 14310 33750 14336 33802
rect 14336 33750 14366 33802
rect 14390 33750 14400 33802
rect 14400 33750 14446 33802
rect 14470 33750 14516 33802
rect 14516 33750 14526 33802
rect 14550 33750 14580 33802
rect 14580 33750 14606 33802
rect 14310 33748 14366 33750
rect 14390 33748 14446 33750
rect 14470 33748 14526 33750
rect 14550 33748 14606 33750
rect 13896 33444 13898 33464
rect 13898 33444 13950 33464
rect 13950 33444 13952 33464
rect 13896 33408 13952 33444
rect 14310 32714 14366 32716
rect 14390 32714 14446 32716
rect 14470 32714 14526 32716
rect 14550 32714 14606 32716
rect 14310 32662 14336 32714
rect 14336 32662 14366 32714
rect 14390 32662 14400 32714
rect 14400 32662 14446 32714
rect 14470 32662 14516 32714
rect 14516 32662 14526 32714
rect 14550 32662 14580 32714
rect 14580 32662 14606 32714
rect 14310 32660 14366 32662
rect 14390 32660 14446 32662
rect 14470 32660 14526 32662
rect 14550 32660 14606 32662
rect 14310 31626 14366 31628
rect 14390 31626 14446 31628
rect 14470 31626 14526 31628
rect 14550 31626 14606 31628
rect 14310 31574 14336 31626
rect 14336 31574 14366 31626
rect 14390 31574 14400 31626
rect 14400 31574 14446 31626
rect 14470 31574 14516 31626
rect 14516 31574 14526 31626
rect 14550 31574 14580 31626
rect 14580 31574 14606 31626
rect 14310 31572 14366 31574
rect 14390 31572 14446 31574
rect 14470 31572 14526 31574
rect 14550 31572 14606 31574
rect 14310 30538 14366 30540
rect 14390 30538 14446 30540
rect 14470 30538 14526 30540
rect 14550 30538 14606 30540
rect 14310 30486 14336 30538
rect 14336 30486 14366 30538
rect 14390 30486 14400 30538
rect 14400 30486 14446 30538
rect 14470 30486 14516 30538
rect 14516 30486 14526 30538
rect 14550 30486 14580 30538
rect 14580 30486 14606 30538
rect 14310 30484 14366 30486
rect 14390 30484 14446 30486
rect 14470 30484 14526 30486
rect 14550 30484 14606 30486
rect 14310 29450 14366 29452
rect 14390 29450 14446 29452
rect 14470 29450 14526 29452
rect 14550 29450 14606 29452
rect 14310 29398 14336 29450
rect 14336 29398 14366 29450
rect 14390 29398 14400 29450
rect 14400 29398 14446 29450
rect 14470 29398 14516 29450
rect 14516 29398 14526 29450
rect 14550 29398 14580 29450
rect 14580 29398 14606 29450
rect 14310 29396 14366 29398
rect 14390 29396 14446 29398
rect 14470 29396 14526 29398
rect 14550 29396 14606 29398
rect 14310 28362 14366 28364
rect 14390 28362 14446 28364
rect 14470 28362 14526 28364
rect 14550 28362 14606 28364
rect 14310 28310 14336 28362
rect 14336 28310 14366 28362
rect 14390 28310 14400 28362
rect 14400 28310 14446 28362
rect 14470 28310 14516 28362
rect 14516 28310 14526 28362
rect 14550 28310 14580 28362
rect 14580 28310 14606 28362
rect 14310 28308 14366 28310
rect 14390 28308 14446 28310
rect 14470 28308 14526 28310
rect 14550 28308 14606 28310
rect 16974 41962 17030 41964
rect 17054 41962 17110 41964
rect 17134 41962 17190 41964
rect 17214 41962 17270 41964
rect 16974 41910 17000 41962
rect 17000 41910 17030 41962
rect 17054 41910 17064 41962
rect 17064 41910 17110 41962
rect 17134 41910 17180 41962
rect 17180 41910 17190 41962
rect 17214 41910 17244 41962
rect 17244 41910 17270 41962
rect 16974 41908 17030 41910
rect 17054 41908 17110 41910
rect 17134 41908 17190 41910
rect 17214 41908 17270 41910
rect 16974 40874 17030 40876
rect 17054 40874 17110 40876
rect 17134 40874 17190 40876
rect 17214 40874 17270 40876
rect 16974 40822 17000 40874
rect 17000 40822 17030 40874
rect 17054 40822 17064 40874
rect 17064 40822 17110 40874
rect 17134 40822 17180 40874
rect 17180 40822 17190 40874
rect 17214 40822 17244 40874
rect 17244 40822 17270 40874
rect 16974 40820 17030 40822
rect 17054 40820 17110 40822
rect 17134 40820 17190 40822
rect 17214 40820 17270 40822
rect 16380 37896 16436 37952
rect 12608 27580 12664 27616
rect 12608 27560 12610 27580
rect 12610 27560 12662 27580
rect 12662 27560 12664 27580
rect 16974 39786 17030 39788
rect 17054 39786 17110 39788
rect 17134 39786 17190 39788
rect 17214 39786 17270 39788
rect 16974 39734 17000 39786
rect 17000 39734 17030 39786
rect 17054 39734 17064 39786
rect 17064 39734 17110 39786
rect 17134 39734 17180 39786
rect 17180 39734 17190 39786
rect 17214 39734 17244 39786
rect 17244 39734 17270 39786
rect 16974 39732 17030 39734
rect 17054 39732 17110 39734
rect 17134 39732 17190 39734
rect 17214 39732 17270 39734
rect 16974 38698 17030 38700
rect 17054 38698 17110 38700
rect 17134 38698 17190 38700
rect 17214 38698 17270 38700
rect 16974 38646 17000 38698
rect 17000 38646 17030 38698
rect 17054 38646 17064 38698
rect 17064 38646 17110 38698
rect 17134 38646 17180 38698
rect 17180 38646 17190 38698
rect 17214 38646 17244 38698
rect 17244 38646 17270 38698
rect 16974 38644 17030 38646
rect 17054 38644 17110 38646
rect 17134 38644 17190 38646
rect 17214 38644 17270 38646
rect 16974 37610 17030 37612
rect 17054 37610 17110 37612
rect 17134 37610 17190 37612
rect 17214 37610 17270 37612
rect 16974 37558 17000 37610
rect 17000 37558 17030 37610
rect 17054 37558 17064 37610
rect 17064 37558 17110 37610
rect 17134 37558 17180 37610
rect 17180 37558 17190 37610
rect 17214 37558 17244 37610
rect 17244 37558 17270 37610
rect 16974 37556 17030 37558
rect 17054 37556 17110 37558
rect 17134 37556 17190 37558
rect 17214 37556 17270 37558
rect 16974 36522 17030 36524
rect 17054 36522 17110 36524
rect 17134 36522 17190 36524
rect 17214 36522 17270 36524
rect 16974 36470 17000 36522
rect 17000 36470 17030 36522
rect 17054 36470 17064 36522
rect 17064 36470 17110 36522
rect 17134 36470 17180 36522
rect 17180 36470 17190 36522
rect 17214 36470 17244 36522
rect 17244 36470 17270 36522
rect 16974 36468 17030 36470
rect 17054 36468 17110 36470
rect 17134 36468 17190 36470
rect 17214 36468 17270 36470
rect 16974 35434 17030 35436
rect 17054 35434 17110 35436
rect 17134 35434 17190 35436
rect 17214 35434 17270 35436
rect 16974 35382 17000 35434
rect 17000 35382 17030 35434
rect 17054 35382 17064 35434
rect 17064 35382 17110 35434
rect 17134 35382 17180 35434
rect 17180 35382 17190 35434
rect 17214 35382 17244 35434
rect 17244 35382 17270 35434
rect 16974 35380 17030 35382
rect 17054 35380 17110 35382
rect 17134 35380 17190 35382
rect 17214 35380 17270 35382
rect 19638 41418 19694 41420
rect 19718 41418 19774 41420
rect 19798 41418 19854 41420
rect 19878 41418 19934 41420
rect 19638 41366 19664 41418
rect 19664 41366 19694 41418
rect 19718 41366 19728 41418
rect 19728 41366 19774 41418
rect 19798 41366 19844 41418
rect 19844 41366 19854 41418
rect 19878 41366 19908 41418
rect 19908 41366 19934 41418
rect 19638 41364 19694 41366
rect 19718 41364 19774 41366
rect 19798 41364 19854 41366
rect 19878 41364 19934 41366
rect 19638 40330 19694 40332
rect 19718 40330 19774 40332
rect 19798 40330 19854 40332
rect 19878 40330 19934 40332
rect 19638 40278 19664 40330
rect 19664 40278 19694 40330
rect 19718 40278 19728 40330
rect 19728 40278 19774 40330
rect 19798 40278 19844 40330
rect 19844 40278 19854 40330
rect 19878 40278 19908 40330
rect 19908 40278 19934 40330
rect 19638 40276 19694 40278
rect 19718 40276 19774 40278
rect 19798 40276 19854 40278
rect 19878 40276 19934 40278
rect 16974 34346 17030 34348
rect 17054 34346 17110 34348
rect 17134 34346 17190 34348
rect 17214 34346 17270 34348
rect 16974 34294 17000 34346
rect 17000 34294 17030 34346
rect 17054 34294 17064 34346
rect 17064 34294 17110 34346
rect 17134 34294 17180 34346
rect 17180 34294 17190 34346
rect 17214 34294 17244 34346
rect 17244 34294 17270 34346
rect 16974 34292 17030 34294
rect 17054 34292 17110 34294
rect 17134 34292 17190 34294
rect 17214 34292 17270 34294
rect 16974 33258 17030 33260
rect 17054 33258 17110 33260
rect 17134 33258 17190 33260
rect 17214 33258 17270 33260
rect 16974 33206 17000 33258
rect 17000 33206 17030 33258
rect 17054 33206 17064 33258
rect 17064 33206 17110 33258
rect 17134 33206 17180 33258
rect 17180 33206 17190 33258
rect 17214 33206 17244 33258
rect 17244 33206 17270 33258
rect 16974 33204 17030 33206
rect 17054 33204 17110 33206
rect 17134 33204 17190 33206
rect 17214 33204 17270 33206
rect 16974 32170 17030 32172
rect 17054 32170 17110 32172
rect 17134 32170 17190 32172
rect 17214 32170 17270 32172
rect 16974 32118 17000 32170
rect 17000 32118 17030 32170
rect 17054 32118 17064 32170
rect 17064 32118 17110 32170
rect 17134 32118 17180 32170
rect 17180 32118 17190 32170
rect 17214 32118 17244 32170
rect 17244 32118 17270 32170
rect 16974 32116 17030 32118
rect 17054 32116 17110 32118
rect 17134 32116 17190 32118
rect 17214 32116 17270 32118
rect 17300 31812 17302 31832
rect 17302 31812 17354 31832
rect 17354 31812 17356 31832
rect 17300 31776 17356 31812
rect 16974 31082 17030 31084
rect 17054 31082 17110 31084
rect 17134 31082 17190 31084
rect 17214 31082 17270 31084
rect 16974 31030 17000 31082
rect 17000 31030 17030 31082
rect 17054 31030 17064 31082
rect 17064 31030 17110 31082
rect 17134 31030 17180 31082
rect 17180 31030 17190 31082
rect 17214 31030 17244 31082
rect 17244 31030 17270 31082
rect 16974 31028 17030 31030
rect 17054 31028 17110 31030
rect 17134 31028 17190 31030
rect 17214 31028 17270 31030
rect 16748 30844 16804 30880
rect 16748 30824 16750 30844
rect 16750 30824 16802 30844
rect 16802 30824 16804 30844
rect 16974 29994 17030 29996
rect 17054 29994 17110 29996
rect 17134 29994 17190 29996
rect 17214 29994 17270 29996
rect 16974 29942 17000 29994
rect 17000 29942 17030 29994
rect 17054 29942 17064 29994
rect 17064 29942 17110 29994
rect 17134 29942 17180 29994
rect 17180 29942 17190 29994
rect 17214 29942 17244 29994
rect 17244 29942 17270 29994
rect 16974 29940 17030 29942
rect 17054 29940 17110 29942
rect 17134 29940 17190 29942
rect 17214 29940 17270 29942
rect 16974 28906 17030 28908
rect 17054 28906 17110 28908
rect 17134 28906 17190 28908
rect 17214 28906 17270 28908
rect 16974 28854 17000 28906
rect 17000 28854 17030 28906
rect 17054 28854 17064 28906
rect 17064 28854 17110 28906
rect 17134 28854 17180 28906
rect 17180 28854 17190 28906
rect 17214 28854 17244 28906
rect 17244 28854 17270 28906
rect 16974 28852 17030 28854
rect 17054 28852 17110 28854
rect 17134 28852 17190 28854
rect 17214 28852 17270 28854
rect 17760 30824 17816 30880
rect 14310 27274 14366 27276
rect 14390 27274 14446 27276
rect 14470 27274 14526 27276
rect 14550 27274 14606 27276
rect 14310 27222 14336 27274
rect 14336 27222 14366 27274
rect 14390 27222 14400 27274
rect 14400 27222 14446 27274
rect 14470 27222 14516 27274
rect 14516 27222 14526 27274
rect 14550 27222 14580 27274
rect 14580 27222 14606 27274
rect 14310 27220 14366 27222
rect 14390 27220 14446 27222
rect 14470 27220 14526 27222
rect 14550 27220 14606 27222
rect 11646 26730 11702 26732
rect 11726 26730 11782 26732
rect 11806 26730 11862 26732
rect 11886 26730 11942 26732
rect 11646 26678 11672 26730
rect 11672 26678 11702 26730
rect 11726 26678 11736 26730
rect 11736 26678 11782 26730
rect 11806 26678 11852 26730
rect 11852 26678 11862 26730
rect 11886 26678 11916 26730
rect 11916 26678 11942 26730
rect 11646 26676 11702 26678
rect 11726 26676 11782 26678
rect 11806 26676 11862 26678
rect 11886 26676 11942 26678
rect 16564 27424 16620 27480
rect 16974 27818 17030 27820
rect 17054 27818 17110 27820
rect 17134 27818 17190 27820
rect 17214 27818 17270 27820
rect 16974 27766 17000 27818
rect 17000 27766 17030 27818
rect 17054 27766 17064 27818
rect 17064 27766 17110 27818
rect 17134 27766 17180 27818
rect 17180 27766 17190 27818
rect 17214 27766 17244 27818
rect 17244 27766 17270 27818
rect 16974 27764 17030 27766
rect 17054 27764 17110 27766
rect 17134 27764 17190 27766
rect 17214 27764 17270 27766
rect 19638 39242 19694 39244
rect 19718 39242 19774 39244
rect 19798 39242 19854 39244
rect 19878 39242 19934 39244
rect 19638 39190 19664 39242
rect 19664 39190 19694 39242
rect 19718 39190 19728 39242
rect 19728 39190 19774 39242
rect 19798 39190 19844 39242
rect 19844 39190 19854 39242
rect 19878 39190 19908 39242
rect 19908 39190 19934 39242
rect 19638 39188 19694 39190
rect 19718 39188 19774 39190
rect 19798 39188 19854 39190
rect 19878 39188 19934 39190
rect 18496 33000 18552 33056
rect 18956 31932 19012 31968
rect 18956 31912 18958 31932
rect 18958 31912 19010 31932
rect 19010 31912 19012 31932
rect 17116 27560 17172 27616
rect 18864 28004 18866 28024
rect 18866 28004 18918 28024
rect 18918 28004 18920 28024
rect 18864 27968 18920 28004
rect 19638 38154 19694 38156
rect 19718 38154 19774 38156
rect 19798 38154 19854 38156
rect 19878 38154 19934 38156
rect 19638 38102 19664 38154
rect 19664 38102 19694 38154
rect 19718 38102 19728 38154
rect 19728 38102 19774 38154
rect 19798 38102 19844 38154
rect 19844 38102 19854 38154
rect 19878 38102 19908 38154
rect 19908 38102 19934 38154
rect 19638 38100 19694 38102
rect 19718 38100 19774 38102
rect 19798 38100 19854 38102
rect 19878 38100 19934 38102
rect 19638 37066 19694 37068
rect 19718 37066 19774 37068
rect 19798 37066 19854 37068
rect 19878 37066 19934 37068
rect 19638 37014 19664 37066
rect 19664 37014 19694 37066
rect 19718 37014 19728 37066
rect 19728 37014 19774 37066
rect 19798 37014 19844 37066
rect 19844 37014 19854 37066
rect 19878 37014 19908 37066
rect 19908 37014 19934 37066
rect 19638 37012 19694 37014
rect 19718 37012 19774 37014
rect 19798 37012 19854 37014
rect 19878 37012 19934 37014
rect 19638 35978 19694 35980
rect 19718 35978 19774 35980
rect 19798 35978 19854 35980
rect 19878 35978 19934 35980
rect 19638 35926 19664 35978
rect 19664 35926 19694 35978
rect 19718 35926 19728 35978
rect 19728 35926 19774 35978
rect 19798 35926 19844 35978
rect 19844 35926 19854 35978
rect 19878 35926 19908 35978
rect 19908 35926 19934 35978
rect 19638 35924 19694 35926
rect 19718 35924 19774 35926
rect 19798 35924 19854 35926
rect 19878 35924 19934 35926
rect 19638 34890 19694 34892
rect 19718 34890 19774 34892
rect 19798 34890 19854 34892
rect 19878 34890 19934 34892
rect 19638 34838 19664 34890
rect 19664 34838 19694 34890
rect 19718 34838 19728 34890
rect 19728 34838 19774 34890
rect 19798 34838 19844 34890
rect 19844 34838 19854 34890
rect 19878 34838 19908 34890
rect 19908 34838 19934 34890
rect 19638 34836 19694 34838
rect 19718 34836 19774 34838
rect 19798 34836 19854 34838
rect 19878 34836 19934 34838
rect 19638 33802 19694 33804
rect 19718 33802 19774 33804
rect 19798 33802 19854 33804
rect 19878 33802 19934 33804
rect 19638 33750 19664 33802
rect 19664 33750 19694 33802
rect 19718 33750 19728 33802
rect 19728 33750 19774 33802
rect 19798 33750 19844 33802
rect 19844 33750 19854 33802
rect 19878 33750 19908 33802
rect 19908 33750 19934 33802
rect 19638 33748 19694 33750
rect 19718 33748 19774 33750
rect 19798 33748 19854 33750
rect 19878 33748 19934 33750
rect 19638 32714 19694 32716
rect 19718 32714 19774 32716
rect 19798 32714 19854 32716
rect 19878 32714 19934 32716
rect 19638 32662 19664 32714
rect 19664 32662 19694 32714
rect 19718 32662 19728 32714
rect 19728 32662 19774 32714
rect 19798 32662 19844 32714
rect 19844 32662 19854 32714
rect 19878 32662 19908 32714
rect 19908 32662 19934 32714
rect 19638 32660 19694 32662
rect 19718 32660 19774 32662
rect 19798 32660 19854 32662
rect 19878 32660 19934 32662
rect 19416 31812 19418 31832
rect 19418 31812 19470 31832
rect 19470 31812 19472 31832
rect 19416 31776 19472 31812
rect 19638 31626 19694 31628
rect 19718 31626 19774 31628
rect 19798 31626 19854 31628
rect 19878 31626 19934 31628
rect 19638 31574 19664 31626
rect 19664 31574 19694 31626
rect 19718 31574 19728 31626
rect 19728 31574 19774 31626
rect 19798 31574 19844 31626
rect 19844 31574 19854 31626
rect 19878 31574 19908 31626
rect 19908 31574 19934 31626
rect 19638 31572 19694 31574
rect 19718 31572 19774 31574
rect 19798 31572 19854 31574
rect 19878 31572 19934 31574
rect 22302 41962 22358 41964
rect 22382 41962 22438 41964
rect 22462 41962 22518 41964
rect 22542 41962 22598 41964
rect 22302 41910 22328 41962
rect 22328 41910 22358 41962
rect 22382 41910 22392 41962
rect 22392 41910 22438 41962
rect 22462 41910 22508 41962
rect 22508 41910 22518 41962
rect 22542 41910 22572 41962
rect 22572 41910 22598 41962
rect 22302 41908 22358 41910
rect 22382 41908 22438 41910
rect 22462 41908 22518 41910
rect 22542 41908 22598 41910
rect 22302 40874 22358 40876
rect 22382 40874 22438 40876
rect 22462 40874 22518 40876
rect 22542 40874 22598 40876
rect 22302 40822 22328 40874
rect 22328 40822 22358 40874
rect 22382 40822 22392 40874
rect 22392 40822 22438 40874
rect 22462 40822 22508 40874
rect 22508 40822 22518 40874
rect 22542 40822 22572 40874
rect 22572 40822 22598 40874
rect 22302 40820 22358 40822
rect 22382 40820 22438 40822
rect 22462 40820 22518 40822
rect 22542 40820 22598 40822
rect 22302 39786 22358 39788
rect 22382 39786 22438 39788
rect 22462 39786 22518 39788
rect 22542 39786 22598 39788
rect 22302 39734 22328 39786
rect 22328 39734 22358 39786
rect 22382 39734 22392 39786
rect 22392 39734 22438 39786
rect 22462 39734 22508 39786
rect 22508 39734 22518 39786
rect 22542 39734 22572 39786
rect 22572 39734 22598 39786
rect 22302 39732 22358 39734
rect 22382 39732 22438 39734
rect 22462 39732 22518 39734
rect 22542 39732 22598 39734
rect 22302 38698 22358 38700
rect 22382 38698 22438 38700
rect 22462 38698 22518 38700
rect 22542 38698 22598 38700
rect 22302 38646 22328 38698
rect 22328 38646 22358 38698
rect 22382 38646 22392 38698
rect 22392 38646 22438 38698
rect 22462 38646 22508 38698
rect 22508 38646 22518 38698
rect 22542 38646 22572 38698
rect 22572 38646 22598 38698
rect 22302 38644 22358 38646
rect 22382 38644 22438 38646
rect 22462 38644 22518 38646
rect 22542 38644 22598 38646
rect 22302 37610 22358 37612
rect 22382 37610 22438 37612
rect 22462 37610 22518 37612
rect 22542 37610 22598 37612
rect 22302 37558 22328 37610
rect 22328 37558 22358 37610
rect 22382 37558 22392 37610
rect 22392 37558 22438 37610
rect 22462 37558 22508 37610
rect 22508 37558 22518 37610
rect 22542 37558 22572 37610
rect 22572 37558 22598 37610
rect 22302 37556 22358 37558
rect 22382 37556 22438 37558
rect 22462 37556 22518 37558
rect 22542 37556 22598 37558
rect 22302 36522 22358 36524
rect 22382 36522 22438 36524
rect 22462 36522 22518 36524
rect 22542 36522 22598 36524
rect 22302 36470 22328 36522
rect 22328 36470 22358 36522
rect 22382 36470 22392 36522
rect 22392 36470 22438 36522
rect 22462 36470 22508 36522
rect 22508 36470 22518 36522
rect 22542 36470 22572 36522
rect 22572 36470 22598 36522
rect 22302 36468 22358 36470
rect 22382 36468 22438 36470
rect 22462 36468 22518 36470
rect 22542 36468 22598 36470
rect 22302 35434 22358 35436
rect 22382 35434 22438 35436
rect 22462 35434 22518 35436
rect 22542 35434 22598 35436
rect 22302 35382 22328 35434
rect 22328 35382 22358 35434
rect 22382 35382 22392 35434
rect 22392 35382 22438 35434
rect 22462 35382 22508 35434
rect 22508 35382 22518 35434
rect 22542 35382 22572 35434
rect 22572 35382 22598 35434
rect 22302 35380 22358 35382
rect 22382 35380 22438 35382
rect 22462 35380 22518 35382
rect 22542 35380 22598 35382
rect 22302 34346 22358 34348
rect 22382 34346 22438 34348
rect 22462 34346 22518 34348
rect 22542 34346 22598 34348
rect 22302 34294 22328 34346
rect 22328 34294 22358 34346
rect 22382 34294 22392 34346
rect 22392 34294 22438 34346
rect 22462 34294 22508 34346
rect 22508 34294 22518 34346
rect 22542 34294 22572 34346
rect 22572 34294 22598 34346
rect 22302 34292 22358 34294
rect 22382 34292 22438 34294
rect 22462 34292 22518 34294
rect 22542 34292 22598 34294
rect 22302 33258 22358 33260
rect 22382 33258 22438 33260
rect 22462 33258 22518 33260
rect 22542 33258 22598 33260
rect 22302 33206 22328 33258
rect 22328 33206 22358 33258
rect 22382 33206 22392 33258
rect 22392 33206 22438 33258
rect 22462 33206 22508 33258
rect 22508 33206 22518 33258
rect 22542 33206 22572 33258
rect 22572 33206 22598 33258
rect 22302 33204 22358 33206
rect 22382 33204 22438 33206
rect 22462 33204 22518 33206
rect 22542 33204 22598 33206
rect 19638 30538 19694 30540
rect 19718 30538 19774 30540
rect 19798 30538 19854 30540
rect 19878 30538 19934 30540
rect 19638 30486 19664 30538
rect 19664 30486 19694 30538
rect 19718 30486 19728 30538
rect 19728 30486 19774 30538
rect 19798 30486 19844 30538
rect 19844 30486 19854 30538
rect 19878 30486 19908 30538
rect 19908 30486 19934 30538
rect 19638 30484 19694 30486
rect 19718 30484 19774 30486
rect 19798 30484 19854 30486
rect 19878 30484 19934 30486
rect 19600 30300 19656 30336
rect 19600 30280 19602 30300
rect 19602 30280 19654 30300
rect 19654 30280 19656 30300
rect 19638 29450 19694 29452
rect 19718 29450 19774 29452
rect 19798 29450 19854 29452
rect 19878 29450 19934 29452
rect 19638 29398 19664 29450
rect 19664 29398 19694 29450
rect 19718 29398 19728 29450
rect 19728 29398 19774 29450
rect 19798 29398 19844 29450
rect 19844 29398 19854 29450
rect 19878 29398 19908 29450
rect 19908 29398 19934 29450
rect 19638 29396 19694 29398
rect 19718 29396 19774 29398
rect 19798 29396 19854 29398
rect 19878 29396 19934 29398
rect 19638 28362 19694 28364
rect 19718 28362 19774 28364
rect 19798 28362 19854 28364
rect 19878 28362 19934 28364
rect 19638 28310 19664 28362
rect 19664 28310 19694 28362
rect 19718 28310 19728 28362
rect 19728 28310 19774 28362
rect 19798 28310 19844 28362
rect 19844 28310 19854 28362
rect 19878 28310 19908 28362
rect 19908 28310 19934 28362
rect 19638 28308 19694 28310
rect 19718 28308 19774 28310
rect 19798 28308 19854 28310
rect 19878 28308 19934 28310
rect 22302 32170 22358 32172
rect 22382 32170 22438 32172
rect 22462 32170 22518 32172
rect 22542 32170 22598 32172
rect 22302 32118 22328 32170
rect 22328 32118 22358 32170
rect 22382 32118 22392 32170
rect 22392 32118 22438 32170
rect 22462 32118 22508 32170
rect 22508 32118 22518 32170
rect 22542 32118 22572 32170
rect 22572 32118 22598 32170
rect 22302 32116 22358 32118
rect 22382 32116 22438 32118
rect 22462 32116 22518 32118
rect 22542 32116 22598 32118
rect 22302 31082 22358 31084
rect 22382 31082 22438 31084
rect 22462 31082 22518 31084
rect 22542 31082 22598 31084
rect 22302 31030 22328 31082
rect 22328 31030 22358 31082
rect 22382 31030 22392 31082
rect 22392 31030 22438 31082
rect 22462 31030 22508 31082
rect 22508 31030 22518 31082
rect 22542 31030 22572 31082
rect 22572 31030 22598 31082
rect 22302 31028 22358 31030
rect 22382 31028 22438 31030
rect 22462 31028 22518 31030
rect 22542 31028 22598 31030
rect 22302 29994 22358 29996
rect 22382 29994 22438 29996
rect 22462 29994 22518 29996
rect 22542 29994 22598 29996
rect 22302 29942 22328 29994
rect 22328 29942 22358 29994
rect 22382 29942 22392 29994
rect 22392 29942 22438 29994
rect 22462 29942 22508 29994
rect 22508 29942 22518 29994
rect 22542 29942 22572 29994
rect 22572 29942 22598 29994
rect 22302 29940 22358 29942
rect 22382 29940 22438 29942
rect 22462 29940 22518 29942
rect 22542 29940 22598 29942
rect 22728 29892 22784 29928
rect 22728 29872 22730 29892
rect 22730 29872 22782 29892
rect 22782 29872 22784 29892
rect 22302 28906 22358 28908
rect 22382 28906 22438 28908
rect 22462 28906 22518 28908
rect 22542 28906 22598 28908
rect 22302 28854 22328 28906
rect 22328 28854 22358 28906
rect 22382 28854 22392 28906
rect 22392 28854 22438 28906
rect 22462 28854 22508 28906
rect 22508 28854 22518 28906
rect 22542 28854 22572 28906
rect 22572 28854 22598 28906
rect 22302 28852 22358 28854
rect 22382 28852 22438 28854
rect 22462 28852 22518 28854
rect 22542 28852 22598 28854
rect 22820 28512 22876 28568
rect 22302 27818 22358 27820
rect 22382 27818 22438 27820
rect 22462 27818 22518 27820
rect 22542 27818 22598 27820
rect 22302 27766 22328 27818
rect 22328 27766 22358 27818
rect 22382 27766 22392 27818
rect 22392 27766 22438 27818
rect 22462 27766 22508 27818
rect 22508 27766 22518 27818
rect 22542 27766 22572 27818
rect 22572 27766 22598 27818
rect 22302 27764 22358 27766
rect 22382 27764 22438 27766
rect 22462 27764 22518 27766
rect 22542 27764 22598 27766
rect 19638 27274 19694 27276
rect 19718 27274 19774 27276
rect 19798 27274 19854 27276
rect 19878 27274 19934 27276
rect 19638 27222 19664 27274
rect 19664 27222 19694 27274
rect 19718 27222 19728 27274
rect 19728 27222 19774 27274
rect 19798 27222 19844 27274
rect 19844 27222 19854 27274
rect 19878 27222 19908 27274
rect 19908 27222 19934 27274
rect 19638 27220 19694 27222
rect 19718 27220 19774 27222
rect 19798 27220 19854 27222
rect 19878 27220 19934 27222
rect 24966 41418 25022 41420
rect 25046 41418 25102 41420
rect 25126 41418 25182 41420
rect 25206 41418 25262 41420
rect 24966 41366 24992 41418
rect 24992 41366 25022 41418
rect 25046 41366 25056 41418
rect 25056 41366 25102 41418
rect 25126 41366 25172 41418
rect 25172 41366 25182 41418
rect 25206 41366 25236 41418
rect 25236 41366 25262 41418
rect 24966 41364 25022 41366
rect 25046 41364 25102 41366
rect 25126 41364 25182 41366
rect 25206 41364 25262 41366
rect 24966 40330 25022 40332
rect 25046 40330 25102 40332
rect 25126 40330 25182 40332
rect 25206 40330 25262 40332
rect 24966 40278 24992 40330
rect 24992 40278 25022 40330
rect 25046 40278 25056 40330
rect 25056 40278 25102 40330
rect 25126 40278 25172 40330
rect 25172 40278 25182 40330
rect 25206 40278 25236 40330
rect 25236 40278 25262 40330
rect 24966 40276 25022 40278
rect 25046 40276 25102 40278
rect 25126 40276 25182 40278
rect 25206 40276 25262 40278
rect 27630 41962 27686 41964
rect 27710 41962 27766 41964
rect 27790 41962 27846 41964
rect 27870 41962 27926 41964
rect 27630 41910 27656 41962
rect 27656 41910 27686 41962
rect 27710 41910 27720 41962
rect 27720 41910 27766 41962
rect 27790 41910 27836 41962
rect 27836 41910 27846 41962
rect 27870 41910 27900 41962
rect 27900 41910 27926 41962
rect 27630 41908 27686 41910
rect 27710 41908 27766 41910
rect 27790 41908 27846 41910
rect 27870 41908 27926 41910
rect 27630 40874 27686 40876
rect 27710 40874 27766 40876
rect 27790 40874 27846 40876
rect 27870 40874 27926 40876
rect 27630 40822 27656 40874
rect 27656 40822 27686 40874
rect 27710 40822 27720 40874
rect 27720 40822 27766 40874
rect 27790 40822 27836 40874
rect 27836 40822 27846 40874
rect 27870 40822 27900 40874
rect 27900 40822 27926 40874
rect 27630 40820 27686 40822
rect 27710 40820 27766 40822
rect 27790 40820 27846 40822
rect 27870 40820 27926 40822
rect 24016 31912 24072 31968
rect 23832 28668 23888 28704
rect 23832 28648 23834 28668
rect 23834 28648 23886 28668
rect 23886 28648 23888 28668
rect 23740 27424 23796 27480
rect 16974 26730 17030 26732
rect 17054 26730 17110 26732
rect 17134 26730 17190 26732
rect 17214 26730 17270 26732
rect 16974 26678 17000 26730
rect 17000 26678 17030 26730
rect 17054 26678 17064 26730
rect 17064 26678 17110 26730
rect 17134 26678 17180 26730
rect 17180 26678 17190 26730
rect 17214 26678 17244 26730
rect 17244 26678 17270 26730
rect 16974 26676 17030 26678
rect 17054 26676 17110 26678
rect 17134 26676 17190 26678
rect 17214 26676 17270 26678
rect 22302 26730 22358 26732
rect 22382 26730 22438 26732
rect 22462 26730 22518 26732
rect 22542 26730 22598 26732
rect 22302 26678 22328 26730
rect 22328 26678 22358 26730
rect 22382 26678 22392 26730
rect 22392 26678 22438 26730
rect 22462 26678 22508 26730
rect 22508 26678 22518 26730
rect 22542 26678 22572 26730
rect 22572 26678 22598 26730
rect 22302 26676 22358 26678
rect 22382 26676 22438 26678
rect 22462 26676 22518 26678
rect 22542 26676 22598 26678
rect 24966 39242 25022 39244
rect 25046 39242 25102 39244
rect 25126 39242 25182 39244
rect 25206 39242 25262 39244
rect 24966 39190 24992 39242
rect 24992 39190 25022 39242
rect 25046 39190 25056 39242
rect 25056 39190 25102 39242
rect 25126 39190 25172 39242
rect 25172 39190 25182 39242
rect 25206 39190 25236 39242
rect 25236 39190 25262 39242
rect 24966 39188 25022 39190
rect 25046 39188 25102 39190
rect 25126 39188 25182 39190
rect 25206 39188 25262 39190
rect 24966 38154 25022 38156
rect 25046 38154 25102 38156
rect 25126 38154 25182 38156
rect 25206 38154 25262 38156
rect 24966 38102 24992 38154
rect 24992 38102 25022 38154
rect 25046 38102 25056 38154
rect 25056 38102 25102 38154
rect 25126 38102 25172 38154
rect 25172 38102 25182 38154
rect 25206 38102 25236 38154
rect 25236 38102 25262 38154
rect 24966 38100 25022 38102
rect 25046 38100 25102 38102
rect 25126 38100 25182 38102
rect 25206 38100 25262 38102
rect 25580 37796 25582 37816
rect 25582 37796 25634 37816
rect 25634 37796 25636 37816
rect 25580 37760 25636 37796
rect 24966 37066 25022 37068
rect 25046 37066 25102 37068
rect 25126 37066 25182 37068
rect 25206 37066 25262 37068
rect 24966 37014 24992 37066
rect 24992 37014 25022 37066
rect 25046 37014 25056 37066
rect 25056 37014 25102 37066
rect 25126 37014 25172 37066
rect 25172 37014 25182 37066
rect 25206 37014 25236 37066
rect 25236 37014 25262 37066
rect 24966 37012 25022 37014
rect 25046 37012 25102 37014
rect 25126 37012 25182 37014
rect 25206 37012 25262 37014
rect 24966 35978 25022 35980
rect 25046 35978 25102 35980
rect 25126 35978 25182 35980
rect 25206 35978 25262 35980
rect 24966 35926 24992 35978
rect 24992 35926 25022 35978
rect 25046 35926 25056 35978
rect 25056 35926 25102 35978
rect 25126 35926 25172 35978
rect 25172 35926 25182 35978
rect 25206 35926 25236 35978
rect 25236 35926 25262 35978
rect 24966 35924 25022 35926
rect 25046 35924 25102 35926
rect 25126 35924 25182 35926
rect 25206 35924 25262 35926
rect 24966 34890 25022 34892
rect 25046 34890 25102 34892
rect 25126 34890 25182 34892
rect 25206 34890 25262 34892
rect 24966 34838 24992 34890
rect 24992 34838 25022 34890
rect 25046 34838 25056 34890
rect 25056 34838 25102 34890
rect 25126 34838 25172 34890
rect 25172 34838 25182 34890
rect 25206 34838 25236 34890
rect 25236 34838 25262 34890
rect 24966 34836 25022 34838
rect 25046 34836 25102 34838
rect 25126 34836 25182 34838
rect 25206 34836 25262 34838
rect 24966 33802 25022 33804
rect 25046 33802 25102 33804
rect 25126 33802 25182 33804
rect 25206 33802 25262 33804
rect 24966 33750 24992 33802
rect 24992 33750 25022 33802
rect 25046 33750 25056 33802
rect 25056 33750 25102 33802
rect 25126 33750 25172 33802
rect 25172 33750 25182 33802
rect 25206 33750 25236 33802
rect 25236 33750 25262 33802
rect 24966 33748 25022 33750
rect 25046 33748 25102 33750
rect 25126 33748 25182 33750
rect 25206 33748 25262 33750
rect 24966 32714 25022 32716
rect 25046 32714 25102 32716
rect 25126 32714 25182 32716
rect 25206 32714 25262 32716
rect 24966 32662 24992 32714
rect 24992 32662 25022 32714
rect 25046 32662 25056 32714
rect 25056 32662 25102 32714
rect 25126 32662 25172 32714
rect 25172 32662 25182 32714
rect 25206 32662 25236 32714
rect 25236 32662 25262 32714
rect 24966 32660 25022 32662
rect 25046 32660 25102 32662
rect 25126 32660 25182 32662
rect 25206 32660 25262 32662
rect 26868 33972 26924 34008
rect 26868 33952 26870 33972
rect 26870 33952 26922 33972
rect 26922 33952 26924 33972
rect 24966 31626 25022 31628
rect 25046 31626 25102 31628
rect 25126 31626 25182 31628
rect 25206 31626 25262 31628
rect 24966 31574 24992 31626
rect 24992 31574 25022 31626
rect 25046 31574 25056 31626
rect 25056 31574 25102 31626
rect 25126 31574 25172 31626
rect 25172 31574 25182 31626
rect 25206 31574 25236 31626
rect 25236 31574 25262 31626
rect 24966 31572 25022 31574
rect 25046 31572 25102 31574
rect 25126 31572 25182 31574
rect 25206 31572 25262 31574
rect 24966 30538 25022 30540
rect 25046 30538 25102 30540
rect 25126 30538 25182 30540
rect 25206 30538 25262 30540
rect 24966 30486 24992 30538
rect 24992 30486 25022 30538
rect 25046 30486 25056 30538
rect 25056 30486 25102 30538
rect 25126 30486 25172 30538
rect 25172 30486 25182 30538
rect 25206 30486 25236 30538
rect 25236 30486 25262 30538
rect 24966 30484 25022 30486
rect 25046 30484 25102 30486
rect 25126 30484 25182 30486
rect 25206 30484 25262 30486
rect 24966 29450 25022 29452
rect 25046 29450 25102 29452
rect 25126 29450 25182 29452
rect 25206 29450 25262 29452
rect 24966 29398 24992 29450
rect 24992 29398 25022 29450
rect 25046 29398 25056 29450
rect 25056 29398 25102 29450
rect 25126 29398 25172 29450
rect 25172 29398 25182 29450
rect 25206 29398 25236 29450
rect 25236 29398 25262 29450
rect 24966 29396 25022 29398
rect 25046 29396 25102 29398
rect 25126 29396 25182 29398
rect 25206 29396 25262 29398
rect 27630 39786 27686 39788
rect 27710 39786 27766 39788
rect 27790 39786 27846 39788
rect 27870 39786 27926 39788
rect 27630 39734 27656 39786
rect 27656 39734 27686 39786
rect 27710 39734 27720 39786
rect 27720 39734 27766 39786
rect 27790 39734 27836 39786
rect 27836 39734 27846 39786
rect 27870 39734 27900 39786
rect 27900 39734 27926 39786
rect 27630 39732 27686 39734
rect 27710 39732 27766 39734
rect 27790 39732 27846 39734
rect 27870 39732 27926 39734
rect 27630 38698 27686 38700
rect 27710 38698 27766 38700
rect 27790 38698 27846 38700
rect 27870 38698 27926 38700
rect 27630 38646 27656 38698
rect 27656 38646 27686 38698
rect 27710 38646 27720 38698
rect 27720 38646 27766 38698
rect 27790 38646 27836 38698
rect 27836 38646 27846 38698
rect 27870 38646 27900 38698
rect 27900 38646 27926 38698
rect 27630 38644 27686 38646
rect 27710 38644 27766 38646
rect 27790 38644 27846 38646
rect 27870 38644 27926 38646
rect 27630 37610 27686 37612
rect 27710 37610 27766 37612
rect 27790 37610 27846 37612
rect 27870 37610 27926 37612
rect 27630 37558 27656 37610
rect 27656 37558 27686 37610
rect 27710 37558 27720 37610
rect 27720 37558 27766 37610
rect 27790 37558 27836 37610
rect 27836 37558 27846 37610
rect 27870 37558 27900 37610
rect 27900 37558 27926 37610
rect 27630 37556 27686 37558
rect 27710 37556 27766 37558
rect 27790 37556 27846 37558
rect 27870 37556 27926 37558
rect 27630 36522 27686 36524
rect 27710 36522 27766 36524
rect 27790 36522 27846 36524
rect 27870 36522 27926 36524
rect 27630 36470 27656 36522
rect 27656 36470 27686 36522
rect 27710 36470 27720 36522
rect 27720 36470 27766 36522
rect 27790 36470 27836 36522
rect 27836 36470 27846 36522
rect 27870 36470 27900 36522
rect 27900 36470 27926 36522
rect 27630 36468 27686 36470
rect 27710 36468 27766 36470
rect 27790 36468 27846 36470
rect 27870 36468 27926 36470
rect 27630 35434 27686 35436
rect 27710 35434 27766 35436
rect 27790 35434 27846 35436
rect 27870 35434 27926 35436
rect 27630 35382 27656 35434
rect 27656 35382 27686 35434
rect 27710 35382 27720 35434
rect 27720 35382 27766 35434
rect 27790 35382 27836 35434
rect 27836 35382 27846 35434
rect 27870 35382 27900 35434
rect 27900 35382 27926 35434
rect 27630 35380 27686 35382
rect 27710 35380 27766 35382
rect 27790 35380 27846 35382
rect 27870 35380 27926 35382
rect 27630 34346 27686 34348
rect 27710 34346 27766 34348
rect 27790 34346 27846 34348
rect 27870 34346 27926 34348
rect 27630 34294 27656 34346
rect 27656 34294 27686 34346
rect 27710 34294 27720 34346
rect 27720 34294 27766 34346
rect 27790 34294 27836 34346
rect 27836 34294 27846 34346
rect 27870 34294 27900 34346
rect 27900 34294 27926 34346
rect 27630 34292 27686 34294
rect 27710 34292 27766 34294
rect 27790 34292 27846 34294
rect 27870 34292 27926 34294
rect 27630 33258 27686 33260
rect 27710 33258 27766 33260
rect 27790 33258 27846 33260
rect 27870 33258 27926 33260
rect 27630 33206 27656 33258
rect 27656 33206 27686 33258
rect 27710 33206 27720 33258
rect 27720 33206 27766 33258
rect 27790 33206 27836 33258
rect 27836 33206 27846 33258
rect 27870 33206 27900 33258
rect 27900 33206 27926 33258
rect 27630 33204 27686 33206
rect 27710 33204 27766 33206
rect 27790 33204 27846 33206
rect 27870 33204 27926 33206
rect 27630 32170 27686 32172
rect 27710 32170 27766 32172
rect 27790 32170 27846 32172
rect 27870 32170 27926 32172
rect 27630 32118 27656 32170
rect 27656 32118 27686 32170
rect 27710 32118 27720 32170
rect 27720 32118 27766 32170
rect 27790 32118 27836 32170
rect 27836 32118 27846 32170
rect 27870 32118 27900 32170
rect 27900 32118 27926 32170
rect 27630 32116 27686 32118
rect 27710 32116 27766 32118
rect 27790 32116 27846 32118
rect 27870 32116 27926 32118
rect 30294 41418 30350 41420
rect 30374 41418 30430 41420
rect 30454 41418 30510 41420
rect 30534 41418 30590 41420
rect 30294 41366 30320 41418
rect 30320 41366 30350 41418
rect 30374 41366 30384 41418
rect 30384 41366 30430 41418
rect 30454 41366 30500 41418
rect 30500 41366 30510 41418
rect 30534 41366 30564 41418
rect 30564 41366 30590 41418
rect 30294 41364 30350 41366
rect 30374 41364 30430 41366
rect 30454 41364 30510 41366
rect 30534 41364 30590 41366
rect 30294 40330 30350 40332
rect 30374 40330 30430 40332
rect 30454 40330 30510 40332
rect 30534 40330 30590 40332
rect 30294 40278 30320 40330
rect 30320 40278 30350 40330
rect 30374 40278 30384 40330
rect 30384 40278 30430 40330
rect 30454 40278 30500 40330
rect 30500 40278 30510 40330
rect 30534 40278 30564 40330
rect 30564 40278 30590 40330
rect 30294 40276 30350 40278
rect 30374 40276 30430 40278
rect 30454 40276 30510 40278
rect 30534 40276 30590 40278
rect 30294 39242 30350 39244
rect 30374 39242 30430 39244
rect 30454 39242 30510 39244
rect 30534 39242 30590 39244
rect 30294 39190 30320 39242
rect 30320 39190 30350 39242
rect 30374 39190 30384 39242
rect 30384 39190 30430 39242
rect 30454 39190 30500 39242
rect 30500 39190 30510 39242
rect 30534 39190 30564 39242
rect 30564 39190 30590 39242
rect 30294 39188 30350 39190
rect 30374 39188 30430 39190
rect 30454 39188 30510 39190
rect 30534 39188 30590 39190
rect 30294 38154 30350 38156
rect 30374 38154 30430 38156
rect 30454 38154 30510 38156
rect 30534 38154 30590 38156
rect 30294 38102 30320 38154
rect 30320 38102 30350 38154
rect 30374 38102 30384 38154
rect 30384 38102 30430 38154
rect 30454 38102 30500 38154
rect 30500 38102 30510 38154
rect 30534 38102 30564 38154
rect 30564 38102 30590 38154
rect 30294 38100 30350 38102
rect 30374 38100 30430 38102
rect 30454 38100 30510 38102
rect 30534 38100 30590 38102
rect 30294 37066 30350 37068
rect 30374 37066 30430 37068
rect 30454 37066 30510 37068
rect 30534 37066 30590 37068
rect 30294 37014 30320 37066
rect 30320 37014 30350 37066
rect 30374 37014 30384 37066
rect 30384 37014 30430 37066
rect 30454 37014 30500 37066
rect 30500 37014 30510 37066
rect 30534 37014 30564 37066
rect 30564 37014 30590 37066
rect 30294 37012 30350 37014
rect 30374 37012 30430 37014
rect 30454 37012 30510 37014
rect 30534 37012 30590 37014
rect 30294 35978 30350 35980
rect 30374 35978 30430 35980
rect 30454 35978 30510 35980
rect 30534 35978 30590 35980
rect 30294 35926 30320 35978
rect 30320 35926 30350 35978
rect 30374 35926 30384 35978
rect 30384 35926 30430 35978
rect 30454 35926 30500 35978
rect 30500 35926 30510 35978
rect 30534 35926 30564 35978
rect 30564 35926 30590 35978
rect 30294 35924 30350 35926
rect 30374 35924 30430 35926
rect 30454 35924 30510 35926
rect 30534 35924 30590 35926
rect 30294 34890 30350 34892
rect 30374 34890 30430 34892
rect 30454 34890 30510 34892
rect 30534 34890 30590 34892
rect 30294 34838 30320 34890
rect 30320 34838 30350 34890
rect 30374 34838 30384 34890
rect 30384 34838 30430 34890
rect 30454 34838 30500 34890
rect 30500 34838 30510 34890
rect 30534 34838 30564 34890
rect 30564 34838 30590 34890
rect 30294 34836 30350 34838
rect 30374 34836 30430 34838
rect 30454 34836 30510 34838
rect 30534 34836 30590 34838
rect 30294 33802 30350 33804
rect 30374 33802 30430 33804
rect 30454 33802 30510 33804
rect 30534 33802 30590 33804
rect 30294 33750 30320 33802
rect 30320 33750 30350 33802
rect 30374 33750 30384 33802
rect 30384 33750 30430 33802
rect 30454 33750 30500 33802
rect 30500 33750 30510 33802
rect 30534 33750 30564 33802
rect 30564 33750 30590 33802
rect 30294 33748 30350 33750
rect 30374 33748 30430 33750
rect 30454 33748 30510 33750
rect 30534 33748 30590 33750
rect 32958 41962 33014 41964
rect 33038 41962 33094 41964
rect 33118 41962 33174 41964
rect 33198 41962 33254 41964
rect 32958 41910 32984 41962
rect 32984 41910 33014 41962
rect 33038 41910 33048 41962
rect 33048 41910 33094 41962
rect 33118 41910 33164 41962
rect 33164 41910 33174 41962
rect 33198 41910 33228 41962
rect 33228 41910 33254 41962
rect 32958 41908 33014 41910
rect 33038 41908 33094 41910
rect 33118 41908 33174 41910
rect 33198 41908 33254 41910
rect 32958 40874 33014 40876
rect 33038 40874 33094 40876
rect 33118 40874 33174 40876
rect 33198 40874 33254 40876
rect 32958 40822 32984 40874
rect 32984 40822 33014 40874
rect 33038 40822 33048 40874
rect 33048 40822 33094 40874
rect 33118 40822 33164 40874
rect 33164 40822 33174 40874
rect 33198 40822 33228 40874
rect 33228 40822 33254 40874
rect 32958 40820 33014 40822
rect 33038 40820 33094 40822
rect 33118 40820 33174 40822
rect 33198 40820 33254 40822
rect 32958 39786 33014 39788
rect 33038 39786 33094 39788
rect 33118 39786 33174 39788
rect 33198 39786 33254 39788
rect 32958 39734 32984 39786
rect 32984 39734 33014 39786
rect 33038 39734 33048 39786
rect 33048 39734 33094 39786
rect 33118 39734 33164 39786
rect 33164 39734 33174 39786
rect 33198 39734 33228 39786
rect 33228 39734 33254 39786
rect 32958 39732 33014 39734
rect 33038 39732 33094 39734
rect 33118 39732 33174 39734
rect 33198 39732 33254 39734
rect 32958 38698 33014 38700
rect 33038 38698 33094 38700
rect 33118 38698 33174 38700
rect 33198 38698 33254 38700
rect 32958 38646 32984 38698
rect 32984 38646 33014 38698
rect 33038 38646 33048 38698
rect 33048 38646 33094 38698
rect 33118 38646 33164 38698
rect 33164 38646 33174 38698
rect 33198 38646 33228 38698
rect 33228 38646 33254 38698
rect 32958 38644 33014 38646
rect 33038 38644 33094 38646
rect 33118 38644 33174 38646
rect 33198 38644 33254 38646
rect 32958 37610 33014 37612
rect 33038 37610 33094 37612
rect 33118 37610 33174 37612
rect 33198 37610 33254 37612
rect 32958 37558 32984 37610
rect 32984 37558 33014 37610
rect 33038 37558 33048 37610
rect 33048 37558 33094 37610
rect 33118 37558 33164 37610
rect 33164 37558 33174 37610
rect 33198 37558 33228 37610
rect 33228 37558 33254 37610
rect 32958 37556 33014 37558
rect 33038 37556 33094 37558
rect 33118 37556 33174 37558
rect 33198 37556 33254 37558
rect 32958 36522 33014 36524
rect 33038 36522 33094 36524
rect 33118 36522 33174 36524
rect 33198 36522 33254 36524
rect 32958 36470 32984 36522
rect 32984 36470 33014 36522
rect 33038 36470 33048 36522
rect 33048 36470 33094 36522
rect 33118 36470 33164 36522
rect 33164 36470 33174 36522
rect 33198 36470 33228 36522
rect 33228 36470 33254 36522
rect 32958 36468 33014 36470
rect 33038 36468 33094 36470
rect 33118 36468 33174 36470
rect 33198 36468 33254 36470
rect 30364 33564 30420 33600
rect 30364 33544 30366 33564
rect 30366 33544 30418 33564
rect 30418 33544 30420 33564
rect 30732 33544 30788 33600
rect 32958 35434 33014 35436
rect 33038 35434 33094 35436
rect 33118 35434 33174 35436
rect 33198 35434 33254 35436
rect 32958 35382 32984 35434
rect 32984 35382 33014 35434
rect 33038 35382 33048 35434
rect 33048 35382 33094 35434
rect 33118 35382 33164 35434
rect 33164 35382 33174 35434
rect 33198 35382 33228 35434
rect 33228 35382 33254 35434
rect 32958 35380 33014 35382
rect 33038 35380 33094 35382
rect 33118 35380 33174 35382
rect 33198 35380 33254 35382
rect 32958 34346 33014 34348
rect 33038 34346 33094 34348
rect 33118 34346 33174 34348
rect 33198 34346 33254 34348
rect 32958 34294 32984 34346
rect 32984 34294 33014 34346
rect 33038 34294 33048 34346
rect 33048 34294 33094 34346
rect 33118 34294 33164 34346
rect 33164 34294 33174 34346
rect 33198 34294 33228 34346
rect 33228 34294 33254 34346
rect 32958 34292 33014 34294
rect 33038 34292 33094 34294
rect 33118 34292 33174 34294
rect 33198 34292 33254 34294
rect 28524 31812 28526 31832
rect 28526 31812 28578 31832
rect 28578 31812 28580 31832
rect 28524 31776 28580 31812
rect 28432 31404 28434 31424
rect 28434 31404 28486 31424
rect 28486 31404 28488 31424
rect 27630 31082 27686 31084
rect 27710 31082 27766 31084
rect 27790 31082 27846 31084
rect 27870 31082 27926 31084
rect 27630 31030 27656 31082
rect 27656 31030 27686 31082
rect 27710 31030 27720 31082
rect 27720 31030 27766 31082
rect 27790 31030 27836 31082
rect 27836 31030 27846 31082
rect 27870 31030 27900 31082
rect 27900 31030 27926 31082
rect 27630 31028 27686 31030
rect 27710 31028 27766 31030
rect 27790 31028 27846 31030
rect 27870 31028 27926 31030
rect 24844 28668 24900 28704
rect 25764 28684 25766 28704
rect 25766 28684 25818 28704
rect 25818 28684 25820 28704
rect 24844 28648 24846 28668
rect 24846 28648 24898 28668
rect 24898 28648 24900 28668
rect 25764 28648 25820 28684
rect 27420 29872 27476 29928
rect 27630 29994 27686 29996
rect 27710 29994 27766 29996
rect 27790 29994 27846 29996
rect 27870 29994 27926 29996
rect 27630 29942 27656 29994
rect 27656 29942 27686 29994
rect 27710 29942 27720 29994
rect 27720 29942 27766 29994
rect 27790 29942 27836 29994
rect 27836 29942 27846 29994
rect 27870 29942 27900 29994
rect 27900 29942 27926 29994
rect 27630 29940 27686 29942
rect 27710 29940 27766 29942
rect 27790 29940 27846 29942
rect 27870 29940 27926 29942
rect 28432 31368 28488 31404
rect 28524 31232 28580 31288
rect 28340 30316 28342 30336
rect 28342 30316 28394 30336
rect 28394 30316 28396 30336
rect 28340 30280 28396 30316
rect 30294 32714 30350 32716
rect 30374 32714 30430 32716
rect 30454 32714 30510 32716
rect 30534 32714 30590 32716
rect 30294 32662 30320 32714
rect 30320 32662 30350 32714
rect 30374 32662 30384 32714
rect 30384 32662 30430 32714
rect 30454 32662 30500 32714
rect 30500 32662 30510 32714
rect 30534 32662 30564 32714
rect 30564 32662 30590 32714
rect 30294 32660 30350 32662
rect 30374 32660 30430 32662
rect 30454 32660 30510 32662
rect 30534 32660 30590 32662
rect 28984 31776 29040 31832
rect 28708 31368 28764 31424
rect 27630 28906 27686 28908
rect 27710 28906 27766 28908
rect 27790 28906 27846 28908
rect 27870 28906 27926 28908
rect 27630 28854 27656 28906
rect 27656 28854 27686 28906
rect 27710 28854 27720 28906
rect 27720 28854 27766 28906
rect 27790 28854 27836 28906
rect 27836 28854 27846 28906
rect 27870 28854 27900 28906
rect 27900 28854 27926 28906
rect 27630 28852 27686 28854
rect 27710 28852 27766 28854
rect 27790 28852 27846 28854
rect 27870 28852 27926 28854
rect 27972 28648 28028 28704
rect 24966 28362 25022 28364
rect 25046 28362 25102 28364
rect 25126 28362 25182 28364
rect 25206 28362 25262 28364
rect 24966 28310 24992 28362
rect 24992 28310 25022 28362
rect 25046 28310 25056 28362
rect 25056 28310 25102 28362
rect 25126 28310 25172 28362
rect 25172 28310 25182 28362
rect 25206 28310 25236 28362
rect 25236 28310 25262 28362
rect 24966 28308 25022 28310
rect 25046 28308 25102 28310
rect 25126 28308 25182 28310
rect 25206 28308 25262 28310
rect 24384 27968 24440 28024
rect 25212 27424 25268 27480
rect 24966 27274 25022 27276
rect 25046 27274 25102 27276
rect 25126 27274 25182 27276
rect 25206 27274 25262 27276
rect 24966 27222 24992 27274
rect 24992 27222 25022 27274
rect 25046 27222 25056 27274
rect 25056 27222 25102 27274
rect 25126 27222 25172 27274
rect 25172 27222 25182 27274
rect 25206 27222 25236 27274
rect 25236 27222 25262 27274
rect 24966 27220 25022 27222
rect 25046 27220 25102 27222
rect 25126 27220 25182 27222
rect 25206 27220 25262 27222
rect 28524 28512 28580 28568
rect 27630 27818 27686 27820
rect 27710 27818 27766 27820
rect 27790 27818 27846 27820
rect 27870 27818 27926 27820
rect 27630 27766 27656 27818
rect 27656 27766 27686 27818
rect 27710 27766 27720 27818
rect 27720 27766 27766 27818
rect 27790 27766 27836 27818
rect 27836 27766 27846 27818
rect 27870 27766 27900 27818
rect 27900 27766 27926 27818
rect 27630 27764 27686 27766
rect 27710 27764 27766 27766
rect 27790 27764 27846 27766
rect 27870 27764 27926 27766
rect 30294 31626 30350 31628
rect 30374 31626 30430 31628
rect 30454 31626 30510 31628
rect 30534 31626 30590 31628
rect 30294 31574 30320 31626
rect 30320 31574 30350 31626
rect 30374 31574 30384 31626
rect 30384 31574 30430 31626
rect 30454 31574 30500 31626
rect 30500 31574 30510 31626
rect 30534 31574 30564 31626
rect 30564 31574 30590 31626
rect 30294 31572 30350 31574
rect 30374 31572 30430 31574
rect 30454 31572 30510 31574
rect 30534 31572 30590 31574
rect 32958 33258 33014 33260
rect 33038 33258 33094 33260
rect 33118 33258 33174 33260
rect 33198 33258 33254 33260
rect 32958 33206 32984 33258
rect 32984 33206 33014 33258
rect 33038 33206 33048 33258
rect 33048 33206 33094 33258
rect 33118 33206 33164 33258
rect 33164 33206 33174 33258
rect 33198 33206 33228 33258
rect 33228 33206 33254 33258
rect 32958 33204 33014 33206
rect 33038 33204 33094 33206
rect 33118 33204 33174 33206
rect 33198 33204 33254 33206
rect 35622 41418 35678 41420
rect 35702 41418 35758 41420
rect 35782 41418 35838 41420
rect 35862 41418 35918 41420
rect 35622 41366 35648 41418
rect 35648 41366 35678 41418
rect 35702 41366 35712 41418
rect 35712 41366 35758 41418
rect 35782 41366 35828 41418
rect 35828 41366 35838 41418
rect 35862 41366 35892 41418
rect 35892 41366 35918 41418
rect 35622 41364 35678 41366
rect 35702 41364 35758 41366
rect 35782 41364 35838 41366
rect 35862 41364 35918 41366
rect 35622 40330 35678 40332
rect 35702 40330 35758 40332
rect 35782 40330 35838 40332
rect 35862 40330 35918 40332
rect 35622 40278 35648 40330
rect 35648 40278 35678 40330
rect 35702 40278 35712 40330
rect 35712 40278 35758 40330
rect 35782 40278 35828 40330
rect 35828 40278 35838 40330
rect 35862 40278 35892 40330
rect 35892 40278 35918 40330
rect 35622 40276 35678 40278
rect 35702 40276 35758 40278
rect 35782 40276 35838 40278
rect 35862 40276 35918 40278
rect 38286 41962 38342 41964
rect 38366 41962 38422 41964
rect 38446 41962 38502 41964
rect 38526 41962 38582 41964
rect 38286 41910 38312 41962
rect 38312 41910 38342 41962
rect 38366 41910 38376 41962
rect 38376 41910 38422 41962
rect 38446 41910 38492 41962
rect 38492 41910 38502 41962
rect 38526 41910 38556 41962
rect 38556 41910 38582 41962
rect 38286 41908 38342 41910
rect 38366 41908 38422 41910
rect 38446 41908 38502 41910
rect 38526 41908 38582 41910
rect 38286 40874 38342 40876
rect 38366 40874 38422 40876
rect 38446 40874 38502 40876
rect 38526 40874 38582 40876
rect 38286 40822 38312 40874
rect 38312 40822 38342 40874
rect 38366 40822 38376 40874
rect 38376 40822 38422 40874
rect 38446 40822 38492 40874
rect 38492 40822 38502 40874
rect 38526 40822 38556 40874
rect 38556 40822 38582 40874
rect 38286 40820 38342 40822
rect 38366 40820 38422 40822
rect 38446 40820 38502 40822
rect 38526 40820 38582 40822
rect 38286 39786 38342 39788
rect 38366 39786 38422 39788
rect 38446 39786 38502 39788
rect 38526 39786 38582 39788
rect 38286 39734 38312 39786
rect 38312 39734 38342 39786
rect 38366 39734 38376 39786
rect 38376 39734 38422 39786
rect 38446 39734 38492 39786
rect 38492 39734 38502 39786
rect 38526 39734 38556 39786
rect 38556 39734 38582 39786
rect 38286 39732 38342 39734
rect 38366 39732 38422 39734
rect 38446 39732 38502 39734
rect 38526 39732 38582 39734
rect 35622 39242 35678 39244
rect 35702 39242 35758 39244
rect 35782 39242 35838 39244
rect 35862 39242 35918 39244
rect 35622 39190 35648 39242
rect 35648 39190 35678 39242
rect 35702 39190 35712 39242
rect 35712 39190 35758 39242
rect 35782 39190 35828 39242
rect 35828 39190 35838 39242
rect 35862 39190 35892 39242
rect 35892 39190 35918 39242
rect 35622 39188 35678 39190
rect 35702 39188 35758 39190
rect 35782 39188 35838 39190
rect 35862 39188 35918 39190
rect 38286 38698 38342 38700
rect 38366 38698 38422 38700
rect 38446 38698 38502 38700
rect 38526 38698 38582 38700
rect 38286 38646 38312 38698
rect 38312 38646 38342 38698
rect 38366 38646 38376 38698
rect 38376 38646 38422 38698
rect 38446 38646 38492 38698
rect 38492 38646 38502 38698
rect 38526 38646 38556 38698
rect 38556 38646 38582 38698
rect 38286 38644 38342 38646
rect 38366 38644 38422 38646
rect 38446 38644 38502 38646
rect 38526 38644 38582 38646
rect 35622 38154 35678 38156
rect 35702 38154 35758 38156
rect 35782 38154 35838 38156
rect 35862 38154 35918 38156
rect 35622 38102 35648 38154
rect 35648 38102 35678 38154
rect 35702 38102 35712 38154
rect 35712 38102 35758 38154
rect 35782 38102 35828 38154
rect 35828 38102 35838 38154
rect 35862 38102 35892 38154
rect 35892 38102 35918 38154
rect 35622 38100 35678 38102
rect 35702 38100 35758 38102
rect 35782 38100 35838 38102
rect 35862 38100 35918 38102
rect 32958 32170 33014 32172
rect 33038 32170 33094 32172
rect 33118 32170 33174 32172
rect 33198 32170 33254 32172
rect 32958 32118 32984 32170
rect 32984 32118 33014 32170
rect 33038 32118 33048 32170
rect 33048 32118 33094 32170
rect 33118 32118 33164 32170
rect 33164 32118 33174 32170
rect 33198 32118 33228 32170
rect 33228 32118 33254 32170
rect 32958 32116 33014 32118
rect 33038 32116 33094 32118
rect 33118 32116 33174 32118
rect 33198 32116 33254 32118
rect 32572 31368 32628 31424
rect 30294 30538 30350 30540
rect 30374 30538 30430 30540
rect 30454 30538 30510 30540
rect 30534 30538 30590 30540
rect 30294 30486 30320 30538
rect 30320 30486 30350 30538
rect 30374 30486 30384 30538
rect 30384 30486 30430 30538
rect 30454 30486 30500 30538
rect 30500 30486 30510 30538
rect 30534 30486 30564 30538
rect 30564 30486 30590 30538
rect 30294 30484 30350 30486
rect 30374 30484 30430 30486
rect 30454 30484 30510 30486
rect 30534 30484 30590 30486
rect 30294 29450 30350 29452
rect 30374 29450 30430 29452
rect 30454 29450 30510 29452
rect 30534 29450 30590 29452
rect 30294 29398 30320 29450
rect 30320 29398 30350 29450
rect 30374 29398 30384 29450
rect 30384 29398 30430 29450
rect 30454 29398 30500 29450
rect 30500 29398 30510 29450
rect 30534 29398 30564 29450
rect 30564 29398 30590 29450
rect 30294 29396 30350 29398
rect 30374 29396 30430 29398
rect 30454 29396 30510 29398
rect 30534 29396 30590 29398
rect 30294 28362 30350 28364
rect 30374 28362 30430 28364
rect 30454 28362 30510 28364
rect 30534 28362 30590 28364
rect 30294 28310 30320 28362
rect 30320 28310 30350 28362
rect 30374 28310 30384 28362
rect 30384 28310 30430 28362
rect 30454 28310 30500 28362
rect 30500 28310 30510 28362
rect 30534 28310 30564 28362
rect 30564 28310 30590 28362
rect 30294 28308 30350 28310
rect 30374 28308 30430 28310
rect 30454 28308 30510 28310
rect 30534 28308 30590 28310
rect 30364 27968 30420 28024
rect 29904 27696 29960 27752
rect 29812 27560 29868 27616
rect 29720 27016 29776 27072
rect 30180 27424 30236 27480
rect 30294 27274 30350 27276
rect 30374 27274 30430 27276
rect 30454 27274 30510 27276
rect 30534 27274 30590 27276
rect 30294 27222 30320 27274
rect 30320 27222 30350 27274
rect 30374 27222 30384 27274
rect 30384 27222 30430 27274
rect 30454 27222 30500 27274
rect 30500 27222 30510 27274
rect 30534 27222 30564 27274
rect 30564 27222 30590 27274
rect 30294 27220 30350 27222
rect 30374 27220 30430 27222
rect 30454 27220 30510 27222
rect 30534 27220 30590 27222
rect 29352 26900 29408 26936
rect 29352 26880 29354 26900
rect 29354 26880 29406 26900
rect 29406 26880 29408 26900
rect 30364 26880 30420 26936
rect 30732 26916 30734 26936
rect 30734 26916 30786 26936
rect 30786 26916 30788 26936
rect 30732 26880 30788 26916
rect 27630 26730 27686 26732
rect 27710 26730 27766 26732
rect 27790 26730 27846 26732
rect 27870 26730 27926 26732
rect 27630 26678 27656 26730
rect 27656 26678 27686 26730
rect 27710 26678 27720 26730
rect 27720 26678 27766 26730
rect 27790 26678 27836 26730
rect 27836 26678 27846 26730
rect 27870 26678 27900 26730
rect 27900 26678 27926 26730
rect 27630 26676 27686 26678
rect 27710 26676 27766 26678
rect 27790 26676 27846 26678
rect 27870 26676 27926 26678
rect 32958 31082 33014 31084
rect 33038 31082 33094 31084
rect 33118 31082 33174 31084
rect 33198 31082 33254 31084
rect 32958 31030 32984 31082
rect 32984 31030 33014 31082
rect 33038 31030 33048 31082
rect 33048 31030 33094 31082
rect 33118 31030 33164 31082
rect 33164 31030 33174 31082
rect 33198 31030 33228 31082
rect 33228 31030 33254 31082
rect 32958 31028 33014 31030
rect 33038 31028 33094 31030
rect 33118 31028 33174 31030
rect 33198 31028 33254 31030
rect 32958 29994 33014 29996
rect 33038 29994 33094 29996
rect 33118 29994 33174 29996
rect 33198 29994 33254 29996
rect 32958 29942 32984 29994
rect 32984 29942 33014 29994
rect 33038 29942 33048 29994
rect 33048 29942 33094 29994
rect 33118 29942 33164 29994
rect 33164 29942 33174 29994
rect 33198 29942 33228 29994
rect 33228 29942 33254 29994
rect 32958 29940 33014 29942
rect 33038 29940 33094 29942
rect 33118 29940 33174 29942
rect 33198 29940 33254 29942
rect 33216 29076 33272 29112
rect 33216 29056 33218 29076
rect 33218 29056 33270 29076
rect 33270 29056 33272 29076
rect 32958 28906 33014 28908
rect 33038 28906 33094 28908
rect 33118 28906 33174 28908
rect 33198 28906 33254 28908
rect 32958 28854 32984 28906
rect 32984 28854 33014 28906
rect 33038 28854 33048 28906
rect 33048 28854 33094 28906
rect 33118 28854 33164 28906
rect 33164 28854 33174 28906
rect 33198 28854 33228 28906
rect 33228 28854 33254 28906
rect 32958 28852 33014 28854
rect 33038 28852 33094 28854
rect 33118 28852 33174 28854
rect 33198 28852 33254 28854
rect 31376 28004 31378 28024
rect 31378 28004 31430 28024
rect 31430 28004 31432 28024
rect 31376 27968 31432 28004
rect 31284 27868 31286 27888
rect 31286 27868 31338 27888
rect 31338 27868 31340 27888
rect 31284 27832 31340 27868
rect 31192 27560 31248 27616
rect 31468 27696 31524 27752
rect 32958 27818 33014 27820
rect 33038 27818 33094 27820
rect 33118 27818 33174 27820
rect 33198 27818 33254 27820
rect 32958 27766 32984 27818
rect 32984 27766 33014 27818
rect 33038 27766 33048 27818
rect 33048 27766 33094 27818
rect 33118 27766 33164 27818
rect 33164 27766 33174 27818
rect 33198 27766 33228 27818
rect 33228 27766 33254 27818
rect 32958 27764 33014 27766
rect 33038 27764 33094 27766
rect 33118 27764 33174 27766
rect 33198 27764 33254 27766
rect 31744 27424 31800 27480
rect 31652 27052 31654 27072
rect 31654 27052 31706 27072
rect 31706 27052 31708 27072
rect 31652 27016 31708 27052
rect 31376 26880 31432 26936
rect 32958 26730 33014 26732
rect 33038 26730 33094 26732
rect 33118 26730 33174 26732
rect 33198 26730 33254 26732
rect 32958 26678 32984 26730
rect 32984 26678 33014 26730
rect 33038 26678 33048 26730
rect 33048 26678 33094 26730
rect 33118 26678 33164 26730
rect 33164 26678 33174 26730
rect 33198 26678 33228 26730
rect 33228 26678 33254 26730
rect 32958 26676 33014 26678
rect 33038 26676 33094 26678
rect 33118 26676 33174 26678
rect 33198 26676 33254 26678
rect 31376 23004 31432 23060
rect 33952 21304 34008 21360
rect 35622 37066 35678 37068
rect 35702 37066 35758 37068
rect 35782 37066 35838 37068
rect 35862 37066 35918 37068
rect 35622 37014 35648 37066
rect 35648 37014 35678 37066
rect 35702 37014 35712 37066
rect 35712 37014 35758 37066
rect 35782 37014 35828 37066
rect 35828 37014 35838 37066
rect 35862 37014 35892 37066
rect 35892 37014 35918 37066
rect 35622 37012 35678 37014
rect 35702 37012 35758 37014
rect 35782 37012 35838 37014
rect 35862 37012 35918 37014
rect 37540 36808 37596 36864
rect 37448 36128 37504 36184
rect 37724 36672 37780 36728
rect 35622 35978 35678 35980
rect 35702 35978 35758 35980
rect 35782 35978 35838 35980
rect 35862 35978 35918 35980
rect 35622 35926 35648 35978
rect 35648 35926 35678 35978
rect 35702 35926 35712 35978
rect 35712 35926 35758 35978
rect 35782 35926 35828 35978
rect 35828 35926 35838 35978
rect 35862 35926 35892 35978
rect 35892 35926 35918 35978
rect 35622 35924 35678 35926
rect 35702 35924 35758 35926
rect 35782 35924 35838 35926
rect 35862 35924 35918 35926
rect 35622 34890 35678 34892
rect 35702 34890 35758 34892
rect 35782 34890 35838 34892
rect 35862 34890 35918 34892
rect 35622 34838 35648 34890
rect 35648 34838 35678 34890
rect 35702 34838 35712 34890
rect 35712 34838 35758 34890
rect 35782 34838 35828 34890
rect 35828 34838 35838 34890
rect 35862 34838 35892 34890
rect 35892 34838 35918 34890
rect 35622 34836 35678 34838
rect 35702 34836 35758 34838
rect 35782 34836 35838 34838
rect 35862 34836 35918 34838
rect 35240 33564 35296 33600
rect 35240 33544 35242 33564
rect 35242 33544 35294 33564
rect 35294 33544 35296 33564
rect 35622 33802 35678 33804
rect 35702 33802 35758 33804
rect 35782 33802 35838 33804
rect 35862 33802 35918 33804
rect 35622 33750 35648 33802
rect 35648 33750 35678 33802
rect 35702 33750 35712 33802
rect 35712 33750 35758 33802
rect 35782 33750 35828 33802
rect 35828 33750 35838 33802
rect 35862 33750 35892 33802
rect 35892 33750 35918 33802
rect 35622 33748 35678 33750
rect 35702 33748 35758 33750
rect 35782 33748 35838 33750
rect 35862 33748 35918 33750
rect 35622 32714 35678 32716
rect 35702 32714 35758 32716
rect 35782 32714 35838 32716
rect 35862 32714 35918 32716
rect 35622 32662 35648 32714
rect 35648 32662 35678 32714
rect 35702 32662 35712 32714
rect 35712 32662 35758 32714
rect 35782 32662 35828 32714
rect 35828 32662 35838 32714
rect 35862 32662 35892 32714
rect 35892 32662 35918 32714
rect 35622 32660 35678 32662
rect 35702 32660 35758 32662
rect 35782 32660 35838 32662
rect 35862 32660 35918 32662
rect 38286 37610 38342 37612
rect 38366 37610 38422 37612
rect 38446 37610 38502 37612
rect 38526 37610 38582 37612
rect 38286 37558 38312 37610
rect 38312 37558 38342 37610
rect 38366 37558 38376 37610
rect 38376 37558 38422 37610
rect 38446 37558 38492 37610
rect 38492 37558 38502 37610
rect 38526 37558 38556 37610
rect 38556 37558 38582 37610
rect 38286 37556 38342 37558
rect 38366 37556 38422 37558
rect 38446 37556 38502 37558
rect 38526 37556 38582 37558
rect 39104 37216 39160 37272
rect 38286 36522 38342 36524
rect 38366 36522 38422 36524
rect 38446 36522 38502 36524
rect 38526 36522 38582 36524
rect 38286 36470 38312 36522
rect 38312 36470 38342 36522
rect 38366 36470 38376 36522
rect 38376 36470 38422 36522
rect 38446 36470 38492 36522
rect 38492 36470 38502 36522
rect 38526 36470 38556 36522
rect 38556 36470 38582 36522
rect 38286 36468 38342 36470
rect 38366 36468 38422 36470
rect 38446 36468 38502 36470
rect 38526 36468 38582 36470
rect 40950 41418 41006 41420
rect 41030 41418 41086 41420
rect 41110 41418 41166 41420
rect 41190 41418 41246 41420
rect 40950 41366 40976 41418
rect 40976 41366 41006 41418
rect 41030 41366 41040 41418
rect 41040 41366 41086 41418
rect 41110 41366 41156 41418
rect 41156 41366 41166 41418
rect 41190 41366 41220 41418
rect 41220 41366 41246 41418
rect 40950 41364 41006 41366
rect 41030 41364 41086 41366
rect 41110 41364 41166 41366
rect 41190 41364 41246 41366
rect 39288 37624 39344 37680
rect 38286 35434 38342 35436
rect 38366 35434 38422 35436
rect 38446 35434 38502 35436
rect 38526 35434 38582 35436
rect 38286 35382 38312 35434
rect 38312 35382 38342 35434
rect 38366 35382 38376 35434
rect 38376 35382 38422 35434
rect 38446 35382 38492 35434
rect 38492 35382 38502 35434
rect 38526 35382 38556 35434
rect 38556 35382 38582 35434
rect 38286 35380 38342 35382
rect 38366 35380 38422 35382
rect 38446 35380 38502 35382
rect 38526 35380 38582 35382
rect 39380 34668 39382 34688
rect 39382 34668 39434 34688
rect 39434 34668 39436 34688
rect 39380 34632 39436 34668
rect 38286 34346 38342 34348
rect 38366 34346 38422 34348
rect 38446 34346 38502 34348
rect 38526 34346 38582 34348
rect 38286 34294 38312 34346
rect 38312 34294 38342 34346
rect 38366 34294 38376 34346
rect 38376 34294 38422 34346
rect 38446 34294 38492 34346
rect 38492 34294 38502 34346
rect 38526 34294 38556 34346
rect 38556 34294 38582 34346
rect 38286 34292 38342 34294
rect 38366 34292 38422 34294
rect 38446 34292 38502 34294
rect 38526 34292 38582 34294
rect 40950 40330 41006 40332
rect 41030 40330 41086 40332
rect 41110 40330 41166 40332
rect 41190 40330 41246 40332
rect 40950 40278 40976 40330
rect 40976 40278 41006 40330
rect 41030 40278 41040 40330
rect 41040 40278 41086 40330
rect 41110 40278 41156 40330
rect 41156 40278 41166 40330
rect 41190 40278 41220 40330
rect 41220 40278 41246 40330
rect 40950 40276 41006 40278
rect 41030 40276 41086 40278
rect 41110 40276 41166 40278
rect 41190 40276 41246 40278
rect 40950 39242 41006 39244
rect 41030 39242 41086 39244
rect 41110 39242 41166 39244
rect 41190 39242 41246 39244
rect 40950 39190 40976 39242
rect 40976 39190 41006 39242
rect 41030 39190 41040 39242
rect 41040 39190 41086 39242
rect 41110 39190 41156 39242
rect 41156 39190 41166 39242
rect 41190 39190 41220 39242
rect 41220 39190 41246 39242
rect 40950 39188 41006 39190
rect 41030 39188 41086 39190
rect 41110 39188 41166 39190
rect 41190 39188 41246 39190
rect 40950 38154 41006 38156
rect 41030 38154 41086 38156
rect 41110 38154 41166 38156
rect 41190 38154 41246 38156
rect 40950 38102 40976 38154
rect 40976 38102 41006 38154
rect 41030 38102 41040 38154
rect 41040 38102 41086 38154
rect 41110 38102 41156 38154
rect 41156 38102 41166 38154
rect 41190 38102 41220 38154
rect 41220 38102 41246 38154
rect 40950 38100 41006 38102
rect 41030 38100 41086 38102
rect 41110 38100 41166 38102
rect 41190 38100 41246 38102
rect 43614 41962 43670 41964
rect 43694 41962 43750 41964
rect 43774 41962 43830 41964
rect 43854 41962 43910 41964
rect 43614 41910 43640 41962
rect 43640 41910 43670 41962
rect 43694 41910 43704 41962
rect 43704 41910 43750 41962
rect 43774 41910 43820 41962
rect 43820 41910 43830 41962
rect 43854 41910 43884 41962
rect 43884 41910 43910 41962
rect 43614 41908 43670 41910
rect 43694 41908 43750 41910
rect 43774 41908 43830 41910
rect 43854 41908 43910 41910
rect 43614 40874 43670 40876
rect 43694 40874 43750 40876
rect 43774 40874 43830 40876
rect 43854 40874 43910 40876
rect 43614 40822 43640 40874
rect 43640 40822 43670 40874
rect 43694 40822 43704 40874
rect 43704 40822 43750 40874
rect 43774 40822 43820 40874
rect 43820 40822 43830 40874
rect 43854 40822 43884 40874
rect 43884 40822 43910 40874
rect 43614 40820 43670 40822
rect 43694 40820 43750 40822
rect 43774 40820 43830 40822
rect 43854 40820 43910 40822
rect 41772 37660 41774 37680
rect 41774 37660 41826 37680
rect 41826 37660 41828 37680
rect 41772 37624 41828 37660
rect 41220 37352 41276 37408
rect 43614 39786 43670 39788
rect 43694 39786 43750 39788
rect 43774 39786 43830 39788
rect 43854 39786 43910 39788
rect 43614 39734 43640 39786
rect 43640 39734 43670 39786
rect 43694 39734 43704 39786
rect 43704 39734 43750 39786
rect 43774 39734 43820 39786
rect 43820 39734 43830 39786
rect 43854 39734 43884 39786
rect 43884 39734 43910 39786
rect 43614 39732 43670 39734
rect 43694 39732 43750 39734
rect 43774 39732 43830 39734
rect 43854 39732 43910 39734
rect 46278 41418 46334 41420
rect 46358 41418 46414 41420
rect 46438 41418 46494 41420
rect 46518 41418 46574 41420
rect 46278 41366 46304 41418
rect 46304 41366 46334 41418
rect 46358 41366 46368 41418
rect 46368 41366 46414 41418
rect 46438 41366 46484 41418
rect 46484 41366 46494 41418
rect 46518 41366 46548 41418
rect 46548 41366 46574 41418
rect 46278 41364 46334 41366
rect 46358 41364 46414 41366
rect 46438 41364 46494 41366
rect 46518 41364 46574 41366
rect 46278 40330 46334 40332
rect 46358 40330 46414 40332
rect 46438 40330 46494 40332
rect 46518 40330 46574 40332
rect 46278 40278 46304 40330
rect 46304 40278 46334 40330
rect 46358 40278 46368 40330
rect 46368 40278 46414 40330
rect 46438 40278 46484 40330
rect 46484 40278 46494 40330
rect 46518 40278 46548 40330
rect 46548 40278 46574 40330
rect 46278 40276 46334 40278
rect 46358 40276 46414 40278
rect 46438 40276 46494 40278
rect 46518 40276 46574 40278
rect 46278 39242 46334 39244
rect 46358 39242 46414 39244
rect 46438 39242 46494 39244
rect 46518 39242 46574 39244
rect 46278 39190 46304 39242
rect 46304 39190 46334 39242
rect 46358 39190 46368 39242
rect 46368 39190 46414 39242
rect 46438 39190 46484 39242
rect 46484 39190 46494 39242
rect 46518 39190 46548 39242
rect 46548 39190 46574 39242
rect 46278 39188 46334 39190
rect 46358 39188 46414 39190
rect 46438 39188 46494 39190
rect 46518 39188 46574 39190
rect 43614 38698 43670 38700
rect 43694 38698 43750 38700
rect 43774 38698 43830 38700
rect 43854 38698 43910 38700
rect 43614 38646 43640 38698
rect 43640 38646 43670 38698
rect 43694 38646 43704 38698
rect 43704 38646 43750 38698
rect 43774 38646 43820 38698
rect 43820 38646 43830 38698
rect 43854 38646 43884 38698
rect 43884 38646 43910 38698
rect 43614 38644 43670 38646
rect 43694 38644 43750 38646
rect 43774 38644 43830 38646
rect 43854 38644 43910 38646
rect 48942 41962 48998 41964
rect 49022 41962 49078 41964
rect 49102 41962 49158 41964
rect 49182 41962 49238 41964
rect 48942 41910 48968 41962
rect 48968 41910 48998 41962
rect 49022 41910 49032 41962
rect 49032 41910 49078 41962
rect 49102 41910 49148 41962
rect 49148 41910 49158 41962
rect 49182 41910 49212 41962
rect 49212 41910 49238 41962
rect 48942 41908 48998 41910
rect 49022 41908 49078 41910
rect 49102 41908 49158 41910
rect 49182 41908 49238 41910
rect 48942 40874 48998 40876
rect 49022 40874 49078 40876
rect 49102 40874 49158 40876
rect 49182 40874 49238 40876
rect 48942 40822 48968 40874
rect 48968 40822 48998 40874
rect 49022 40822 49032 40874
rect 49032 40822 49078 40874
rect 49102 40822 49148 40874
rect 49148 40822 49158 40874
rect 49182 40822 49212 40874
rect 49212 40822 49238 40874
rect 48942 40820 48998 40822
rect 49022 40820 49078 40822
rect 49102 40820 49158 40822
rect 49182 40820 49238 40822
rect 48942 39786 48998 39788
rect 49022 39786 49078 39788
rect 49102 39786 49158 39788
rect 49182 39786 49238 39788
rect 48942 39734 48968 39786
rect 48968 39734 48998 39786
rect 49022 39734 49032 39786
rect 49032 39734 49078 39786
rect 49102 39734 49148 39786
rect 49148 39734 49158 39786
rect 49182 39734 49212 39786
rect 49212 39734 49238 39786
rect 48942 39732 48998 39734
rect 49022 39732 49078 39734
rect 49102 39732 49158 39734
rect 49182 39732 49238 39734
rect 50328 38984 50384 39040
rect 43614 37610 43670 37612
rect 43694 37610 43750 37612
rect 43774 37610 43830 37612
rect 43854 37610 43910 37612
rect 43614 37558 43640 37610
rect 43640 37558 43670 37610
rect 43694 37558 43704 37610
rect 43704 37558 43750 37610
rect 43774 37558 43820 37610
rect 43820 37558 43830 37610
rect 43854 37558 43884 37610
rect 43884 37558 43910 37610
rect 43614 37556 43670 37558
rect 43694 37556 43750 37558
rect 43774 37556 43830 37558
rect 43854 37556 43910 37558
rect 40950 37066 41006 37068
rect 41030 37066 41086 37068
rect 41110 37066 41166 37068
rect 41190 37066 41246 37068
rect 40950 37014 40976 37066
rect 40976 37014 41006 37066
rect 41030 37014 41040 37066
rect 41040 37014 41086 37066
rect 41110 37014 41156 37066
rect 41156 37014 41166 37066
rect 41190 37014 41220 37066
rect 41220 37014 41246 37066
rect 40950 37012 41006 37014
rect 41030 37012 41086 37014
rect 41110 37012 41166 37014
rect 41190 37012 41246 37014
rect 43612 37372 43668 37408
rect 43612 37352 43614 37372
rect 43614 37352 43666 37372
rect 43666 37352 43668 37372
rect 43704 36672 43760 36728
rect 43614 36522 43670 36524
rect 43694 36522 43750 36524
rect 43774 36522 43830 36524
rect 43854 36522 43910 36524
rect 43614 36470 43640 36522
rect 43640 36470 43670 36522
rect 43694 36470 43704 36522
rect 43704 36470 43750 36522
rect 43774 36470 43820 36522
rect 43820 36470 43830 36522
rect 43854 36470 43884 36522
rect 43884 36470 43910 36522
rect 43614 36468 43670 36470
rect 43694 36468 43750 36470
rect 43774 36468 43830 36470
rect 43854 36468 43910 36470
rect 38286 33258 38342 33260
rect 38366 33258 38422 33260
rect 38446 33258 38502 33260
rect 38526 33258 38582 33260
rect 38286 33206 38312 33258
rect 38312 33206 38342 33258
rect 38366 33206 38376 33258
rect 38376 33206 38422 33258
rect 38446 33206 38492 33258
rect 38492 33206 38502 33258
rect 38526 33206 38556 33258
rect 38556 33206 38582 33258
rect 38286 33204 38342 33206
rect 38366 33204 38422 33206
rect 38446 33204 38502 33206
rect 38526 33204 38582 33206
rect 35622 31626 35678 31628
rect 35702 31626 35758 31628
rect 35782 31626 35838 31628
rect 35862 31626 35918 31628
rect 35622 31574 35648 31626
rect 35648 31574 35678 31626
rect 35702 31574 35712 31626
rect 35712 31574 35758 31626
rect 35782 31574 35828 31626
rect 35828 31574 35838 31626
rect 35862 31574 35892 31626
rect 35892 31574 35918 31626
rect 35622 31572 35678 31574
rect 35702 31572 35758 31574
rect 35782 31572 35838 31574
rect 35862 31572 35918 31574
rect 35622 30538 35678 30540
rect 35702 30538 35758 30540
rect 35782 30538 35838 30540
rect 35862 30538 35918 30540
rect 35622 30486 35648 30538
rect 35648 30486 35678 30538
rect 35702 30486 35712 30538
rect 35712 30486 35758 30538
rect 35782 30486 35828 30538
rect 35828 30486 35838 30538
rect 35862 30486 35892 30538
rect 35892 30486 35918 30538
rect 35622 30484 35678 30486
rect 35702 30484 35758 30486
rect 35782 30484 35838 30486
rect 35862 30484 35918 30486
rect 35622 29450 35678 29452
rect 35702 29450 35758 29452
rect 35782 29450 35838 29452
rect 35862 29450 35918 29452
rect 35622 29398 35648 29450
rect 35648 29398 35678 29450
rect 35702 29398 35712 29450
rect 35712 29398 35758 29450
rect 35782 29398 35828 29450
rect 35828 29398 35838 29450
rect 35862 29398 35892 29450
rect 35892 29398 35918 29450
rect 35622 29396 35678 29398
rect 35702 29396 35758 29398
rect 35782 29396 35838 29398
rect 35862 29396 35918 29398
rect 35622 28362 35678 28364
rect 35702 28362 35758 28364
rect 35782 28362 35838 28364
rect 35862 28362 35918 28364
rect 35622 28310 35648 28362
rect 35648 28310 35678 28362
rect 35702 28310 35712 28362
rect 35712 28310 35758 28362
rect 35782 28310 35828 28362
rect 35828 28310 35838 28362
rect 35862 28310 35892 28362
rect 35892 28310 35918 28362
rect 35622 28308 35678 28310
rect 35702 28308 35758 28310
rect 35782 28308 35838 28310
rect 35862 28308 35918 28310
rect 34320 23480 34376 23536
rect 34780 22428 34782 22448
rect 34782 22428 34834 22448
rect 34834 22428 34836 22448
rect 34780 22392 34836 22428
rect 34412 20252 34414 20272
rect 34414 20252 34466 20272
rect 34466 20252 34468 20272
rect 34412 20216 34468 20252
rect 34412 19164 34414 19184
rect 34414 19164 34466 19184
rect 34466 19164 34468 19184
rect 34412 19128 34468 19164
rect 34780 21340 34782 21360
rect 34782 21340 34834 21360
rect 34834 21340 34836 21360
rect 34780 21304 34836 21340
rect 36712 27988 36768 28024
rect 36712 27968 36714 27988
rect 36714 27968 36766 27988
rect 36766 27968 36768 27988
rect 35622 27274 35678 27276
rect 35702 27274 35758 27276
rect 35782 27274 35838 27276
rect 35862 27274 35918 27276
rect 35622 27222 35648 27274
rect 35648 27222 35678 27274
rect 35702 27222 35712 27274
rect 35712 27222 35758 27274
rect 35782 27222 35828 27274
rect 35828 27222 35838 27274
rect 35862 27222 35892 27274
rect 35892 27222 35918 27274
rect 35622 27220 35678 27222
rect 35702 27220 35758 27222
rect 35782 27220 35838 27222
rect 35862 27220 35918 27222
rect 35622 26186 35678 26188
rect 35702 26186 35758 26188
rect 35782 26186 35838 26188
rect 35862 26186 35918 26188
rect 35622 26134 35648 26186
rect 35648 26134 35678 26186
rect 35702 26134 35712 26186
rect 35712 26134 35758 26186
rect 35782 26134 35828 26186
rect 35828 26134 35838 26186
rect 35862 26134 35892 26186
rect 35892 26134 35918 26186
rect 35622 26132 35678 26134
rect 35702 26132 35758 26134
rect 35782 26132 35838 26134
rect 35862 26132 35918 26134
rect 35622 25098 35678 25100
rect 35702 25098 35758 25100
rect 35782 25098 35838 25100
rect 35862 25098 35918 25100
rect 35622 25046 35648 25098
rect 35648 25046 35678 25098
rect 35702 25046 35712 25098
rect 35712 25046 35758 25098
rect 35782 25046 35828 25098
rect 35828 25046 35838 25098
rect 35862 25046 35892 25098
rect 35892 25046 35918 25098
rect 35622 25044 35678 25046
rect 35702 25044 35758 25046
rect 35782 25044 35838 25046
rect 35862 25044 35918 25046
rect 35622 24010 35678 24012
rect 35702 24010 35758 24012
rect 35782 24010 35838 24012
rect 35862 24010 35918 24012
rect 35622 23958 35648 24010
rect 35648 23958 35678 24010
rect 35702 23958 35712 24010
rect 35712 23958 35758 24010
rect 35782 23958 35828 24010
rect 35828 23958 35838 24010
rect 35862 23958 35892 24010
rect 35892 23958 35918 24010
rect 35622 23956 35678 23958
rect 35702 23956 35758 23958
rect 35782 23956 35838 23958
rect 35862 23956 35918 23958
rect 35622 22922 35678 22924
rect 35702 22922 35758 22924
rect 35782 22922 35838 22924
rect 35862 22922 35918 22924
rect 35622 22870 35648 22922
rect 35648 22870 35678 22922
rect 35702 22870 35712 22922
rect 35712 22870 35758 22922
rect 35782 22870 35828 22922
rect 35828 22870 35838 22922
rect 35862 22870 35892 22922
rect 35892 22870 35918 22922
rect 35622 22868 35678 22870
rect 35702 22868 35758 22870
rect 35782 22868 35838 22870
rect 35862 22868 35918 22870
rect 35622 21834 35678 21836
rect 35702 21834 35758 21836
rect 35782 21834 35838 21836
rect 35862 21834 35918 21836
rect 35622 21782 35648 21834
rect 35648 21782 35678 21834
rect 35702 21782 35712 21834
rect 35712 21782 35758 21834
rect 35782 21782 35828 21834
rect 35828 21782 35838 21834
rect 35862 21782 35892 21834
rect 35892 21782 35918 21834
rect 35622 21780 35678 21782
rect 35702 21780 35758 21782
rect 35782 21780 35838 21782
rect 35862 21780 35918 21782
rect 35622 20746 35678 20748
rect 35702 20746 35758 20748
rect 35782 20746 35838 20748
rect 35862 20746 35918 20748
rect 35622 20694 35648 20746
rect 35648 20694 35678 20746
rect 35702 20694 35712 20746
rect 35712 20694 35758 20746
rect 35782 20694 35828 20746
rect 35828 20694 35838 20746
rect 35862 20694 35892 20746
rect 35892 20694 35918 20746
rect 35622 20692 35678 20694
rect 35702 20692 35758 20694
rect 35782 20692 35838 20694
rect 35862 20692 35918 20694
rect 35622 19658 35678 19660
rect 35702 19658 35758 19660
rect 35782 19658 35838 19660
rect 35862 19658 35918 19660
rect 35622 19606 35648 19658
rect 35648 19606 35678 19658
rect 35702 19606 35712 19658
rect 35712 19606 35758 19658
rect 35782 19606 35828 19658
rect 35828 19606 35838 19658
rect 35862 19606 35892 19658
rect 35892 19606 35918 19658
rect 35622 19604 35678 19606
rect 35702 19604 35758 19606
rect 35782 19604 35838 19606
rect 35862 19604 35918 19606
rect 35622 18570 35678 18572
rect 35702 18570 35758 18572
rect 35782 18570 35838 18572
rect 35862 18570 35918 18572
rect 35622 18518 35648 18570
rect 35648 18518 35678 18570
rect 35702 18518 35712 18570
rect 35712 18518 35758 18570
rect 35782 18518 35828 18570
rect 35828 18518 35838 18570
rect 35862 18518 35892 18570
rect 35892 18518 35918 18570
rect 35622 18516 35678 18518
rect 35702 18516 35758 18518
rect 35782 18516 35838 18518
rect 35862 18516 35918 18518
rect 34412 18076 34414 18096
rect 34414 18076 34466 18096
rect 34466 18076 34468 18096
rect 34412 18040 34468 18076
rect 35622 17482 35678 17484
rect 35702 17482 35758 17484
rect 35782 17482 35838 17484
rect 35862 17482 35918 17484
rect 35622 17430 35648 17482
rect 35648 17430 35678 17482
rect 35702 17430 35712 17482
rect 35712 17430 35758 17482
rect 35782 17430 35828 17482
rect 35828 17430 35838 17482
rect 35862 17430 35892 17482
rect 35892 17430 35918 17482
rect 35622 17428 35678 17430
rect 35702 17428 35758 17430
rect 35782 17428 35838 17430
rect 35862 17428 35918 17430
rect 34412 16988 34414 17008
rect 34414 16988 34466 17008
rect 34466 16988 34468 17008
rect 34412 16952 34468 16988
rect 36988 21440 37044 21496
rect 36344 16544 36400 16600
rect 35622 16394 35678 16396
rect 35702 16394 35758 16396
rect 35782 16394 35838 16396
rect 35862 16394 35918 16396
rect 35622 16342 35648 16394
rect 35648 16342 35678 16394
rect 35702 16342 35712 16394
rect 35712 16342 35758 16394
rect 35782 16342 35828 16394
rect 35828 16342 35838 16394
rect 35862 16342 35892 16394
rect 35892 16342 35918 16394
rect 35622 16340 35678 16342
rect 35702 16340 35758 16342
rect 35782 16340 35838 16342
rect 35862 16340 35918 16342
rect 37816 29056 37872 29112
rect 38286 32170 38342 32172
rect 38366 32170 38422 32172
rect 38446 32170 38502 32172
rect 38526 32170 38582 32172
rect 38286 32118 38312 32170
rect 38312 32118 38342 32170
rect 38366 32118 38376 32170
rect 38376 32118 38422 32170
rect 38446 32118 38492 32170
rect 38492 32118 38502 32170
rect 38526 32118 38556 32170
rect 38556 32118 38582 32170
rect 38286 32116 38342 32118
rect 38366 32116 38422 32118
rect 38446 32116 38502 32118
rect 38526 32116 38582 32118
rect 40950 35978 41006 35980
rect 41030 35978 41086 35980
rect 41110 35978 41166 35980
rect 41190 35978 41246 35980
rect 40950 35926 40976 35978
rect 40976 35926 41006 35978
rect 41030 35926 41040 35978
rect 41040 35926 41086 35978
rect 41110 35926 41156 35978
rect 41156 35926 41166 35978
rect 41190 35926 41220 35978
rect 41220 35926 41246 35978
rect 40950 35924 41006 35926
rect 41030 35924 41086 35926
rect 41110 35924 41166 35926
rect 41190 35924 41246 35926
rect 40116 32864 40172 32920
rect 43614 35434 43670 35436
rect 43694 35434 43750 35436
rect 43774 35434 43830 35436
rect 43854 35434 43910 35436
rect 43614 35382 43640 35434
rect 43640 35382 43670 35434
rect 43694 35382 43704 35434
rect 43704 35382 43750 35434
rect 43774 35382 43820 35434
rect 43820 35382 43830 35434
rect 43854 35382 43884 35434
rect 43884 35382 43910 35434
rect 43614 35380 43670 35382
rect 43694 35380 43750 35382
rect 43774 35380 43830 35382
rect 43854 35380 43910 35382
rect 44256 36672 44312 36728
rect 45452 36808 45508 36864
rect 44256 36128 44312 36184
rect 40950 34890 41006 34892
rect 41030 34890 41086 34892
rect 41110 34890 41166 34892
rect 41190 34890 41246 34892
rect 40950 34838 40976 34890
rect 40976 34838 41006 34890
rect 41030 34838 41040 34890
rect 41040 34838 41086 34890
rect 41110 34838 41156 34890
rect 41156 34838 41166 34890
rect 41190 34838 41220 34890
rect 41220 34838 41246 34890
rect 40950 34836 41006 34838
rect 41030 34836 41086 34838
rect 41110 34836 41166 34838
rect 41190 34836 41246 34838
rect 40950 33802 41006 33804
rect 41030 33802 41086 33804
rect 41110 33802 41166 33804
rect 41190 33802 41246 33804
rect 40950 33750 40976 33802
rect 40976 33750 41006 33802
rect 41030 33750 41040 33802
rect 41040 33750 41086 33802
rect 41110 33750 41156 33802
rect 41156 33750 41166 33802
rect 41190 33750 41220 33802
rect 41220 33750 41246 33802
rect 40950 33748 41006 33750
rect 41030 33748 41086 33750
rect 41110 33748 41166 33750
rect 41190 33748 41246 33750
rect 40950 32714 41006 32716
rect 41030 32714 41086 32716
rect 41110 32714 41166 32716
rect 41190 32714 41246 32716
rect 40950 32662 40976 32714
rect 40976 32662 41006 32714
rect 41030 32662 41040 32714
rect 41040 32662 41086 32714
rect 41110 32662 41156 32714
rect 41156 32662 41166 32714
rect 41190 32662 41220 32714
rect 41220 32662 41246 32714
rect 40950 32660 41006 32662
rect 41030 32660 41086 32662
rect 41110 32660 41166 32662
rect 41190 32660 41246 32662
rect 41772 32320 41828 32376
rect 40950 31626 41006 31628
rect 41030 31626 41086 31628
rect 41110 31626 41166 31628
rect 41190 31626 41246 31628
rect 40950 31574 40976 31626
rect 40976 31574 41006 31626
rect 41030 31574 41040 31626
rect 41040 31574 41086 31626
rect 41110 31574 41156 31626
rect 41156 31574 41166 31626
rect 41190 31574 41220 31626
rect 41220 31574 41246 31626
rect 40950 31572 41006 31574
rect 41030 31572 41086 31574
rect 41110 31572 41166 31574
rect 41190 31572 41246 31574
rect 40852 31268 40854 31288
rect 40854 31268 40906 31288
rect 40906 31268 40908 31288
rect 40852 31232 40908 31268
rect 38286 31082 38342 31084
rect 38366 31082 38422 31084
rect 38446 31082 38502 31084
rect 38526 31082 38582 31084
rect 38286 31030 38312 31082
rect 38312 31030 38342 31082
rect 38366 31030 38376 31082
rect 38376 31030 38422 31082
rect 38446 31030 38492 31082
rect 38492 31030 38502 31082
rect 38526 31030 38556 31082
rect 38556 31030 38582 31082
rect 38286 31028 38342 31030
rect 38366 31028 38422 31030
rect 38446 31028 38502 31030
rect 38526 31028 38582 31030
rect 40950 30538 41006 30540
rect 41030 30538 41086 30540
rect 41110 30538 41166 30540
rect 41190 30538 41246 30540
rect 40950 30486 40976 30538
rect 40976 30486 41006 30538
rect 41030 30486 41040 30538
rect 41040 30486 41086 30538
rect 41110 30486 41156 30538
rect 41156 30486 41166 30538
rect 41190 30486 41220 30538
rect 41220 30486 41246 30538
rect 40950 30484 41006 30486
rect 41030 30484 41086 30486
rect 41110 30484 41166 30486
rect 41190 30484 41246 30486
rect 38286 29994 38342 29996
rect 38366 29994 38422 29996
rect 38446 29994 38502 29996
rect 38526 29994 38582 29996
rect 38286 29942 38312 29994
rect 38312 29942 38342 29994
rect 38366 29942 38376 29994
rect 38376 29942 38422 29994
rect 38446 29942 38492 29994
rect 38492 29942 38502 29994
rect 38526 29942 38556 29994
rect 38556 29942 38582 29994
rect 38286 29940 38342 29942
rect 38366 29940 38422 29942
rect 38446 29940 38502 29942
rect 38526 29940 38582 29942
rect 38276 29076 38332 29112
rect 38276 29056 38278 29076
rect 38278 29056 38330 29076
rect 38330 29056 38332 29076
rect 38286 28906 38342 28908
rect 38366 28906 38422 28908
rect 38446 28906 38502 28908
rect 38526 28906 38582 28908
rect 38286 28854 38312 28906
rect 38312 28854 38342 28906
rect 38366 28854 38376 28906
rect 38376 28854 38422 28906
rect 38446 28854 38492 28906
rect 38492 28854 38502 28906
rect 38526 28854 38556 28906
rect 38556 28854 38582 28906
rect 38286 28852 38342 28854
rect 38366 28852 38422 28854
rect 38446 28852 38502 28854
rect 38526 28852 38582 28854
rect 38286 27818 38342 27820
rect 38366 27818 38422 27820
rect 38446 27818 38502 27820
rect 38526 27818 38582 27820
rect 38286 27766 38312 27818
rect 38312 27766 38342 27818
rect 38366 27766 38376 27818
rect 38376 27766 38422 27818
rect 38446 27766 38492 27818
rect 38492 27766 38502 27818
rect 38526 27766 38556 27818
rect 38556 27766 38582 27818
rect 38286 27764 38342 27766
rect 38366 27764 38422 27766
rect 38446 27764 38502 27766
rect 38526 27764 38582 27766
rect 38286 26730 38342 26732
rect 38366 26730 38422 26732
rect 38446 26730 38502 26732
rect 38526 26730 38582 26732
rect 38286 26678 38312 26730
rect 38312 26678 38342 26730
rect 38366 26678 38376 26730
rect 38376 26678 38422 26730
rect 38446 26678 38492 26730
rect 38492 26678 38502 26730
rect 38526 26678 38556 26730
rect 38556 26678 38582 26730
rect 38286 26676 38342 26678
rect 38366 26676 38422 26678
rect 38446 26676 38502 26678
rect 38526 26676 38582 26678
rect 38286 25642 38342 25644
rect 38366 25642 38422 25644
rect 38446 25642 38502 25644
rect 38526 25642 38582 25644
rect 38286 25590 38312 25642
rect 38312 25590 38342 25642
rect 38366 25590 38376 25642
rect 38376 25590 38422 25642
rect 38446 25590 38492 25642
rect 38492 25590 38502 25642
rect 38526 25590 38556 25642
rect 38556 25590 38582 25642
rect 38286 25588 38342 25590
rect 38366 25588 38422 25590
rect 38446 25588 38502 25590
rect 38526 25588 38582 25590
rect 38286 24554 38342 24556
rect 38366 24554 38422 24556
rect 38446 24554 38502 24556
rect 38526 24554 38582 24556
rect 38286 24502 38312 24554
rect 38312 24502 38342 24554
rect 38366 24502 38376 24554
rect 38376 24502 38422 24554
rect 38446 24502 38492 24554
rect 38492 24502 38502 24554
rect 38526 24502 38556 24554
rect 38556 24502 38582 24554
rect 38286 24500 38342 24502
rect 38366 24500 38422 24502
rect 38446 24500 38502 24502
rect 38526 24500 38582 24502
rect 38286 23466 38342 23468
rect 38366 23466 38422 23468
rect 38446 23466 38502 23468
rect 38526 23466 38582 23468
rect 38286 23414 38312 23466
rect 38312 23414 38342 23466
rect 38366 23414 38376 23466
rect 38376 23414 38422 23466
rect 38446 23414 38492 23466
rect 38492 23414 38502 23466
rect 38526 23414 38556 23466
rect 38556 23414 38582 23466
rect 38286 23412 38342 23414
rect 38366 23412 38422 23414
rect 38446 23412 38502 23414
rect 38526 23412 38582 23414
rect 38286 22378 38342 22380
rect 38366 22378 38422 22380
rect 38446 22378 38502 22380
rect 38526 22378 38582 22380
rect 38286 22326 38312 22378
rect 38312 22326 38342 22378
rect 38366 22326 38376 22378
rect 38376 22326 38422 22378
rect 38446 22326 38492 22378
rect 38492 22326 38502 22378
rect 38526 22326 38556 22378
rect 38556 22326 38582 22378
rect 38286 22324 38342 22326
rect 38366 22324 38422 22326
rect 38446 22324 38502 22326
rect 38526 22324 38582 22326
rect 38286 21290 38342 21292
rect 38366 21290 38422 21292
rect 38446 21290 38502 21292
rect 38526 21290 38582 21292
rect 38286 21238 38312 21290
rect 38312 21238 38342 21290
rect 38366 21238 38376 21290
rect 38376 21238 38422 21290
rect 38446 21238 38492 21290
rect 38492 21238 38502 21290
rect 38526 21238 38556 21290
rect 38556 21238 38582 21290
rect 38286 21236 38342 21238
rect 38366 21236 38422 21238
rect 38446 21236 38502 21238
rect 38526 21236 38582 21238
rect 38286 20202 38342 20204
rect 38366 20202 38422 20204
rect 38446 20202 38502 20204
rect 38526 20202 38582 20204
rect 38286 20150 38312 20202
rect 38312 20150 38342 20202
rect 38366 20150 38376 20202
rect 38376 20150 38422 20202
rect 38446 20150 38492 20202
rect 38492 20150 38502 20202
rect 38526 20150 38556 20202
rect 38556 20150 38582 20202
rect 38286 20148 38342 20150
rect 38366 20148 38422 20150
rect 38446 20148 38502 20150
rect 38526 20148 38582 20150
rect 38286 19114 38342 19116
rect 38366 19114 38422 19116
rect 38446 19114 38502 19116
rect 38526 19114 38582 19116
rect 38286 19062 38312 19114
rect 38312 19062 38342 19114
rect 38366 19062 38376 19114
rect 38376 19062 38422 19114
rect 38446 19062 38492 19114
rect 38492 19062 38502 19114
rect 38526 19062 38556 19114
rect 38556 19062 38582 19114
rect 38286 19060 38342 19062
rect 38366 19060 38422 19062
rect 38446 19060 38502 19062
rect 38526 19060 38582 19062
rect 38286 18026 38342 18028
rect 38366 18026 38422 18028
rect 38446 18026 38502 18028
rect 38526 18026 38582 18028
rect 38286 17974 38312 18026
rect 38312 17974 38342 18026
rect 38366 17974 38376 18026
rect 38376 17974 38422 18026
rect 38446 17974 38492 18026
rect 38492 17974 38502 18026
rect 38526 17974 38556 18026
rect 38556 17974 38582 18026
rect 38286 17972 38342 17974
rect 38366 17972 38422 17974
rect 38446 17972 38502 17974
rect 38526 17972 38582 17974
rect 40950 29450 41006 29452
rect 41030 29450 41086 29452
rect 41110 29450 41166 29452
rect 41190 29450 41246 29452
rect 40950 29398 40976 29450
rect 40976 29398 41006 29450
rect 41030 29398 41040 29450
rect 41040 29398 41086 29450
rect 41110 29398 41156 29450
rect 41156 29398 41166 29450
rect 41190 29398 41220 29450
rect 41220 29398 41246 29450
rect 40950 29396 41006 29398
rect 41030 29396 41086 29398
rect 41110 29396 41166 29398
rect 41190 29396 41246 29398
rect 40950 28362 41006 28364
rect 41030 28362 41086 28364
rect 41110 28362 41166 28364
rect 41190 28362 41246 28364
rect 40950 28310 40976 28362
rect 40976 28310 41006 28362
rect 41030 28310 41040 28362
rect 41040 28310 41086 28362
rect 41110 28310 41156 28362
rect 41156 28310 41166 28362
rect 41190 28310 41220 28362
rect 41220 28310 41246 28362
rect 40950 28308 41006 28310
rect 41030 28308 41086 28310
rect 41110 28308 41166 28310
rect 41190 28308 41246 28310
rect 40950 27274 41006 27276
rect 41030 27274 41086 27276
rect 41110 27274 41166 27276
rect 41190 27274 41246 27276
rect 40950 27222 40976 27274
rect 40976 27222 41006 27274
rect 41030 27222 41040 27274
rect 41040 27222 41086 27274
rect 41110 27222 41156 27274
rect 41156 27222 41166 27274
rect 41190 27222 41220 27274
rect 41220 27222 41246 27274
rect 40950 27220 41006 27222
rect 41030 27220 41086 27222
rect 41110 27220 41166 27222
rect 41190 27220 41246 27222
rect 40950 26186 41006 26188
rect 41030 26186 41086 26188
rect 41110 26186 41166 26188
rect 41190 26186 41246 26188
rect 40950 26134 40976 26186
rect 40976 26134 41006 26186
rect 41030 26134 41040 26186
rect 41040 26134 41086 26186
rect 41110 26134 41156 26186
rect 41156 26134 41166 26186
rect 41190 26134 41220 26186
rect 41220 26134 41246 26186
rect 40950 26132 41006 26134
rect 41030 26132 41086 26134
rect 41110 26132 41166 26134
rect 41190 26132 41246 26134
rect 40950 25098 41006 25100
rect 41030 25098 41086 25100
rect 41110 25098 41166 25100
rect 41190 25098 41246 25100
rect 40950 25046 40976 25098
rect 40976 25046 41006 25098
rect 41030 25046 41040 25098
rect 41040 25046 41086 25098
rect 41110 25046 41156 25098
rect 41156 25046 41166 25098
rect 41190 25046 41220 25098
rect 41220 25046 41246 25098
rect 40950 25044 41006 25046
rect 41030 25044 41086 25046
rect 41110 25044 41166 25046
rect 41190 25044 41246 25046
rect 40950 24010 41006 24012
rect 41030 24010 41086 24012
rect 41110 24010 41166 24012
rect 41190 24010 41246 24012
rect 40950 23958 40976 24010
rect 40976 23958 41006 24010
rect 41030 23958 41040 24010
rect 41040 23958 41086 24010
rect 41110 23958 41156 24010
rect 41156 23958 41166 24010
rect 41190 23958 41220 24010
rect 41220 23958 41246 24010
rect 40950 23956 41006 23958
rect 41030 23956 41086 23958
rect 41110 23956 41166 23958
rect 41190 23956 41246 23958
rect 40950 22922 41006 22924
rect 41030 22922 41086 22924
rect 41110 22922 41166 22924
rect 41190 22922 41246 22924
rect 40950 22870 40976 22922
rect 40976 22870 41006 22922
rect 41030 22870 41040 22922
rect 41040 22870 41086 22922
rect 41110 22870 41156 22922
rect 41156 22870 41166 22922
rect 41190 22870 41220 22922
rect 41220 22870 41246 22922
rect 40950 22868 41006 22870
rect 41030 22868 41086 22870
rect 41110 22868 41166 22870
rect 41190 22868 41246 22870
rect 43060 22428 43062 22448
rect 43062 22428 43114 22448
rect 43114 22428 43116 22448
rect 43060 22392 43116 22428
rect 40950 21834 41006 21836
rect 41030 21834 41086 21836
rect 41110 21834 41166 21836
rect 41190 21834 41246 21836
rect 40950 21782 40976 21834
rect 40976 21782 41006 21834
rect 41030 21782 41040 21834
rect 41040 21782 41086 21834
rect 41110 21782 41156 21834
rect 41156 21782 41166 21834
rect 41190 21782 41220 21834
rect 41220 21782 41246 21834
rect 40950 21780 41006 21782
rect 41030 21780 41086 21782
rect 41110 21780 41166 21782
rect 41190 21780 41246 21782
rect 43060 21340 43062 21360
rect 43062 21340 43114 21360
rect 43114 21340 43116 21360
rect 43060 21304 43116 21340
rect 40950 20746 41006 20748
rect 41030 20746 41086 20748
rect 41110 20746 41166 20748
rect 41190 20746 41246 20748
rect 40950 20694 40976 20746
rect 40976 20694 41006 20746
rect 41030 20694 41040 20746
rect 41040 20694 41086 20746
rect 41110 20694 41156 20746
rect 41156 20694 41166 20746
rect 41190 20694 41220 20746
rect 41220 20694 41246 20746
rect 40950 20692 41006 20694
rect 41030 20692 41086 20694
rect 41110 20692 41166 20694
rect 41190 20692 41246 20694
rect 41496 19944 41552 20000
rect 43060 20252 43062 20272
rect 43062 20252 43114 20272
rect 43114 20252 43116 20272
rect 43060 20216 43116 20252
rect 40950 19658 41006 19660
rect 41030 19658 41086 19660
rect 41110 19658 41166 19660
rect 41190 19658 41246 19660
rect 40950 19606 40976 19658
rect 40976 19606 41006 19658
rect 41030 19606 41040 19658
rect 41040 19606 41086 19658
rect 41110 19606 41156 19658
rect 41156 19606 41166 19658
rect 41190 19606 41220 19658
rect 41220 19606 41246 19658
rect 40950 19604 41006 19606
rect 41030 19604 41086 19606
rect 41110 19604 41166 19606
rect 41190 19604 41246 19606
rect 42324 19128 42380 19184
rect 43614 34346 43670 34348
rect 43694 34346 43750 34348
rect 43774 34346 43830 34348
rect 43854 34346 43910 34348
rect 43614 34294 43640 34346
rect 43640 34294 43670 34346
rect 43694 34294 43704 34346
rect 43704 34294 43750 34346
rect 43774 34294 43820 34346
rect 43820 34294 43830 34346
rect 43854 34294 43884 34346
rect 43884 34294 43910 34346
rect 43614 34292 43670 34294
rect 43694 34292 43750 34294
rect 43774 34292 43830 34294
rect 43854 34292 43910 34294
rect 43614 33258 43670 33260
rect 43694 33258 43750 33260
rect 43774 33258 43830 33260
rect 43854 33258 43910 33260
rect 43614 33206 43640 33258
rect 43640 33206 43670 33258
rect 43694 33206 43704 33258
rect 43704 33206 43750 33258
rect 43774 33206 43820 33258
rect 43820 33206 43830 33258
rect 43854 33206 43884 33258
rect 43884 33206 43910 33258
rect 43614 33204 43670 33206
rect 43694 33204 43750 33206
rect 43774 33204 43830 33206
rect 43854 33204 43910 33206
rect 43614 32170 43670 32172
rect 43694 32170 43750 32172
rect 43774 32170 43830 32172
rect 43854 32170 43910 32172
rect 43614 32118 43640 32170
rect 43640 32118 43670 32170
rect 43694 32118 43704 32170
rect 43704 32118 43750 32170
rect 43774 32118 43820 32170
rect 43820 32118 43830 32170
rect 43854 32118 43884 32170
rect 43884 32118 43910 32170
rect 43614 32116 43670 32118
rect 43694 32116 43750 32118
rect 43774 32116 43830 32118
rect 43854 32116 43910 32118
rect 43614 31082 43670 31084
rect 43694 31082 43750 31084
rect 43774 31082 43830 31084
rect 43854 31082 43910 31084
rect 43614 31030 43640 31082
rect 43640 31030 43670 31082
rect 43694 31030 43704 31082
rect 43704 31030 43750 31082
rect 43774 31030 43820 31082
rect 43820 31030 43830 31082
rect 43854 31030 43884 31082
rect 43884 31030 43910 31082
rect 43614 31028 43670 31030
rect 43694 31028 43750 31030
rect 43774 31028 43830 31030
rect 43854 31028 43910 31030
rect 44992 33272 45048 33328
rect 44900 32884 44956 32920
rect 44900 32864 44902 32884
rect 44902 32864 44954 32884
rect 44954 32864 44956 32884
rect 46278 38154 46334 38156
rect 46358 38154 46414 38156
rect 46438 38154 46494 38156
rect 46518 38154 46574 38156
rect 46278 38102 46304 38154
rect 46304 38102 46334 38154
rect 46358 38102 46368 38154
rect 46368 38102 46414 38154
rect 46438 38102 46484 38154
rect 46484 38102 46494 38154
rect 46518 38102 46548 38154
rect 46548 38102 46574 38154
rect 46278 38100 46334 38102
rect 46358 38100 46414 38102
rect 46438 38100 46494 38102
rect 46518 38100 46574 38102
rect 46278 37066 46334 37068
rect 46358 37066 46414 37068
rect 46438 37066 46494 37068
rect 46518 37066 46574 37068
rect 46278 37014 46304 37066
rect 46304 37014 46334 37066
rect 46358 37014 46368 37066
rect 46368 37014 46414 37066
rect 46438 37014 46484 37066
rect 46484 37014 46494 37066
rect 46518 37014 46548 37066
rect 46548 37014 46574 37066
rect 46278 37012 46334 37014
rect 46358 37012 46414 37014
rect 46438 37012 46494 37014
rect 46518 37012 46574 37014
rect 51606 41418 51662 41420
rect 51686 41418 51742 41420
rect 51766 41418 51822 41420
rect 51846 41418 51902 41420
rect 51606 41366 51632 41418
rect 51632 41366 51662 41418
rect 51686 41366 51696 41418
rect 51696 41366 51742 41418
rect 51766 41366 51812 41418
rect 51812 41366 51822 41418
rect 51846 41366 51876 41418
rect 51876 41366 51902 41418
rect 51606 41364 51662 41366
rect 51686 41364 51742 41366
rect 51766 41364 51822 41366
rect 51846 41364 51902 41366
rect 54270 41962 54326 41964
rect 54350 41962 54406 41964
rect 54430 41962 54486 41964
rect 54510 41962 54566 41964
rect 54270 41910 54296 41962
rect 54296 41910 54326 41962
rect 54350 41910 54360 41962
rect 54360 41910 54406 41962
rect 54430 41910 54476 41962
rect 54476 41910 54486 41962
rect 54510 41910 54540 41962
rect 54540 41910 54566 41962
rect 54270 41908 54326 41910
rect 54350 41908 54406 41910
rect 54430 41908 54486 41910
rect 54510 41908 54566 41910
rect 48942 38698 48998 38700
rect 49022 38698 49078 38700
rect 49102 38698 49158 38700
rect 49182 38698 49238 38700
rect 48942 38646 48968 38698
rect 48968 38646 48998 38698
rect 49022 38646 49032 38698
rect 49032 38646 49078 38698
rect 49102 38646 49148 38698
rect 49148 38646 49158 38698
rect 49182 38646 49212 38698
rect 49212 38646 49238 38698
rect 48942 38644 48998 38646
rect 49022 38644 49078 38646
rect 49102 38644 49158 38646
rect 49182 38644 49238 38646
rect 54270 40874 54326 40876
rect 54350 40874 54406 40876
rect 54430 40874 54486 40876
rect 54510 40874 54566 40876
rect 54270 40822 54296 40874
rect 54296 40822 54326 40874
rect 54350 40822 54360 40874
rect 54360 40822 54406 40874
rect 54430 40822 54476 40874
rect 54476 40822 54486 40874
rect 54510 40822 54540 40874
rect 54540 40822 54566 40874
rect 54270 40820 54326 40822
rect 54350 40820 54406 40822
rect 54430 40820 54486 40822
rect 54510 40820 54566 40822
rect 51606 40330 51662 40332
rect 51686 40330 51742 40332
rect 51766 40330 51822 40332
rect 51846 40330 51902 40332
rect 51606 40278 51632 40330
rect 51632 40278 51662 40330
rect 51686 40278 51696 40330
rect 51696 40278 51742 40330
rect 51766 40278 51812 40330
rect 51812 40278 51822 40330
rect 51846 40278 51876 40330
rect 51876 40278 51902 40330
rect 51606 40276 51662 40278
rect 51686 40276 51742 40278
rect 51766 40276 51822 40278
rect 51846 40276 51902 40278
rect 56934 41418 56990 41420
rect 57014 41418 57070 41420
rect 57094 41418 57150 41420
rect 57174 41418 57230 41420
rect 56934 41366 56960 41418
rect 56960 41366 56990 41418
rect 57014 41366 57024 41418
rect 57024 41366 57070 41418
rect 57094 41366 57140 41418
rect 57140 41366 57150 41418
rect 57174 41366 57204 41418
rect 57204 41366 57230 41418
rect 56934 41364 56990 41366
rect 57014 41364 57070 41366
rect 57094 41364 57150 41366
rect 57174 41364 57230 41366
rect 54270 39786 54326 39788
rect 54350 39786 54406 39788
rect 54430 39786 54486 39788
rect 54510 39786 54566 39788
rect 54270 39734 54296 39786
rect 54296 39734 54326 39786
rect 54350 39734 54360 39786
rect 54360 39734 54406 39786
rect 54430 39734 54476 39786
rect 54476 39734 54486 39786
rect 54510 39734 54540 39786
rect 54540 39734 54566 39786
rect 54270 39732 54326 39734
rect 54350 39732 54406 39734
rect 54430 39732 54486 39734
rect 54510 39732 54566 39734
rect 51606 39242 51662 39244
rect 51686 39242 51742 39244
rect 51766 39242 51822 39244
rect 51846 39242 51902 39244
rect 51606 39190 51632 39242
rect 51632 39190 51662 39242
rect 51686 39190 51696 39242
rect 51696 39190 51742 39242
rect 51766 39190 51812 39242
rect 51812 39190 51822 39242
rect 51846 39190 51876 39242
rect 51876 39190 51902 39242
rect 51606 39188 51662 39190
rect 51686 39188 51742 39190
rect 51766 39188 51822 39190
rect 51846 39188 51902 39190
rect 46924 37216 46980 37272
rect 51606 38154 51662 38156
rect 51686 38154 51742 38156
rect 51766 38154 51822 38156
rect 51846 38154 51902 38156
rect 51606 38102 51632 38154
rect 51632 38102 51662 38154
rect 51686 38102 51696 38154
rect 51696 38102 51742 38154
rect 51766 38102 51812 38154
rect 51812 38102 51822 38154
rect 51846 38102 51876 38154
rect 51876 38102 51902 38154
rect 51606 38100 51662 38102
rect 51686 38100 51742 38102
rect 51766 38100 51822 38102
rect 51846 38100 51902 38102
rect 48942 37610 48998 37612
rect 49022 37610 49078 37612
rect 49102 37610 49158 37612
rect 49182 37610 49238 37612
rect 48942 37558 48968 37610
rect 48968 37558 48998 37610
rect 49022 37558 49032 37610
rect 49032 37558 49078 37610
rect 49102 37558 49148 37610
rect 49148 37558 49158 37610
rect 49182 37558 49212 37610
rect 49212 37558 49238 37610
rect 48942 37556 48998 37558
rect 49022 37556 49078 37558
rect 49102 37556 49158 37558
rect 49182 37556 49238 37558
rect 46278 35978 46334 35980
rect 46358 35978 46414 35980
rect 46438 35978 46494 35980
rect 46518 35978 46574 35980
rect 46278 35926 46304 35978
rect 46304 35926 46334 35978
rect 46358 35926 46368 35978
rect 46368 35926 46414 35978
rect 46438 35926 46484 35978
rect 46484 35926 46494 35978
rect 46518 35926 46548 35978
rect 46548 35926 46574 35978
rect 46278 35924 46334 35926
rect 46358 35924 46414 35926
rect 46438 35924 46494 35926
rect 46518 35924 46574 35926
rect 46278 34890 46334 34892
rect 46358 34890 46414 34892
rect 46438 34890 46494 34892
rect 46518 34890 46574 34892
rect 46278 34838 46304 34890
rect 46304 34838 46334 34890
rect 46358 34838 46368 34890
rect 46368 34838 46414 34890
rect 46438 34838 46484 34890
rect 46484 34838 46494 34890
rect 46518 34838 46548 34890
rect 46548 34838 46574 34890
rect 46278 34836 46334 34838
rect 46358 34836 46414 34838
rect 46438 34836 46494 34838
rect 46518 34836 46574 34838
rect 46278 33802 46334 33804
rect 46358 33802 46414 33804
rect 46438 33802 46494 33804
rect 46518 33802 46574 33804
rect 46278 33750 46304 33802
rect 46304 33750 46334 33802
rect 46358 33750 46368 33802
rect 46368 33750 46414 33802
rect 46438 33750 46484 33802
rect 46484 33750 46494 33802
rect 46518 33750 46548 33802
rect 46548 33750 46574 33802
rect 46278 33748 46334 33750
rect 46358 33748 46414 33750
rect 46438 33748 46494 33750
rect 46518 33748 46574 33750
rect 47016 34632 47072 34688
rect 47660 36708 47662 36728
rect 47662 36708 47714 36728
rect 47714 36708 47716 36728
rect 47660 36672 47716 36708
rect 50420 37236 50476 37272
rect 50420 37216 50422 37236
rect 50422 37216 50474 37236
rect 50474 37216 50476 37236
rect 54270 38698 54326 38700
rect 54350 38698 54406 38700
rect 54430 38698 54486 38700
rect 54510 38698 54566 38700
rect 54270 38646 54296 38698
rect 54296 38646 54326 38698
rect 54350 38646 54360 38698
rect 54360 38646 54406 38698
rect 54430 38646 54476 38698
rect 54476 38646 54486 38698
rect 54510 38646 54540 38698
rect 54540 38646 54566 38698
rect 54270 38644 54326 38646
rect 54350 38644 54406 38646
rect 54430 38644 54486 38646
rect 54510 38644 54566 38646
rect 51606 37066 51662 37068
rect 51686 37066 51742 37068
rect 51766 37066 51822 37068
rect 51846 37066 51902 37068
rect 51606 37014 51632 37066
rect 51632 37014 51662 37066
rect 51686 37014 51696 37066
rect 51696 37014 51742 37066
rect 51766 37014 51812 37066
rect 51812 37014 51822 37066
rect 51846 37014 51876 37066
rect 51876 37014 51902 37066
rect 51606 37012 51662 37014
rect 51686 37012 51742 37014
rect 51766 37012 51822 37014
rect 51846 37012 51902 37014
rect 50420 36536 50476 36592
rect 48942 36522 48998 36524
rect 49022 36522 49078 36524
rect 49102 36522 49158 36524
rect 49182 36522 49238 36524
rect 48942 36470 48968 36522
rect 48968 36470 48998 36522
rect 49022 36470 49032 36522
rect 49032 36470 49078 36522
rect 49102 36470 49148 36522
rect 49148 36470 49158 36522
rect 49182 36470 49212 36522
rect 49212 36470 49238 36522
rect 48942 36468 48998 36470
rect 49022 36468 49078 36470
rect 49102 36468 49158 36470
rect 49182 36468 49238 36470
rect 51800 36808 51856 36864
rect 51432 36672 51488 36728
rect 48942 35434 48998 35436
rect 49022 35434 49078 35436
rect 49102 35434 49158 35436
rect 49182 35434 49238 35436
rect 48942 35382 48968 35434
rect 48968 35382 48998 35434
rect 49022 35382 49032 35434
rect 49032 35382 49078 35434
rect 49102 35382 49148 35434
rect 49148 35382 49158 35434
rect 49182 35382 49212 35434
rect 49212 35382 49238 35434
rect 48942 35380 48998 35382
rect 49022 35380 49078 35382
rect 49102 35380 49158 35382
rect 49182 35380 49238 35382
rect 52352 36808 52408 36864
rect 54270 37610 54326 37612
rect 54350 37610 54406 37612
rect 54430 37610 54486 37612
rect 54510 37610 54566 37612
rect 54270 37558 54296 37610
rect 54296 37558 54326 37610
rect 54350 37558 54360 37610
rect 54360 37558 54406 37610
rect 54430 37558 54476 37610
rect 54476 37558 54486 37610
rect 54510 37558 54540 37610
rect 54540 37558 54566 37610
rect 54270 37556 54326 37558
rect 54350 37556 54406 37558
rect 54430 37556 54486 37558
rect 54510 37556 54566 37558
rect 56934 40330 56990 40332
rect 57014 40330 57070 40332
rect 57094 40330 57150 40332
rect 57174 40330 57230 40332
rect 56934 40278 56960 40330
rect 56960 40278 56990 40330
rect 57014 40278 57024 40330
rect 57024 40278 57070 40330
rect 57094 40278 57140 40330
rect 57140 40278 57150 40330
rect 57174 40278 57204 40330
rect 57204 40278 57230 40330
rect 56934 40276 56990 40278
rect 57014 40276 57070 40278
rect 57094 40276 57150 40278
rect 57174 40276 57230 40278
rect 55480 39020 55482 39040
rect 55482 39020 55534 39040
rect 55534 39020 55536 39040
rect 55480 38984 55536 39020
rect 52536 37216 52592 37272
rect 53456 36672 53512 36728
rect 52720 36536 52776 36592
rect 54270 36522 54326 36524
rect 54350 36522 54406 36524
rect 54430 36522 54486 36524
rect 54510 36522 54566 36524
rect 54270 36470 54296 36522
rect 54296 36470 54326 36522
rect 54350 36470 54360 36522
rect 54360 36470 54406 36522
rect 54430 36470 54476 36522
rect 54476 36470 54486 36522
rect 54510 36470 54540 36522
rect 54540 36470 54566 36522
rect 54270 36468 54326 36470
rect 54350 36468 54406 36470
rect 54430 36468 54486 36470
rect 54510 36468 54566 36470
rect 51606 35978 51662 35980
rect 51686 35978 51742 35980
rect 51766 35978 51822 35980
rect 51846 35978 51902 35980
rect 51606 35926 51632 35978
rect 51632 35926 51662 35978
rect 51686 35926 51696 35978
rect 51696 35926 51742 35978
rect 51766 35926 51812 35978
rect 51812 35926 51822 35978
rect 51846 35926 51876 35978
rect 51876 35926 51902 35978
rect 51606 35924 51662 35926
rect 51686 35924 51742 35926
rect 51766 35924 51822 35926
rect 51846 35924 51902 35926
rect 51524 35720 51580 35776
rect 51606 34890 51662 34892
rect 51686 34890 51742 34892
rect 51766 34890 51822 34892
rect 51846 34890 51902 34892
rect 51606 34838 51632 34890
rect 51632 34838 51662 34890
rect 51686 34838 51696 34890
rect 51696 34838 51742 34890
rect 51766 34838 51812 34890
rect 51812 34838 51822 34890
rect 51846 34838 51876 34890
rect 51876 34838 51902 34890
rect 51606 34836 51662 34838
rect 51686 34836 51742 34838
rect 51766 34836 51822 34838
rect 51846 34836 51902 34838
rect 48942 34346 48998 34348
rect 49022 34346 49078 34348
rect 49102 34346 49158 34348
rect 49182 34346 49238 34348
rect 48942 34294 48968 34346
rect 48968 34294 48998 34346
rect 49022 34294 49032 34346
rect 49032 34294 49078 34346
rect 49102 34294 49148 34346
rect 49148 34294 49158 34346
rect 49182 34294 49212 34346
rect 49212 34294 49238 34346
rect 48942 34292 48998 34294
rect 49022 34292 49078 34294
rect 49102 34292 49158 34294
rect 49182 34292 49238 34294
rect 46740 32764 46742 32784
rect 46742 32764 46794 32784
rect 46794 32764 46796 32784
rect 46740 32728 46796 32764
rect 46278 32714 46334 32716
rect 46358 32714 46414 32716
rect 46438 32714 46494 32716
rect 46518 32714 46574 32716
rect 46278 32662 46304 32714
rect 46304 32662 46334 32714
rect 46358 32662 46368 32714
rect 46368 32662 46414 32714
rect 46438 32662 46484 32714
rect 46484 32662 46494 32714
rect 46518 32662 46548 32714
rect 46548 32662 46574 32714
rect 46278 32660 46334 32662
rect 46358 32660 46414 32662
rect 46438 32660 46494 32662
rect 46518 32660 46574 32662
rect 46464 32184 46520 32240
rect 47108 33272 47164 33328
rect 51606 33802 51662 33804
rect 51686 33802 51742 33804
rect 51766 33802 51822 33804
rect 51846 33802 51902 33804
rect 51606 33750 51632 33802
rect 51632 33750 51662 33802
rect 51686 33750 51696 33802
rect 51696 33750 51742 33802
rect 51766 33750 51812 33802
rect 51812 33750 51822 33802
rect 51846 33750 51876 33802
rect 51876 33750 51902 33802
rect 51606 33748 51662 33750
rect 51686 33748 51742 33750
rect 51766 33748 51822 33750
rect 51846 33748 51902 33750
rect 47292 32900 47294 32920
rect 47294 32900 47346 32920
rect 47346 32900 47348 32920
rect 47292 32864 47348 32900
rect 47384 32728 47440 32784
rect 47568 32764 47570 32784
rect 47570 32764 47622 32784
rect 47622 32764 47624 32784
rect 47568 32728 47624 32764
rect 47200 32356 47202 32376
rect 47202 32356 47254 32376
rect 47254 32356 47256 32376
rect 46278 31626 46334 31628
rect 46358 31626 46414 31628
rect 46438 31626 46494 31628
rect 46518 31626 46574 31628
rect 46278 31574 46304 31626
rect 46304 31574 46334 31626
rect 46358 31574 46368 31626
rect 46368 31574 46414 31626
rect 46438 31574 46484 31626
rect 46484 31574 46494 31626
rect 46518 31574 46548 31626
rect 46548 31574 46574 31626
rect 46278 31572 46334 31574
rect 46358 31572 46414 31574
rect 46438 31572 46494 31574
rect 46518 31572 46574 31574
rect 46464 31388 46520 31424
rect 46464 31368 46466 31388
rect 46466 31368 46518 31388
rect 46518 31368 46520 31388
rect 47200 32320 47256 32356
rect 48396 32492 48398 32512
rect 48398 32492 48450 32512
rect 48450 32492 48452 32512
rect 48396 32456 48452 32492
rect 48942 33258 48998 33260
rect 49022 33258 49078 33260
rect 49102 33258 49158 33260
rect 49182 33258 49238 33260
rect 48942 33206 48968 33258
rect 48968 33206 48998 33258
rect 49022 33206 49032 33258
rect 49032 33206 49078 33258
rect 49102 33206 49148 33258
rect 49148 33206 49158 33258
rect 49182 33206 49212 33258
rect 49212 33206 49238 33258
rect 48942 33204 48998 33206
rect 49022 33204 49078 33206
rect 49102 33204 49158 33206
rect 49182 33204 49238 33206
rect 47568 32220 47570 32240
rect 47570 32220 47622 32240
rect 47622 32220 47624 32240
rect 47568 32184 47624 32220
rect 47936 32320 47992 32376
rect 43614 29994 43670 29996
rect 43694 29994 43750 29996
rect 43774 29994 43830 29996
rect 43854 29994 43910 29996
rect 43614 29942 43640 29994
rect 43640 29942 43670 29994
rect 43694 29942 43704 29994
rect 43704 29942 43750 29994
rect 43774 29942 43820 29994
rect 43820 29942 43830 29994
rect 43854 29942 43884 29994
rect 43884 29942 43910 29994
rect 43614 29940 43670 29942
rect 43694 29940 43750 29942
rect 43774 29940 43830 29942
rect 43854 29940 43910 29942
rect 43614 28906 43670 28908
rect 43694 28906 43750 28908
rect 43774 28906 43830 28908
rect 43854 28906 43910 28908
rect 43614 28854 43640 28906
rect 43640 28854 43670 28906
rect 43694 28854 43704 28906
rect 43704 28854 43750 28906
rect 43774 28854 43820 28906
rect 43820 28854 43830 28906
rect 43854 28854 43884 28906
rect 43884 28854 43910 28906
rect 43614 28852 43670 28854
rect 43694 28852 43750 28854
rect 43774 28852 43830 28854
rect 43854 28852 43910 28854
rect 43614 27818 43670 27820
rect 43694 27818 43750 27820
rect 43774 27818 43830 27820
rect 43854 27818 43910 27820
rect 43614 27766 43640 27818
rect 43640 27766 43670 27818
rect 43694 27766 43704 27818
rect 43704 27766 43750 27818
rect 43774 27766 43820 27818
rect 43820 27766 43830 27818
rect 43854 27766 43884 27818
rect 43884 27766 43910 27818
rect 43614 27764 43670 27766
rect 43694 27764 43750 27766
rect 43774 27764 43830 27766
rect 43854 27764 43910 27766
rect 46278 30538 46334 30540
rect 46358 30538 46414 30540
rect 46438 30538 46494 30540
rect 46518 30538 46574 30540
rect 46278 30486 46304 30538
rect 46304 30486 46334 30538
rect 46358 30486 46368 30538
rect 46368 30486 46414 30538
rect 46438 30486 46484 30538
rect 46484 30486 46494 30538
rect 46518 30486 46548 30538
rect 46548 30486 46574 30538
rect 46278 30484 46334 30486
rect 46358 30484 46414 30486
rect 46438 30484 46494 30486
rect 46518 30484 46574 30486
rect 46278 29450 46334 29452
rect 46358 29450 46414 29452
rect 46438 29450 46494 29452
rect 46518 29450 46574 29452
rect 46278 29398 46304 29450
rect 46304 29398 46334 29450
rect 46358 29398 46368 29450
rect 46368 29398 46414 29450
rect 46438 29398 46484 29450
rect 46484 29398 46494 29450
rect 46518 29398 46548 29450
rect 46548 29398 46574 29450
rect 46278 29396 46334 29398
rect 46358 29396 46414 29398
rect 46438 29396 46494 29398
rect 46518 29396 46574 29398
rect 46004 29056 46060 29112
rect 46278 28362 46334 28364
rect 46358 28362 46414 28364
rect 46438 28362 46494 28364
rect 46518 28362 46574 28364
rect 46278 28310 46304 28362
rect 46304 28310 46334 28362
rect 46358 28310 46368 28362
rect 46368 28310 46414 28362
rect 46438 28310 46484 28362
rect 46484 28310 46494 28362
rect 46518 28310 46548 28362
rect 46548 28310 46574 28362
rect 46278 28308 46334 28310
rect 46358 28308 46414 28310
rect 46438 28308 46494 28310
rect 46518 28308 46574 28310
rect 43614 26730 43670 26732
rect 43694 26730 43750 26732
rect 43774 26730 43830 26732
rect 43854 26730 43910 26732
rect 43614 26678 43640 26730
rect 43640 26678 43670 26730
rect 43694 26678 43704 26730
rect 43704 26678 43750 26730
rect 43774 26678 43820 26730
rect 43820 26678 43830 26730
rect 43854 26678 43884 26730
rect 43884 26678 43910 26730
rect 43614 26676 43670 26678
rect 43694 26676 43750 26678
rect 43774 26676 43830 26678
rect 43854 26676 43910 26678
rect 48942 32170 48998 32172
rect 49022 32170 49078 32172
rect 49102 32170 49158 32172
rect 49182 32170 49238 32172
rect 48942 32118 48968 32170
rect 48968 32118 48998 32170
rect 49022 32118 49032 32170
rect 49032 32118 49078 32170
rect 49102 32118 49148 32170
rect 49148 32118 49158 32170
rect 49182 32118 49212 32170
rect 49212 32118 49238 32170
rect 48942 32116 48998 32118
rect 49022 32116 49078 32118
rect 49102 32116 49158 32118
rect 49182 32116 49238 32118
rect 51606 32714 51662 32716
rect 51686 32714 51742 32716
rect 51766 32714 51822 32716
rect 51846 32714 51902 32716
rect 51606 32662 51632 32714
rect 51632 32662 51662 32714
rect 51686 32662 51696 32714
rect 51696 32662 51742 32714
rect 51766 32662 51812 32714
rect 51812 32662 51822 32714
rect 51846 32662 51876 32714
rect 51876 32662 51902 32714
rect 51606 32660 51662 32662
rect 51686 32660 51742 32662
rect 51766 32660 51822 32662
rect 51846 32660 51902 32662
rect 52812 32456 52868 32512
rect 51606 31626 51662 31628
rect 51686 31626 51742 31628
rect 51766 31626 51822 31628
rect 51846 31626 51902 31628
rect 51606 31574 51632 31626
rect 51632 31574 51662 31626
rect 51686 31574 51696 31626
rect 51696 31574 51742 31626
rect 51766 31574 51812 31626
rect 51812 31574 51822 31626
rect 51846 31574 51876 31626
rect 51876 31574 51902 31626
rect 51606 31572 51662 31574
rect 51686 31572 51742 31574
rect 51766 31572 51822 31574
rect 51846 31572 51902 31574
rect 48942 31082 48998 31084
rect 49022 31082 49078 31084
rect 49102 31082 49158 31084
rect 49182 31082 49238 31084
rect 48942 31030 48968 31082
rect 48968 31030 48998 31082
rect 49022 31030 49032 31082
rect 49032 31030 49078 31082
rect 49102 31030 49148 31082
rect 49148 31030 49158 31082
rect 49182 31030 49212 31082
rect 49212 31030 49238 31082
rect 48942 31028 48998 31030
rect 49022 31028 49078 31030
rect 49102 31028 49158 31030
rect 49182 31028 49238 31030
rect 48212 27968 48268 28024
rect 48396 27424 48452 27480
rect 46278 27274 46334 27276
rect 46358 27274 46414 27276
rect 46438 27274 46494 27276
rect 46518 27274 46574 27276
rect 46278 27222 46304 27274
rect 46304 27222 46334 27274
rect 46358 27222 46368 27274
rect 46368 27222 46414 27274
rect 46438 27222 46484 27274
rect 46484 27222 46494 27274
rect 46518 27222 46548 27274
rect 46548 27222 46574 27274
rect 46278 27220 46334 27222
rect 46358 27220 46414 27222
rect 46438 27220 46494 27222
rect 46518 27220 46574 27222
rect 48942 29994 48998 29996
rect 49022 29994 49078 29996
rect 49102 29994 49158 29996
rect 49182 29994 49238 29996
rect 48942 29942 48968 29994
rect 48968 29942 48998 29994
rect 49022 29942 49032 29994
rect 49032 29942 49078 29994
rect 49102 29942 49148 29994
rect 49148 29942 49158 29994
rect 49182 29942 49212 29994
rect 49212 29942 49238 29994
rect 48942 29940 48998 29942
rect 49022 29940 49078 29942
rect 49102 29940 49158 29942
rect 49182 29940 49238 29942
rect 48942 28906 48998 28908
rect 49022 28906 49078 28908
rect 49102 28906 49158 28908
rect 49182 28906 49238 28908
rect 48942 28854 48968 28906
rect 48968 28854 48998 28906
rect 49022 28854 49032 28906
rect 49032 28854 49078 28906
rect 49102 28854 49148 28906
rect 49148 28854 49158 28906
rect 49182 28854 49212 28906
rect 49212 28854 49238 28906
rect 48942 28852 48998 28854
rect 49022 28852 49078 28854
rect 49102 28852 49158 28854
rect 49182 28852 49238 28854
rect 48942 27818 48998 27820
rect 49022 27818 49078 27820
rect 49102 27818 49158 27820
rect 49182 27818 49238 27820
rect 48942 27766 48968 27818
rect 48968 27766 48998 27818
rect 49022 27766 49032 27818
rect 49032 27766 49078 27818
rect 49102 27766 49148 27818
rect 49148 27766 49158 27818
rect 49182 27766 49212 27818
rect 49212 27766 49238 27818
rect 48942 27764 48998 27766
rect 49022 27764 49078 27766
rect 49102 27764 49158 27766
rect 49182 27764 49238 27766
rect 51606 30538 51662 30540
rect 51686 30538 51742 30540
rect 51766 30538 51822 30540
rect 51846 30538 51902 30540
rect 51606 30486 51632 30538
rect 51632 30486 51662 30538
rect 51686 30486 51696 30538
rect 51696 30486 51742 30538
rect 51766 30486 51812 30538
rect 51812 30486 51822 30538
rect 51846 30486 51876 30538
rect 51876 30486 51902 30538
rect 51606 30484 51662 30486
rect 51686 30484 51742 30486
rect 51766 30484 51822 30486
rect 51846 30484 51902 30486
rect 52168 30860 52170 30880
rect 52170 30860 52222 30880
rect 52222 30860 52224 30880
rect 52168 30824 52224 30860
rect 54270 35434 54326 35436
rect 54350 35434 54406 35436
rect 54430 35434 54486 35436
rect 54510 35434 54566 35436
rect 54270 35382 54296 35434
rect 54296 35382 54326 35434
rect 54350 35382 54360 35434
rect 54360 35382 54406 35434
rect 54430 35382 54476 35434
rect 54476 35382 54486 35434
rect 54510 35382 54540 35434
rect 54540 35382 54566 35434
rect 54270 35380 54326 35382
rect 54350 35380 54406 35382
rect 54430 35380 54486 35382
rect 54510 35380 54566 35382
rect 54270 34346 54326 34348
rect 54350 34346 54406 34348
rect 54430 34346 54486 34348
rect 54510 34346 54566 34348
rect 54270 34294 54296 34346
rect 54296 34294 54326 34346
rect 54350 34294 54360 34346
rect 54360 34294 54406 34346
rect 54430 34294 54476 34346
rect 54476 34294 54486 34346
rect 54510 34294 54540 34346
rect 54540 34294 54566 34346
rect 54270 34292 54326 34294
rect 54350 34292 54406 34294
rect 54430 34292 54486 34294
rect 54510 34292 54566 34294
rect 54270 33258 54326 33260
rect 54350 33258 54406 33260
rect 54430 33258 54486 33260
rect 54510 33258 54566 33260
rect 54270 33206 54296 33258
rect 54296 33206 54326 33258
rect 54350 33206 54360 33258
rect 54360 33206 54406 33258
rect 54430 33206 54476 33258
rect 54476 33206 54486 33258
rect 54510 33206 54540 33258
rect 54540 33206 54566 33258
rect 54270 33204 54326 33206
rect 54350 33204 54406 33206
rect 54430 33204 54486 33206
rect 54510 33204 54566 33206
rect 56934 39242 56990 39244
rect 57014 39242 57070 39244
rect 57094 39242 57150 39244
rect 57174 39242 57230 39244
rect 56934 39190 56960 39242
rect 56960 39190 56990 39242
rect 57014 39190 57024 39242
rect 57024 39190 57070 39242
rect 57094 39190 57140 39242
rect 57140 39190 57150 39242
rect 57174 39190 57204 39242
rect 57204 39190 57230 39242
rect 56934 39188 56990 39190
rect 57014 39188 57070 39190
rect 57094 39188 57150 39190
rect 57174 39188 57230 39190
rect 56934 38154 56990 38156
rect 57014 38154 57070 38156
rect 57094 38154 57150 38156
rect 57174 38154 57230 38156
rect 56934 38102 56960 38154
rect 56960 38102 56990 38154
rect 57014 38102 57024 38154
rect 57024 38102 57070 38154
rect 57094 38102 57140 38154
rect 57140 38102 57150 38154
rect 57174 38102 57204 38154
rect 57204 38102 57230 38154
rect 56934 38100 56990 38102
rect 57014 38100 57070 38102
rect 57094 38100 57150 38102
rect 57174 38100 57230 38102
rect 56934 37066 56990 37068
rect 57014 37066 57070 37068
rect 57094 37066 57150 37068
rect 57174 37066 57230 37068
rect 56934 37014 56960 37066
rect 56960 37014 56990 37066
rect 57014 37014 57024 37066
rect 57024 37014 57070 37066
rect 57094 37014 57140 37066
rect 57140 37014 57150 37066
rect 57174 37014 57204 37066
rect 57204 37014 57230 37066
rect 56934 37012 56990 37014
rect 57014 37012 57070 37014
rect 57094 37012 57150 37014
rect 57174 37012 57230 37014
rect 56934 35978 56990 35980
rect 57014 35978 57070 35980
rect 57094 35978 57150 35980
rect 57174 35978 57230 35980
rect 56934 35926 56960 35978
rect 56960 35926 56990 35978
rect 57014 35926 57024 35978
rect 57024 35926 57070 35978
rect 57094 35926 57140 35978
rect 57140 35926 57150 35978
rect 57174 35926 57204 35978
rect 57204 35926 57230 35978
rect 56934 35924 56990 35926
rect 57014 35924 57070 35926
rect 57094 35924 57150 35926
rect 57174 35924 57230 35926
rect 56676 35720 56732 35776
rect 56934 34890 56990 34892
rect 57014 34890 57070 34892
rect 57094 34890 57150 34892
rect 57174 34890 57230 34892
rect 56934 34838 56960 34890
rect 56960 34838 56990 34890
rect 57014 34838 57024 34890
rect 57024 34838 57070 34890
rect 57094 34838 57140 34890
rect 57140 34838 57150 34890
rect 57174 34838 57204 34890
rect 57204 34838 57230 34890
rect 56934 34836 56990 34838
rect 57014 34836 57070 34838
rect 57094 34836 57150 34838
rect 57174 34836 57230 34838
rect 56934 33802 56990 33804
rect 57014 33802 57070 33804
rect 57094 33802 57150 33804
rect 57174 33802 57230 33804
rect 56934 33750 56960 33802
rect 56960 33750 56990 33802
rect 57014 33750 57024 33802
rect 57024 33750 57070 33802
rect 57094 33750 57140 33802
rect 57140 33750 57150 33802
rect 57174 33750 57204 33802
rect 57204 33750 57230 33802
rect 56934 33748 56990 33750
rect 57014 33748 57070 33750
rect 57094 33748 57150 33750
rect 57174 33748 57230 33750
rect 59598 41962 59654 41964
rect 59678 41962 59734 41964
rect 59758 41962 59814 41964
rect 59838 41962 59894 41964
rect 59598 41910 59624 41962
rect 59624 41910 59654 41962
rect 59678 41910 59688 41962
rect 59688 41910 59734 41962
rect 59758 41910 59804 41962
rect 59804 41910 59814 41962
rect 59838 41910 59868 41962
rect 59868 41910 59894 41962
rect 59598 41908 59654 41910
rect 59678 41908 59734 41910
rect 59758 41908 59814 41910
rect 59838 41908 59894 41910
rect 62262 41418 62318 41420
rect 62342 41418 62398 41420
rect 62422 41418 62478 41420
rect 62502 41418 62558 41420
rect 62262 41366 62288 41418
rect 62288 41366 62318 41418
rect 62342 41366 62352 41418
rect 62352 41366 62398 41418
rect 62422 41366 62468 41418
rect 62468 41366 62478 41418
rect 62502 41366 62532 41418
rect 62532 41366 62558 41418
rect 62262 41364 62318 41366
rect 62342 41364 62398 41366
rect 62422 41364 62478 41366
rect 62502 41364 62558 41366
rect 59598 40874 59654 40876
rect 59678 40874 59734 40876
rect 59758 40874 59814 40876
rect 59838 40874 59894 40876
rect 59598 40822 59624 40874
rect 59624 40822 59654 40874
rect 59678 40822 59688 40874
rect 59688 40822 59734 40874
rect 59758 40822 59804 40874
rect 59804 40822 59814 40874
rect 59838 40822 59868 40874
rect 59868 40822 59894 40874
rect 59598 40820 59654 40822
rect 59678 40820 59734 40822
rect 59758 40820 59814 40822
rect 59838 40820 59894 40822
rect 59598 39786 59654 39788
rect 59678 39786 59734 39788
rect 59758 39786 59814 39788
rect 59838 39786 59894 39788
rect 59598 39734 59624 39786
rect 59624 39734 59654 39786
rect 59678 39734 59688 39786
rect 59688 39734 59734 39786
rect 59758 39734 59804 39786
rect 59804 39734 59814 39786
rect 59838 39734 59868 39786
rect 59868 39734 59894 39786
rect 59598 39732 59654 39734
rect 59678 39732 59734 39734
rect 59758 39732 59814 39734
rect 59838 39732 59894 39734
rect 59598 38698 59654 38700
rect 59678 38698 59734 38700
rect 59758 38698 59814 38700
rect 59838 38698 59894 38700
rect 59598 38646 59624 38698
rect 59624 38646 59654 38698
rect 59678 38646 59688 38698
rect 59688 38646 59734 38698
rect 59758 38646 59804 38698
rect 59804 38646 59814 38698
rect 59838 38646 59868 38698
rect 59868 38646 59894 38698
rect 59598 38644 59654 38646
rect 59678 38644 59734 38646
rect 59758 38644 59814 38646
rect 59838 38644 59894 38646
rect 57872 37760 57928 37816
rect 57780 37080 57836 37136
rect 57688 36692 57744 36728
rect 57688 36672 57690 36692
rect 57690 36672 57742 36692
rect 57742 36672 57744 36692
rect 57964 37236 58020 37272
rect 57964 37216 57966 37236
rect 57966 37216 58018 37236
rect 58018 37216 58020 37236
rect 58424 36692 58480 36728
rect 58424 36672 58426 36692
rect 58426 36672 58478 36692
rect 58478 36672 58480 36692
rect 59598 37610 59654 37612
rect 59678 37610 59734 37612
rect 59758 37610 59814 37612
rect 59838 37610 59894 37612
rect 59598 37558 59624 37610
rect 59624 37558 59654 37610
rect 59678 37558 59688 37610
rect 59688 37558 59734 37610
rect 59758 37558 59804 37610
rect 59804 37558 59814 37610
rect 59838 37558 59868 37610
rect 59868 37558 59894 37610
rect 59598 37556 59654 37558
rect 59678 37556 59734 37558
rect 59758 37556 59814 37558
rect 59838 37556 59894 37558
rect 62262 40330 62318 40332
rect 62342 40330 62398 40332
rect 62422 40330 62478 40332
rect 62502 40330 62558 40332
rect 62262 40278 62288 40330
rect 62288 40278 62318 40330
rect 62342 40278 62352 40330
rect 62352 40278 62398 40330
rect 62422 40278 62468 40330
rect 62468 40278 62478 40330
rect 62502 40278 62532 40330
rect 62532 40278 62558 40330
rect 62262 40276 62318 40278
rect 62342 40276 62398 40278
rect 62422 40276 62478 40278
rect 62502 40276 62558 40278
rect 62262 39242 62318 39244
rect 62342 39242 62398 39244
rect 62422 39242 62478 39244
rect 62502 39242 62558 39244
rect 62262 39190 62288 39242
rect 62288 39190 62318 39242
rect 62342 39190 62352 39242
rect 62352 39190 62398 39242
rect 62422 39190 62468 39242
rect 62468 39190 62478 39242
rect 62502 39190 62532 39242
rect 62532 39190 62558 39242
rect 62262 39188 62318 39190
rect 62342 39188 62398 39190
rect 62422 39188 62478 39190
rect 62502 39188 62558 39190
rect 62262 38154 62318 38156
rect 62342 38154 62398 38156
rect 62422 38154 62478 38156
rect 62502 38154 62558 38156
rect 62262 38102 62288 38154
rect 62288 38102 62318 38154
rect 62342 38102 62352 38154
rect 62352 38102 62398 38154
rect 62422 38102 62468 38154
rect 62468 38102 62478 38154
rect 62502 38102 62532 38154
rect 62532 38102 62558 38154
rect 62262 38100 62318 38102
rect 62342 38100 62398 38102
rect 62422 38100 62478 38102
rect 62502 38100 62558 38102
rect 59620 37252 59622 37272
rect 59622 37252 59674 37272
rect 59674 37252 59676 37272
rect 59620 37216 59676 37252
rect 62104 37116 62106 37136
rect 62106 37116 62158 37136
rect 62158 37116 62160 37136
rect 62104 37080 62160 37116
rect 62262 37066 62318 37068
rect 62342 37066 62398 37068
rect 62422 37066 62478 37068
rect 62502 37066 62558 37068
rect 62262 37014 62288 37066
rect 62288 37014 62318 37066
rect 62342 37014 62352 37066
rect 62352 37014 62398 37066
rect 62422 37014 62468 37066
rect 62468 37014 62478 37066
rect 62502 37014 62532 37066
rect 62532 37014 62558 37066
rect 62262 37012 62318 37014
rect 62342 37012 62398 37014
rect 62422 37012 62478 37014
rect 62502 37012 62558 37014
rect 59598 36522 59654 36524
rect 59678 36522 59734 36524
rect 59758 36522 59814 36524
rect 59838 36522 59894 36524
rect 59598 36470 59624 36522
rect 59624 36470 59654 36522
rect 59678 36470 59688 36522
rect 59688 36470 59734 36522
rect 59758 36470 59804 36522
rect 59804 36470 59814 36522
rect 59838 36470 59868 36522
rect 59868 36470 59894 36522
rect 59598 36468 59654 36470
rect 59678 36468 59734 36470
rect 59758 36468 59814 36470
rect 59838 36468 59894 36470
rect 57872 35740 57928 35776
rect 57872 35720 57874 35740
rect 57874 35720 57926 35740
rect 57926 35720 57928 35740
rect 62564 36148 62620 36184
rect 62564 36128 62566 36148
rect 62566 36128 62618 36148
rect 62618 36128 62620 36148
rect 62262 35978 62318 35980
rect 62342 35978 62398 35980
rect 62422 35978 62478 35980
rect 62502 35978 62558 35980
rect 62262 35926 62288 35978
rect 62288 35926 62318 35978
rect 62342 35926 62352 35978
rect 62352 35926 62398 35978
rect 62422 35926 62468 35978
rect 62468 35926 62478 35978
rect 62502 35926 62532 35978
rect 62532 35926 62558 35978
rect 62262 35924 62318 35926
rect 62342 35924 62398 35926
rect 62422 35924 62478 35926
rect 62502 35924 62558 35926
rect 59598 35434 59654 35436
rect 59678 35434 59734 35436
rect 59758 35434 59814 35436
rect 59838 35434 59894 35436
rect 59598 35382 59624 35434
rect 59624 35382 59654 35434
rect 59678 35382 59688 35434
rect 59688 35382 59734 35434
rect 59758 35382 59804 35434
rect 59804 35382 59814 35434
rect 59838 35382 59868 35434
rect 59868 35382 59894 35434
rect 59598 35380 59654 35382
rect 59678 35380 59734 35382
rect 59758 35380 59814 35382
rect 59838 35380 59894 35382
rect 58424 34532 58426 34552
rect 58426 34532 58478 34552
rect 58478 34532 58480 34552
rect 58424 34496 58480 34532
rect 59598 34346 59654 34348
rect 59678 34346 59734 34348
rect 59758 34346 59814 34348
rect 59838 34346 59894 34348
rect 59598 34294 59624 34346
rect 59624 34294 59654 34346
rect 59678 34294 59688 34346
rect 59688 34294 59734 34346
rect 59758 34294 59804 34346
rect 59804 34294 59814 34346
rect 59838 34294 59868 34346
rect 59868 34294 59894 34346
rect 59598 34292 59654 34294
rect 59678 34292 59734 34294
rect 59758 34292 59814 34294
rect 59838 34292 59894 34294
rect 56934 32714 56990 32716
rect 57014 32714 57070 32716
rect 57094 32714 57150 32716
rect 57174 32714 57230 32716
rect 56934 32662 56960 32714
rect 56960 32662 56990 32714
rect 57014 32662 57024 32714
rect 57024 32662 57070 32714
rect 57094 32662 57140 32714
rect 57140 32662 57150 32714
rect 57174 32662 57204 32714
rect 57204 32662 57230 32714
rect 56934 32660 56990 32662
rect 57014 32660 57070 32662
rect 57094 32660 57150 32662
rect 57174 32660 57230 32662
rect 57872 32592 57928 32648
rect 58792 32864 58848 32920
rect 60816 35312 60872 35368
rect 59598 33258 59654 33260
rect 59678 33258 59734 33260
rect 59758 33258 59814 33260
rect 59838 33258 59894 33260
rect 59598 33206 59624 33258
rect 59624 33206 59654 33258
rect 59678 33206 59688 33258
rect 59688 33206 59734 33258
rect 59758 33206 59804 33258
rect 59804 33206 59814 33258
rect 59838 33206 59868 33258
rect 59868 33206 59894 33258
rect 59598 33204 59654 33206
rect 59678 33204 59734 33206
rect 59758 33204 59814 33206
rect 59838 33204 59894 33206
rect 60908 33544 60964 33600
rect 62380 35448 62436 35504
rect 62262 34890 62318 34892
rect 62342 34890 62398 34892
rect 62422 34890 62478 34892
rect 62502 34890 62558 34892
rect 62262 34838 62288 34890
rect 62288 34838 62318 34890
rect 62342 34838 62352 34890
rect 62352 34838 62398 34890
rect 62422 34838 62468 34890
rect 62468 34838 62478 34890
rect 62502 34838 62532 34890
rect 62532 34838 62558 34890
rect 62262 34836 62318 34838
rect 62342 34836 62398 34838
rect 62422 34836 62478 34838
rect 62502 34836 62558 34838
rect 62262 33802 62318 33804
rect 62342 33802 62398 33804
rect 62422 33802 62478 33804
rect 62502 33802 62558 33804
rect 62262 33750 62288 33802
rect 62288 33750 62318 33802
rect 62342 33750 62352 33802
rect 62352 33750 62398 33802
rect 62422 33750 62468 33802
rect 62468 33750 62478 33802
rect 62502 33750 62532 33802
rect 62532 33750 62558 33802
rect 62262 33748 62318 33750
rect 62342 33748 62398 33750
rect 62422 33748 62478 33750
rect 62502 33748 62558 33750
rect 62656 33680 62712 33736
rect 59804 32456 59860 32512
rect 58424 32220 58426 32240
rect 58426 32220 58478 32240
rect 58478 32220 58480 32240
rect 58424 32184 58480 32220
rect 54270 32170 54326 32172
rect 54350 32170 54406 32172
rect 54430 32170 54486 32172
rect 54510 32170 54566 32172
rect 54270 32118 54296 32170
rect 54296 32118 54326 32170
rect 54350 32118 54360 32170
rect 54360 32118 54406 32170
rect 54430 32118 54476 32170
rect 54476 32118 54486 32170
rect 54510 32118 54540 32170
rect 54540 32118 54566 32170
rect 54270 32116 54326 32118
rect 54350 32116 54406 32118
rect 54430 32116 54486 32118
rect 54510 32116 54566 32118
rect 58700 32184 58756 32240
rect 60080 32184 60136 32240
rect 59598 32170 59654 32172
rect 59678 32170 59734 32172
rect 59758 32170 59814 32172
rect 59838 32170 59894 32172
rect 59598 32118 59624 32170
rect 59624 32118 59654 32170
rect 59678 32118 59688 32170
rect 59688 32118 59734 32170
rect 59758 32118 59804 32170
rect 59804 32118 59814 32170
rect 59838 32118 59868 32170
rect 59868 32118 59894 32170
rect 59598 32116 59654 32118
rect 59678 32116 59734 32118
rect 59758 32116 59814 32118
rect 59838 32116 59894 32118
rect 58608 31948 58610 31968
rect 58610 31948 58662 31968
rect 58662 31948 58664 31968
rect 58608 31912 58664 31948
rect 62262 32714 62318 32716
rect 62342 32714 62398 32716
rect 62422 32714 62478 32716
rect 62502 32714 62558 32716
rect 62262 32662 62288 32714
rect 62288 32662 62318 32714
rect 62342 32662 62352 32714
rect 62352 32662 62398 32714
rect 62422 32662 62468 32714
rect 62468 32662 62478 32714
rect 62502 32662 62532 32714
rect 62532 32662 62558 32714
rect 62262 32660 62318 32662
rect 62342 32660 62398 32662
rect 62422 32660 62478 32662
rect 62502 32660 62558 32662
rect 62012 32592 62068 32648
rect 57596 31776 57652 31832
rect 56934 31626 56990 31628
rect 57014 31626 57070 31628
rect 57094 31626 57150 31628
rect 57174 31626 57230 31628
rect 56934 31574 56960 31626
rect 56960 31574 56990 31626
rect 57014 31574 57024 31626
rect 57024 31574 57070 31626
rect 57094 31574 57140 31626
rect 57140 31574 57150 31626
rect 57174 31574 57204 31626
rect 57204 31574 57230 31626
rect 56934 31572 56990 31574
rect 57014 31572 57070 31574
rect 57094 31572 57150 31574
rect 57174 31572 57230 31574
rect 50420 27832 50476 27888
rect 52260 29620 52316 29656
rect 52260 29600 52262 29620
rect 52262 29600 52314 29620
rect 52314 29600 52316 29620
rect 51606 29450 51662 29452
rect 51686 29450 51742 29452
rect 51766 29450 51822 29452
rect 51846 29450 51902 29452
rect 51606 29398 51632 29450
rect 51632 29398 51662 29450
rect 51686 29398 51696 29450
rect 51696 29398 51742 29450
rect 51766 29398 51812 29450
rect 51812 29398 51822 29450
rect 51846 29398 51876 29450
rect 51876 29398 51902 29450
rect 51606 29396 51662 29398
rect 51686 29396 51742 29398
rect 51766 29396 51822 29398
rect 51846 29396 51902 29398
rect 52076 28668 52132 28704
rect 52076 28648 52078 28668
rect 52078 28648 52130 28668
rect 52130 28648 52132 28668
rect 51606 28362 51662 28364
rect 51686 28362 51742 28364
rect 51766 28362 51822 28364
rect 51846 28362 51902 28364
rect 51606 28310 51632 28362
rect 51632 28310 51662 28362
rect 51686 28310 51696 28362
rect 51696 28310 51742 28362
rect 51766 28310 51812 28362
rect 51812 28310 51822 28362
rect 51846 28310 51876 28362
rect 51876 28310 51902 28362
rect 51606 28308 51662 28310
rect 51686 28308 51742 28310
rect 51766 28308 51822 28310
rect 51846 28308 51902 28310
rect 51524 27968 51580 28024
rect 51156 27832 51212 27888
rect 51064 27016 51120 27072
rect 51606 27274 51662 27276
rect 51686 27274 51742 27276
rect 51766 27274 51822 27276
rect 51846 27274 51902 27276
rect 51606 27222 51632 27274
rect 51632 27222 51662 27274
rect 51686 27222 51696 27274
rect 51696 27222 51742 27274
rect 51766 27222 51812 27274
rect 51812 27222 51822 27274
rect 51846 27222 51876 27274
rect 51876 27222 51902 27274
rect 51606 27220 51662 27222
rect 51686 27220 51742 27222
rect 51766 27220 51822 27222
rect 51846 27220 51902 27222
rect 53916 30824 53972 30880
rect 54744 31388 54800 31424
rect 54744 31368 54746 31388
rect 54746 31368 54798 31388
rect 54798 31368 54800 31388
rect 57504 31268 57506 31288
rect 57506 31268 57558 31288
rect 57558 31268 57560 31288
rect 57504 31232 57560 31268
rect 54270 31082 54326 31084
rect 54350 31082 54406 31084
rect 54430 31082 54486 31084
rect 54510 31082 54566 31084
rect 54270 31030 54296 31082
rect 54296 31030 54326 31082
rect 54350 31030 54360 31082
rect 54360 31030 54406 31082
rect 54430 31030 54476 31082
rect 54476 31030 54486 31082
rect 54510 31030 54540 31082
rect 54540 31030 54566 31082
rect 54270 31028 54326 31030
rect 54350 31028 54406 31030
rect 54430 31028 54486 31030
rect 54510 31028 54566 31030
rect 52628 29076 52684 29112
rect 52628 29056 52630 29076
rect 52630 29056 52682 29076
rect 52682 29056 52684 29076
rect 52996 28648 53052 28704
rect 54270 29994 54326 29996
rect 54350 29994 54406 29996
rect 54430 29994 54486 29996
rect 54510 29994 54566 29996
rect 54270 29942 54296 29994
rect 54296 29942 54326 29994
rect 54350 29942 54360 29994
rect 54360 29942 54406 29994
rect 54430 29942 54476 29994
rect 54476 29942 54486 29994
rect 54510 29942 54540 29994
rect 54540 29942 54566 29994
rect 54270 29940 54326 29942
rect 54350 29940 54406 29942
rect 54430 29940 54486 29942
rect 54510 29940 54566 29942
rect 58884 31776 58940 31832
rect 56934 30538 56990 30540
rect 57014 30538 57070 30540
rect 57094 30538 57150 30540
rect 57174 30538 57230 30540
rect 56934 30486 56960 30538
rect 56960 30486 56990 30538
rect 57014 30486 57024 30538
rect 57024 30486 57070 30538
rect 57094 30486 57140 30538
rect 57140 30486 57150 30538
rect 57174 30486 57204 30538
rect 57204 30486 57230 30538
rect 56934 30484 56990 30486
rect 57014 30484 57070 30486
rect 57094 30484 57150 30486
rect 57174 30484 57230 30486
rect 54468 29620 54524 29656
rect 54468 29600 54470 29620
rect 54470 29600 54522 29620
rect 54522 29600 54524 29620
rect 54270 28906 54326 28908
rect 54350 28906 54406 28908
rect 54430 28906 54486 28908
rect 54510 28906 54566 28908
rect 54270 28854 54296 28906
rect 54296 28854 54326 28906
rect 54350 28854 54360 28906
rect 54360 28854 54406 28906
rect 54430 28854 54476 28906
rect 54476 28854 54486 28906
rect 54510 28854 54540 28906
rect 54540 28854 54566 28906
rect 54270 28852 54326 28854
rect 54350 28852 54406 28854
rect 54430 28852 54486 28854
rect 54510 28852 54566 28854
rect 56934 29450 56990 29452
rect 57014 29450 57070 29452
rect 57094 29450 57150 29452
rect 57174 29450 57230 29452
rect 56934 29398 56960 29450
rect 56960 29398 56990 29450
rect 57014 29398 57024 29450
rect 57024 29398 57070 29450
rect 57094 29398 57140 29450
rect 57140 29398 57150 29450
rect 57174 29398 57204 29450
rect 57204 29398 57230 29450
rect 56934 29396 56990 29398
rect 57014 29396 57070 29398
rect 57094 29396 57150 29398
rect 57174 29396 57230 29398
rect 56584 29056 56640 29112
rect 52904 27424 52960 27480
rect 52904 27052 52906 27072
rect 52906 27052 52958 27072
rect 52958 27052 52960 27072
rect 52904 27016 52960 27052
rect 54008 27832 54064 27888
rect 54270 27818 54326 27820
rect 54350 27818 54406 27820
rect 54430 27818 54486 27820
rect 54510 27818 54566 27820
rect 54270 27766 54296 27818
rect 54296 27766 54326 27818
rect 54350 27766 54360 27818
rect 54360 27766 54406 27818
rect 54430 27766 54476 27818
rect 54476 27766 54486 27818
rect 54510 27766 54540 27818
rect 54540 27766 54566 27818
rect 54270 27764 54326 27766
rect 54350 27764 54406 27766
rect 54430 27764 54486 27766
rect 54510 27764 54566 27766
rect 56934 28362 56990 28364
rect 57014 28362 57070 28364
rect 57094 28362 57150 28364
rect 57174 28362 57230 28364
rect 56934 28310 56960 28362
rect 56960 28310 56990 28362
rect 57014 28310 57024 28362
rect 57024 28310 57070 28362
rect 57094 28310 57140 28362
rect 57140 28310 57150 28362
rect 57174 28310 57204 28362
rect 57204 28310 57230 28362
rect 56934 28308 56990 28310
rect 57014 28308 57070 28310
rect 57094 28308 57150 28310
rect 57174 28308 57230 28310
rect 56934 27274 56990 27276
rect 57014 27274 57070 27276
rect 57094 27274 57150 27276
rect 57174 27274 57230 27276
rect 56934 27222 56960 27274
rect 56960 27222 56990 27274
rect 57014 27222 57024 27274
rect 57024 27222 57070 27274
rect 57094 27222 57140 27274
rect 57140 27222 57150 27274
rect 57174 27222 57204 27274
rect 57204 27222 57230 27274
rect 56934 27220 56990 27222
rect 57014 27220 57070 27222
rect 57094 27220 57150 27222
rect 57174 27220 57230 27222
rect 63024 36128 63080 36184
rect 64926 41962 64982 41964
rect 65006 41962 65062 41964
rect 65086 41962 65142 41964
rect 65166 41962 65222 41964
rect 64926 41910 64952 41962
rect 64952 41910 64982 41962
rect 65006 41910 65016 41962
rect 65016 41910 65062 41962
rect 65086 41910 65132 41962
rect 65132 41910 65142 41962
rect 65166 41910 65196 41962
rect 65196 41910 65222 41962
rect 64926 41908 64982 41910
rect 65006 41908 65062 41910
rect 65086 41908 65142 41910
rect 65166 41908 65222 41910
rect 64926 40874 64982 40876
rect 65006 40874 65062 40876
rect 65086 40874 65142 40876
rect 65166 40874 65222 40876
rect 64926 40822 64952 40874
rect 64952 40822 64982 40874
rect 65006 40822 65016 40874
rect 65016 40822 65062 40874
rect 65086 40822 65132 40874
rect 65132 40822 65142 40874
rect 65166 40822 65196 40874
rect 65196 40822 65222 40874
rect 64926 40820 64982 40822
rect 65006 40820 65062 40822
rect 65086 40820 65142 40822
rect 65166 40820 65222 40822
rect 64926 39786 64982 39788
rect 65006 39786 65062 39788
rect 65086 39786 65142 39788
rect 65166 39786 65222 39788
rect 64926 39734 64952 39786
rect 64952 39734 64982 39786
rect 65006 39734 65016 39786
rect 65016 39734 65062 39786
rect 65086 39734 65132 39786
rect 65132 39734 65142 39786
rect 65166 39734 65196 39786
rect 65196 39734 65222 39786
rect 64926 39732 64982 39734
rect 65006 39732 65062 39734
rect 65086 39732 65142 39734
rect 65166 39732 65222 39734
rect 67590 41418 67646 41420
rect 67670 41418 67726 41420
rect 67750 41418 67806 41420
rect 67830 41418 67886 41420
rect 67590 41366 67616 41418
rect 67616 41366 67646 41418
rect 67670 41366 67680 41418
rect 67680 41366 67726 41418
rect 67750 41366 67796 41418
rect 67796 41366 67806 41418
rect 67830 41366 67860 41418
rect 67860 41366 67886 41418
rect 67590 41364 67646 41366
rect 67670 41364 67726 41366
rect 67750 41364 67806 41366
rect 67830 41364 67886 41366
rect 67590 40330 67646 40332
rect 67670 40330 67726 40332
rect 67750 40330 67806 40332
rect 67830 40330 67886 40332
rect 67590 40278 67616 40330
rect 67616 40278 67646 40330
rect 67670 40278 67680 40330
rect 67680 40278 67726 40330
rect 67750 40278 67796 40330
rect 67796 40278 67806 40330
rect 67830 40278 67860 40330
rect 67860 40278 67886 40330
rect 67590 40276 67646 40278
rect 67670 40276 67726 40278
rect 67750 40276 67806 40278
rect 67830 40276 67886 40278
rect 67808 39548 67864 39584
rect 67808 39528 67810 39548
rect 67810 39528 67862 39548
rect 67862 39528 67864 39548
rect 67590 39242 67646 39244
rect 67670 39242 67726 39244
rect 67750 39242 67806 39244
rect 67830 39242 67886 39244
rect 67590 39190 67616 39242
rect 67616 39190 67646 39242
rect 67670 39190 67680 39242
rect 67680 39190 67726 39242
rect 67750 39190 67796 39242
rect 67796 39190 67806 39242
rect 67830 39190 67860 39242
rect 67860 39190 67886 39242
rect 67590 39188 67646 39190
rect 67670 39188 67726 39190
rect 67750 39188 67806 39190
rect 67830 39188 67886 39190
rect 64926 38698 64982 38700
rect 65006 38698 65062 38700
rect 65086 38698 65142 38700
rect 65166 38698 65222 38700
rect 64926 38646 64952 38698
rect 64952 38646 64982 38698
rect 65006 38646 65016 38698
rect 65016 38646 65062 38698
rect 65086 38646 65132 38698
rect 65132 38646 65142 38698
rect 65166 38646 65196 38698
rect 65196 38646 65222 38698
rect 64926 38644 64982 38646
rect 65006 38644 65062 38646
rect 65086 38644 65142 38646
rect 65166 38644 65222 38646
rect 67590 38154 67646 38156
rect 67670 38154 67726 38156
rect 67750 38154 67806 38156
rect 67830 38154 67886 38156
rect 67590 38102 67616 38154
rect 67616 38102 67646 38154
rect 67670 38102 67680 38154
rect 67680 38102 67726 38154
rect 67750 38102 67796 38154
rect 67796 38102 67806 38154
rect 67830 38102 67860 38154
rect 67860 38102 67886 38154
rect 67590 38100 67646 38102
rect 67670 38100 67726 38102
rect 67750 38100 67806 38102
rect 67830 38100 67886 38102
rect 64926 37610 64982 37612
rect 65006 37610 65062 37612
rect 65086 37610 65142 37612
rect 65166 37610 65222 37612
rect 64926 37558 64952 37610
rect 64952 37558 64982 37610
rect 65006 37558 65016 37610
rect 65016 37558 65062 37610
rect 65086 37558 65132 37610
rect 65132 37558 65142 37610
rect 65166 37558 65196 37610
rect 65196 37558 65222 37610
rect 64926 37556 64982 37558
rect 65006 37556 65062 37558
rect 65086 37556 65142 37558
rect 65166 37556 65222 37558
rect 67590 37066 67646 37068
rect 67670 37066 67726 37068
rect 67750 37066 67806 37068
rect 67830 37066 67886 37068
rect 67590 37014 67616 37066
rect 67616 37014 67646 37066
rect 67670 37014 67680 37066
rect 67680 37014 67726 37066
rect 67750 37014 67796 37066
rect 67796 37014 67806 37066
rect 67830 37014 67860 37066
rect 67860 37014 67886 37066
rect 67590 37012 67646 37014
rect 67670 37012 67726 37014
rect 67750 37012 67806 37014
rect 67830 37012 67886 37014
rect 64926 36522 64982 36524
rect 65006 36522 65062 36524
rect 65086 36522 65142 36524
rect 65166 36522 65222 36524
rect 64926 36470 64952 36522
rect 64952 36470 64982 36522
rect 65006 36470 65016 36522
rect 65016 36470 65062 36522
rect 65086 36470 65132 36522
rect 65132 36470 65142 36522
rect 65166 36470 65196 36522
rect 65196 36470 65222 36522
rect 64926 36468 64982 36470
rect 65006 36468 65062 36470
rect 65086 36468 65142 36470
rect 65166 36468 65222 36470
rect 63300 35312 63356 35368
rect 63944 35448 64000 35504
rect 64926 35434 64982 35436
rect 65006 35434 65062 35436
rect 65086 35434 65142 35436
rect 65166 35434 65222 35436
rect 64926 35382 64952 35434
rect 64952 35382 64982 35434
rect 65006 35382 65016 35434
rect 65016 35382 65062 35434
rect 65086 35382 65132 35434
rect 65132 35382 65142 35434
rect 65166 35382 65196 35434
rect 65196 35382 65222 35434
rect 64926 35380 64982 35382
rect 65006 35380 65062 35382
rect 65086 35380 65142 35382
rect 65166 35380 65222 35382
rect 63208 32728 63264 32784
rect 63392 32592 63448 32648
rect 60172 31268 60174 31288
rect 60174 31268 60226 31288
rect 60226 31268 60228 31288
rect 60172 31232 60228 31268
rect 59598 31082 59654 31084
rect 59678 31082 59734 31084
rect 59758 31082 59814 31084
rect 59838 31082 59894 31084
rect 59598 31030 59624 31082
rect 59624 31030 59654 31082
rect 59678 31030 59688 31082
rect 59688 31030 59734 31082
rect 59758 31030 59804 31082
rect 59804 31030 59814 31082
rect 59838 31030 59868 31082
rect 59868 31030 59894 31082
rect 59598 31028 59654 31030
rect 59678 31028 59734 31030
rect 59758 31028 59814 31030
rect 59838 31028 59894 31030
rect 59988 30180 59990 30200
rect 59990 30180 60042 30200
rect 60042 30180 60044 30200
rect 59988 30144 60044 30180
rect 59598 29994 59654 29996
rect 59678 29994 59734 29996
rect 59758 29994 59814 29996
rect 59838 29994 59894 29996
rect 59598 29942 59624 29994
rect 59624 29942 59654 29994
rect 59678 29942 59688 29994
rect 59688 29942 59734 29994
rect 59758 29942 59804 29994
rect 59804 29942 59814 29994
rect 59838 29942 59868 29994
rect 59868 29942 59894 29994
rect 59598 29940 59654 29942
rect 59678 29940 59734 29942
rect 59758 29940 59814 29942
rect 59838 29940 59894 29942
rect 60356 29192 60412 29248
rect 59598 28906 59654 28908
rect 59678 28906 59734 28908
rect 59758 28906 59814 28908
rect 59838 28906 59894 28908
rect 59598 28854 59624 28906
rect 59624 28854 59654 28906
rect 59678 28854 59688 28906
rect 59688 28854 59734 28906
rect 59758 28854 59804 28906
rect 59804 28854 59814 28906
rect 59838 28854 59868 28906
rect 59868 28854 59894 28906
rect 59598 28852 59654 28854
rect 59678 28852 59734 28854
rect 59758 28852 59814 28854
rect 59838 28852 59894 28854
rect 63300 32048 63356 32104
rect 64128 34496 64184 34552
rect 64926 34346 64982 34348
rect 65006 34346 65062 34348
rect 65086 34346 65142 34348
rect 65166 34346 65222 34348
rect 64926 34294 64952 34346
rect 64952 34294 64982 34346
rect 65006 34294 65016 34346
rect 65016 34294 65062 34346
rect 65086 34294 65132 34346
rect 65132 34294 65142 34346
rect 65166 34294 65196 34346
rect 65196 34294 65222 34346
rect 64926 34292 64982 34294
rect 65006 34292 65062 34294
rect 65086 34292 65142 34294
rect 65166 34292 65222 34294
rect 64926 33258 64982 33260
rect 65006 33258 65062 33260
rect 65086 33258 65142 33260
rect 65166 33258 65222 33260
rect 64926 33206 64952 33258
rect 64952 33206 64982 33258
rect 65006 33206 65016 33258
rect 65016 33206 65062 33258
rect 65086 33206 65132 33258
rect 65132 33206 65142 33258
rect 65166 33206 65196 33258
rect 65196 33206 65222 33258
rect 64926 33204 64982 33206
rect 65006 33204 65062 33206
rect 65086 33204 65142 33206
rect 65166 33204 65222 33206
rect 64680 32884 64736 32920
rect 64680 32864 64682 32884
rect 64682 32864 64734 32884
rect 64734 32864 64736 32884
rect 64128 32728 64184 32784
rect 64680 32592 64736 32648
rect 64496 32184 64552 32240
rect 64680 32048 64736 32104
rect 62262 31626 62318 31628
rect 62342 31626 62398 31628
rect 62422 31626 62478 31628
rect 62502 31626 62558 31628
rect 62262 31574 62288 31626
rect 62288 31574 62318 31626
rect 62342 31574 62352 31626
rect 62352 31574 62398 31626
rect 62422 31574 62468 31626
rect 62468 31574 62478 31626
rect 62502 31574 62532 31626
rect 62532 31574 62558 31626
rect 62262 31572 62318 31574
rect 62342 31572 62398 31574
rect 62422 31572 62478 31574
rect 62502 31572 62558 31574
rect 62262 30538 62318 30540
rect 62342 30538 62398 30540
rect 62422 30538 62478 30540
rect 62502 30538 62558 30540
rect 62262 30486 62288 30538
rect 62288 30486 62318 30538
rect 62342 30486 62352 30538
rect 62352 30486 62398 30538
rect 62422 30486 62468 30538
rect 62468 30486 62478 30538
rect 62502 30486 62532 30538
rect 62532 30486 62558 30538
rect 62262 30484 62318 30486
rect 62342 30484 62398 30486
rect 62422 30484 62478 30486
rect 62502 30484 62558 30486
rect 62104 30280 62160 30336
rect 62262 29450 62318 29452
rect 62342 29450 62398 29452
rect 62422 29450 62478 29452
rect 62502 29450 62558 29452
rect 62262 29398 62288 29450
rect 62288 29398 62318 29450
rect 62342 29398 62352 29450
rect 62352 29398 62398 29450
rect 62422 29398 62468 29450
rect 62468 29398 62478 29450
rect 62502 29398 62532 29450
rect 62532 29398 62558 29450
rect 62262 29396 62318 29398
rect 62342 29396 62398 29398
rect 62422 29396 62478 29398
rect 62502 29396 62558 29398
rect 59598 27818 59654 27820
rect 59678 27818 59734 27820
rect 59758 27818 59814 27820
rect 59838 27818 59894 27820
rect 59598 27766 59624 27818
rect 59624 27766 59654 27818
rect 59678 27766 59688 27818
rect 59688 27766 59734 27818
rect 59758 27766 59804 27818
rect 59804 27766 59814 27818
rect 59838 27766 59868 27818
rect 59868 27766 59894 27818
rect 59598 27764 59654 27766
rect 59678 27764 59734 27766
rect 59758 27764 59814 27766
rect 59838 27764 59894 27766
rect 62262 28362 62318 28364
rect 62342 28362 62398 28364
rect 62422 28362 62478 28364
rect 62502 28362 62558 28364
rect 62262 28310 62288 28362
rect 62288 28310 62318 28362
rect 62342 28310 62352 28362
rect 62352 28310 62398 28362
rect 62422 28310 62468 28362
rect 62468 28310 62478 28362
rect 62502 28310 62532 28362
rect 62532 28310 62558 28362
rect 62262 28308 62318 28310
rect 62342 28308 62398 28310
rect 62422 28308 62478 28310
rect 62502 28308 62558 28310
rect 64496 29192 64552 29248
rect 64926 32170 64982 32172
rect 65006 32170 65062 32172
rect 65086 32170 65142 32172
rect 65166 32170 65222 32172
rect 64926 32118 64952 32170
rect 64952 32118 64982 32170
rect 65006 32118 65016 32170
rect 65016 32118 65062 32170
rect 65086 32118 65132 32170
rect 65132 32118 65142 32170
rect 65166 32118 65196 32170
rect 65196 32118 65222 32170
rect 64926 32116 64982 32118
rect 65006 32116 65062 32118
rect 65086 32116 65142 32118
rect 65166 32116 65222 32118
rect 65508 31912 65564 31968
rect 65968 33700 66024 33736
rect 65968 33680 65970 33700
rect 65970 33680 66022 33700
rect 66022 33680 66024 33700
rect 67590 35978 67646 35980
rect 67670 35978 67726 35980
rect 67750 35978 67806 35980
rect 67830 35978 67886 35980
rect 67590 35926 67616 35978
rect 67616 35926 67646 35978
rect 67670 35926 67680 35978
rect 67680 35926 67726 35978
rect 67750 35926 67796 35978
rect 67796 35926 67806 35978
rect 67830 35926 67860 35978
rect 67860 35926 67886 35978
rect 67590 35924 67646 35926
rect 67670 35924 67726 35926
rect 67750 35924 67806 35926
rect 67830 35924 67886 35926
rect 66704 32764 66706 32784
rect 66706 32764 66758 32784
rect 66758 32764 66760 32784
rect 66704 32728 66760 32764
rect 64926 31082 64982 31084
rect 65006 31082 65062 31084
rect 65086 31082 65142 31084
rect 65166 31082 65222 31084
rect 64926 31030 64952 31082
rect 64952 31030 64982 31082
rect 65006 31030 65016 31082
rect 65016 31030 65062 31082
rect 65086 31030 65132 31082
rect 65132 31030 65142 31082
rect 65166 31030 65196 31082
rect 65196 31030 65222 31082
rect 64926 31028 64982 31030
rect 65006 31028 65062 31030
rect 65086 31028 65142 31030
rect 65166 31028 65222 31030
rect 65416 30280 65472 30336
rect 64926 29994 64982 29996
rect 65006 29994 65062 29996
rect 65086 29994 65142 29996
rect 65166 29994 65222 29996
rect 64926 29942 64952 29994
rect 64952 29942 64982 29994
rect 65006 29942 65016 29994
rect 65016 29942 65062 29994
rect 65086 29942 65132 29994
rect 65132 29942 65142 29994
rect 65166 29942 65196 29994
rect 65196 29942 65222 29994
rect 64926 29940 64982 29942
rect 65006 29940 65062 29942
rect 65086 29940 65142 29942
rect 65166 29940 65222 29942
rect 64926 28906 64982 28908
rect 65006 28906 65062 28908
rect 65086 28906 65142 28908
rect 65166 28906 65222 28908
rect 64926 28854 64952 28906
rect 64952 28854 64982 28906
rect 65006 28854 65016 28906
rect 65016 28854 65062 28906
rect 65086 28854 65132 28906
rect 65132 28854 65142 28906
rect 65166 28854 65196 28906
rect 65196 28854 65222 28906
rect 64926 28852 64982 28854
rect 65006 28852 65062 28854
rect 65086 28852 65142 28854
rect 65166 28852 65222 28854
rect 68176 37352 68232 37408
rect 70254 41962 70310 41964
rect 70334 41962 70390 41964
rect 70414 41962 70470 41964
rect 70494 41962 70550 41964
rect 70254 41910 70280 41962
rect 70280 41910 70310 41962
rect 70334 41910 70344 41962
rect 70344 41910 70390 41962
rect 70414 41910 70460 41962
rect 70460 41910 70470 41962
rect 70494 41910 70524 41962
rect 70524 41910 70550 41962
rect 70254 41908 70310 41910
rect 70334 41908 70390 41910
rect 70414 41908 70470 41910
rect 70494 41908 70550 41910
rect 70254 40874 70310 40876
rect 70334 40874 70390 40876
rect 70414 40874 70470 40876
rect 70494 40874 70550 40876
rect 70254 40822 70280 40874
rect 70280 40822 70310 40874
rect 70334 40822 70344 40874
rect 70344 40822 70390 40874
rect 70414 40822 70460 40874
rect 70460 40822 70470 40874
rect 70494 40822 70524 40874
rect 70524 40822 70550 40874
rect 70254 40820 70310 40822
rect 70334 40820 70390 40822
rect 70414 40820 70470 40822
rect 70494 40820 70550 40822
rect 70254 39786 70310 39788
rect 70334 39786 70390 39788
rect 70414 39786 70470 39788
rect 70494 39786 70550 39788
rect 70254 39734 70280 39786
rect 70280 39734 70310 39786
rect 70334 39734 70344 39786
rect 70344 39734 70390 39786
rect 70414 39734 70460 39786
rect 70460 39734 70470 39786
rect 70494 39734 70524 39786
rect 70524 39734 70550 39786
rect 70254 39732 70310 39734
rect 70334 39732 70390 39734
rect 70414 39732 70470 39734
rect 70494 39732 70550 39734
rect 72918 41418 72974 41420
rect 72998 41418 73054 41420
rect 73078 41418 73134 41420
rect 73158 41418 73214 41420
rect 72918 41366 72944 41418
rect 72944 41366 72974 41418
rect 72998 41366 73008 41418
rect 73008 41366 73054 41418
rect 73078 41366 73124 41418
rect 73124 41366 73134 41418
rect 73158 41366 73188 41418
rect 73188 41366 73214 41418
rect 72918 41364 72974 41366
rect 72998 41364 73054 41366
rect 73078 41364 73134 41366
rect 73158 41364 73214 41366
rect 72918 40330 72974 40332
rect 72998 40330 73054 40332
rect 73078 40330 73134 40332
rect 73158 40330 73214 40332
rect 72918 40278 72944 40330
rect 72944 40278 72974 40330
rect 72998 40278 73008 40330
rect 73008 40278 73054 40330
rect 73078 40278 73124 40330
rect 73124 40278 73134 40330
rect 73158 40278 73188 40330
rect 73188 40278 73214 40330
rect 72918 40276 72974 40278
rect 72998 40276 73054 40278
rect 73078 40276 73134 40278
rect 73158 40276 73214 40278
rect 70254 38698 70310 38700
rect 70334 38698 70390 38700
rect 70414 38698 70470 38700
rect 70494 38698 70550 38700
rect 70254 38646 70280 38698
rect 70280 38646 70310 38698
rect 70334 38646 70344 38698
rect 70344 38646 70390 38698
rect 70414 38646 70460 38698
rect 70460 38646 70470 38698
rect 70494 38646 70524 38698
rect 70524 38646 70550 38698
rect 70254 38644 70310 38646
rect 70334 38644 70390 38646
rect 70414 38644 70470 38646
rect 70494 38644 70550 38646
rect 70254 37610 70310 37612
rect 70334 37610 70390 37612
rect 70414 37610 70470 37612
rect 70494 37610 70550 37612
rect 70254 37558 70280 37610
rect 70280 37558 70310 37610
rect 70334 37558 70344 37610
rect 70344 37558 70390 37610
rect 70414 37558 70460 37610
rect 70460 37558 70470 37610
rect 70494 37558 70524 37610
rect 70524 37558 70550 37610
rect 70254 37556 70310 37558
rect 70334 37556 70390 37558
rect 70414 37556 70470 37558
rect 70494 37556 70550 37558
rect 69280 37372 69336 37408
rect 69280 37352 69282 37372
rect 69282 37352 69334 37372
rect 69334 37352 69336 37372
rect 69188 37216 69244 37272
rect 68912 36692 68968 36728
rect 68912 36672 68914 36692
rect 68914 36672 68966 36692
rect 68966 36672 68968 36692
rect 67992 35720 68048 35776
rect 67590 34890 67646 34892
rect 67670 34890 67726 34892
rect 67750 34890 67806 34892
rect 67830 34890 67886 34892
rect 67590 34838 67616 34890
rect 67616 34838 67646 34890
rect 67670 34838 67680 34890
rect 67680 34838 67726 34890
rect 67750 34838 67796 34890
rect 67796 34838 67806 34890
rect 67830 34838 67860 34890
rect 67860 34838 67886 34890
rect 67590 34836 67646 34838
rect 67670 34836 67726 34838
rect 67750 34836 67806 34838
rect 67830 34836 67886 34838
rect 67590 33802 67646 33804
rect 67670 33802 67726 33804
rect 67750 33802 67806 33804
rect 67830 33802 67886 33804
rect 67590 33750 67616 33802
rect 67616 33750 67646 33802
rect 67670 33750 67680 33802
rect 67680 33750 67726 33802
rect 67750 33750 67796 33802
rect 67796 33750 67806 33802
rect 67830 33750 67860 33802
rect 67860 33750 67886 33802
rect 67590 33748 67646 33750
rect 67670 33748 67726 33750
rect 67750 33748 67806 33750
rect 67830 33748 67886 33750
rect 67072 32864 67128 32920
rect 67440 32864 67496 32920
rect 67590 32714 67646 32716
rect 67670 32714 67726 32716
rect 67750 32714 67806 32716
rect 67830 32714 67886 32716
rect 67590 32662 67616 32714
rect 67616 32662 67646 32714
rect 67670 32662 67680 32714
rect 67680 32662 67726 32714
rect 67750 32662 67796 32714
rect 67796 32662 67806 32714
rect 67830 32662 67860 32714
rect 67860 32662 67886 32714
rect 67590 32660 67646 32662
rect 67670 32660 67726 32662
rect 67750 32660 67806 32662
rect 67830 32660 67886 32662
rect 66612 30144 66668 30200
rect 64926 27818 64982 27820
rect 65006 27818 65062 27820
rect 65086 27818 65142 27820
rect 65166 27818 65222 27820
rect 64926 27766 64952 27818
rect 64952 27766 64982 27818
rect 65006 27766 65016 27818
rect 65016 27766 65062 27818
rect 65086 27766 65132 27818
rect 65132 27766 65142 27818
rect 65166 27766 65196 27818
rect 65196 27766 65222 27818
rect 64926 27764 64982 27766
rect 65006 27764 65062 27766
rect 65086 27764 65142 27766
rect 65166 27764 65222 27766
rect 62262 27274 62318 27276
rect 62342 27274 62398 27276
rect 62422 27274 62478 27276
rect 62502 27274 62558 27276
rect 62262 27222 62288 27274
rect 62288 27222 62318 27274
rect 62342 27222 62352 27274
rect 62352 27222 62398 27274
rect 62422 27222 62468 27274
rect 62468 27222 62478 27274
rect 62502 27222 62532 27274
rect 62532 27222 62558 27274
rect 62262 27220 62318 27222
rect 62342 27220 62398 27222
rect 62422 27220 62478 27222
rect 62502 27220 62558 27222
rect 67900 32456 67956 32512
rect 67164 32320 67220 32376
rect 67590 31626 67646 31628
rect 67670 31626 67726 31628
rect 67750 31626 67806 31628
rect 67830 31626 67886 31628
rect 67590 31574 67616 31626
rect 67616 31574 67646 31626
rect 67670 31574 67680 31626
rect 67680 31574 67726 31626
rect 67750 31574 67796 31626
rect 67796 31574 67806 31626
rect 67830 31574 67860 31626
rect 67860 31574 67886 31626
rect 67590 31572 67646 31574
rect 67670 31572 67726 31574
rect 67750 31572 67806 31574
rect 67830 31572 67886 31574
rect 67590 30538 67646 30540
rect 67670 30538 67726 30540
rect 67750 30538 67806 30540
rect 67830 30538 67886 30540
rect 67590 30486 67616 30538
rect 67616 30486 67646 30538
rect 67670 30486 67680 30538
rect 67680 30486 67726 30538
rect 67750 30486 67796 30538
rect 67796 30486 67806 30538
rect 67830 30486 67860 30538
rect 67860 30486 67886 30538
rect 67590 30484 67646 30486
rect 67670 30484 67726 30486
rect 67750 30484 67806 30486
rect 67830 30484 67886 30486
rect 67590 29450 67646 29452
rect 67670 29450 67726 29452
rect 67750 29450 67806 29452
rect 67830 29450 67886 29452
rect 67590 29398 67616 29450
rect 67616 29398 67646 29450
rect 67670 29398 67680 29450
rect 67680 29398 67726 29450
rect 67750 29398 67796 29450
rect 67796 29398 67806 29450
rect 67830 29398 67860 29450
rect 67860 29398 67886 29450
rect 67590 29396 67646 29398
rect 67670 29396 67726 29398
rect 67750 29396 67806 29398
rect 67830 29396 67886 29398
rect 69740 33000 69796 33056
rect 68360 32320 68416 32376
rect 67590 28362 67646 28364
rect 67670 28362 67726 28364
rect 67750 28362 67806 28364
rect 67830 28362 67886 28364
rect 67590 28310 67616 28362
rect 67616 28310 67646 28362
rect 67670 28310 67680 28362
rect 67680 28310 67726 28362
rect 67750 28310 67796 28362
rect 67796 28310 67806 28362
rect 67830 28310 67860 28362
rect 67860 28310 67886 28362
rect 67590 28308 67646 28310
rect 67670 28308 67726 28310
rect 67750 28308 67806 28310
rect 67830 28308 67886 28310
rect 68176 28104 68232 28160
rect 67590 27274 67646 27276
rect 67670 27274 67726 27276
rect 67750 27274 67806 27276
rect 67830 27274 67886 27276
rect 67590 27222 67616 27274
rect 67616 27222 67646 27274
rect 67670 27222 67680 27274
rect 67680 27222 67726 27274
rect 67750 27222 67796 27274
rect 67796 27222 67806 27274
rect 67830 27222 67860 27274
rect 67860 27222 67886 27274
rect 67590 27220 67646 27222
rect 67670 27220 67726 27222
rect 67750 27220 67806 27222
rect 67830 27220 67886 27222
rect 48942 26730 48998 26732
rect 49022 26730 49078 26732
rect 49102 26730 49158 26732
rect 49182 26730 49238 26732
rect 48942 26678 48968 26730
rect 48968 26678 48998 26730
rect 49022 26678 49032 26730
rect 49032 26678 49078 26730
rect 49102 26678 49148 26730
rect 49148 26678 49158 26730
rect 49182 26678 49212 26730
rect 49212 26678 49238 26730
rect 48942 26676 48998 26678
rect 49022 26676 49078 26678
rect 49102 26676 49158 26678
rect 49182 26676 49238 26678
rect 54270 26730 54326 26732
rect 54350 26730 54406 26732
rect 54430 26730 54486 26732
rect 54510 26730 54566 26732
rect 54270 26678 54296 26730
rect 54296 26678 54326 26730
rect 54350 26678 54360 26730
rect 54360 26678 54406 26730
rect 54430 26678 54476 26730
rect 54476 26678 54486 26730
rect 54510 26678 54540 26730
rect 54540 26678 54566 26730
rect 54270 26676 54326 26678
rect 54350 26676 54406 26678
rect 54430 26676 54486 26678
rect 54510 26676 54566 26678
rect 59598 26730 59654 26732
rect 59678 26730 59734 26732
rect 59758 26730 59814 26732
rect 59838 26730 59894 26732
rect 59598 26678 59624 26730
rect 59624 26678 59654 26730
rect 59678 26678 59688 26730
rect 59688 26678 59734 26730
rect 59758 26678 59804 26730
rect 59804 26678 59814 26730
rect 59838 26678 59868 26730
rect 59868 26678 59894 26730
rect 59598 26676 59654 26678
rect 59678 26676 59734 26678
rect 59758 26676 59814 26678
rect 59838 26676 59894 26678
rect 64926 26730 64982 26732
rect 65006 26730 65062 26732
rect 65086 26730 65142 26732
rect 65166 26730 65222 26732
rect 64926 26678 64952 26730
rect 64952 26678 64982 26730
rect 65006 26678 65016 26730
rect 65016 26678 65062 26730
rect 65086 26678 65132 26730
rect 65132 26678 65142 26730
rect 65166 26678 65196 26730
rect 65196 26678 65222 26730
rect 64926 26676 64982 26678
rect 65006 26676 65062 26678
rect 65086 26676 65142 26678
rect 65166 26676 65222 26678
rect 46096 23548 46152 23604
rect 43520 22936 43576 22992
rect 67164 21304 67220 21360
rect 67072 20624 67128 20680
rect 40950 18570 41006 18572
rect 41030 18570 41086 18572
rect 41110 18570 41166 18572
rect 41190 18570 41246 18572
rect 40950 18518 40976 18570
rect 40976 18518 41006 18570
rect 41030 18518 41040 18570
rect 41040 18518 41086 18570
rect 41110 18518 41156 18570
rect 41156 18518 41166 18570
rect 41190 18518 41220 18570
rect 41220 18518 41246 18570
rect 40950 18516 41006 18518
rect 41030 18516 41086 18518
rect 41110 18516 41166 18518
rect 41190 18516 41246 18518
rect 42048 17924 42104 17960
rect 42048 17904 42050 17924
rect 42050 17904 42102 17924
rect 42102 17904 42104 17924
rect 40950 17482 41006 17484
rect 41030 17482 41086 17484
rect 41110 17482 41166 17484
rect 41190 17482 41246 17484
rect 40950 17430 40976 17482
rect 40976 17430 41006 17482
rect 41030 17430 41040 17482
rect 41040 17430 41086 17482
rect 41110 17430 41156 17482
rect 41156 17430 41166 17482
rect 41190 17430 41220 17482
rect 41220 17430 41246 17482
rect 40950 17428 41006 17430
rect 41030 17428 41086 17430
rect 41110 17428 41166 17430
rect 41190 17428 41246 17430
rect 38286 16938 38342 16940
rect 38366 16938 38422 16940
rect 38446 16938 38502 16940
rect 38526 16938 38582 16940
rect 38286 16886 38312 16938
rect 38312 16886 38342 16938
rect 38366 16886 38376 16938
rect 38376 16886 38422 16938
rect 38446 16886 38492 16938
rect 38492 16886 38502 16938
rect 38526 16886 38556 16938
rect 38556 16886 38582 16938
rect 38286 16884 38342 16886
rect 38366 16884 38422 16886
rect 38446 16884 38502 16886
rect 38526 16884 38582 16886
rect 38828 17108 38884 17144
rect 38828 17088 38830 17108
rect 38830 17088 38882 17108
rect 38882 17088 38884 17108
rect 40760 17124 40762 17144
rect 40762 17124 40814 17144
rect 40814 17124 40816 17144
rect 40760 17088 40816 17124
rect 35622 15306 35678 15308
rect 35702 15306 35758 15308
rect 35782 15306 35838 15308
rect 35862 15306 35918 15308
rect 35622 15254 35648 15306
rect 35648 15254 35678 15306
rect 35702 15254 35712 15306
rect 35712 15254 35758 15306
rect 35782 15254 35828 15306
rect 35828 15254 35838 15306
rect 35862 15254 35892 15306
rect 35892 15254 35918 15306
rect 35622 15252 35678 15254
rect 35702 15252 35758 15254
rect 35782 15252 35838 15254
rect 35862 15252 35918 15254
rect 38286 15850 38342 15852
rect 38366 15850 38422 15852
rect 38446 15850 38502 15852
rect 38526 15850 38582 15852
rect 38286 15798 38312 15850
rect 38312 15798 38342 15850
rect 38366 15798 38376 15850
rect 38376 15798 38422 15850
rect 38446 15798 38492 15850
rect 38492 15798 38502 15850
rect 38526 15798 38556 15850
rect 38556 15798 38582 15850
rect 38286 15796 38342 15798
rect 38366 15796 38422 15798
rect 38446 15796 38502 15798
rect 38526 15796 38582 15798
rect 41680 16580 41682 16600
rect 41682 16580 41734 16600
rect 41734 16580 41736 16600
rect 41680 16544 41736 16580
rect 40950 16394 41006 16396
rect 41030 16394 41086 16396
rect 41110 16394 41166 16396
rect 41190 16394 41246 16396
rect 40950 16342 40976 16394
rect 40976 16342 41006 16394
rect 41030 16342 41040 16394
rect 41040 16342 41086 16394
rect 41110 16342 41156 16394
rect 41156 16342 41166 16394
rect 41190 16342 41220 16394
rect 41220 16342 41246 16394
rect 40950 16340 41006 16342
rect 41030 16340 41086 16342
rect 41110 16340 41166 16342
rect 41190 16340 41246 16342
rect 40950 15306 41006 15308
rect 41030 15306 41086 15308
rect 41110 15306 41166 15308
rect 41190 15306 41246 15308
rect 40950 15254 40976 15306
rect 40976 15254 41006 15306
rect 41030 15254 41040 15306
rect 41040 15254 41086 15306
rect 41110 15254 41156 15306
rect 41156 15254 41166 15306
rect 41190 15254 41220 15306
rect 41220 15254 41246 15306
rect 40950 15252 41006 15254
rect 41030 15252 41086 15254
rect 41110 15252 41166 15254
rect 41190 15252 41246 15254
rect 34412 14812 34414 14832
rect 34414 14812 34466 14832
rect 34466 14812 34468 14832
rect 34412 14776 34468 14812
rect 38286 14762 38342 14764
rect 38366 14762 38422 14764
rect 38446 14762 38502 14764
rect 38526 14762 38582 14764
rect 38286 14710 38312 14762
rect 38312 14710 38342 14762
rect 38366 14710 38376 14762
rect 38376 14710 38422 14762
rect 38446 14710 38492 14762
rect 38492 14710 38502 14762
rect 38526 14710 38556 14762
rect 38556 14710 38582 14762
rect 38286 14708 38342 14710
rect 38366 14708 38422 14710
rect 38446 14708 38502 14710
rect 38526 14708 38582 14710
rect 35622 14218 35678 14220
rect 35702 14218 35758 14220
rect 35782 14218 35838 14220
rect 35862 14218 35918 14220
rect 35622 14166 35648 14218
rect 35648 14166 35678 14218
rect 35702 14166 35712 14218
rect 35712 14166 35758 14218
rect 35782 14166 35828 14218
rect 35828 14166 35838 14218
rect 35862 14166 35892 14218
rect 35892 14166 35918 14218
rect 35622 14164 35678 14166
rect 35702 14164 35758 14166
rect 35782 14164 35838 14166
rect 35862 14164 35918 14166
rect 38286 13674 38342 13676
rect 38366 13674 38422 13676
rect 38446 13674 38502 13676
rect 38526 13674 38582 13676
rect 38286 13622 38312 13674
rect 38312 13622 38342 13674
rect 38366 13622 38376 13674
rect 38376 13622 38422 13674
rect 38446 13622 38492 13674
rect 38492 13622 38502 13674
rect 38526 13622 38556 13674
rect 38556 13622 38582 13674
rect 38286 13620 38342 13622
rect 38366 13620 38422 13622
rect 38446 13620 38502 13622
rect 38526 13620 38582 13622
rect 35622 13130 35678 13132
rect 35702 13130 35758 13132
rect 35782 13130 35838 13132
rect 35862 13130 35918 13132
rect 35622 13078 35648 13130
rect 35648 13078 35678 13130
rect 35702 13078 35712 13130
rect 35712 13078 35758 13130
rect 35782 13078 35828 13130
rect 35828 13078 35838 13130
rect 35862 13078 35892 13130
rect 35892 13078 35918 13130
rect 35622 13076 35678 13078
rect 35702 13076 35758 13078
rect 35782 13076 35838 13078
rect 35862 13076 35918 13078
rect 38286 12586 38342 12588
rect 38366 12586 38422 12588
rect 38446 12586 38502 12588
rect 38526 12586 38582 12588
rect 38286 12534 38312 12586
rect 38312 12534 38342 12586
rect 38366 12534 38376 12586
rect 38376 12534 38422 12586
rect 38446 12534 38492 12586
rect 38492 12534 38502 12586
rect 38526 12534 38556 12586
rect 38556 12534 38582 12586
rect 38286 12532 38342 12534
rect 38366 12532 38422 12534
rect 38446 12532 38502 12534
rect 38526 12532 38582 12534
rect 35622 12042 35678 12044
rect 35702 12042 35758 12044
rect 35782 12042 35838 12044
rect 35862 12042 35918 12044
rect 35622 11990 35648 12042
rect 35648 11990 35678 12042
rect 35702 11990 35712 12042
rect 35712 11990 35758 12042
rect 35782 11990 35828 12042
rect 35828 11990 35838 12042
rect 35862 11990 35892 12042
rect 35892 11990 35918 12042
rect 35622 11988 35678 11990
rect 35702 11988 35758 11990
rect 35782 11988 35838 11990
rect 35862 11988 35918 11990
rect 40950 14218 41006 14220
rect 41030 14218 41086 14220
rect 41110 14218 41166 14220
rect 41190 14218 41246 14220
rect 40950 14166 40976 14218
rect 40976 14166 41006 14218
rect 41030 14166 41040 14218
rect 41040 14166 41086 14218
rect 41110 14166 41156 14218
rect 41156 14166 41166 14218
rect 41190 14166 41220 14218
rect 41220 14166 41246 14218
rect 40950 14164 41006 14166
rect 41030 14164 41086 14166
rect 41110 14164 41166 14166
rect 41190 14164 41246 14166
rect 40950 13130 41006 13132
rect 41030 13130 41086 13132
rect 41110 13130 41166 13132
rect 41190 13130 41246 13132
rect 40950 13078 40976 13130
rect 40976 13078 41006 13130
rect 41030 13078 41040 13130
rect 41040 13078 41086 13130
rect 41110 13078 41156 13130
rect 41156 13078 41166 13130
rect 41190 13078 41220 13130
rect 41220 13078 41246 13130
rect 40950 13076 41006 13078
rect 41030 13076 41086 13078
rect 41110 13076 41166 13078
rect 41190 13076 41246 13078
rect 40950 12042 41006 12044
rect 41030 12042 41086 12044
rect 41110 12042 41166 12044
rect 41190 12042 41246 12044
rect 40950 11990 40976 12042
rect 40976 11990 41006 12042
rect 41030 11990 41040 12042
rect 41040 11990 41086 12042
rect 41110 11990 41156 12042
rect 41156 11990 41166 12042
rect 41190 11990 41220 12042
rect 41220 11990 41246 12042
rect 40950 11988 41006 11990
rect 41030 11988 41086 11990
rect 41110 11988 41166 11990
rect 41190 11988 41246 11990
rect 38286 11498 38342 11500
rect 38366 11498 38422 11500
rect 38446 11498 38502 11500
rect 38526 11498 38582 11500
rect 38286 11446 38312 11498
rect 38312 11446 38342 11498
rect 38366 11446 38376 11498
rect 38376 11446 38422 11498
rect 38446 11446 38492 11498
rect 38492 11446 38502 11498
rect 38526 11446 38556 11498
rect 38556 11446 38582 11498
rect 38286 11444 38342 11446
rect 38366 11444 38422 11446
rect 38446 11444 38502 11446
rect 38526 11444 38582 11446
rect 35622 10954 35678 10956
rect 35702 10954 35758 10956
rect 35782 10954 35838 10956
rect 35862 10954 35918 10956
rect 35622 10902 35648 10954
rect 35648 10902 35678 10954
rect 35702 10902 35712 10954
rect 35712 10902 35758 10954
rect 35782 10902 35828 10954
rect 35828 10902 35838 10954
rect 35862 10902 35892 10954
rect 35892 10902 35918 10954
rect 35622 10900 35678 10902
rect 35702 10900 35758 10902
rect 35782 10900 35838 10902
rect 35862 10900 35918 10902
rect 40950 10954 41006 10956
rect 41030 10954 41086 10956
rect 41110 10954 41166 10956
rect 41190 10954 41246 10956
rect 40950 10902 40976 10954
rect 40976 10902 41006 10954
rect 41030 10902 41040 10954
rect 41040 10902 41086 10954
rect 41110 10902 41156 10954
rect 41156 10902 41166 10954
rect 41190 10902 41220 10954
rect 41220 10902 41246 10954
rect 40950 10900 41006 10902
rect 41030 10900 41086 10902
rect 41110 10900 41166 10902
rect 41190 10900 41246 10902
rect 34412 10460 34414 10480
rect 34414 10460 34466 10480
rect 34466 10460 34468 10480
rect 34412 10424 34468 10460
rect 38286 10410 38342 10412
rect 38366 10410 38422 10412
rect 38446 10410 38502 10412
rect 38526 10410 38582 10412
rect 38286 10358 38312 10410
rect 38312 10358 38342 10410
rect 38366 10358 38376 10410
rect 38376 10358 38422 10410
rect 38446 10358 38492 10410
rect 38492 10358 38502 10410
rect 38526 10358 38556 10410
rect 38556 10358 38582 10410
rect 38286 10356 38342 10358
rect 38366 10356 38422 10358
rect 38446 10356 38502 10358
rect 38526 10356 38582 10358
rect 3654 9866 3710 9868
rect 3734 9866 3790 9868
rect 3814 9866 3870 9868
rect 3894 9866 3950 9868
rect 3654 9814 3680 9866
rect 3680 9814 3710 9866
rect 3734 9814 3744 9866
rect 3744 9814 3790 9866
rect 3814 9814 3860 9866
rect 3860 9814 3870 9866
rect 3894 9814 3924 9866
rect 3924 9814 3950 9866
rect 3654 9812 3710 9814
rect 3734 9812 3790 9814
rect 3814 9812 3870 9814
rect 3894 9812 3950 9814
rect 6318 9322 6374 9324
rect 6398 9322 6454 9324
rect 6478 9322 6534 9324
rect 6558 9322 6614 9324
rect 6318 9270 6344 9322
rect 6344 9270 6374 9322
rect 6398 9270 6408 9322
rect 6408 9270 6454 9322
rect 6478 9270 6524 9322
rect 6524 9270 6534 9322
rect 6558 9270 6588 9322
rect 6588 9270 6614 9322
rect 6318 9268 6374 9270
rect 6398 9268 6454 9270
rect 6478 9268 6534 9270
rect 6558 9268 6614 9270
rect 3654 8778 3710 8780
rect 3734 8778 3790 8780
rect 3814 8778 3870 8780
rect 3894 8778 3950 8780
rect 3654 8726 3680 8778
rect 3680 8726 3710 8778
rect 3734 8726 3744 8778
rect 3744 8726 3790 8778
rect 3814 8726 3860 8778
rect 3860 8726 3870 8778
rect 3894 8726 3924 8778
rect 3924 8726 3950 8778
rect 3654 8724 3710 8726
rect 3734 8724 3790 8726
rect 3814 8724 3870 8726
rect 3894 8724 3950 8726
rect 6318 8234 6374 8236
rect 6398 8234 6454 8236
rect 6478 8234 6534 8236
rect 6558 8234 6614 8236
rect 6318 8182 6344 8234
rect 6344 8182 6374 8234
rect 6398 8182 6408 8234
rect 6408 8182 6454 8234
rect 6478 8182 6524 8234
rect 6524 8182 6534 8234
rect 6558 8182 6588 8234
rect 6588 8182 6614 8234
rect 6318 8180 6374 8182
rect 6398 8180 6454 8182
rect 6478 8180 6534 8182
rect 6558 8180 6614 8182
rect 3654 7690 3710 7692
rect 3734 7690 3790 7692
rect 3814 7690 3870 7692
rect 3894 7690 3950 7692
rect 3654 7638 3680 7690
rect 3680 7638 3710 7690
rect 3734 7638 3744 7690
rect 3744 7638 3790 7690
rect 3814 7638 3860 7690
rect 3860 7638 3870 7690
rect 3894 7638 3924 7690
rect 3924 7638 3950 7690
rect 3654 7636 3710 7638
rect 3734 7636 3790 7638
rect 3814 7636 3870 7638
rect 3894 7636 3950 7638
rect 6318 7146 6374 7148
rect 6398 7146 6454 7148
rect 6478 7146 6534 7148
rect 6558 7146 6614 7148
rect 6318 7094 6344 7146
rect 6344 7094 6374 7146
rect 6398 7094 6408 7146
rect 6408 7094 6454 7146
rect 6478 7094 6524 7146
rect 6524 7094 6534 7146
rect 6558 7094 6588 7146
rect 6588 7094 6614 7146
rect 6318 7092 6374 7094
rect 6398 7092 6454 7094
rect 6478 7092 6534 7094
rect 6558 7092 6614 7094
rect 3654 6602 3710 6604
rect 3734 6602 3790 6604
rect 3814 6602 3870 6604
rect 3894 6602 3950 6604
rect 3654 6550 3680 6602
rect 3680 6550 3710 6602
rect 3734 6550 3744 6602
rect 3744 6550 3790 6602
rect 3814 6550 3860 6602
rect 3860 6550 3870 6602
rect 3894 6550 3924 6602
rect 3924 6550 3950 6602
rect 3654 6548 3710 6550
rect 3734 6548 3790 6550
rect 3814 6548 3870 6550
rect 3894 6548 3950 6550
rect 6318 6058 6374 6060
rect 6398 6058 6454 6060
rect 6478 6058 6534 6060
rect 6558 6058 6614 6060
rect 6318 6006 6344 6058
rect 6344 6006 6374 6058
rect 6398 6006 6408 6058
rect 6408 6006 6454 6058
rect 6478 6006 6524 6058
rect 6524 6006 6534 6058
rect 6558 6006 6588 6058
rect 6588 6006 6614 6058
rect 6318 6004 6374 6006
rect 6398 6004 6454 6006
rect 6478 6004 6534 6006
rect 6558 6004 6614 6006
rect 3654 5514 3710 5516
rect 3734 5514 3790 5516
rect 3814 5514 3870 5516
rect 3894 5514 3950 5516
rect 3654 5462 3680 5514
rect 3680 5462 3710 5514
rect 3734 5462 3744 5514
rect 3744 5462 3790 5514
rect 3814 5462 3860 5514
rect 3860 5462 3870 5514
rect 3894 5462 3924 5514
rect 3924 5462 3950 5514
rect 3654 5460 3710 5462
rect 3734 5460 3790 5462
rect 3814 5460 3870 5462
rect 3894 5460 3950 5462
rect 6318 4970 6374 4972
rect 6398 4970 6454 4972
rect 6478 4970 6534 4972
rect 6558 4970 6614 4972
rect 6318 4918 6344 4970
rect 6344 4918 6374 4970
rect 6398 4918 6408 4970
rect 6408 4918 6454 4970
rect 6478 4918 6524 4970
rect 6524 4918 6534 4970
rect 6558 4918 6588 4970
rect 6588 4918 6614 4970
rect 6318 4916 6374 4918
rect 6398 4916 6454 4918
rect 6478 4916 6534 4918
rect 6558 4916 6614 4918
rect 3654 4426 3710 4428
rect 3734 4426 3790 4428
rect 3814 4426 3870 4428
rect 3894 4426 3950 4428
rect 3654 4374 3680 4426
rect 3680 4374 3710 4426
rect 3734 4374 3744 4426
rect 3744 4374 3790 4426
rect 3814 4374 3860 4426
rect 3860 4374 3870 4426
rect 3894 4374 3924 4426
rect 3924 4374 3950 4426
rect 3654 4372 3710 4374
rect 3734 4372 3790 4374
rect 3814 4372 3870 4374
rect 3894 4372 3950 4374
rect 6318 3882 6374 3884
rect 6398 3882 6454 3884
rect 6478 3882 6534 3884
rect 6558 3882 6614 3884
rect 6318 3830 6344 3882
rect 6344 3830 6374 3882
rect 6398 3830 6408 3882
rect 6408 3830 6454 3882
rect 6478 3830 6524 3882
rect 6524 3830 6534 3882
rect 6558 3830 6588 3882
rect 6588 3830 6614 3882
rect 6318 3828 6374 3830
rect 6398 3828 6454 3830
rect 6478 3828 6534 3830
rect 6558 3828 6614 3830
rect 3654 3338 3710 3340
rect 3734 3338 3790 3340
rect 3814 3338 3870 3340
rect 3894 3338 3950 3340
rect 3654 3286 3680 3338
rect 3680 3286 3710 3338
rect 3734 3286 3744 3338
rect 3744 3286 3790 3338
rect 3814 3286 3860 3338
rect 3860 3286 3870 3338
rect 3894 3286 3924 3338
rect 3924 3286 3950 3338
rect 3654 3284 3710 3286
rect 3734 3284 3790 3286
rect 3814 3284 3870 3286
rect 3894 3284 3950 3286
rect 6318 2794 6374 2796
rect 6398 2794 6454 2796
rect 6478 2794 6534 2796
rect 6558 2794 6614 2796
rect 6318 2742 6344 2794
rect 6344 2742 6374 2794
rect 6398 2742 6408 2794
rect 6408 2742 6454 2794
rect 6478 2742 6524 2794
rect 6524 2742 6534 2794
rect 6558 2742 6588 2794
rect 6588 2742 6614 2794
rect 6318 2740 6374 2742
rect 6398 2740 6454 2742
rect 6478 2740 6534 2742
rect 6558 2740 6614 2742
rect 3654 2250 3710 2252
rect 3734 2250 3790 2252
rect 3814 2250 3870 2252
rect 3894 2250 3950 2252
rect 3654 2198 3680 2250
rect 3680 2198 3710 2250
rect 3734 2198 3744 2250
rect 3744 2198 3790 2250
rect 3814 2198 3860 2250
rect 3860 2198 3870 2250
rect 3894 2198 3924 2250
rect 3924 2198 3950 2250
rect 3654 2196 3710 2198
rect 3734 2196 3790 2198
rect 3814 2196 3870 2198
rect 3894 2196 3950 2198
rect 35622 9866 35678 9868
rect 35702 9866 35758 9868
rect 35782 9866 35838 9868
rect 35862 9866 35918 9868
rect 35622 9814 35648 9866
rect 35648 9814 35678 9866
rect 35702 9814 35712 9866
rect 35712 9814 35758 9866
rect 35782 9814 35828 9866
rect 35828 9814 35838 9866
rect 35862 9814 35892 9866
rect 35892 9814 35918 9866
rect 35622 9812 35678 9814
rect 35702 9812 35758 9814
rect 35782 9812 35838 9814
rect 35862 9812 35918 9814
rect 40950 9866 41006 9868
rect 41030 9866 41086 9868
rect 41110 9866 41166 9868
rect 41190 9866 41246 9868
rect 40950 9814 40976 9866
rect 40976 9814 41006 9866
rect 41030 9814 41040 9866
rect 41040 9814 41086 9866
rect 41110 9814 41156 9866
rect 41156 9814 41166 9866
rect 41190 9814 41220 9866
rect 41220 9814 41246 9866
rect 40950 9812 41006 9814
rect 41030 9812 41086 9814
rect 41110 9812 41166 9814
rect 41190 9812 41246 9814
rect 38286 9322 38342 9324
rect 38366 9322 38422 9324
rect 38446 9322 38502 9324
rect 38526 9322 38582 9324
rect 38286 9270 38312 9322
rect 38312 9270 38342 9322
rect 38366 9270 38376 9322
rect 38376 9270 38422 9322
rect 38446 9270 38492 9322
rect 38492 9270 38502 9322
rect 38526 9270 38556 9322
rect 38556 9270 38582 9322
rect 38286 9268 38342 9270
rect 38366 9268 38422 9270
rect 38446 9268 38502 9270
rect 38526 9268 38582 9270
rect 35622 8778 35678 8780
rect 35702 8778 35758 8780
rect 35782 8778 35838 8780
rect 35862 8778 35918 8780
rect 35622 8726 35648 8778
rect 35648 8726 35678 8778
rect 35702 8726 35712 8778
rect 35712 8726 35758 8778
rect 35782 8726 35828 8778
rect 35828 8726 35838 8778
rect 35862 8726 35892 8778
rect 35892 8726 35918 8778
rect 35622 8724 35678 8726
rect 35702 8724 35758 8726
rect 35782 8724 35838 8726
rect 35862 8724 35918 8726
rect 40950 8778 41006 8780
rect 41030 8778 41086 8780
rect 41110 8778 41166 8780
rect 41190 8778 41246 8780
rect 40950 8726 40976 8778
rect 40976 8726 41006 8778
rect 41030 8726 41040 8778
rect 41040 8726 41086 8778
rect 41110 8726 41156 8778
rect 41156 8726 41166 8778
rect 41190 8726 41220 8778
rect 41220 8726 41246 8778
rect 40950 8724 41006 8726
rect 41030 8724 41086 8726
rect 41110 8724 41166 8726
rect 41190 8724 41246 8726
rect 38286 8234 38342 8236
rect 38366 8234 38422 8236
rect 38446 8234 38502 8236
rect 38526 8234 38582 8236
rect 38286 8182 38312 8234
rect 38312 8182 38342 8234
rect 38366 8182 38376 8234
rect 38376 8182 38422 8234
rect 38446 8182 38492 8234
rect 38492 8182 38502 8234
rect 38526 8182 38556 8234
rect 38556 8182 38582 8234
rect 38286 8180 38342 8182
rect 38366 8180 38422 8182
rect 38446 8180 38502 8182
rect 38526 8180 38582 8182
rect 35622 7690 35678 7692
rect 35702 7690 35758 7692
rect 35782 7690 35838 7692
rect 35862 7690 35918 7692
rect 35622 7638 35648 7690
rect 35648 7638 35678 7690
rect 35702 7638 35712 7690
rect 35712 7638 35758 7690
rect 35782 7638 35828 7690
rect 35828 7638 35838 7690
rect 35862 7638 35892 7690
rect 35892 7638 35918 7690
rect 35622 7636 35678 7638
rect 35702 7636 35758 7638
rect 35782 7636 35838 7638
rect 35862 7636 35918 7638
rect 40950 7690 41006 7692
rect 41030 7690 41086 7692
rect 41110 7690 41166 7692
rect 41190 7690 41246 7692
rect 40950 7638 40976 7690
rect 40976 7638 41006 7690
rect 41030 7638 41040 7690
rect 41040 7638 41086 7690
rect 41110 7638 41156 7690
rect 41156 7638 41166 7690
rect 41190 7638 41220 7690
rect 41220 7638 41246 7690
rect 40950 7636 41006 7638
rect 41030 7636 41086 7638
rect 41110 7636 41166 7638
rect 41190 7636 41246 7638
rect 38286 7146 38342 7148
rect 38366 7146 38422 7148
rect 38446 7146 38502 7148
rect 38526 7146 38582 7148
rect 38286 7094 38312 7146
rect 38312 7094 38342 7146
rect 38366 7094 38376 7146
rect 38376 7094 38422 7146
rect 38446 7094 38492 7146
rect 38492 7094 38502 7146
rect 38526 7094 38556 7146
rect 38556 7094 38582 7146
rect 38286 7092 38342 7094
rect 38366 7092 38422 7094
rect 38446 7092 38502 7094
rect 38526 7092 38582 7094
rect 35622 6602 35678 6604
rect 35702 6602 35758 6604
rect 35782 6602 35838 6604
rect 35862 6602 35918 6604
rect 35622 6550 35648 6602
rect 35648 6550 35678 6602
rect 35702 6550 35712 6602
rect 35712 6550 35758 6602
rect 35782 6550 35828 6602
rect 35828 6550 35838 6602
rect 35862 6550 35892 6602
rect 35892 6550 35918 6602
rect 35622 6548 35678 6550
rect 35702 6548 35758 6550
rect 35782 6548 35838 6550
rect 35862 6548 35918 6550
rect 40950 6602 41006 6604
rect 41030 6602 41086 6604
rect 41110 6602 41166 6604
rect 41190 6602 41246 6604
rect 40950 6550 40976 6602
rect 40976 6550 41006 6602
rect 41030 6550 41040 6602
rect 41040 6550 41086 6602
rect 41110 6550 41156 6602
rect 41156 6550 41166 6602
rect 41190 6550 41220 6602
rect 41220 6550 41246 6602
rect 40950 6548 41006 6550
rect 41030 6548 41086 6550
rect 41110 6548 41166 6550
rect 41190 6548 41246 6550
rect 38286 6058 38342 6060
rect 38366 6058 38422 6060
rect 38446 6058 38502 6060
rect 38526 6058 38582 6060
rect 38286 6006 38312 6058
rect 38312 6006 38342 6058
rect 38366 6006 38376 6058
rect 38376 6006 38422 6058
rect 38446 6006 38492 6058
rect 38492 6006 38502 6058
rect 38526 6006 38556 6058
rect 38556 6006 38582 6058
rect 38286 6004 38342 6006
rect 38366 6004 38422 6006
rect 38446 6004 38502 6006
rect 38526 6004 38582 6006
rect 35622 5514 35678 5516
rect 35702 5514 35758 5516
rect 35782 5514 35838 5516
rect 35862 5514 35918 5516
rect 35622 5462 35648 5514
rect 35648 5462 35678 5514
rect 35702 5462 35712 5514
rect 35712 5462 35758 5514
rect 35782 5462 35828 5514
rect 35828 5462 35838 5514
rect 35862 5462 35892 5514
rect 35892 5462 35918 5514
rect 35622 5460 35678 5462
rect 35702 5460 35758 5462
rect 35782 5460 35838 5462
rect 35862 5460 35918 5462
rect 40950 5514 41006 5516
rect 41030 5514 41086 5516
rect 41110 5514 41166 5516
rect 41190 5514 41246 5516
rect 40950 5462 40976 5514
rect 40976 5462 41006 5514
rect 41030 5462 41040 5514
rect 41040 5462 41086 5514
rect 41110 5462 41156 5514
rect 41156 5462 41166 5514
rect 41190 5462 41220 5514
rect 41220 5462 41246 5514
rect 40950 5460 41006 5462
rect 41030 5460 41086 5462
rect 41110 5460 41166 5462
rect 41190 5460 41246 5462
rect 38286 4970 38342 4972
rect 38366 4970 38422 4972
rect 38446 4970 38502 4972
rect 38526 4970 38582 4972
rect 38286 4918 38312 4970
rect 38312 4918 38342 4970
rect 38366 4918 38376 4970
rect 38376 4918 38422 4970
rect 38446 4918 38492 4970
rect 38492 4918 38502 4970
rect 38526 4918 38556 4970
rect 38556 4918 38582 4970
rect 38286 4916 38342 4918
rect 38366 4916 38422 4918
rect 38446 4916 38502 4918
rect 38526 4916 38582 4918
rect 35622 4426 35678 4428
rect 35702 4426 35758 4428
rect 35782 4426 35838 4428
rect 35862 4426 35918 4428
rect 35622 4374 35648 4426
rect 35648 4374 35678 4426
rect 35702 4374 35712 4426
rect 35712 4374 35758 4426
rect 35782 4374 35828 4426
rect 35828 4374 35838 4426
rect 35862 4374 35892 4426
rect 35892 4374 35918 4426
rect 35622 4372 35678 4374
rect 35702 4372 35758 4374
rect 35782 4372 35838 4374
rect 35862 4372 35918 4374
rect 40950 4426 41006 4428
rect 41030 4426 41086 4428
rect 41110 4426 41166 4428
rect 41190 4426 41246 4428
rect 40950 4374 40976 4426
rect 40976 4374 41006 4426
rect 41030 4374 41040 4426
rect 41040 4374 41086 4426
rect 41110 4374 41156 4426
rect 41156 4374 41166 4426
rect 41190 4374 41220 4426
rect 41220 4374 41246 4426
rect 40950 4372 41006 4374
rect 41030 4372 41086 4374
rect 41110 4372 41166 4374
rect 41190 4372 41246 4374
rect 38286 3882 38342 3884
rect 38366 3882 38422 3884
rect 38446 3882 38502 3884
rect 38526 3882 38582 3884
rect 38286 3830 38312 3882
rect 38312 3830 38342 3882
rect 38366 3830 38376 3882
rect 38376 3830 38422 3882
rect 38446 3830 38492 3882
rect 38492 3830 38502 3882
rect 38526 3830 38556 3882
rect 38556 3830 38582 3882
rect 38286 3828 38342 3830
rect 38366 3828 38422 3830
rect 38446 3828 38502 3830
rect 38526 3828 38582 3830
rect 35622 3338 35678 3340
rect 35702 3338 35758 3340
rect 35782 3338 35838 3340
rect 35862 3338 35918 3340
rect 35622 3286 35648 3338
rect 35648 3286 35678 3338
rect 35702 3286 35712 3338
rect 35712 3286 35758 3338
rect 35782 3286 35828 3338
rect 35828 3286 35838 3338
rect 35862 3286 35892 3338
rect 35892 3286 35918 3338
rect 35622 3284 35678 3286
rect 35702 3284 35758 3286
rect 35782 3284 35838 3286
rect 35862 3284 35918 3286
rect 40950 3338 41006 3340
rect 41030 3338 41086 3340
rect 41110 3338 41166 3340
rect 41190 3338 41246 3340
rect 40950 3286 40976 3338
rect 40976 3286 41006 3338
rect 41030 3286 41040 3338
rect 41040 3286 41086 3338
rect 41110 3286 41156 3338
rect 41156 3286 41166 3338
rect 41190 3286 41220 3338
rect 41220 3286 41246 3338
rect 40950 3284 41006 3286
rect 41030 3284 41086 3286
rect 41110 3284 41166 3286
rect 41190 3284 41246 3286
rect 38286 2794 38342 2796
rect 38366 2794 38422 2796
rect 38446 2794 38502 2796
rect 38526 2794 38582 2796
rect 38286 2742 38312 2794
rect 38312 2742 38342 2794
rect 38366 2742 38376 2794
rect 38376 2742 38422 2794
rect 38446 2742 38492 2794
rect 38492 2742 38502 2794
rect 38526 2742 38556 2794
rect 38556 2742 38582 2794
rect 38286 2740 38342 2742
rect 38366 2740 38422 2742
rect 38446 2740 38502 2742
rect 38526 2740 38582 2742
rect 69004 31932 69060 31968
rect 69004 31912 69006 31932
rect 69006 31912 69058 31932
rect 69058 31912 69060 31932
rect 69648 31948 69650 31968
rect 69650 31948 69702 31968
rect 69702 31948 69704 31968
rect 69648 31912 69704 31948
rect 72918 39242 72974 39244
rect 72998 39242 73054 39244
rect 73078 39242 73134 39244
rect 73158 39242 73214 39244
rect 72918 39190 72944 39242
rect 72944 39190 72974 39242
rect 72998 39190 73008 39242
rect 73008 39190 73054 39242
rect 73078 39190 73124 39242
rect 73124 39190 73134 39242
rect 73158 39190 73188 39242
rect 73188 39190 73214 39242
rect 72918 39188 72974 39190
rect 72998 39188 73054 39190
rect 73078 39188 73134 39190
rect 73158 39188 73214 39190
rect 72918 38154 72974 38156
rect 72998 38154 73054 38156
rect 73078 38154 73134 38156
rect 73158 38154 73214 38156
rect 72918 38102 72944 38154
rect 72944 38102 72974 38154
rect 72998 38102 73008 38154
rect 73008 38102 73054 38154
rect 73078 38102 73124 38154
rect 73124 38102 73134 38154
rect 73158 38102 73188 38154
rect 73188 38102 73214 38154
rect 72918 38100 72974 38102
rect 72998 38100 73054 38102
rect 73078 38100 73134 38102
rect 73158 38100 73214 38102
rect 72918 37066 72974 37068
rect 72998 37066 73054 37068
rect 73078 37066 73134 37068
rect 73158 37066 73214 37068
rect 72918 37014 72944 37066
rect 72944 37014 72974 37066
rect 72998 37014 73008 37066
rect 73008 37014 73054 37066
rect 73078 37014 73124 37066
rect 73124 37014 73134 37066
rect 73158 37014 73188 37066
rect 73188 37014 73214 37066
rect 72918 37012 72974 37014
rect 72998 37012 73054 37014
rect 73078 37012 73134 37014
rect 73158 37012 73214 37014
rect 70254 36522 70310 36524
rect 70334 36522 70390 36524
rect 70414 36522 70470 36524
rect 70494 36522 70550 36524
rect 70254 36470 70280 36522
rect 70280 36470 70310 36522
rect 70334 36470 70344 36522
rect 70344 36470 70390 36522
rect 70414 36470 70460 36522
rect 70460 36470 70470 36522
rect 70494 36470 70524 36522
rect 70524 36470 70550 36522
rect 70254 36468 70310 36470
rect 70334 36468 70390 36470
rect 70414 36468 70470 36470
rect 70494 36468 70550 36470
rect 75582 41962 75638 41964
rect 75662 41962 75718 41964
rect 75742 41962 75798 41964
rect 75822 41962 75878 41964
rect 75582 41910 75608 41962
rect 75608 41910 75638 41962
rect 75662 41910 75672 41962
rect 75672 41910 75718 41962
rect 75742 41910 75788 41962
rect 75788 41910 75798 41962
rect 75822 41910 75852 41962
rect 75852 41910 75878 41962
rect 75582 41908 75638 41910
rect 75662 41908 75718 41910
rect 75742 41908 75798 41910
rect 75822 41908 75878 41910
rect 75582 40874 75638 40876
rect 75662 40874 75718 40876
rect 75742 40874 75798 40876
rect 75822 40874 75878 40876
rect 75582 40822 75608 40874
rect 75608 40822 75638 40874
rect 75662 40822 75672 40874
rect 75672 40822 75718 40874
rect 75742 40822 75788 40874
rect 75788 40822 75798 40874
rect 75822 40822 75852 40874
rect 75852 40822 75878 40874
rect 75582 40820 75638 40822
rect 75662 40820 75718 40822
rect 75742 40820 75798 40822
rect 75822 40820 75878 40822
rect 78246 41418 78302 41420
rect 78326 41418 78382 41420
rect 78406 41418 78462 41420
rect 78486 41418 78542 41420
rect 78246 41366 78272 41418
rect 78272 41366 78302 41418
rect 78326 41366 78336 41418
rect 78336 41366 78382 41418
rect 78406 41366 78452 41418
rect 78452 41366 78462 41418
rect 78486 41366 78516 41418
rect 78516 41366 78542 41418
rect 78246 41364 78302 41366
rect 78326 41364 78382 41366
rect 78406 41364 78462 41366
rect 78486 41364 78542 41366
rect 75582 39786 75638 39788
rect 75662 39786 75718 39788
rect 75742 39786 75798 39788
rect 75822 39786 75878 39788
rect 75582 39734 75608 39786
rect 75608 39734 75638 39786
rect 75662 39734 75672 39786
rect 75672 39734 75718 39786
rect 75742 39734 75788 39786
rect 75788 39734 75798 39786
rect 75822 39734 75852 39786
rect 75852 39734 75878 39786
rect 75582 39732 75638 39734
rect 75662 39732 75718 39734
rect 75742 39732 75798 39734
rect 75822 39732 75878 39734
rect 75444 39528 75500 39584
rect 75582 38698 75638 38700
rect 75662 38698 75718 38700
rect 75742 38698 75798 38700
rect 75822 38698 75878 38700
rect 75582 38646 75608 38698
rect 75608 38646 75638 38698
rect 75662 38646 75672 38698
rect 75672 38646 75718 38698
rect 75742 38646 75788 38698
rect 75788 38646 75798 38698
rect 75822 38646 75852 38698
rect 75852 38646 75878 38698
rect 75582 38644 75638 38646
rect 75662 38644 75718 38646
rect 75742 38644 75798 38646
rect 75822 38644 75878 38646
rect 72918 35978 72974 35980
rect 72998 35978 73054 35980
rect 73078 35978 73134 35980
rect 73158 35978 73214 35980
rect 72918 35926 72944 35978
rect 72944 35926 72974 35978
rect 72998 35926 73008 35978
rect 73008 35926 73054 35978
rect 73078 35926 73124 35978
rect 73124 35926 73134 35978
rect 73158 35926 73188 35978
rect 73188 35926 73214 35978
rect 72918 35924 72974 35926
rect 72998 35924 73054 35926
rect 73078 35924 73134 35926
rect 73158 35924 73214 35926
rect 70254 35434 70310 35436
rect 70334 35434 70390 35436
rect 70414 35434 70470 35436
rect 70494 35434 70550 35436
rect 70254 35382 70280 35434
rect 70280 35382 70310 35434
rect 70334 35382 70344 35434
rect 70344 35382 70390 35434
rect 70414 35382 70460 35434
rect 70460 35382 70470 35434
rect 70494 35382 70524 35434
rect 70524 35382 70550 35434
rect 70254 35380 70310 35382
rect 70334 35380 70390 35382
rect 70414 35380 70470 35382
rect 70494 35380 70550 35382
rect 72918 34890 72974 34892
rect 72998 34890 73054 34892
rect 73078 34890 73134 34892
rect 73158 34890 73214 34892
rect 72918 34838 72944 34890
rect 72944 34838 72974 34890
rect 72998 34838 73008 34890
rect 73008 34838 73054 34890
rect 73078 34838 73124 34890
rect 73124 34838 73134 34890
rect 73158 34838 73188 34890
rect 73188 34838 73214 34890
rect 72918 34836 72974 34838
rect 72998 34836 73054 34838
rect 73078 34836 73134 34838
rect 73158 34836 73214 34838
rect 70254 34346 70310 34348
rect 70334 34346 70390 34348
rect 70414 34346 70470 34348
rect 70494 34346 70550 34348
rect 70254 34294 70280 34346
rect 70280 34294 70310 34346
rect 70334 34294 70344 34346
rect 70344 34294 70390 34346
rect 70414 34294 70460 34346
rect 70460 34294 70470 34346
rect 70494 34294 70524 34346
rect 70524 34294 70550 34346
rect 70254 34292 70310 34294
rect 70334 34292 70390 34294
rect 70414 34292 70470 34294
rect 70494 34292 70550 34294
rect 72918 33802 72974 33804
rect 72998 33802 73054 33804
rect 73078 33802 73134 33804
rect 73158 33802 73214 33804
rect 72918 33750 72944 33802
rect 72944 33750 72974 33802
rect 72998 33750 73008 33802
rect 73008 33750 73054 33802
rect 73078 33750 73124 33802
rect 73124 33750 73134 33802
rect 73158 33750 73188 33802
rect 73188 33750 73214 33802
rect 72918 33748 72974 33750
rect 72998 33748 73054 33750
rect 73078 33748 73134 33750
rect 73158 33748 73214 33750
rect 74156 37216 74212 37272
rect 74248 36672 74304 36728
rect 74064 33988 74066 34008
rect 74066 33988 74118 34008
rect 74118 33988 74120 34008
rect 74064 33952 74120 33988
rect 70254 33258 70310 33260
rect 70334 33258 70390 33260
rect 70414 33258 70470 33260
rect 70494 33258 70550 33260
rect 70254 33206 70280 33258
rect 70280 33206 70310 33258
rect 70334 33206 70344 33258
rect 70344 33206 70390 33258
rect 70414 33206 70460 33258
rect 70460 33206 70470 33258
rect 70494 33206 70524 33258
rect 70524 33206 70550 33258
rect 70254 33204 70310 33206
rect 70334 33204 70390 33206
rect 70414 33204 70470 33206
rect 70494 33204 70550 33206
rect 70254 32170 70310 32172
rect 70334 32170 70390 32172
rect 70414 32170 70470 32172
rect 70494 32170 70550 32172
rect 70254 32118 70280 32170
rect 70280 32118 70310 32170
rect 70334 32118 70344 32170
rect 70344 32118 70390 32170
rect 70414 32118 70460 32170
rect 70460 32118 70470 32170
rect 70494 32118 70524 32170
rect 70524 32118 70550 32170
rect 70254 32116 70310 32118
rect 70334 32116 70390 32118
rect 70414 32116 70470 32118
rect 70494 32116 70550 32118
rect 70254 31082 70310 31084
rect 70334 31082 70390 31084
rect 70414 31082 70470 31084
rect 70494 31082 70550 31084
rect 70254 31030 70280 31082
rect 70280 31030 70310 31082
rect 70334 31030 70344 31082
rect 70344 31030 70390 31082
rect 70414 31030 70460 31082
rect 70460 31030 70470 31082
rect 70494 31030 70524 31082
rect 70524 31030 70550 31082
rect 70254 31028 70310 31030
rect 70334 31028 70390 31030
rect 70414 31028 70470 31030
rect 70494 31028 70550 31030
rect 72918 32714 72974 32716
rect 72998 32714 73054 32716
rect 73078 32714 73134 32716
rect 73158 32714 73214 32716
rect 72918 32662 72944 32714
rect 72944 32662 72974 32714
rect 72998 32662 73008 32714
rect 73008 32662 73054 32714
rect 73078 32662 73124 32714
rect 73124 32662 73134 32714
rect 73158 32662 73188 32714
rect 73188 32662 73214 32714
rect 72918 32660 72974 32662
rect 72998 32660 73054 32662
rect 73078 32660 73134 32662
rect 73158 32660 73214 32662
rect 73696 32356 73698 32376
rect 73698 32356 73750 32376
rect 73750 32356 73752 32376
rect 73696 32320 73752 32356
rect 69832 30300 69888 30336
rect 69832 30280 69834 30300
rect 69834 30280 69886 30300
rect 69886 30280 69888 30300
rect 70254 29994 70310 29996
rect 70334 29994 70390 29996
rect 70414 29994 70470 29996
rect 70494 29994 70550 29996
rect 70254 29942 70280 29994
rect 70280 29942 70310 29994
rect 70334 29942 70344 29994
rect 70344 29942 70390 29994
rect 70414 29942 70460 29994
rect 70460 29942 70470 29994
rect 70494 29942 70524 29994
rect 70524 29942 70550 29994
rect 70254 29940 70310 29942
rect 70334 29940 70390 29942
rect 70414 29940 70470 29942
rect 70494 29940 70550 29942
rect 68176 20216 68232 20272
rect 67164 19980 67166 20000
rect 67166 19980 67218 20000
rect 67218 19980 67220 20000
rect 67164 19944 67220 19980
rect 68360 23480 68416 23536
rect 68268 19128 68324 19184
rect 68268 18448 68324 18504
rect 43520 18040 43576 18096
rect 67072 18040 67128 18096
rect 68268 17904 68324 17960
rect 43336 16952 43392 17008
rect 43520 14776 43576 14832
rect 68360 16544 68416 16600
rect 43520 10424 43576 10480
rect 68268 10424 68324 10480
rect 70254 28906 70310 28908
rect 70334 28906 70390 28908
rect 70414 28906 70470 28908
rect 70494 28906 70550 28908
rect 70254 28854 70280 28906
rect 70280 28854 70310 28906
rect 70334 28854 70344 28906
rect 70344 28854 70390 28906
rect 70414 28854 70460 28906
rect 70460 28854 70470 28906
rect 70494 28854 70524 28906
rect 70524 28854 70550 28906
rect 70254 28852 70310 28854
rect 70334 28852 70390 28854
rect 70414 28852 70470 28854
rect 70494 28852 70550 28854
rect 70254 27818 70310 27820
rect 70334 27818 70390 27820
rect 70414 27818 70470 27820
rect 70494 27818 70550 27820
rect 70254 27766 70280 27818
rect 70280 27766 70310 27818
rect 70334 27766 70344 27818
rect 70344 27766 70390 27818
rect 70414 27766 70460 27818
rect 70460 27766 70470 27818
rect 70494 27766 70524 27818
rect 70524 27766 70550 27818
rect 70254 27764 70310 27766
rect 70334 27764 70390 27766
rect 70414 27764 70470 27766
rect 70494 27764 70550 27766
rect 72918 31626 72974 31628
rect 72998 31626 73054 31628
rect 73078 31626 73134 31628
rect 73158 31626 73214 31628
rect 72918 31574 72944 31626
rect 72944 31574 72974 31626
rect 72998 31574 73008 31626
rect 73008 31574 73054 31626
rect 73078 31574 73124 31626
rect 73124 31574 73134 31626
rect 73158 31574 73188 31626
rect 73188 31574 73214 31626
rect 72918 31572 72974 31574
rect 72998 31572 73054 31574
rect 73078 31572 73134 31574
rect 73158 31572 73214 31574
rect 72918 30538 72974 30540
rect 72998 30538 73054 30540
rect 73078 30538 73134 30540
rect 73158 30538 73214 30540
rect 72918 30486 72944 30538
rect 72944 30486 72974 30538
rect 72998 30486 73008 30538
rect 73008 30486 73054 30538
rect 73078 30486 73124 30538
rect 73124 30486 73134 30538
rect 73158 30486 73188 30538
rect 73188 30486 73214 30538
rect 72918 30484 72974 30486
rect 72998 30484 73054 30486
rect 73078 30484 73134 30486
rect 73158 30484 73214 30486
rect 75582 37610 75638 37612
rect 75662 37610 75718 37612
rect 75742 37610 75798 37612
rect 75822 37610 75878 37612
rect 75582 37558 75608 37610
rect 75608 37558 75638 37610
rect 75662 37558 75672 37610
rect 75672 37558 75718 37610
rect 75742 37558 75788 37610
rect 75788 37558 75798 37610
rect 75822 37558 75852 37610
rect 75852 37558 75878 37610
rect 75582 37556 75638 37558
rect 75662 37556 75718 37558
rect 75742 37556 75798 37558
rect 75822 37556 75878 37558
rect 75582 36522 75638 36524
rect 75662 36522 75718 36524
rect 75742 36522 75798 36524
rect 75822 36522 75878 36524
rect 75582 36470 75608 36522
rect 75608 36470 75638 36522
rect 75662 36470 75672 36522
rect 75672 36470 75718 36522
rect 75742 36470 75788 36522
rect 75788 36470 75798 36522
rect 75822 36470 75852 36522
rect 75852 36470 75878 36522
rect 75582 36468 75638 36470
rect 75662 36468 75718 36470
rect 75742 36468 75798 36470
rect 75822 36468 75878 36470
rect 75582 35434 75638 35436
rect 75662 35434 75718 35436
rect 75742 35434 75798 35436
rect 75822 35434 75878 35436
rect 75582 35382 75608 35434
rect 75608 35382 75638 35434
rect 75662 35382 75672 35434
rect 75672 35382 75718 35434
rect 75742 35382 75788 35434
rect 75788 35382 75798 35434
rect 75822 35382 75852 35434
rect 75852 35382 75878 35434
rect 75582 35380 75638 35382
rect 75662 35380 75718 35382
rect 75742 35380 75798 35382
rect 75822 35380 75878 35382
rect 75582 34346 75638 34348
rect 75662 34346 75718 34348
rect 75742 34346 75798 34348
rect 75822 34346 75878 34348
rect 75582 34294 75608 34346
rect 75608 34294 75638 34346
rect 75662 34294 75672 34346
rect 75672 34294 75718 34346
rect 75742 34294 75788 34346
rect 75788 34294 75798 34346
rect 75822 34294 75852 34346
rect 75852 34294 75878 34346
rect 75582 34292 75638 34294
rect 75662 34292 75718 34294
rect 75742 34292 75798 34294
rect 75822 34292 75878 34294
rect 75582 33258 75638 33260
rect 75662 33258 75718 33260
rect 75742 33258 75798 33260
rect 75822 33258 75878 33260
rect 75582 33206 75608 33258
rect 75608 33206 75638 33258
rect 75662 33206 75672 33258
rect 75672 33206 75718 33258
rect 75742 33206 75788 33258
rect 75788 33206 75798 33258
rect 75822 33206 75852 33258
rect 75852 33206 75878 33258
rect 75582 33204 75638 33206
rect 75662 33204 75718 33206
rect 75742 33204 75798 33206
rect 75822 33204 75878 33206
rect 74616 32320 74672 32376
rect 78246 40330 78302 40332
rect 78326 40330 78382 40332
rect 78406 40330 78462 40332
rect 78486 40330 78542 40332
rect 78246 40278 78272 40330
rect 78272 40278 78302 40330
rect 78326 40278 78336 40330
rect 78336 40278 78382 40330
rect 78406 40278 78452 40330
rect 78452 40278 78462 40330
rect 78486 40278 78516 40330
rect 78516 40278 78542 40330
rect 78246 40276 78302 40278
rect 78326 40276 78382 40278
rect 78406 40276 78462 40278
rect 78486 40276 78542 40278
rect 80910 41962 80966 41964
rect 80990 41962 81046 41964
rect 81070 41962 81126 41964
rect 81150 41962 81206 41964
rect 80910 41910 80936 41962
rect 80936 41910 80966 41962
rect 80990 41910 81000 41962
rect 81000 41910 81046 41962
rect 81070 41910 81116 41962
rect 81116 41910 81126 41962
rect 81150 41910 81180 41962
rect 81180 41910 81206 41962
rect 80910 41908 80966 41910
rect 80990 41908 81046 41910
rect 81070 41908 81126 41910
rect 81150 41908 81206 41910
rect 80910 40874 80966 40876
rect 80990 40874 81046 40876
rect 81070 40874 81126 40876
rect 81150 40874 81206 40876
rect 80910 40822 80936 40874
rect 80936 40822 80966 40874
rect 80990 40822 81000 40874
rect 81000 40822 81046 40874
rect 81070 40822 81116 40874
rect 81116 40822 81126 40874
rect 81150 40822 81180 40874
rect 81180 40822 81206 40874
rect 80910 40820 80966 40822
rect 80990 40820 81046 40822
rect 81070 40820 81126 40822
rect 81150 40820 81206 40822
rect 80910 39786 80966 39788
rect 80990 39786 81046 39788
rect 81070 39786 81126 39788
rect 81150 39786 81206 39788
rect 80910 39734 80936 39786
rect 80936 39734 80966 39786
rect 80990 39734 81000 39786
rect 81000 39734 81046 39786
rect 81070 39734 81116 39786
rect 81116 39734 81126 39786
rect 81150 39734 81180 39786
rect 81180 39734 81206 39786
rect 80910 39732 80966 39734
rect 80990 39732 81046 39734
rect 81070 39732 81126 39734
rect 81150 39732 81206 39734
rect 78246 39242 78302 39244
rect 78326 39242 78382 39244
rect 78406 39242 78462 39244
rect 78486 39242 78542 39244
rect 78246 39190 78272 39242
rect 78272 39190 78302 39242
rect 78326 39190 78336 39242
rect 78336 39190 78382 39242
rect 78406 39190 78452 39242
rect 78452 39190 78462 39242
rect 78486 39190 78516 39242
rect 78516 39190 78542 39242
rect 78246 39188 78302 39190
rect 78326 39188 78382 39190
rect 78406 39188 78462 39190
rect 78486 39188 78542 39190
rect 78246 38154 78302 38156
rect 78326 38154 78382 38156
rect 78406 38154 78462 38156
rect 78486 38154 78542 38156
rect 78246 38102 78272 38154
rect 78272 38102 78302 38154
rect 78326 38102 78336 38154
rect 78336 38102 78382 38154
rect 78406 38102 78452 38154
rect 78452 38102 78462 38154
rect 78486 38102 78516 38154
rect 78516 38102 78542 38154
rect 78246 38100 78302 38102
rect 78326 38100 78382 38102
rect 78406 38100 78462 38102
rect 78486 38100 78542 38102
rect 78246 37066 78302 37068
rect 78326 37066 78382 37068
rect 78406 37066 78462 37068
rect 78486 37066 78542 37068
rect 78246 37014 78272 37066
rect 78272 37014 78302 37066
rect 78326 37014 78336 37066
rect 78336 37014 78382 37066
rect 78406 37014 78452 37066
rect 78452 37014 78462 37066
rect 78486 37014 78516 37066
rect 78516 37014 78542 37066
rect 78246 37012 78302 37014
rect 78326 37012 78382 37014
rect 78406 37012 78462 37014
rect 78486 37012 78542 37014
rect 78246 35978 78302 35980
rect 78326 35978 78382 35980
rect 78406 35978 78462 35980
rect 78486 35978 78542 35980
rect 78246 35926 78272 35978
rect 78272 35926 78302 35978
rect 78326 35926 78336 35978
rect 78336 35926 78382 35978
rect 78406 35926 78452 35978
rect 78452 35926 78462 35978
rect 78486 35926 78516 35978
rect 78516 35926 78542 35978
rect 78246 35924 78302 35926
rect 78326 35924 78382 35926
rect 78406 35924 78462 35926
rect 78486 35924 78542 35926
rect 78246 34890 78302 34892
rect 78326 34890 78382 34892
rect 78406 34890 78462 34892
rect 78486 34890 78542 34892
rect 78246 34838 78272 34890
rect 78272 34838 78302 34890
rect 78326 34838 78336 34890
rect 78336 34838 78382 34890
rect 78406 34838 78452 34890
rect 78452 34838 78462 34890
rect 78486 34838 78516 34890
rect 78516 34838 78542 34890
rect 78246 34836 78302 34838
rect 78326 34836 78382 34838
rect 78406 34836 78462 34838
rect 78486 34836 78542 34838
rect 78246 33802 78302 33804
rect 78326 33802 78382 33804
rect 78406 33802 78462 33804
rect 78486 33802 78542 33804
rect 78246 33750 78272 33802
rect 78272 33750 78302 33802
rect 78326 33750 78336 33802
rect 78336 33750 78382 33802
rect 78406 33750 78452 33802
rect 78452 33750 78462 33802
rect 78486 33750 78516 33802
rect 78516 33750 78542 33802
rect 78246 33748 78302 33750
rect 78326 33748 78382 33750
rect 78406 33748 78462 33750
rect 78486 33748 78542 33750
rect 78246 32714 78302 32716
rect 78326 32714 78382 32716
rect 78406 32714 78462 32716
rect 78486 32714 78542 32716
rect 78246 32662 78272 32714
rect 78272 32662 78302 32714
rect 78326 32662 78336 32714
rect 78336 32662 78382 32714
rect 78406 32662 78452 32714
rect 78452 32662 78462 32714
rect 78486 32662 78516 32714
rect 78516 32662 78542 32714
rect 78246 32660 78302 32662
rect 78326 32660 78382 32662
rect 78406 32660 78462 32662
rect 78486 32660 78542 32662
rect 75582 32170 75638 32172
rect 75662 32170 75718 32172
rect 75742 32170 75798 32172
rect 75822 32170 75878 32172
rect 75582 32118 75608 32170
rect 75608 32118 75638 32170
rect 75662 32118 75672 32170
rect 75672 32118 75718 32170
rect 75742 32118 75788 32170
rect 75788 32118 75798 32170
rect 75822 32118 75852 32170
rect 75852 32118 75878 32170
rect 75582 32116 75638 32118
rect 75662 32116 75718 32118
rect 75742 32116 75798 32118
rect 75822 32116 75878 32118
rect 74524 30280 74580 30336
rect 75582 31082 75638 31084
rect 75662 31082 75718 31084
rect 75742 31082 75798 31084
rect 75822 31082 75878 31084
rect 75582 31030 75608 31082
rect 75608 31030 75638 31082
rect 75662 31030 75672 31082
rect 75672 31030 75718 31082
rect 75742 31030 75788 31082
rect 75788 31030 75798 31082
rect 75822 31030 75852 31082
rect 75852 31030 75878 31082
rect 75582 31028 75638 31030
rect 75662 31028 75718 31030
rect 75742 31028 75798 31030
rect 75822 31028 75878 31030
rect 74984 29756 75040 29792
rect 74984 29736 74986 29756
rect 74986 29736 75038 29756
rect 75038 29736 75040 29756
rect 72918 29450 72974 29452
rect 72998 29450 73054 29452
rect 73078 29450 73134 29452
rect 73158 29450 73214 29452
rect 72918 29398 72944 29450
rect 72944 29398 72974 29450
rect 72998 29398 73008 29450
rect 73008 29398 73054 29450
rect 73078 29398 73124 29450
rect 73124 29398 73134 29450
rect 73158 29398 73188 29450
rect 73188 29398 73214 29450
rect 72918 29396 72974 29398
rect 72998 29396 73054 29398
rect 73078 29396 73134 29398
rect 73158 29396 73214 29398
rect 75582 29994 75638 29996
rect 75662 29994 75718 29996
rect 75742 29994 75798 29996
rect 75822 29994 75878 29996
rect 75582 29942 75608 29994
rect 75608 29942 75638 29994
rect 75662 29942 75672 29994
rect 75672 29942 75718 29994
rect 75742 29942 75788 29994
rect 75788 29942 75798 29994
rect 75822 29942 75852 29994
rect 75852 29942 75878 29994
rect 75582 29940 75638 29942
rect 75662 29940 75718 29942
rect 75742 29940 75798 29942
rect 75822 29940 75878 29942
rect 72918 28362 72974 28364
rect 72998 28362 73054 28364
rect 73078 28362 73134 28364
rect 73158 28362 73214 28364
rect 72918 28310 72944 28362
rect 72944 28310 72974 28362
rect 72998 28310 73008 28362
rect 73008 28310 73054 28362
rect 73078 28310 73124 28362
rect 73124 28310 73134 28362
rect 73158 28310 73188 28362
rect 73188 28310 73214 28362
rect 72918 28308 72974 28310
rect 72998 28308 73054 28310
rect 73078 28308 73134 28310
rect 73158 28308 73214 28310
rect 72918 27274 72974 27276
rect 72998 27274 73054 27276
rect 73078 27274 73134 27276
rect 73158 27274 73214 27276
rect 72918 27222 72944 27274
rect 72944 27222 72974 27274
rect 72998 27222 73008 27274
rect 73008 27222 73054 27274
rect 73078 27222 73124 27274
rect 73124 27222 73134 27274
rect 73158 27222 73188 27274
rect 73188 27222 73214 27274
rect 72918 27220 72974 27222
rect 72998 27220 73054 27222
rect 73078 27220 73134 27222
rect 73158 27220 73214 27222
rect 75582 28906 75638 28908
rect 75662 28906 75718 28908
rect 75742 28906 75798 28908
rect 75822 28906 75878 28908
rect 75582 28854 75608 28906
rect 75608 28854 75638 28906
rect 75662 28854 75672 28906
rect 75672 28854 75718 28906
rect 75742 28854 75788 28906
rect 75788 28854 75798 28906
rect 75822 28854 75852 28906
rect 75852 28854 75878 28906
rect 75582 28852 75638 28854
rect 75662 28852 75718 28854
rect 75742 28852 75798 28854
rect 75822 28852 75878 28854
rect 75582 27818 75638 27820
rect 75662 27818 75718 27820
rect 75742 27818 75798 27820
rect 75822 27818 75878 27820
rect 75582 27766 75608 27818
rect 75608 27766 75638 27818
rect 75662 27766 75672 27818
rect 75672 27766 75718 27818
rect 75742 27766 75788 27818
rect 75788 27766 75798 27818
rect 75822 27766 75852 27818
rect 75852 27766 75878 27818
rect 75582 27764 75638 27766
rect 75662 27764 75718 27766
rect 75742 27764 75798 27766
rect 75822 27764 75878 27766
rect 76640 29736 76696 29792
rect 78246 31626 78302 31628
rect 78326 31626 78382 31628
rect 78406 31626 78462 31628
rect 78486 31626 78542 31628
rect 78246 31574 78272 31626
rect 78272 31574 78302 31626
rect 78326 31574 78336 31626
rect 78336 31574 78382 31626
rect 78406 31574 78452 31626
rect 78452 31574 78462 31626
rect 78486 31574 78516 31626
rect 78516 31574 78542 31626
rect 78246 31572 78302 31574
rect 78326 31572 78382 31574
rect 78406 31572 78462 31574
rect 78486 31572 78542 31574
rect 78246 30538 78302 30540
rect 78326 30538 78382 30540
rect 78406 30538 78462 30540
rect 78486 30538 78542 30540
rect 78246 30486 78272 30538
rect 78272 30486 78302 30538
rect 78326 30486 78336 30538
rect 78336 30486 78382 30538
rect 78406 30486 78452 30538
rect 78452 30486 78462 30538
rect 78486 30486 78516 30538
rect 78516 30486 78542 30538
rect 78246 30484 78302 30486
rect 78326 30484 78382 30486
rect 78406 30484 78462 30486
rect 78486 30484 78542 30486
rect 78246 29450 78302 29452
rect 78326 29450 78382 29452
rect 78406 29450 78462 29452
rect 78486 29450 78542 29452
rect 78246 29398 78272 29450
rect 78272 29398 78302 29450
rect 78326 29398 78336 29450
rect 78336 29398 78382 29450
rect 78406 29398 78452 29450
rect 78452 29398 78462 29450
rect 78486 29398 78516 29450
rect 78516 29398 78542 29450
rect 78246 29396 78302 29398
rect 78326 29396 78382 29398
rect 78406 29396 78462 29398
rect 78486 29396 78542 29398
rect 78246 28362 78302 28364
rect 78326 28362 78382 28364
rect 78406 28362 78462 28364
rect 78486 28362 78542 28364
rect 78246 28310 78272 28362
rect 78272 28310 78302 28362
rect 78326 28310 78336 28362
rect 78336 28310 78382 28362
rect 78406 28310 78452 28362
rect 78452 28310 78462 28362
rect 78486 28310 78516 28362
rect 78516 28310 78542 28362
rect 78246 28308 78302 28310
rect 78326 28308 78382 28310
rect 78406 28308 78462 28310
rect 78486 28308 78542 28310
rect 80910 38698 80966 38700
rect 80990 38698 81046 38700
rect 81070 38698 81126 38700
rect 81150 38698 81206 38700
rect 80910 38646 80936 38698
rect 80936 38646 80966 38698
rect 80990 38646 81000 38698
rect 81000 38646 81046 38698
rect 81070 38646 81116 38698
rect 81116 38646 81126 38698
rect 81150 38646 81180 38698
rect 81180 38646 81206 38698
rect 80910 38644 80966 38646
rect 80990 38644 81046 38646
rect 81070 38644 81126 38646
rect 81150 38644 81206 38646
rect 80910 37610 80966 37612
rect 80990 37610 81046 37612
rect 81070 37610 81126 37612
rect 81150 37610 81206 37612
rect 80910 37558 80936 37610
rect 80936 37558 80966 37610
rect 80990 37558 81000 37610
rect 81000 37558 81046 37610
rect 81070 37558 81116 37610
rect 81116 37558 81126 37610
rect 81150 37558 81180 37610
rect 81180 37558 81206 37610
rect 80910 37556 80966 37558
rect 80990 37556 81046 37558
rect 81070 37556 81126 37558
rect 81150 37556 81206 37558
rect 80910 36522 80966 36524
rect 80990 36522 81046 36524
rect 81070 36522 81126 36524
rect 81150 36522 81206 36524
rect 80910 36470 80936 36522
rect 80936 36470 80966 36522
rect 80990 36470 81000 36522
rect 81000 36470 81046 36522
rect 81070 36470 81116 36522
rect 81116 36470 81126 36522
rect 81150 36470 81180 36522
rect 81180 36470 81206 36522
rect 80910 36468 80966 36470
rect 80990 36468 81046 36470
rect 81070 36468 81126 36470
rect 81150 36468 81206 36470
rect 80910 35434 80966 35436
rect 80990 35434 81046 35436
rect 81070 35434 81126 35436
rect 81150 35434 81206 35436
rect 80910 35382 80936 35434
rect 80936 35382 80966 35434
rect 80990 35382 81000 35434
rect 81000 35382 81046 35434
rect 81070 35382 81116 35434
rect 81116 35382 81126 35434
rect 81150 35382 81180 35434
rect 81180 35382 81206 35434
rect 80910 35380 80966 35382
rect 80990 35380 81046 35382
rect 81070 35380 81126 35382
rect 81150 35380 81206 35382
rect 80910 34346 80966 34348
rect 80990 34346 81046 34348
rect 81070 34346 81126 34348
rect 81150 34346 81206 34348
rect 80910 34294 80936 34346
rect 80936 34294 80966 34346
rect 80990 34294 81000 34346
rect 81000 34294 81046 34346
rect 81070 34294 81116 34346
rect 81116 34294 81126 34346
rect 81150 34294 81180 34346
rect 81180 34294 81206 34346
rect 80910 34292 80966 34294
rect 80990 34292 81046 34294
rect 81070 34292 81126 34294
rect 81150 34292 81206 34294
rect 80910 33258 80966 33260
rect 80990 33258 81046 33260
rect 81070 33258 81126 33260
rect 81150 33258 81206 33260
rect 80910 33206 80936 33258
rect 80936 33206 80966 33258
rect 80990 33206 81000 33258
rect 81000 33206 81046 33258
rect 81070 33206 81116 33258
rect 81116 33206 81126 33258
rect 81150 33206 81180 33258
rect 81180 33206 81206 33258
rect 80910 33204 80966 33206
rect 80990 33204 81046 33206
rect 81070 33204 81126 33206
rect 81150 33204 81206 33206
rect 83574 41418 83630 41420
rect 83654 41418 83710 41420
rect 83734 41418 83790 41420
rect 83814 41418 83870 41420
rect 83574 41366 83600 41418
rect 83600 41366 83630 41418
rect 83654 41366 83664 41418
rect 83664 41366 83710 41418
rect 83734 41366 83780 41418
rect 83780 41366 83790 41418
rect 83814 41366 83844 41418
rect 83844 41366 83870 41418
rect 83574 41364 83630 41366
rect 83654 41364 83710 41366
rect 83734 41364 83790 41366
rect 83814 41364 83870 41366
rect 83574 40330 83630 40332
rect 83654 40330 83710 40332
rect 83734 40330 83790 40332
rect 83814 40330 83870 40332
rect 83574 40278 83600 40330
rect 83600 40278 83630 40330
rect 83654 40278 83664 40330
rect 83664 40278 83710 40330
rect 83734 40278 83780 40330
rect 83780 40278 83790 40330
rect 83814 40278 83844 40330
rect 83844 40278 83870 40330
rect 83574 40276 83630 40278
rect 83654 40276 83710 40278
rect 83734 40276 83790 40278
rect 83814 40276 83870 40278
rect 83574 39242 83630 39244
rect 83654 39242 83710 39244
rect 83734 39242 83790 39244
rect 83814 39242 83870 39244
rect 83574 39190 83600 39242
rect 83600 39190 83630 39242
rect 83654 39190 83664 39242
rect 83664 39190 83710 39242
rect 83734 39190 83780 39242
rect 83780 39190 83790 39242
rect 83814 39190 83844 39242
rect 83844 39190 83870 39242
rect 83574 39188 83630 39190
rect 83654 39188 83710 39190
rect 83734 39188 83790 39190
rect 83814 39188 83870 39190
rect 83574 38154 83630 38156
rect 83654 38154 83710 38156
rect 83734 38154 83790 38156
rect 83814 38154 83870 38156
rect 83574 38102 83600 38154
rect 83600 38102 83630 38154
rect 83654 38102 83664 38154
rect 83664 38102 83710 38154
rect 83734 38102 83780 38154
rect 83780 38102 83790 38154
rect 83814 38102 83844 38154
rect 83844 38102 83870 38154
rect 83574 38100 83630 38102
rect 83654 38100 83710 38102
rect 83734 38100 83790 38102
rect 83814 38100 83870 38102
rect 83574 37066 83630 37068
rect 83654 37066 83710 37068
rect 83734 37066 83790 37068
rect 83814 37066 83870 37068
rect 83574 37014 83600 37066
rect 83600 37014 83630 37066
rect 83654 37014 83664 37066
rect 83664 37014 83710 37066
rect 83734 37014 83780 37066
rect 83780 37014 83790 37066
rect 83814 37014 83844 37066
rect 83844 37014 83870 37066
rect 83574 37012 83630 37014
rect 83654 37012 83710 37014
rect 83734 37012 83790 37014
rect 83814 37012 83870 37014
rect 83574 35978 83630 35980
rect 83654 35978 83710 35980
rect 83734 35978 83790 35980
rect 83814 35978 83870 35980
rect 83574 35926 83600 35978
rect 83600 35926 83630 35978
rect 83654 35926 83664 35978
rect 83664 35926 83710 35978
rect 83734 35926 83780 35978
rect 83780 35926 83790 35978
rect 83814 35926 83844 35978
rect 83844 35926 83870 35978
rect 83574 35924 83630 35926
rect 83654 35924 83710 35926
rect 83734 35924 83790 35926
rect 83814 35924 83870 35926
rect 80910 32170 80966 32172
rect 80990 32170 81046 32172
rect 81070 32170 81126 32172
rect 81150 32170 81206 32172
rect 80910 32118 80936 32170
rect 80936 32118 80966 32170
rect 80990 32118 81000 32170
rect 81000 32118 81046 32170
rect 81070 32118 81116 32170
rect 81116 32118 81126 32170
rect 81150 32118 81180 32170
rect 81180 32118 81206 32170
rect 80910 32116 80966 32118
rect 80990 32116 81046 32118
rect 81070 32116 81126 32118
rect 81150 32116 81206 32118
rect 83574 34890 83630 34892
rect 83654 34890 83710 34892
rect 83734 34890 83790 34892
rect 83814 34890 83870 34892
rect 83574 34838 83600 34890
rect 83600 34838 83630 34890
rect 83654 34838 83664 34890
rect 83664 34838 83710 34890
rect 83734 34838 83780 34890
rect 83780 34838 83790 34890
rect 83814 34838 83844 34890
rect 83844 34838 83870 34890
rect 83574 34836 83630 34838
rect 83654 34836 83710 34838
rect 83734 34836 83790 34838
rect 83814 34836 83870 34838
rect 83574 33802 83630 33804
rect 83654 33802 83710 33804
rect 83734 33802 83790 33804
rect 83814 33802 83870 33804
rect 83574 33750 83600 33802
rect 83600 33750 83630 33802
rect 83654 33750 83664 33802
rect 83664 33750 83710 33802
rect 83734 33750 83780 33802
rect 83780 33750 83790 33802
rect 83814 33750 83844 33802
rect 83844 33750 83870 33802
rect 83574 33748 83630 33750
rect 83654 33748 83710 33750
rect 83734 33748 83790 33750
rect 83814 33748 83870 33750
rect 86238 41962 86294 41964
rect 86318 41962 86374 41964
rect 86398 41962 86454 41964
rect 86478 41962 86534 41964
rect 86238 41910 86264 41962
rect 86264 41910 86294 41962
rect 86318 41910 86328 41962
rect 86328 41910 86374 41962
rect 86398 41910 86444 41962
rect 86444 41910 86454 41962
rect 86478 41910 86508 41962
rect 86508 41910 86534 41962
rect 86238 41908 86294 41910
rect 86318 41908 86374 41910
rect 86398 41908 86454 41910
rect 86478 41908 86534 41910
rect 88902 41418 88958 41420
rect 88982 41418 89038 41420
rect 89062 41418 89118 41420
rect 89142 41418 89198 41420
rect 88902 41366 88928 41418
rect 88928 41366 88958 41418
rect 88982 41366 88992 41418
rect 88992 41366 89038 41418
rect 89062 41366 89108 41418
rect 89108 41366 89118 41418
rect 89142 41366 89172 41418
rect 89172 41366 89198 41418
rect 88902 41364 88958 41366
rect 88982 41364 89038 41366
rect 89062 41364 89118 41366
rect 89142 41364 89198 41366
rect 86238 40874 86294 40876
rect 86318 40874 86374 40876
rect 86398 40874 86454 40876
rect 86478 40874 86534 40876
rect 86238 40822 86264 40874
rect 86264 40822 86294 40874
rect 86318 40822 86328 40874
rect 86328 40822 86374 40874
rect 86398 40822 86444 40874
rect 86444 40822 86454 40874
rect 86478 40822 86508 40874
rect 86508 40822 86534 40874
rect 86238 40820 86294 40822
rect 86318 40820 86374 40822
rect 86398 40820 86454 40822
rect 86478 40820 86534 40822
rect 86238 39786 86294 39788
rect 86318 39786 86374 39788
rect 86398 39786 86454 39788
rect 86478 39786 86534 39788
rect 86238 39734 86264 39786
rect 86264 39734 86294 39786
rect 86318 39734 86328 39786
rect 86328 39734 86374 39786
rect 86398 39734 86444 39786
rect 86444 39734 86454 39786
rect 86478 39734 86508 39786
rect 86508 39734 86534 39786
rect 86238 39732 86294 39734
rect 86318 39732 86374 39734
rect 86398 39732 86454 39734
rect 86478 39732 86534 39734
rect 86238 38698 86294 38700
rect 86318 38698 86374 38700
rect 86398 38698 86454 38700
rect 86478 38698 86534 38700
rect 86238 38646 86264 38698
rect 86264 38646 86294 38698
rect 86318 38646 86328 38698
rect 86328 38646 86374 38698
rect 86398 38646 86444 38698
rect 86444 38646 86454 38698
rect 86478 38646 86508 38698
rect 86508 38646 86534 38698
rect 86238 38644 86294 38646
rect 86318 38644 86374 38646
rect 86398 38644 86454 38646
rect 86478 38644 86534 38646
rect 86238 37610 86294 37612
rect 86318 37610 86374 37612
rect 86398 37610 86454 37612
rect 86478 37610 86534 37612
rect 86238 37558 86264 37610
rect 86264 37558 86294 37610
rect 86318 37558 86328 37610
rect 86328 37558 86374 37610
rect 86398 37558 86444 37610
rect 86444 37558 86454 37610
rect 86478 37558 86508 37610
rect 86508 37558 86534 37610
rect 86238 37556 86294 37558
rect 86318 37556 86374 37558
rect 86398 37556 86454 37558
rect 86478 37556 86534 37558
rect 86238 36522 86294 36524
rect 86318 36522 86374 36524
rect 86398 36522 86454 36524
rect 86478 36522 86534 36524
rect 86238 36470 86264 36522
rect 86264 36470 86294 36522
rect 86318 36470 86328 36522
rect 86328 36470 86374 36522
rect 86398 36470 86444 36522
rect 86444 36470 86454 36522
rect 86478 36470 86508 36522
rect 86508 36470 86534 36522
rect 86238 36468 86294 36470
rect 86318 36468 86374 36470
rect 86398 36468 86454 36470
rect 86478 36468 86534 36470
rect 88902 40330 88958 40332
rect 88982 40330 89038 40332
rect 89062 40330 89118 40332
rect 89142 40330 89198 40332
rect 88902 40278 88928 40330
rect 88928 40278 88958 40330
rect 88982 40278 88992 40330
rect 88992 40278 89038 40330
rect 89062 40278 89108 40330
rect 89108 40278 89118 40330
rect 89142 40278 89172 40330
rect 89172 40278 89198 40330
rect 88902 40276 88958 40278
rect 88982 40276 89038 40278
rect 89062 40276 89118 40278
rect 89142 40276 89198 40278
rect 88902 39242 88958 39244
rect 88982 39242 89038 39244
rect 89062 39242 89118 39244
rect 89142 39242 89198 39244
rect 88902 39190 88928 39242
rect 88928 39190 88958 39242
rect 88982 39190 88992 39242
rect 88992 39190 89038 39242
rect 89062 39190 89108 39242
rect 89108 39190 89118 39242
rect 89142 39190 89172 39242
rect 89172 39190 89198 39242
rect 88902 39188 88958 39190
rect 88982 39188 89038 39190
rect 89062 39188 89118 39190
rect 89142 39188 89198 39190
rect 88902 38154 88958 38156
rect 88982 38154 89038 38156
rect 89062 38154 89118 38156
rect 89142 38154 89198 38156
rect 88902 38102 88928 38154
rect 88928 38102 88958 38154
rect 88982 38102 88992 38154
rect 88992 38102 89038 38154
rect 89062 38102 89108 38154
rect 89108 38102 89118 38154
rect 89142 38102 89172 38154
rect 89172 38102 89198 38154
rect 88902 38100 88958 38102
rect 88982 38100 89038 38102
rect 89062 38100 89118 38102
rect 89142 38100 89198 38102
rect 88902 37066 88958 37068
rect 88982 37066 89038 37068
rect 89062 37066 89118 37068
rect 89142 37066 89198 37068
rect 88902 37014 88928 37066
rect 88928 37014 88958 37066
rect 88982 37014 88992 37066
rect 88992 37014 89038 37066
rect 89062 37014 89108 37066
rect 89108 37014 89118 37066
rect 89142 37014 89172 37066
rect 89172 37014 89198 37066
rect 88902 37012 88958 37014
rect 88982 37012 89038 37014
rect 89062 37012 89118 37014
rect 89142 37012 89198 37014
rect 88902 35978 88958 35980
rect 88982 35978 89038 35980
rect 89062 35978 89118 35980
rect 89142 35978 89198 35980
rect 88902 35926 88928 35978
rect 88928 35926 88958 35978
rect 88982 35926 88992 35978
rect 88992 35926 89038 35978
rect 89062 35926 89108 35978
rect 89108 35926 89118 35978
rect 89142 35926 89172 35978
rect 89172 35926 89198 35978
rect 88902 35924 88958 35926
rect 88982 35924 89038 35926
rect 89062 35924 89118 35926
rect 89142 35924 89198 35926
rect 86238 35434 86294 35436
rect 86318 35434 86374 35436
rect 86398 35434 86454 35436
rect 86478 35434 86534 35436
rect 86238 35382 86264 35434
rect 86264 35382 86294 35434
rect 86318 35382 86328 35434
rect 86328 35382 86374 35434
rect 86398 35382 86444 35434
rect 86444 35382 86454 35434
rect 86478 35382 86508 35434
rect 86508 35382 86534 35434
rect 86238 35380 86294 35382
rect 86318 35380 86374 35382
rect 86398 35380 86454 35382
rect 86478 35380 86534 35382
rect 86238 34346 86294 34348
rect 86318 34346 86374 34348
rect 86398 34346 86454 34348
rect 86478 34346 86534 34348
rect 86238 34294 86264 34346
rect 86264 34294 86294 34346
rect 86318 34294 86328 34346
rect 86328 34294 86374 34346
rect 86398 34294 86444 34346
rect 86444 34294 86454 34346
rect 86478 34294 86508 34346
rect 86508 34294 86534 34346
rect 86238 34292 86294 34294
rect 86318 34292 86374 34294
rect 86398 34292 86454 34294
rect 86478 34292 86534 34294
rect 84368 33408 84424 33464
rect 86024 33444 86026 33464
rect 86026 33444 86078 33464
rect 86078 33444 86080 33464
rect 86024 33408 86080 33444
rect 83574 32714 83630 32716
rect 83654 32714 83710 32716
rect 83734 32714 83790 32716
rect 83814 32714 83870 32716
rect 83574 32662 83600 32714
rect 83600 32662 83630 32714
rect 83654 32662 83664 32714
rect 83664 32662 83710 32714
rect 83734 32662 83780 32714
rect 83780 32662 83790 32714
rect 83814 32662 83844 32714
rect 83844 32662 83870 32714
rect 83574 32660 83630 32662
rect 83654 32660 83710 32662
rect 83734 32660 83790 32662
rect 83814 32660 83870 32662
rect 83574 31626 83630 31628
rect 83654 31626 83710 31628
rect 83734 31626 83790 31628
rect 83814 31626 83870 31628
rect 83574 31574 83600 31626
rect 83600 31574 83630 31626
rect 83654 31574 83664 31626
rect 83664 31574 83710 31626
rect 83734 31574 83780 31626
rect 83780 31574 83790 31626
rect 83814 31574 83844 31626
rect 83844 31574 83870 31626
rect 83574 31572 83630 31574
rect 83654 31572 83710 31574
rect 83734 31572 83790 31574
rect 83814 31572 83870 31574
rect 80320 30824 80376 30880
rect 78246 27274 78302 27276
rect 78326 27274 78382 27276
rect 78406 27274 78462 27276
rect 78486 27274 78542 27276
rect 78246 27222 78272 27274
rect 78272 27222 78302 27274
rect 78326 27222 78336 27274
rect 78336 27222 78382 27274
rect 78406 27222 78452 27274
rect 78452 27222 78462 27274
rect 78486 27222 78516 27274
rect 78516 27222 78542 27274
rect 78246 27220 78302 27222
rect 78326 27220 78382 27222
rect 78406 27220 78462 27222
rect 78486 27220 78542 27222
rect 80910 31082 80966 31084
rect 80990 31082 81046 31084
rect 81070 31082 81126 31084
rect 81150 31082 81206 31084
rect 80910 31030 80936 31082
rect 80936 31030 80966 31082
rect 80990 31030 81000 31082
rect 81000 31030 81046 31082
rect 81070 31030 81116 31082
rect 81116 31030 81126 31082
rect 81150 31030 81180 31082
rect 81180 31030 81206 31082
rect 80910 31028 80966 31030
rect 80990 31028 81046 31030
rect 81070 31028 81126 31030
rect 81150 31028 81206 31030
rect 80964 30844 81020 30880
rect 80964 30824 80966 30844
rect 80966 30824 81018 30844
rect 81018 30824 81020 30844
rect 83574 30538 83630 30540
rect 83654 30538 83710 30540
rect 83734 30538 83790 30540
rect 83814 30538 83870 30540
rect 83574 30486 83600 30538
rect 83600 30486 83630 30538
rect 83654 30486 83664 30538
rect 83664 30486 83710 30538
rect 83734 30486 83780 30538
rect 83780 30486 83790 30538
rect 83814 30486 83844 30538
rect 83844 30486 83870 30538
rect 83574 30484 83630 30486
rect 83654 30484 83710 30486
rect 83734 30484 83790 30486
rect 83814 30484 83870 30486
rect 80910 29994 80966 29996
rect 80990 29994 81046 29996
rect 81070 29994 81126 29996
rect 81150 29994 81206 29996
rect 80910 29942 80936 29994
rect 80936 29942 80966 29994
rect 80990 29942 81000 29994
rect 81000 29942 81046 29994
rect 81070 29942 81116 29994
rect 81116 29942 81126 29994
rect 81150 29942 81180 29994
rect 81180 29942 81206 29994
rect 80910 29940 80966 29942
rect 80990 29940 81046 29942
rect 81070 29940 81126 29942
rect 81150 29940 81206 29942
rect 86238 33258 86294 33260
rect 86318 33258 86374 33260
rect 86398 33258 86454 33260
rect 86478 33258 86534 33260
rect 86238 33206 86264 33258
rect 86264 33206 86294 33258
rect 86318 33206 86328 33258
rect 86328 33206 86374 33258
rect 86398 33206 86444 33258
rect 86444 33206 86454 33258
rect 86478 33206 86508 33258
rect 86508 33206 86534 33258
rect 86238 33204 86294 33206
rect 86318 33204 86374 33206
rect 86398 33204 86454 33206
rect 86478 33204 86534 33206
rect 88902 34890 88958 34892
rect 88982 34890 89038 34892
rect 89062 34890 89118 34892
rect 89142 34890 89198 34892
rect 88902 34838 88928 34890
rect 88928 34838 88958 34890
rect 88982 34838 88992 34890
rect 88992 34838 89038 34890
rect 89062 34838 89108 34890
rect 89108 34838 89118 34890
rect 89142 34838 89172 34890
rect 89172 34838 89198 34890
rect 88902 34836 88958 34838
rect 88982 34836 89038 34838
rect 89062 34836 89118 34838
rect 89142 34836 89198 34838
rect 86238 32170 86294 32172
rect 86318 32170 86374 32172
rect 86398 32170 86454 32172
rect 86478 32170 86534 32172
rect 86238 32118 86264 32170
rect 86264 32118 86294 32170
rect 86318 32118 86328 32170
rect 86328 32118 86374 32170
rect 86398 32118 86444 32170
rect 86444 32118 86454 32170
rect 86478 32118 86508 32170
rect 86508 32118 86534 32170
rect 86238 32116 86294 32118
rect 86318 32116 86374 32118
rect 86398 32116 86454 32118
rect 86478 32116 86534 32118
rect 86238 31082 86294 31084
rect 86318 31082 86374 31084
rect 86398 31082 86454 31084
rect 86478 31082 86534 31084
rect 86238 31030 86264 31082
rect 86264 31030 86294 31082
rect 86318 31030 86328 31082
rect 86328 31030 86374 31082
rect 86398 31030 86444 31082
rect 86444 31030 86454 31082
rect 86478 31030 86508 31082
rect 86508 31030 86534 31082
rect 86238 31028 86294 31030
rect 86318 31028 86374 31030
rect 86398 31028 86454 31030
rect 86478 31028 86534 31030
rect 80910 28906 80966 28908
rect 80990 28906 81046 28908
rect 81070 28906 81126 28908
rect 81150 28906 81206 28908
rect 80910 28854 80936 28906
rect 80936 28854 80966 28906
rect 80990 28854 81000 28906
rect 81000 28854 81046 28906
rect 81070 28854 81116 28906
rect 81116 28854 81126 28906
rect 81150 28854 81180 28906
rect 81180 28854 81206 28906
rect 80910 28852 80966 28854
rect 80990 28852 81046 28854
rect 81070 28852 81126 28854
rect 81150 28852 81206 28854
rect 80910 27818 80966 27820
rect 80990 27818 81046 27820
rect 81070 27818 81126 27820
rect 81150 27818 81206 27820
rect 80910 27766 80936 27818
rect 80936 27766 80966 27818
rect 80990 27766 81000 27818
rect 81000 27766 81046 27818
rect 81070 27766 81116 27818
rect 81116 27766 81126 27818
rect 81150 27766 81180 27818
rect 81180 27766 81206 27818
rect 80910 27764 80966 27766
rect 80990 27764 81046 27766
rect 81070 27764 81126 27766
rect 81150 27764 81206 27766
rect 83574 29450 83630 29452
rect 83654 29450 83710 29452
rect 83734 29450 83790 29452
rect 83814 29450 83870 29452
rect 83574 29398 83600 29450
rect 83600 29398 83630 29450
rect 83654 29398 83664 29450
rect 83664 29398 83710 29450
rect 83734 29398 83780 29450
rect 83780 29398 83790 29450
rect 83814 29398 83844 29450
rect 83844 29398 83870 29450
rect 83574 29396 83630 29398
rect 83654 29396 83710 29398
rect 83734 29396 83790 29398
rect 83814 29396 83870 29398
rect 83574 28362 83630 28364
rect 83654 28362 83710 28364
rect 83734 28362 83790 28364
rect 83814 28362 83870 28364
rect 83574 28310 83600 28362
rect 83600 28310 83630 28362
rect 83654 28310 83664 28362
rect 83664 28310 83710 28362
rect 83734 28310 83780 28362
rect 83780 28310 83790 28362
rect 83814 28310 83844 28362
rect 83844 28310 83870 28362
rect 83574 28308 83630 28310
rect 83654 28308 83710 28310
rect 83734 28308 83790 28310
rect 83814 28308 83870 28310
rect 86238 29994 86294 29996
rect 86318 29994 86374 29996
rect 86398 29994 86454 29996
rect 86478 29994 86534 29996
rect 86238 29942 86264 29994
rect 86264 29942 86294 29994
rect 86318 29942 86328 29994
rect 86328 29942 86374 29994
rect 86398 29942 86444 29994
rect 86444 29942 86454 29994
rect 86478 29942 86508 29994
rect 86508 29942 86534 29994
rect 86238 29940 86294 29942
rect 86318 29940 86374 29942
rect 86398 29940 86454 29942
rect 86478 29940 86534 29942
rect 88902 33802 88958 33804
rect 88982 33802 89038 33804
rect 89062 33802 89118 33804
rect 89142 33802 89198 33804
rect 88902 33750 88928 33802
rect 88928 33750 88958 33802
rect 88982 33750 88992 33802
rect 88992 33750 89038 33802
rect 89062 33750 89108 33802
rect 89108 33750 89118 33802
rect 89142 33750 89172 33802
rect 89172 33750 89198 33802
rect 88902 33748 88958 33750
rect 88982 33748 89038 33750
rect 89062 33748 89118 33750
rect 89142 33748 89198 33750
rect 88902 32714 88958 32716
rect 88982 32714 89038 32716
rect 89062 32714 89118 32716
rect 89142 32714 89198 32716
rect 88902 32662 88928 32714
rect 88928 32662 88958 32714
rect 88982 32662 88992 32714
rect 88992 32662 89038 32714
rect 89062 32662 89108 32714
rect 89108 32662 89118 32714
rect 89142 32662 89172 32714
rect 89172 32662 89198 32714
rect 88902 32660 88958 32662
rect 88982 32660 89038 32662
rect 89062 32660 89118 32662
rect 89142 32660 89198 32662
rect 88902 31626 88958 31628
rect 88982 31626 89038 31628
rect 89062 31626 89118 31628
rect 89142 31626 89198 31628
rect 88902 31574 88928 31626
rect 88928 31574 88958 31626
rect 88982 31574 88992 31626
rect 88992 31574 89038 31626
rect 89062 31574 89108 31626
rect 89108 31574 89118 31626
rect 89142 31574 89172 31626
rect 89172 31574 89198 31626
rect 88902 31572 88958 31574
rect 88982 31572 89038 31574
rect 89062 31572 89118 31574
rect 89142 31572 89198 31574
rect 86238 28906 86294 28908
rect 86318 28906 86374 28908
rect 86398 28906 86454 28908
rect 86478 28906 86534 28908
rect 86238 28854 86264 28906
rect 86264 28854 86294 28906
rect 86318 28854 86328 28906
rect 86328 28854 86374 28906
rect 86398 28854 86444 28906
rect 86444 28854 86454 28906
rect 86478 28854 86508 28906
rect 86508 28854 86534 28906
rect 86238 28852 86294 28854
rect 86318 28852 86374 28854
rect 86398 28852 86454 28854
rect 86478 28852 86534 28854
rect 83574 27274 83630 27276
rect 83654 27274 83710 27276
rect 83734 27274 83790 27276
rect 83814 27274 83870 27276
rect 83574 27222 83600 27274
rect 83600 27222 83630 27274
rect 83654 27222 83664 27274
rect 83664 27222 83710 27274
rect 83734 27222 83780 27274
rect 83780 27222 83790 27274
rect 83814 27222 83844 27274
rect 83844 27222 83870 27274
rect 83574 27220 83630 27222
rect 83654 27220 83710 27222
rect 83734 27220 83790 27222
rect 83814 27220 83870 27222
rect 88902 30538 88958 30540
rect 88982 30538 89038 30540
rect 89062 30538 89118 30540
rect 89142 30538 89198 30540
rect 88902 30486 88928 30538
rect 88928 30486 88958 30538
rect 88982 30486 88992 30538
rect 88992 30486 89038 30538
rect 89062 30486 89108 30538
rect 89108 30486 89118 30538
rect 89142 30486 89172 30538
rect 89172 30486 89198 30538
rect 88902 30484 88958 30486
rect 88982 30484 89038 30486
rect 89062 30484 89118 30486
rect 89142 30484 89198 30486
rect 88902 29450 88958 29452
rect 88982 29450 89038 29452
rect 89062 29450 89118 29452
rect 89142 29450 89198 29452
rect 88902 29398 88928 29450
rect 88928 29398 88958 29450
rect 88982 29398 88992 29450
rect 88992 29398 89038 29450
rect 89062 29398 89108 29450
rect 89108 29398 89118 29450
rect 89142 29398 89172 29450
rect 89172 29398 89198 29450
rect 88902 29396 88958 29398
rect 88982 29396 89038 29398
rect 89062 29396 89118 29398
rect 89142 29396 89198 29398
rect 88902 28362 88958 28364
rect 88982 28362 89038 28364
rect 89062 28362 89118 28364
rect 89142 28362 89198 28364
rect 88902 28310 88928 28362
rect 88928 28310 88958 28362
rect 88982 28310 88992 28362
rect 88992 28310 89038 28362
rect 89062 28310 89108 28362
rect 89108 28310 89118 28362
rect 89142 28310 89172 28362
rect 89172 28310 89198 28362
rect 88902 28308 88958 28310
rect 88982 28308 89038 28310
rect 89062 28308 89118 28310
rect 89142 28308 89198 28310
rect 86238 27818 86294 27820
rect 86318 27818 86374 27820
rect 86398 27818 86454 27820
rect 86478 27818 86534 27820
rect 86238 27766 86264 27818
rect 86264 27766 86294 27818
rect 86318 27766 86328 27818
rect 86328 27766 86374 27818
rect 86398 27766 86444 27818
rect 86444 27766 86454 27818
rect 86478 27766 86508 27818
rect 86508 27766 86534 27818
rect 86238 27764 86294 27766
rect 86318 27764 86374 27766
rect 86398 27764 86454 27766
rect 86478 27764 86534 27766
rect 88902 27274 88958 27276
rect 88982 27274 89038 27276
rect 89062 27274 89118 27276
rect 89142 27274 89198 27276
rect 88902 27222 88928 27274
rect 88928 27222 88958 27274
rect 88982 27222 88992 27274
rect 88992 27222 89038 27274
rect 89062 27222 89108 27274
rect 89108 27222 89118 27274
rect 89142 27222 89172 27274
rect 89172 27222 89198 27274
rect 88902 27220 88958 27222
rect 88982 27220 89038 27222
rect 89062 27220 89118 27222
rect 89142 27220 89198 27222
rect 91566 41962 91622 41964
rect 91646 41962 91702 41964
rect 91726 41962 91782 41964
rect 91806 41962 91862 41964
rect 91566 41910 91592 41962
rect 91592 41910 91622 41962
rect 91646 41910 91656 41962
rect 91656 41910 91702 41962
rect 91726 41910 91772 41962
rect 91772 41910 91782 41962
rect 91806 41910 91836 41962
rect 91836 41910 91862 41962
rect 91566 41908 91622 41910
rect 91646 41908 91702 41910
rect 91726 41908 91782 41910
rect 91806 41908 91862 41910
rect 91566 40874 91622 40876
rect 91646 40874 91702 40876
rect 91726 40874 91782 40876
rect 91806 40874 91862 40876
rect 91566 40822 91592 40874
rect 91592 40822 91622 40874
rect 91646 40822 91656 40874
rect 91656 40822 91702 40874
rect 91726 40822 91772 40874
rect 91772 40822 91782 40874
rect 91806 40822 91836 40874
rect 91836 40822 91862 40874
rect 91566 40820 91622 40822
rect 91646 40820 91702 40822
rect 91726 40820 91782 40822
rect 91806 40820 91862 40822
rect 91566 39786 91622 39788
rect 91646 39786 91702 39788
rect 91726 39786 91782 39788
rect 91806 39786 91862 39788
rect 91566 39734 91592 39786
rect 91592 39734 91622 39786
rect 91646 39734 91656 39786
rect 91656 39734 91702 39786
rect 91726 39734 91772 39786
rect 91772 39734 91782 39786
rect 91806 39734 91836 39786
rect 91836 39734 91862 39786
rect 91566 39732 91622 39734
rect 91646 39732 91702 39734
rect 91726 39732 91782 39734
rect 91806 39732 91862 39734
rect 91566 38698 91622 38700
rect 91646 38698 91702 38700
rect 91726 38698 91782 38700
rect 91806 38698 91862 38700
rect 91566 38646 91592 38698
rect 91592 38646 91622 38698
rect 91646 38646 91656 38698
rect 91656 38646 91702 38698
rect 91726 38646 91772 38698
rect 91772 38646 91782 38698
rect 91806 38646 91836 38698
rect 91836 38646 91862 38698
rect 91566 38644 91622 38646
rect 91646 38644 91702 38646
rect 91726 38644 91782 38646
rect 91806 38644 91862 38646
rect 91566 37610 91622 37612
rect 91646 37610 91702 37612
rect 91726 37610 91782 37612
rect 91806 37610 91862 37612
rect 91566 37558 91592 37610
rect 91592 37558 91622 37610
rect 91646 37558 91656 37610
rect 91656 37558 91702 37610
rect 91726 37558 91772 37610
rect 91772 37558 91782 37610
rect 91806 37558 91836 37610
rect 91836 37558 91862 37610
rect 91566 37556 91622 37558
rect 91646 37556 91702 37558
rect 91726 37556 91782 37558
rect 91806 37556 91862 37558
rect 91566 36522 91622 36524
rect 91646 36522 91702 36524
rect 91726 36522 91782 36524
rect 91806 36522 91862 36524
rect 91566 36470 91592 36522
rect 91592 36470 91622 36522
rect 91646 36470 91656 36522
rect 91656 36470 91702 36522
rect 91726 36470 91772 36522
rect 91772 36470 91782 36522
rect 91806 36470 91836 36522
rect 91836 36470 91862 36522
rect 91566 36468 91622 36470
rect 91646 36468 91702 36470
rect 91726 36468 91782 36470
rect 91806 36468 91862 36470
rect 91566 35434 91622 35436
rect 91646 35434 91702 35436
rect 91726 35434 91782 35436
rect 91806 35434 91862 35436
rect 91566 35382 91592 35434
rect 91592 35382 91622 35434
rect 91646 35382 91656 35434
rect 91656 35382 91702 35434
rect 91726 35382 91772 35434
rect 91772 35382 91782 35434
rect 91806 35382 91836 35434
rect 91836 35382 91862 35434
rect 91566 35380 91622 35382
rect 91646 35380 91702 35382
rect 91726 35380 91782 35382
rect 91806 35380 91862 35382
rect 91268 35176 91324 35232
rect 91566 34346 91622 34348
rect 91646 34346 91702 34348
rect 91726 34346 91782 34348
rect 91806 34346 91862 34348
rect 91566 34294 91592 34346
rect 91592 34294 91622 34346
rect 91646 34294 91656 34346
rect 91656 34294 91702 34346
rect 91726 34294 91772 34346
rect 91772 34294 91782 34346
rect 91806 34294 91836 34346
rect 91836 34294 91862 34346
rect 91566 34292 91622 34294
rect 91646 34292 91702 34294
rect 91726 34292 91782 34294
rect 91806 34292 91862 34294
rect 91360 33544 91416 33600
rect 91566 33258 91622 33260
rect 91646 33258 91702 33260
rect 91726 33258 91782 33260
rect 91806 33258 91862 33260
rect 91566 33206 91592 33258
rect 91592 33206 91622 33258
rect 91646 33206 91656 33258
rect 91656 33206 91702 33258
rect 91726 33206 91772 33258
rect 91772 33206 91782 33258
rect 91806 33206 91836 33258
rect 91836 33206 91862 33258
rect 91566 33204 91622 33206
rect 91646 33204 91702 33206
rect 91726 33204 91782 33206
rect 91806 33204 91862 33206
rect 91084 32592 91140 32648
rect 91566 32170 91622 32172
rect 91646 32170 91702 32172
rect 91726 32170 91782 32172
rect 91806 32170 91862 32172
rect 91566 32118 91592 32170
rect 91592 32118 91622 32170
rect 91646 32118 91656 32170
rect 91656 32118 91702 32170
rect 91726 32118 91772 32170
rect 91772 32118 91782 32170
rect 91806 32118 91836 32170
rect 91836 32118 91862 32170
rect 91566 32116 91622 32118
rect 91646 32116 91702 32118
rect 91726 32116 91782 32118
rect 91806 32116 91862 32118
rect 91566 31082 91622 31084
rect 91646 31082 91702 31084
rect 91726 31082 91782 31084
rect 91806 31082 91862 31084
rect 91566 31030 91592 31082
rect 91592 31030 91622 31082
rect 91646 31030 91656 31082
rect 91656 31030 91702 31082
rect 91726 31030 91772 31082
rect 91772 31030 91782 31082
rect 91806 31030 91836 31082
rect 91836 31030 91862 31082
rect 91566 31028 91622 31030
rect 91646 31028 91702 31030
rect 91726 31028 91782 31030
rect 91806 31028 91862 31030
rect 91566 29994 91622 29996
rect 91646 29994 91702 29996
rect 91726 29994 91782 29996
rect 91806 29994 91862 29996
rect 91566 29942 91592 29994
rect 91592 29942 91622 29994
rect 91646 29942 91656 29994
rect 91656 29942 91702 29994
rect 91726 29942 91772 29994
rect 91772 29942 91782 29994
rect 91806 29942 91836 29994
rect 91836 29942 91862 29994
rect 91566 29940 91622 29942
rect 91646 29940 91702 29942
rect 91726 29940 91782 29942
rect 91806 29940 91862 29942
rect 91566 28906 91622 28908
rect 91646 28906 91702 28908
rect 91726 28906 91782 28908
rect 91806 28906 91862 28908
rect 91566 28854 91592 28906
rect 91592 28854 91622 28906
rect 91646 28854 91656 28906
rect 91656 28854 91702 28906
rect 91726 28854 91772 28906
rect 91772 28854 91782 28906
rect 91806 28854 91836 28906
rect 91836 28854 91862 28906
rect 91566 28852 91622 28854
rect 91646 28852 91702 28854
rect 91726 28852 91782 28854
rect 91806 28852 91862 28854
rect 91566 27818 91622 27820
rect 91646 27818 91702 27820
rect 91726 27818 91782 27820
rect 91806 27818 91862 27820
rect 91566 27766 91592 27818
rect 91592 27766 91622 27818
rect 91646 27766 91656 27818
rect 91656 27766 91702 27818
rect 91726 27766 91772 27818
rect 91772 27766 91782 27818
rect 91806 27766 91836 27818
rect 91836 27766 91862 27818
rect 91566 27764 91622 27766
rect 91646 27764 91702 27766
rect 91726 27764 91782 27766
rect 91806 27764 91862 27766
rect 70254 26730 70310 26732
rect 70334 26730 70390 26732
rect 70414 26730 70470 26732
rect 70494 26730 70550 26732
rect 70254 26678 70280 26730
rect 70280 26678 70310 26730
rect 70334 26678 70344 26730
rect 70344 26678 70390 26730
rect 70414 26678 70460 26730
rect 70460 26678 70470 26730
rect 70494 26678 70524 26730
rect 70524 26678 70550 26730
rect 70254 26676 70310 26678
rect 70334 26676 70390 26678
rect 70414 26676 70470 26678
rect 70494 26676 70550 26678
rect 70016 22936 70072 22992
rect 70200 22460 70256 22516
rect 70384 18448 70440 18504
rect 70476 17020 70532 17076
rect 75582 26730 75638 26732
rect 75662 26730 75718 26732
rect 75742 26730 75798 26732
rect 75822 26730 75878 26732
rect 75582 26678 75608 26730
rect 75608 26678 75638 26730
rect 75662 26678 75672 26730
rect 75672 26678 75718 26730
rect 75742 26678 75788 26730
rect 75788 26678 75798 26730
rect 75822 26678 75852 26730
rect 75852 26678 75878 26730
rect 75582 26676 75638 26678
rect 75662 26676 75718 26678
rect 75742 26676 75798 26678
rect 75822 26676 75878 26678
rect 80910 26730 80966 26732
rect 80990 26730 81046 26732
rect 81070 26730 81126 26732
rect 81150 26730 81206 26732
rect 80910 26678 80936 26730
rect 80936 26678 80966 26730
rect 80990 26678 81000 26730
rect 81000 26678 81046 26730
rect 81070 26678 81116 26730
rect 81116 26678 81126 26730
rect 81150 26678 81180 26730
rect 81180 26678 81206 26730
rect 80910 26676 80966 26678
rect 80990 26676 81046 26678
rect 81070 26676 81126 26678
rect 81150 26676 81206 26678
rect 86238 26730 86294 26732
rect 86318 26730 86374 26732
rect 86398 26730 86454 26732
rect 86478 26730 86534 26732
rect 86238 26678 86264 26730
rect 86264 26678 86294 26730
rect 86318 26678 86328 26730
rect 86328 26678 86374 26730
rect 86398 26678 86444 26730
rect 86444 26678 86454 26730
rect 86478 26678 86508 26730
rect 86508 26678 86534 26730
rect 86238 26676 86294 26678
rect 86318 26676 86374 26678
rect 86398 26676 86454 26678
rect 86478 26676 86534 26678
rect 70476 14844 70532 14900
rect 91566 26730 91622 26732
rect 91646 26730 91702 26732
rect 91726 26730 91782 26732
rect 91806 26730 91862 26732
rect 91566 26678 91592 26730
rect 91592 26678 91622 26730
rect 91646 26678 91656 26730
rect 91656 26678 91702 26730
rect 91726 26678 91772 26730
rect 91772 26678 91782 26730
rect 91806 26678 91836 26730
rect 91836 26678 91862 26730
rect 91566 26676 91622 26678
rect 91646 26676 91702 26678
rect 91726 26676 91782 26678
rect 91806 26676 91862 26678
rect 91176 9472 91232 9528
rect 31376 2300 31378 2320
rect 31378 2300 31430 2320
rect 31430 2300 31432 2320
rect 31376 2264 31432 2300
rect 35622 2250 35678 2252
rect 35702 2250 35758 2252
rect 35782 2250 35838 2252
rect 35862 2250 35918 2252
rect 35622 2198 35648 2250
rect 35648 2198 35678 2250
rect 35702 2198 35712 2250
rect 35712 2198 35758 2250
rect 35782 2198 35828 2250
rect 35828 2198 35838 2250
rect 35862 2198 35892 2250
rect 35892 2198 35918 2250
rect 35622 2196 35678 2198
rect 35702 2196 35758 2198
rect 35782 2196 35838 2198
rect 35862 2196 35918 2198
rect 43244 2264 43300 2320
rect 69740 2264 69796 2320
rect 40950 2250 41006 2252
rect 41030 2250 41086 2252
rect 41110 2250 41166 2252
rect 41190 2250 41246 2252
rect 40950 2198 40976 2250
rect 40976 2198 41006 2250
rect 41030 2198 41040 2250
rect 41040 2198 41086 2250
rect 41110 2198 41156 2250
rect 41156 2198 41166 2250
rect 41190 2198 41220 2250
rect 41220 2198 41246 2250
rect 40950 2196 41006 2198
rect 41030 2196 41086 2198
rect 41110 2196 41166 2198
rect 41190 2196 41246 2198
rect 6318 1706 6374 1708
rect 6398 1706 6454 1708
rect 6478 1706 6534 1708
rect 6558 1706 6614 1708
rect 6318 1654 6344 1706
rect 6344 1654 6374 1706
rect 6398 1654 6408 1706
rect 6408 1654 6454 1706
rect 6478 1654 6524 1706
rect 6524 1654 6534 1706
rect 6558 1654 6588 1706
rect 6588 1654 6614 1706
rect 6318 1652 6374 1654
rect 6398 1652 6454 1654
rect 6478 1652 6534 1654
rect 6558 1652 6614 1654
rect 38286 1706 38342 1708
rect 38366 1706 38422 1708
rect 38446 1706 38502 1708
rect 38526 1706 38582 1708
rect 38286 1654 38312 1706
rect 38312 1654 38342 1706
rect 38366 1654 38376 1706
rect 38376 1654 38422 1706
rect 38446 1654 38492 1706
rect 38492 1654 38502 1706
rect 38526 1654 38556 1706
rect 38556 1654 38582 1706
rect 38286 1652 38342 1654
rect 38366 1652 38422 1654
rect 38446 1652 38502 1654
rect 38526 1652 38582 1654
rect 3654 1162 3710 1164
rect 3734 1162 3790 1164
rect 3814 1162 3870 1164
rect 3894 1162 3950 1164
rect 3654 1110 3680 1162
rect 3680 1110 3710 1162
rect 3734 1110 3744 1162
rect 3744 1110 3790 1162
rect 3814 1110 3860 1162
rect 3860 1110 3870 1162
rect 3894 1110 3924 1162
rect 3924 1110 3950 1162
rect 3654 1108 3710 1110
rect 3734 1108 3790 1110
rect 3814 1108 3870 1110
rect 3894 1108 3950 1110
rect 35622 1162 35678 1164
rect 35702 1162 35758 1164
rect 35782 1162 35838 1164
rect 35862 1162 35918 1164
rect 35622 1110 35648 1162
rect 35648 1110 35678 1162
rect 35702 1110 35712 1162
rect 35712 1110 35758 1162
rect 35782 1110 35828 1162
rect 35828 1110 35838 1162
rect 35862 1110 35892 1162
rect 35892 1110 35918 1162
rect 35622 1108 35678 1110
rect 35702 1108 35758 1110
rect 35782 1108 35838 1110
rect 35862 1108 35918 1110
rect 40950 1162 41006 1164
rect 41030 1162 41086 1164
rect 41110 1162 41166 1164
rect 41190 1162 41246 1164
rect 40950 1110 40976 1162
rect 40976 1110 41006 1162
rect 41030 1110 41040 1162
rect 41040 1110 41086 1162
rect 41110 1110 41156 1162
rect 41156 1110 41166 1162
rect 41190 1110 41220 1162
rect 41220 1110 41246 1162
rect 40950 1108 41006 1110
rect 41030 1108 41086 1110
rect 41110 1108 41166 1110
rect 41190 1108 41246 1110
rect 6318 618 6374 620
rect 6398 618 6454 620
rect 6478 618 6534 620
rect 6558 618 6614 620
rect 6318 566 6344 618
rect 6344 566 6374 618
rect 6398 566 6408 618
rect 6408 566 6454 618
rect 6478 566 6524 618
rect 6524 566 6534 618
rect 6558 566 6588 618
rect 6588 566 6614 618
rect 6318 564 6374 566
rect 6398 564 6454 566
rect 6478 564 6534 566
rect 6558 564 6614 566
rect 38286 618 38342 620
rect 38366 618 38422 620
rect 38446 618 38502 620
rect 38526 618 38582 620
rect 38286 566 38312 618
rect 38312 566 38342 618
rect 38366 566 38376 618
rect 38376 566 38422 618
rect 38446 566 38492 618
rect 38492 566 38502 618
rect 38526 566 38556 618
rect 38556 566 38582 618
rect 38286 564 38342 566
rect 38366 564 38422 566
rect 38446 564 38502 566
rect 38526 564 38582 566
rect 3654 74 3710 76
rect 3734 74 3790 76
rect 3814 74 3870 76
rect 3894 74 3950 76
rect 3654 22 3680 74
rect 3680 22 3710 74
rect 3734 22 3744 74
rect 3744 22 3790 74
rect 3814 22 3860 74
rect 3860 22 3870 74
rect 3894 22 3924 74
rect 3924 22 3950 74
rect 3654 20 3710 22
rect 3734 20 3790 22
rect 3814 20 3870 22
rect 3894 20 3950 22
rect 35622 74 35678 76
rect 35702 74 35758 76
rect 35782 74 35838 76
rect 35862 74 35918 76
rect 35622 22 35648 74
rect 35648 22 35678 74
rect 35702 22 35712 74
rect 35712 22 35758 74
rect 35782 22 35828 74
rect 35828 22 35838 74
rect 35862 22 35892 74
rect 35892 22 35918 74
rect 35622 20 35678 22
rect 35702 20 35758 22
rect 35782 20 35838 22
rect 35862 20 35918 22
rect 40950 74 41006 76
rect 41030 74 41086 76
rect 41110 74 41166 76
rect 41190 74 41246 76
rect 40950 22 40976 74
rect 40976 22 41006 74
rect 41030 22 41040 74
rect 41040 22 41086 74
rect 41110 22 41156 74
rect 41156 22 41166 74
rect 41190 22 41220 74
rect 41220 22 41246 74
rect 40950 20 41006 22
rect 41030 20 41086 22
rect 41110 20 41166 22
rect 41190 20 41246 22
<< metal3 >>
rect 6306 41968 6626 41969
rect 6306 41904 6314 41968
rect 6378 41904 6394 41968
rect 6458 41904 6474 41968
rect 6538 41904 6554 41968
rect 6618 41904 6626 41968
rect 6306 41903 6626 41904
rect 11634 41968 11954 41969
rect 11634 41904 11642 41968
rect 11706 41904 11722 41968
rect 11786 41904 11802 41968
rect 11866 41904 11882 41968
rect 11946 41904 11954 41968
rect 11634 41903 11954 41904
rect 16962 41968 17282 41969
rect 16962 41904 16970 41968
rect 17034 41904 17050 41968
rect 17114 41904 17130 41968
rect 17194 41904 17210 41968
rect 17274 41904 17282 41968
rect 16962 41903 17282 41904
rect 22290 41968 22610 41969
rect 22290 41904 22298 41968
rect 22362 41904 22378 41968
rect 22442 41904 22458 41968
rect 22522 41904 22538 41968
rect 22602 41904 22610 41968
rect 22290 41903 22610 41904
rect 27618 41968 27938 41969
rect 27618 41904 27626 41968
rect 27690 41904 27706 41968
rect 27770 41904 27786 41968
rect 27850 41904 27866 41968
rect 27930 41904 27938 41968
rect 27618 41903 27938 41904
rect 32946 41968 33266 41969
rect 32946 41904 32954 41968
rect 33018 41904 33034 41968
rect 33098 41904 33114 41968
rect 33178 41904 33194 41968
rect 33258 41904 33266 41968
rect 32946 41903 33266 41904
rect 38274 41968 38594 41969
rect 38274 41904 38282 41968
rect 38346 41904 38362 41968
rect 38426 41904 38442 41968
rect 38506 41904 38522 41968
rect 38586 41904 38594 41968
rect 38274 41903 38594 41904
rect 43602 41968 43922 41969
rect 43602 41904 43610 41968
rect 43674 41904 43690 41968
rect 43754 41904 43770 41968
rect 43834 41904 43850 41968
rect 43914 41904 43922 41968
rect 43602 41903 43922 41904
rect 48930 41968 49250 41969
rect 48930 41904 48938 41968
rect 49002 41904 49018 41968
rect 49082 41904 49098 41968
rect 49162 41904 49178 41968
rect 49242 41904 49250 41968
rect 48930 41903 49250 41904
rect 54258 41968 54578 41969
rect 54258 41904 54266 41968
rect 54330 41904 54346 41968
rect 54410 41904 54426 41968
rect 54490 41904 54506 41968
rect 54570 41904 54578 41968
rect 54258 41903 54578 41904
rect 59586 41968 59906 41969
rect 59586 41904 59594 41968
rect 59658 41904 59674 41968
rect 59738 41904 59754 41968
rect 59818 41904 59834 41968
rect 59898 41904 59906 41968
rect 59586 41903 59906 41904
rect 64914 41968 65234 41969
rect 64914 41904 64922 41968
rect 64986 41904 65002 41968
rect 65066 41904 65082 41968
rect 65146 41904 65162 41968
rect 65226 41904 65234 41968
rect 64914 41903 65234 41904
rect 70242 41968 70562 41969
rect 70242 41904 70250 41968
rect 70314 41904 70330 41968
rect 70394 41904 70410 41968
rect 70474 41904 70490 41968
rect 70554 41904 70562 41968
rect 70242 41903 70562 41904
rect 75570 41968 75890 41969
rect 75570 41904 75578 41968
rect 75642 41904 75658 41968
rect 75722 41904 75738 41968
rect 75802 41904 75818 41968
rect 75882 41904 75890 41968
rect 75570 41903 75890 41904
rect 80898 41968 81218 41969
rect 80898 41904 80906 41968
rect 80970 41904 80986 41968
rect 81050 41904 81066 41968
rect 81130 41904 81146 41968
rect 81210 41904 81218 41968
rect 80898 41903 81218 41904
rect 86226 41968 86546 41969
rect 86226 41904 86234 41968
rect 86298 41904 86314 41968
rect 86378 41904 86394 41968
rect 86458 41904 86474 41968
rect 86538 41904 86546 41968
rect 86226 41903 86546 41904
rect 91554 41968 91874 41969
rect 91554 41904 91562 41968
rect 91626 41904 91642 41968
rect 91706 41904 91722 41968
rect 91786 41904 91802 41968
rect 91866 41904 91874 41968
rect 91554 41903 91874 41904
rect 3642 41424 3962 41425
rect 3642 41360 3650 41424
rect 3714 41360 3730 41424
rect 3794 41360 3810 41424
rect 3874 41360 3890 41424
rect 3954 41360 3962 41424
rect 3642 41359 3962 41360
rect 8970 41424 9290 41425
rect 8970 41360 8978 41424
rect 9042 41360 9058 41424
rect 9122 41360 9138 41424
rect 9202 41360 9218 41424
rect 9282 41360 9290 41424
rect 8970 41359 9290 41360
rect 14298 41424 14618 41425
rect 14298 41360 14306 41424
rect 14370 41360 14386 41424
rect 14450 41360 14466 41424
rect 14530 41360 14546 41424
rect 14610 41360 14618 41424
rect 14298 41359 14618 41360
rect 19626 41424 19946 41425
rect 19626 41360 19634 41424
rect 19698 41360 19714 41424
rect 19778 41360 19794 41424
rect 19858 41360 19874 41424
rect 19938 41360 19946 41424
rect 19626 41359 19946 41360
rect 24954 41424 25274 41425
rect 24954 41360 24962 41424
rect 25026 41360 25042 41424
rect 25106 41360 25122 41424
rect 25186 41360 25202 41424
rect 25266 41360 25274 41424
rect 24954 41359 25274 41360
rect 30282 41424 30602 41425
rect 30282 41360 30290 41424
rect 30354 41360 30370 41424
rect 30434 41360 30450 41424
rect 30514 41360 30530 41424
rect 30594 41360 30602 41424
rect 30282 41359 30602 41360
rect 35610 41424 35930 41425
rect 35610 41360 35618 41424
rect 35682 41360 35698 41424
rect 35762 41360 35778 41424
rect 35842 41360 35858 41424
rect 35922 41360 35930 41424
rect 35610 41359 35930 41360
rect 40938 41424 41258 41425
rect 40938 41360 40946 41424
rect 41010 41360 41026 41424
rect 41090 41360 41106 41424
rect 41170 41360 41186 41424
rect 41250 41360 41258 41424
rect 40938 41359 41258 41360
rect 46266 41424 46586 41425
rect 46266 41360 46274 41424
rect 46338 41360 46354 41424
rect 46418 41360 46434 41424
rect 46498 41360 46514 41424
rect 46578 41360 46586 41424
rect 46266 41359 46586 41360
rect 51594 41424 51914 41425
rect 51594 41360 51602 41424
rect 51666 41360 51682 41424
rect 51746 41360 51762 41424
rect 51826 41360 51842 41424
rect 51906 41360 51914 41424
rect 51594 41359 51914 41360
rect 56922 41424 57242 41425
rect 56922 41360 56930 41424
rect 56994 41360 57010 41424
rect 57074 41360 57090 41424
rect 57154 41360 57170 41424
rect 57234 41360 57242 41424
rect 56922 41359 57242 41360
rect 62250 41424 62570 41425
rect 62250 41360 62258 41424
rect 62322 41360 62338 41424
rect 62402 41360 62418 41424
rect 62482 41360 62498 41424
rect 62562 41360 62570 41424
rect 62250 41359 62570 41360
rect 67578 41424 67898 41425
rect 67578 41360 67586 41424
rect 67650 41360 67666 41424
rect 67730 41360 67746 41424
rect 67810 41360 67826 41424
rect 67890 41360 67898 41424
rect 67578 41359 67898 41360
rect 72906 41424 73226 41425
rect 72906 41360 72914 41424
rect 72978 41360 72994 41424
rect 73058 41360 73074 41424
rect 73138 41360 73154 41424
rect 73218 41360 73226 41424
rect 72906 41359 73226 41360
rect 78234 41424 78554 41425
rect 78234 41360 78242 41424
rect 78306 41360 78322 41424
rect 78386 41360 78402 41424
rect 78466 41360 78482 41424
rect 78546 41360 78554 41424
rect 78234 41359 78554 41360
rect 83562 41424 83882 41425
rect 83562 41360 83570 41424
rect 83634 41360 83650 41424
rect 83714 41360 83730 41424
rect 83794 41360 83810 41424
rect 83874 41360 83882 41424
rect 83562 41359 83882 41360
rect 88890 41424 89210 41425
rect 88890 41360 88898 41424
rect 88962 41360 88978 41424
rect 89042 41360 89058 41424
rect 89122 41360 89138 41424
rect 89202 41360 89210 41424
rect 88890 41359 89210 41360
rect 6306 40880 6626 40881
rect 6306 40816 6314 40880
rect 6378 40816 6394 40880
rect 6458 40816 6474 40880
rect 6538 40816 6554 40880
rect 6618 40816 6626 40880
rect 6306 40815 6626 40816
rect 11634 40880 11954 40881
rect 11634 40816 11642 40880
rect 11706 40816 11722 40880
rect 11786 40816 11802 40880
rect 11866 40816 11882 40880
rect 11946 40816 11954 40880
rect 11634 40815 11954 40816
rect 16962 40880 17282 40881
rect 16962 40816 16970 40880
rect 17034 40816 17050 40880
rect 17114 40816 17130 40880
rect 17194 40816 17210 40880
rect 17274 40816 17282 40880
rect 16962 40815 17282 40816
rect 22290 40880 22610 40881
rect 22290 40816 22298 40880
rect 22362 40816 22378 40880
rect 22442 40816 22458 40880
rect 22522 40816 22538 40880
rect 22602 40816 22610 40880
rect 22290 40815 22610 40816
rect 27618 40880 27938 40881
rect 27618 40816 27626 40880
rect 27690 40816 27706 40880
rect 27770 40816 27786 40880
rect 27850 40816 27866 40880
rect 27930 40816 27938 40880
rect 27618 40815 27938 40816
rect 32946 40880 33266 40881
rect 32946 40816 32954 40880
rect 33018 40816 33034 40880
rect 33098 40816 33114 40880
rect 33178 40816 33194 40880
rect 33258 40816 33266 40880
rect 32946 40815 33266 40816
rect 38274 40880 38594 40881
rect 38274 40816 38282 40880
rect 38346 40816 38362 40880
rect 38426 40816 38442 40880
rect 38506 40816 38522 40880
rect 38586 40816 38594 40880
rect 38274 40815 38594 40816
rect 43602 40880 43922 40881
rect 43602 40816 43610 40880
rect 43674 40816 43690 40880
rect 43754 40816 43770 40880
rect 43834 40816 43850 40880
rect 43914 40816 43922 40880
rect 43602 40815 43922 40816
rect 48930 40880 49250 40881
rect 48930 40816 48938 40880
rect 49002 40816 49018 40880
rect 49082 40816 49098 40880
rect 49162 40816 49178 40880
rect 49242 40816 49250 40880
rect 48930 40815 49250 40816
rect 54258 40880 54578 40881
rect 54258 40816 54266 40880
rect 54330 40816 54346 40880
rect 54410 40816 54426 40880
rect 54490 40816 54506 40880
rect 54570 40816 54578 40880
rect 54258 40815 54578 40816
rect 59586 40880 59906 40881
rect 59586 40816 59594 40880
rect 59658 40816 59674 40880
rect 59738 40816 59754 40880
rect 59818 40816 59834 40880
rect 59898 40816 59906 40880
rect 59586 40815 59906 40816
rect 64914 40880 65234 40881
rect 64914 40816 64922 40880
rect 64986 40816 65002 40880
rect 65066 40816 65082 40880
rect 65146 40816 65162 40880
rect 65226 40816 65234 40880
rect 64914 40815 65234 40816
rect 70242 40880 70562 40881
rect 70242 40816 70250 40880
rect 70314 40816 70330 40880
rect 70394 40816 70410 40880
rect 70474 40816 70490 40880
rect 70554 40816 70562 40880
rect 70242 40815 70562 40816
rect 75570 40880 75890 40881
rect 75570 40816 75578 40880
rect 75642 40816 75658 40880
rect 75722 40816 75738 40880
rect 75802 40816 75818 40880
rect 75882 40816 75890 40880
rect 75570 40815 75890 40816
rect 80898 40880 81218 40881
rect 80898 40816 80906 40880
rect 80970 40816 80986 40880
rect 81050 40816 81066 40880
rect 81130 40816 81146 40880
rect 81210 40816 81218 40880
rect 80898 40815 81218 40816
rect 86226 40880 86546 40881
rect 86226 40816 86234 40880
rect 86298 40816 86314 40880
rect 86378 40816 86394 40880
rect 86458 40816 86474 40880
rect 86538 40816 86546 40880
rect 86226 40815 86546 40816
rect 91554 40880 91874 40881
rect 91554 40816 91562 40880
rect 91626 40816 91642 40880
rect 91706 40816 91722 40880
rect 91786 40816 91802 40880
rect 91866 40816 91874 40880
rect 91554 40815 91874 40816
rect 3642 40336 3962 40337
rect 3642 40272 3650 40336
rect 3714 40272 3730 40336
rect 3794 40272 3810 40336
rect 3874 40272 3890 40336
rect 3954 40272 3962 40336
rect 3642 40271 3962 40272
rect 8970 40336 9290 40337
rect 8970 40272 8978 40336
rect 9042 40272 9058 40336
rect 9122 40272 9138 40336
rect 9202 40272 9218 40336
rect 9282 40272 9290 40336
rect 8970 40271 9290 40272
rect 14298 40336 14618 40337
rect 14298 40272 14306 40336
rect 14370 40272 14386 40336
rect 14450 40272 14466 40336
rect 14530 40272 14546 40336
rect 14610 40272 14618 40336
rect 14298 40271 14618 40272
rect 19626 40336 19946 40337
rect 19626 40272 19634 40336
rect 19698 40272 19714 40336
rect 19778 40272 19794 40336
rect 19858 40272 19874 40336
rect 19938 40272 19946 40336
rect 19626 40271 19946 40272
rect 24954 40336 25274 40337
rect 24954 40272 24962 40336
rect 25026 40272 25042 40336
rect 25106 40272 25122 40336
rect 25186 40272 25202 40336
rect 25266 40272 25274 40336
rect 24954 40271 25274 40272
rect 30282 40336 30602 40337
rect 30282 40272 30290 40336
rect 30354 40272 30370 40336
rect 30434 40272 30450 40336
rect 30514 40272 30530 40336
rect 30594 40272 30602 40336
rect 30282 40271 30602 40272
rect 35610 40336 35930 40337
rect 35610 40272 35618 40336
rect 35682 40272 35698 40336
rect 35762 40272 35778 40336
rect 35842 40272 35858 40336
rect 35922 40272 35930 40336
rect 35610 40271 35930 40272
rect 40938 40336 41258 40337
rect 40938 40272 40946 40336
rect 41010 40272 41026 40336
rect 41090 40272 41106 40336
rect 41170 40272 41186 40336
rect 41250 40272 41258 40336
rect 40938 40271 41258 40272
rect 46266 40336 46586 40337
rect 46266 40272 46274 40336
rect 46338 40272 46354 40336
rect 46418 40272 46434 40336
rect 46498 40272 46514 40336
rect 46578 40272 46586 40336
rect 46266 40271 46586 40272
rect 51594 40336 51914 40337
rect 51594 40272 51602 40336
rect 51666 40272 51682 40336
rect 51746 40272 51762 40336
rect 51826 40272 51842 40336
rect 51906 40272 51914 40336
rect 51594 40271 51914 40272
rect 56922 40336 57242 40337
rect 56922 40272 56930 40336
rect 56994 40272 57010 40336
rect 57074 40272 57090 40336
rect 57154 40272 57170 40336
rect 57234 40272 57242 40336
rect 56922 40271 57242 40272
rect 62250 40336 62570 40337
rect 62250 40272 62258 40336
rect 62322 40272 62338 40336
rect 62402 40272 62418 40336
rect 62482 40272 62498 40336
rect 62562 40272 62570 40336
rect 62250 40271 62570 40272
rect 67578 40336 67898 40337
rect 67578 40272 67586 40336
rect 67650 40272 67666 40336
rect 67730 40272 67746 40336
rect 67810 40272 67826 40336
rect 67890 40272 67898 40336
rect 67578 40271 67898 40272
rect 72906 40336 73226 40337
rect 72906 40272 72914 40336
rect 72978 40272 72994 40336
rect 73058 40272 73074 40336
rect 73138 40272 73154 40336
rect 73218 40272 73226 40336
rect 72906 40271 73226 40272
rect 78234 40336 78554 40337
rect 78234 40272 78242 40336
rect 78306 40272 78322 40336
rect 78386 40272 78402 40336
rect 78466 40272 78482 40336
rect 78546 40272 78554 40336
rect 78234 40271 78554 40272
rect 83562 40336 83882 40337
rect 83562 40272 83570 40336
rect 83634 40272 83650 40336
rect 83714 40272 83730 40336
rect 83794 40272 83810 40336
rect 83874 40272 83882 40336
rect 83562 40271 83882 40272
rect 88890 40336 89210 40337
rect 88890 40272 88898 40336
rect 88962 40272 88978 40336
rect 89042 40272 89058 40336
rect 89122 40272 89138 40336
rect 89202 40272 89210 40336
rect 88890 40271 89210 40272
rect 6306 39792 6626 39793
rect 6306 39728 6314 39792
rect 6378 39728 6394 39792
rect 6458 39728 6474 39792
rect 6538 39728 6554 39792
rect 6618 39728 6626 39792
rect 6306 39727 6626 39728
rect 11634 39792 11954 39793
rect 11634 39728 11642 39792
rect 11706 39728 11722 39792
rect 11786 39728 11802 39792
rect 11866 39728 11882 39792
rect 11946 39728 11954 39792
rect 11634 39727 11954 39728
rect 16962 39792 17282 39793
rect 16962 39728 16970 39792
rect 17034 39728 17050 39792
rect 17114 39728 17130 39792
rect 17194 39728 17210 39792
rect 17274 39728 17282 39792
rect 16962 39727 17282 39728
rect 22290 39792 22610 39793
rect 22290 39728 22298 39792
rect 22362 39728 22378 39792
rect 22442 39728 22458 39792
rect 22522 39728 22538 39792
rect 22602 39728 22610 39792
rect 22290 39727 22610 39728
rect 27618 39792 27938 39793
rect 27618 39728 27626 39792
rect 27690 39728 27706 39792
rect 27770 39728 27786 39792
rect 27850 39728 27866 39792
rect 27930 39728 27938 39792
rect 27618 39727 27938 39728
rect 32946 39792 33266 39793
rect 32946 39728 32954 39792
rect 33018 39728 33034 39792
rect 33098 39728 33114 39792
rect 33178 39728 33194 39792
rect 33258 39728 33266 39792
rect 32946 39727 33266 39728
rect 38274 39792 38594 39793
rect 38274 39728 38282 39792
rect 38346 39728 38362 39792
rect 38426 39728 38442 39792
rect 38506 39728 38522 39792
rect 38586 39728 38594 39792
rect 38274 39727 38594 39728
rect 43602 39792 43922 39793
rect 43602 39728 43610 39792
rect 43674 39728 43690 39792
rect 43754 39728 43770 39792
rect 43834 39728 43850 39792
rect 43914 39728 43922 39792
rect 43602 39727 43922 39728
rect 48930 39792 49250 39793
rect 48930 39728 48938 39792
rect 49002 39728 49018 39792
rect 49082 39728 49098 39792
rect 49162 39728 49178 39792
rect 49242 39728 49250 39792
rect 48930 39727 49250 39728
rect 54258 39792 54578 39793
rect 54258 39728 54266 39792
rect 54330 39728 54346 39792
rect 54410 39728 54426 39792
rect 54490 39728 54506 39792
rect 54570 39728 54578 39792
rect 54258 39727 54578 39728
rect 59586 39792 59906 39793
rect 59586 39728 59594 39792
rect 59658 39728 59674 39792
rect 59738 39728 59754 39792
rect 59818 39728 59834 39792
rect 59898 39728 59906 39792
rect 59586 39727 59906 39728
rect 64914 39792 65234 39793
rect 64914 39728 64922 39792
rect 64986 39728 65002 39792
rect 65066 39728 65082 39792
rect 65146 39728 65162 39792
rect 65226 39728 65234 39792
rect 64914 39727 65234 39728
rect 70242 39792 70562 39793
rect 70242 39728 70250 39792
rect 70314 39728 70330 39792
rect 70394 39728 70410 39792
rect 70474 39728 70490 39792
rect 70554 39728 70562 39792
rect 70242 39727 70562 39728
rect 75570 39792 75890 39793
rect 75570 39728 75578 39792
rect 75642 39728 75658 39792
rect 75722 39728 75738 39792
rect 75802 39728 75818 39792
rect 75882 39728 75890 39792
rect 75570 39727 75890 39728
rect 80898 39792 81218 39793
rect 80898 39728 80906 39792
rect 80970 39728 80986 39792
rect 81050 39728 81066 39792
rect 81130 39728 81146 39792
rect 81210 39728 81218 39792
rect 80898 39727 81218 39728
rect 86226 39792 86546 39793
rect 86226 39728 86234 39792
rect 86298 39728 86314 39792
rect 86378 39728 86394 39792
rect 86458 39728 86474 39792
rect 86538 39728 86546 39792
rect 86226 39727 86546 39728
rect 91554 39792 91874 39793
rect 91554 39728 91562 39792
rect 91626 39728 91642 39792
rect 91706 39728 91722 39792
rect 91786 39728 91802 39792
rect 91866 39728 91874 39792
rect 91554 39727 91874 39728
rect 67803 39586 67869 39589
rect 75439 39586 75505 39589
rect 67803 39584 75505 39586
rect 67803 39528 67808 39584
rect 67864 39528 75444 39584
rect 75500 39528 75505 39584
rect 67803 39526 75505 39528
rect 67803 39523 67869 39526
rect 75439 39523 75505 39526
rect 3642 39248 3962 39249
rect 3642 39184 3650 39248
rect 3714 39184 3730 39248
rect 3794 39184 3810 39248
rect 3874 39184 3890 39248
rect 3954 39184 3962 39248
rect 3642 39183 3962 39184
rect 8970 39248 9290 39249
rect 8970 39184 8978 39248
rect 9042 39184 9058 39248
rect 9122 39184 9138 39248
rect 9202 39184 9218 39248
rect 9282 39184 9290 39248
rect 8970 39183 9290 39184
rect 14298 39248 14618 39249
rect 14298 39184 14306 39248
rect 14370 39184 14386 39248
rect 14450 39184 14466 39248
rect 14530 39184 14546 39248
rect 14610 39184 14618 39248
rect 14298 39183 14618 39184
rect 19626 39248 19946 39249
rect 19626 39184 19634 39248
rect 19698 39184 19714 39248
rect 19778 39184 19794 39248
rect 19858 39184 19874 39248
rect 19938 39184 19946 39248
rect 19626 39183 19946 39184
rect 24954 39248 25274 39249
rect 24954 39184 24962 39248
rect 25026 39184 25042 39248
rect 25106 39184 25122 39248
rect 25186 39184 25202 39248
rect 25266 39184 25274 39248
rect 24954 39183 25274 39184
rect 30282 39248 30602 39249
rect 30282 39184 30290 39248
rect 30354 39184 30370 39248
rect 30434 39184 30450 39248
rect 30514 39184 30530 39248
rect 30594 39184 30602 39248
rect 30282 39183 30602 39184
rect 35610 39248 35930 39249
rect 35610 39184 35618 39248
rect 35682 39184 35698 39248
rect 35762 39184 35778 39248
rect 35842 39184 35858 39248
rect 35922 39184 35930 39248
rect 35610 39183 35930 39184
rect 40938 39248 41258 39249
rect 40938 39184 40946 39248
rect 41010 39184 41026 39248
rect 41090 39184 41106 39248
rect 41170 39184 41186 39248
rect 41250 39184 41258 39248
rect 40938 39183 41258 39184
rect 46266 39248 46586 39249
rect 46266 39184 46274 39248
rect 46338 39184 46354 39248
rect 46418 39184 46434 39248
rect 46498 39184 46514 39248
rect 46578 39184 46586 39248
rect 46266 39183 46586 39184
rect 51594 39248 51914 39249
rect 51594 39184 51602 39248
rect 51666 39184 51682 39248
rect 51746 39184 51762 39248
rect 51826 39184 51842 39248
rect 51906 39184 51914 39248
rect 51594 39183 51914 39184
rect 56922 39248 57242 39249
rect 56922 39184 56930 39248
rect 56994 39184 57010 39248
rect 57074 39184 57090 39248
rect 57154 39184 57170 39248
rect 57234 39184 57242 39248
rect 56922 39183 57242 39184
rect 62250 39248 62570 39249
rect 62250 39184 62258 39248
rect 62322 39184 62338 39248
rect 62402 39184 62418 39248
rect 62482 39184 62498 39248
rect 62562 39184 62570 39248
rect 62250 39183 62570 39184
rect 67578 39248 67898 39249
rect 67578 39184 67586 39248
rect 67650 39184 67666 39248
rect 67730 39184 67746 39248
rect 67810 39184 67826 39248
rect 67890 39184 67898 39248
rect 67578 39183 67898 39184
rect 72906 39248 73226 39249
rect 72906 39184 72914 39248
rect 72978 39184 72994 39248
rect 73058 39184 73074 39248
rect 73138 39184 73154 39248
rect 73218 39184 73226 39248
rect 72906 39183 73226 39184
rect 78234 39248 78554 39249
rect 78234 39184 78242 39248
rect 78306 39184 78322 39248
rect 78386 39184 78402 39248
rect 78466 39184 78482 39248
rect 78546 39184 78554 39248
rect 78234 39183 78554 39184
rect 83562 39248 83882 39249
rect 83562 39184 83570 39248
rect 83634 39184 83650 39248
rect 83714 39184 83730 39248
rect 83794 39184 83810 39248
rect 83874 39184 83882 39248
rect 83562 39183 83882 39184
rect 88890 39248 89210 39249
rect 88890 39184 88898 39248
rect 88962 39184 88978 39248
rect 89042 39184 89058 39248
rect 89122 39184 89138 39248
rect 89202 39184 89210 39248
rect 88890 39183 89210 39184
rect 50323 39042 50389 39045
rect 55475 39042 55541 39045
rect 50323 39040 55541 39042
rect 50323 38984 50328 39040
rect 50384 38984 55480 39040
rect 55536 38984 55541 39040
rect 50323 38982 55541 38984
rect 50323 38979 50389 38982
rect 55475 38979 55541 38982
rect 6306 38704 6626 38705
rect 6306 38640 6314 38704
rect 6378 38640 6394 38704
rect 6458 38640 6474 38704
rect 6538 38640 6554 38704
rect 6618 38640 6626 38704
rect 6306 38639 6626 38640
rect 11634 38704 11954 38705
rect 11634 38640 11642 38704
rect 11706 38640 11722 38704
rect 11786 38640 11802 38704
rect 11866 38640 11882 38704
rect 11946 38640 11954 38704
rect 11634 38639 11954 38640
rect 16962 38704 17282 38705
rect 16962 38640 16970 38704
rect 17034 38640 17050 38704
rect 17114 38640 17130 38704
rect 17194 38640 17210 38704
rect 17274 38640 17282 38704
rect 16962 38639 17282 38640
rect 22290 38704 22610 38705
rect 22290 38640 22298 38704
rect 22362 38640 22378 38704
rect 22442 38640 22458 38704
rect 22522 38640 22538 38704
rect 22602 38640 22610 38704
rect 22290 38639 22610 38640
rect 27618 38704 27938 38705
rect 27618 38640 27626 38704
rect 27690 38640 27706 38704
rect 27770 38640 27786 38704
rect 27850 38640 27866 38704
rect 27930 38640 27938 38704
rect 27618 38639 27938 38640
rect 32946 38704 33266 38705
rect 32946 38640 32954 38704
rect 33018 38640 33034 38704
rect 33098 38640 33114 38704
rect 33178 38640 33194 38704
rect 33258 38640 33266 38704
rect 32946 38639 33266 38640
rect 38274 38704 38594 38705
rect 38274 38640 38282 38704
rect 38346 38640 38362 38704
rect 38426 38640 38442 38704
rect 38506 38640 38522 38704
rect 38586 38640 38594 38704
rect 38274 38639 38594 38640
rect 43602 38704 43922 38705
rect 43602 38640 43610 38704
rect 43674 38640 43690 38704
rect 43754 38640 43770 38704
rect 43834 38640 43850 38704
rect 43914 38640 43922 38704
rect 43602 38639 43922 38640
rect 48930 38704 49250 38705
rect 48930 38640 48938 38704
rect 49002 38640 49018 38704
rect 49082 38640 49098 38704
rect 49162 38640 49178 38704
rect 49242 38640 49250 38704
rect 48930 38639 49250 38640
rect 54258 38704 54578 38705
rect 54258 38640 54266 38704
rect 54330 38640 54346 38704
rect 54410 38640 54426 38704
rect 54490 38640 54506 38704
rect 54570 38640 54578 38704
rect 54258 38639 54578 38640
rect 59586 38704 59906 38705
rect 59586 38640 59594 38704
rect 59658 38640 59674 38704
rect 59738 38640 59754 38704
rect 59818 38640 59834 38704
rect 59898 38640 59906 38704
rect 59586 38639 59906 38640
rect 64914 38704 65234 38705
rect 64914 38640 64922 38704
rect 64986 38640 65002 38704
rect 65066 38640 65082 38704
rect 65146 38640 65162 38704
rect 65226 38640 65234 38704
rect 64914 38639 65234 38640
rect 70242 38704 70562 38705
rect 70242 38640 70250 38704
rect 70314 38640 70330 38704
rect 70394 38640 70410 38704
rect 70474 38640 70490 38704
rect 70554 38640 70562 38704
rect 70242 38639 70562 38640
rect 75570 38704 75890 38705
rect 75570 38640 75578 38704
rect 75642 38640 75658 38704
rect 75722 38640 75738 38704
rect 75802 38640 75818 38704
rect 75882 38640 75890 38704
rect 75570 38639 75890 38640
rect 80898 38704 81218 38705
rect 80898 38640 80906 38704
rect 80970 38640 80986 38704
rect 81050 38640 81066 38704
rect 81130 38640 81146 38704
rect 81210 38640 81218 38704
rect 80898 38639 81218 38640
rect 86226 38704 86546 38705
rect 86226 38640 86234 38704
rect 86298 38640 86314 38704
rect 86378 38640 86394 38704
rect 86458 38640 86474 38704
rect 86538 38640 86546 38704
rect 86226 38639 86546 38640
rect 91554 38704 91874 38705
rect 91554 38640 91562 38704
rect 91626 38640 91642 38704
rect 91706 38640 91722 38704
rect 91786 38640 91802 38704
rect 91866 38640 91874 38704
rect 91554 38639 91874 38640
rect 3642 38160 3962 38161
rect 3642 38096 3650 38160
rect 3714 38096 3730 38160
rect 3794 38096 3810 38160
rect 3874 38096 3890 38160
rect 3954 38096 3962 38160
rect 3642 38095 3962 38096
rect 8970 38160 9290 38161
rect 8970 38096 8978 38160
rect 9042 38096 9058 38160
rect 9122 38096 9138 38160
rect 9202 38096 9218 38160
rect 9282 38096 9290 38160
rect 8970 38095 9290 38096
rect 14298 38160 14618 38161
rect 14298 38096 14306 38160
rect 14370 38096 14386 38160
rect 14450 38096 14466 38160
rect 14530 38096 14546 38160
rect 14610 38096 14618 38160
rect 14298 38095 14618 38096
rect 19626 38160 19946 38161
rect 19626 38096 19634 38160
rect 19698 38096 19714 38160
rect 19778 38096 19794 38160
rect 19858 38096 19874 38160
rect 19938 38096 19946 38160
rect 19626 38095 19946 38096
rect 24954 38160 25274 38161
rect 24954 38096 24962 38160
rect 25026 38096 25042 38160
rect 25106 38096 25122 38160
rect 25186 38096 25202 38160
rect 25266 38096 25274 38160
rect 24954 38095 25274 38096
rect 30282 38160 30602 38161
rect 30282 38096 30290 38160
rect 30354 38096 30370 38160
rect 30434 38096 30450 38160
rect 30514 38096 30530 38160
rect 30594 38096 30602 38160
rect 30282 38095 30602 38096
rect 35610 38160 35930 38161
rect 35610 38096 35618 38160
rect 35682 38096 35698 38160
rect 35762 38096 35778 38160
rect 35842 38096 35858 38160
rect 35922 38096 35930 38160
rect 35610 38095 35930 38096
rect 40938 38160 41258 38161
rect 40938 38096 40946 38160
rect 41010 38096 41026 38160
rect 41090 38096 41106 38160
rect 41170 38096 41186 38160
rect 41250 38096 41258 38160
rect 40938 38095 41258 38096
rect 46266 38160 46586 38161
rect 46266 38096 46274 38160
rect 46338 38096 46354 38160
rect 46418 38096 46434 38160
rect 46498 38096 46514 38160
rect 46578 38096 46586 38160
rect 46266 38095 46586 38096
rect 51594 38160 51914 38161
rect 51594 38096 51602 38160
rect 51666 38096 51682 38160
rect 51746 38096 51762 38160
rect 51826 38096 51842 38160
rect 51906 38096 51914 38160
rect 51594 38095 51914 38096
rect 56922 38160 57242 38161
rect 56922 38096 56930 38160
rect 56994 38096 57010 38160
rect 57074 38096 57090 38160
rect 57154 38096 57170 38160
rect 57234 38096 57242 38160
rect 56922 38095 57242 38096
rect 62250 38160 62570 38161
rect 62250 38096 62258 38160
rect 62322 38096 62338 38160
rect 62402 38096 62418 38160
rect 62482 38096 62498 38160
rect 62562 38096 62570 38160
rect 62250 38095 62570 38096
rect 67578 38160 67898 38161
rect 67578 38096 67586 38160
rect 67650 38096 67666 38160
rect 67730 38096 67746 38160
rect 67810 38096 67826 38160
rect 67890 38096 67898 38160
rect 67578 38095 67898 38096
rect 72906 38160 73226 38161
rect 72906 38096 72914 38160
rect 72978 38096 72994 38160
rect 73058 38096 73074 38160
rect 73138 38096 73154 38160
rect 73218 38096 73226 38160
rect 72906 38095 73226 38096
rect 78234 38160 78554 38161
rect 78234 38096 78242 38160
rect 78306 38096 78322 38160
rect 78386 38096 78402 38160
rect 78466 38096 78482 38160
rect 78546 38096 78554 38160
rect 78234 38095 78554 38096
rect 83562 38160 83882 38161
rect 83562 38096 83570 38160
rect 83634 38096 83650 38160
rect 83714 38096 83730 38160
rect 83794 38096 83810 38160
rect 83874 38096 83882 38160
rect 83562 38095 83882 38096
rect 88890 38160 89210 38161
rect 88890 38096 88898 38160
rect 88962 38096 88978 38160
rect 89042 38096 89058 38160
rect 89122 38096 89138 38160
rect 89202 38096 89210 38160
rect 88890 38095 89210 38096
rect 9107 37954 9173 37957
rect 16375 37954 16441 37957
rect 9107 37952 16441 37954
rect 9107 37896 9112 37952
rect 9168 37896 16380 37952
rect 16436 37896 16441 37952
rect 9107 37894 16441 37896
rect 9107 37891 9173 37894
rect 16375 37891 16441 37894
rect 25575 37818 25641 37821
rect 57867 37818 57933 37821
rect 25575 37816 57933 37818
rect 25575 37760 25580 37816
rect 25636 37760 57872 37816
rect 57928 37760 57933 37816
rect 25575 37758 57933 37760
rect 25575 37755 25641 37758
rect 57867 37755 57933 37758
rect 39283 37682 39349 37685
rect 41767 37682 41833 37685
rect 39283 37680 41833 37682
rect 39283 37624 39288 37680
rect 39344 37624 41772 37680
rect 41828 37624 41833 37680
rect 39283 37622 41833 37624
rect 39283 37619 39349 37622
rect 41767 37619 41833 37622
rect 6306 37616 6626 37617
rect 6306 37552 6314 37616
rect 6378 37552 6394 37616
rect 6458 37552 6474 37616
rect 6538 37552 6554 37616
rect 6618 37552 6626 37616
rect 6306 37551 6626 37552
rect 11634 37616 11954 37617
rect 11634 37552 11642 37616
rect 11706 37552 11722 37616
rect 11786 37552 11802 37616
rect 11866 37552 11882 37616
rect 11946 37552 11954 37616
rect 11634 37551 11954 37552
rect 16962 37616 17282 37617
rect 16962 37552 16970 37616
rect 17034 37552 17050 37616
rect 17114 37552 17130 37616
rect 17194 37552 17210 37616
rect 17274 37552 17282 37616
rect 16962 37551 17282 37552
rect 22290 37616 22610 37617
rect 22290 37552 22298 37616
rect 22362 37552 22378 37616
rect 22442 37552 22458 37616
rect 22522 37552 22538 37616
rect 22602 37552 22610 37616
rect 22290 37551 22610 37552
rect 27618 37616 27938 37617
rect 27618 37552 27626 37616
rect 27690 37552 27706 37616
rect 27770 37552 27786 37616
rect 27850 37552 27866 37616
rect 27930 37552 27938 37616
rect 27618 37551 27938 37552
rect 32946 37616 33266 37617
rect 32946 37552 32954 37616
rect 33018 37552 33034 37616
rect 33098 37552 33114 37616
rect 33178 37552 33194 37616
rect 33258 37552 33266 37616
rect 32946 37551 33266 37552
rect 38274 37616 38594 37617
rect 38274 37552 38282 37616
rect 38346 37552 38362 37616
rect 38426 37552 38442 37616
rect 38506 37552 38522 37616
rect 38586 37552 38594 37616
rect 38274 37551 38594 37552
rect 43602 37616 43922 37617
rect 43602 37552 43610 37616
rect 43674 37552 43690 37616
rect 43754 37552 43770 37616
rect 43834 37552 43850 37616
rect 43914 37552 43922 37616
rect 43602 37551 43922 37552
rect 48930 37616 49250 37617
rect 48930 37552 48938 37616
rect 49002 37552 49018 37616
rect 49082 37552 49098 37616
rect 49162 37552 49178 37616
rect 49242 37552 49250 37616
rect 48930 37551 49250 37552
rect 54258 37616 54578 37617
rect 54258 37552 54266 37616
rect 54330 37552 54346 37616
rect 54410 37552 54426 37616
rect 54490 37552 54506 37616
rect 54570 37552 54578 37616
rect 54258 37551 54578 37552
rect 59586 37616 59906 37617
rect 59586 37552 59594 37616
rect 59658 37552 59674 37616
rect 59738 37552 59754 37616
rect 59818 37552 59834 37616
rect 59898 37552 59906 37616
rect 59586 37551 59906 37552
rect 64914 37616 65234 37617
rect 64914 37552 64922 37616
rect 64986 37552 65002 37616
rect 65066 37552 65082 37616
rect 65146 37552 65162 37616
rect 65226 37552 65234 37616
rect 64914 37551 65234 37552
rect 70242 37616 70562 37617
rect 70242 37552 70250 37616
rect 70314 37552 70330 37616
rect 70394 37552 70410 37616
rect 70474 37552 70490 37616
rect 70554 37552 70562 37616
rect 70242 37551 70562 37552
rect 75570 37616 75890 37617
rect 75570 37552 75578 37616
rect 75642 37552 75658 37616
rect 75722 37552 75738 37616
rect 75802 37552 75818 37616
rect 75882 37552 75890 37616
rect 75570 37551 75890 37552
rect 80898 37616 81218 37617
rect 80898 37552 80906 37616
rect 80970 37552 80986 37616
rect 81050 37552 81066 37616
rect 81130 37552 81146 37616
rect 81210 37552 81218 37616
rect 80898 37551 81218 37552
rect 86226 37616 86546 37617
rect 86226 37552 86234 37616
rect 86298 37552 86314 37616
rect 86378 37552 86394 37616
rect 86458 37552 86474 37616
rect 86538 37552 86546 37616
rect 86226 37551 86546 37552
rect 91554 37616 91874 37617
rect 91554 37552 91562 37616
rect 91626 37552 91642 37616
rect 91706 37552 91722 37616
rect 91786 37552 91802 37616
rect 91866 37552 91874 37616
rect 91554 37551 91874 37552
rect 41215 37410 41281 37413
rect 43607 37410 43673 37413
rect 41215 37408 43673 37410
rect 41215 37352 41220 37408
rect 41276 37352 43612 37408
rect 43668 37352 43673 37408
rect 41215 37350 43673 37352
rect 41215 37347 41281 37350
rect 43607 37347 43673 37350
rect 68171 37410 68237 37413
rect 69275 37410 69341 37413
rect 68171 37408 69341 37410
rect 68171 37352 68176 37408
rect 68232 37352 69280 37408
rect 69336 37352 69341 37408
rect 68171 37350 69341 37352
rect 68171 37347 68237 37350
rect 69275 37347 69341 37350
rect 39099 37274 39165 37277
rect 46919 37274 46985 37277
rect 39099 37272 46985 37274
rect 39099 37216 39104 37272
rect 39160 37216 46924 37272
rect 46980 37216 46985 37272
rect 39099 37214 46985 37216
rect 39099 37211 39165 37214
rect 46919 37211 46985 37214
rect 50415 37274 50481 37277
rect 52531 37274 52597 37277
rect 50415 37272 52597 37274
rect 50415 37216 50420 37272
rect 50476 37216 52536 37272
rect 52592 37216 52597 37272
rect 50415 37214 52597 37216
rect 50415 37211 50481 37214
rect 52531 37211 52597 37214
rect 57959 37274 58025 37277
rect 59615 37274 59681 37277
rect 57959 37272 59681 37274
rect 57959 37216 57964 37272
rect 58020 37216 59620 37272
rect 59676 37216 59681 37272
rect 57959 37214 59681 37216
rect 57959 37211 58025 37214
rect 59615 37211 59681 37214
rect 69183 37274 69249 37277
rect 74151 37274 74217 37277
rect 69183 37272 74217 37274
rect 69183 37216 69188 37272
rect 69244 37216 74156 37272
rect 74212 37216 74217 37272
rect 69183 37214 74217 37216
rect 69183 37211 69249 37214
rect 74151 37211 74217 37214
rect 57775 37138 57841 37141
rect 62099 37138 62165 37141
rect 57775 37136 62165 37138
rect 57775 37080 57780 37136
rect 57836 37080 62104 37136
rect 62160 37080 62165 37136
rect 57775 37078 62165 37080
rect 57775 37075 57841 37078
rect 62099 37075 62165 37078
rect 3642 37072 3962 37073
rect 3642 37008 3650 37072
rect 3714 37008 3730 37072
rect 3794 37008 3810 37072
rect 3874 37008 3890 37072
rect 3954 37008 3962 37072
rect 3642 37007 3962 37008
rect 8970 37072 9290 37073
rect 8970 37008 8978 37072
rect 9042 37008 9058 37072
rect 9122 37008 9138 37072
rect 9202 37008 9218 37072
rect 9282 37008 9290 37072
rect 8970 37007 9290 37008
rect 14298 37072 14618 37073
rect 14298 37008 14306 37072
rect 14370 37008 14386 37072
rect 14450 37008 14466 37072
rect 14530 37008 14546 37072
rect 14610 37008 14618 37072
rect 14298 37007 14618 37008
rect 19626 37072 19946 37073
rect 19626 37008 19634 37072
rect 19698 37008 19714 37072
rect 19778 37008 19794 37072
rect 19858 37008 19874 37072
rect 19938 37008 19946 37072
rect 19626 37007 19946 37008
rect 24954 37072 25274 37073
rect 24954 37008 24962 37072
rect 25026 37008 25042 37072
rect 25106 37008 25122 37072
rect 25186 37008 25202 37072
rect 25266 37008 25274 37072
rect 24954 37007 25274 37008
rect 30282 37072 30602 37073
rect 30282 37008 30290 37072
rect 30354 37008 30370 37072
rect 30434 37008 30450 37072
rect 30514 37008 30530 37072
rect 30594 37008 30602 37072
rect 30282 37007 30602 37008
rect 35610 37072 35930 37073
rect 35610 37008 35618 37072
rect 35682 37008 35698 37072
rect 35762 37008 35778 37072
rect 35842 37008 35858 37072
rect 35922 37008 35930 37072
rect 35610 37007 35930 37008
rect 40938 37072 41258 37073
rect 40938 37008 40946 37072
rect 41010 37008 41026 37072
rect 41090 37008 41106 37072
rect 41170 37008 41186 37072
rect 41250 37008 41258 37072
rect 40938 37007 41258 37008
rect 46266 37072 46586 37073
rect 46266 37008 46274 37072
rect 46338 37008 46354 37072
rect 46418 37008 46434 37072
rect 46498 37008 46514 37072
rect 46578 37008 46586 37072
rect 46266 37007 46586 37008
rect 51594 37072 51914 37073
rect 51594 37008 51602 37072
rect 51666 37008 51682 37072
rect 51746 37008 51762 37072
rect 51826 37008 51842 37072
rect 51906 37008 51914 37072
rect 51594 37007 51914 37008
rect 56922 37072 57242 37073
rect 56922 37008 56930 37072
rect 56994 37008 57010 37072
rect 57074 37008 57090 37072
rect 57154 37008 57170 37072
rect 57234 37008 57242 37072
rect 56922 37007 57242 37008
rect 62250 37072 62570 37073
rect 62250 37008 62258 37072
rect 62322 37008 62338 37072
rect 62402 37008 62418 37072
rect 62482 37008 62498 37072
rect 62562 37008 62570 37072
rect 62250 37007 62570 37008
rect 67578 37072 67898 37073
rect 67578 37008 67586 37072
rect 67650 37008 67666 37072
rect 67730 37008 67746 37072
rect 67810 37008 67826 37072
rect 67890 37008 67898 37072
rect 67578 37007 67898 37008
rect 72906 37072 73226 37073
rect 72906 37008 72914 37072
rect 72978 37008 72994 37072
rect 73058 37008 73074 37072
rect 73138 37008 73154 37072
rect 73218 37008 73226 37072
rect 72906 37007 73226 37008
rect 78234 37072 78554 37073
rect 78234 37008 78242 37072
rect 78306 37008 78322 37072
rect 78386 37008 78402 37072
rect 78466 37008 78482 37072
rect 78546 37008 78554 37072
rect 78234 37007 78554 37008
rect 83562 37072 83882 37073
rect 83562 37008 83570 37072
rect 83634 37008 83650 37072
rect 83714 37008 83730 37072
rect 83794 37008 83810 37072
rect 83874 37008 83882 37072
rect 83562 37007 83882 37008
rect 88890 37072 89210 37073
rect 88890 37008 88898 37072
rect 88962 37008 88978 37072
rect 89042 37008 89058 37072
rect 89122 37008 89138 37072
rect 89202 37008 89210 37072
rect 88890 37007 89210 37008
rect 37535 36866 37601 36869
rect 45447 36866 45513 36869
rect 37535 36864 45513 36866
rect 37535 36808 37540 36864
rect 37596 36808 45452 36864
rect 45508 36808 45513 36864
rect 37535 36806 45513 36808
rect 37535 36803 37601 36806
rect 45447 36803 45513 36806
rect 51795 36866 51861 36869
rect 52347 36866 52413 36869
rect 51795 36864 52413 36866
rect 51795 36808 51800 36864
rect 51856 36808 52352 36864
rect 52408 36808 52413 36864
rect 51795 36806 52413 36808
rect 51795 36803 51861 36806
rect 52347 36803 52413 36806
rect 37719 36730 37785 36733
rect 43699 36730 43765 36733
rect 37719 36728 43765 36730
rect 37719 36672 37724 36728
rect 37780 36672 43704 36728
rect 43760 36672 43765 36728
rect 37719 36670 43765 36672
rect 37719 36667 37785 36670
rect 43699 36667 43765 36670
rect 44251 36730 44317 36733
rect 47655 36730 47721 36733
rect 44251 36728 47721 36730
rect 44251 36672 44256 36728
rect 44312 36672 47660 36728
rect 47716 36672 47721 36728
rect 44251 36670 47721 36672
rect 44251 36667 44317 36670
rect 47655 36667 47721 36670
rect 51427 36730 51493 36733
rect 53451 36730 53517 36733
rect 51427 36728 53517 36730
rect 51427 36672 51432 36728
rect 51488 36672 53456 36728
rect 53512 36672 53517 36728
rect 51427 36670 53517 36672
rect 51427 36667 51493 36670
rect 53451 36667 53517 36670
rect 57683 36730 57749 36733
rect 58419 36730 58485 36733
rect 57683 36728 58485 36730
rect 57683 36672 57688 36728
rect 57744 36672 58424 36728
rect 58480 36672 58485 36728
rect 57683 36670 58485 36672
rect 57683 36667 57749 36670
rect 58419 36667 58485 36670
rect 68907 36730 68973 36733
rect 74243 36730 74309 36733
rect 68907 36728 74309 36730
rect 68907 36672 68912 36728
rect 68968 36672 74248 36728
rect 74304 36672 74309 36728
rect 68907 36670 74309 36672
rect 68907 36667 68973 36670
rect 74243 36667 74309 36670
rect 50415 36594 50481 36597
rect 52715 36594 52781 36597
rect 50415 36592 52781 36594
rect 50415 36536 50420 36592
rect 50476 36536 52720 36592
rect 52776 36536 52781 36592
rect 50415 36534 52781 36536
rect 50415 36531 50481 36534
rect 52715 36531 52781 36534
rect 6306 36528 6626 36529
rect 6306 36464 6314 36528
rect 6378 36464 6394 36528
rect 6458 36464 6474 36528
rect 6538 36464 6554 36528
rect 6618 36464 6626 36528
rect 6306 36463 6626 36464
rect 11634 36528 11954 36529
rect 11634 36464 11642 36528
rect 11706 36464 11722 36528
rect 11786 36464 11802 36528
rect 11866 36464 11882 36528
rect 11946 36464 11954 36528
rect 11634 36463 11954 36464
rect 16962 36528 17282 36529
rect 16962 36464 16970 36528
rect 17034 36464 17050 36528
rect 17114 36464 17130 36528
rect 17194 36464 17210 36528
rect 17274 36464 17282 36528
rect 16962 36463 17282 36464
rect 22290 36528 22610 36529
rect 22290 36464 22298 36528
rect 22362 36464 22378 36528
rect 22442 36464 22458 36528
rect 22522 36464 22538 36528
rect 22602 36464 22610 36528
rect 22290 36463 22610 36464
rect 27618 36528 27938 36529
rect 27618 36464 27626 36528
rect 27690 36464 27706 36528
rect 27770 36464 27786 36528
rect 27850 36464 27866 36528
rect 27930 36464 27938 36528
rect 27618 36463 27938 36464
rect 32946 36528 33266 36529
rect 32946 36464 32954 36528
rect 33018 36464 33034 36528
rect 33098 36464 33114 36528
rect 33178 36464 33194 36528
rect 33258 36464 33266 36528
rect 32946 36463 33266 36464
rect 38274 36528 38594 36529
rect 38274 36464 38282 36528
rect 38346 36464 38362 36528
rect 38426 36464 38442 36528
rect 38506 36464 38522 36528
rect 38586 36464 38594 36528
rect 38274 36463 38594 36464
rect 43602 36528 43922 36529
rect 43602 36464 43610 36528
rect 43674 36464 43690 36528
rect 43754 36464 43770 36528
rect 43834 36464 43850 36528
rect 43914 36464 43922 36528
rect 43602 36463 43922 36464
rect 48930 36528 49250 36529
rect 48930 36464 48938 36528
rect 49002 36464 49018 36528
rect 49082 36464 49098 36528
rect 49162 36464 49178 36528
rect 49242 36464 49250 36528
rect 48930 36463 49250 36464
rect 54258 36528 54578 36529
rect 54258 36464 54266 36528
rect 54330 36464 54346 36528
rect 54410 36464 54426 36528
rect 54490 36464 54506 36528
rect 54570 36464 54578 36528
rect 54258 36463 54578 36464
rect 59586 36528 59906 36529
rect 59586 36464 59594 36528
rect 59658 36464 59674 36528
rect 59738 36464 59754 36528
rect 59818 36464 59834 36528
rect 59898 36464 59906 36528
rect 59586 36463 59906 36464
rect 64914 36528 65234 36529
rect 64914 36464 64922 36528
rect 64986 36464 65002 36528
rect 65066 36464 65082 36528
rect 65146 36464 65162 36528
rect 65226 36464 65234 36528
rect 64914 36463 65234 36464
rect 70242 36528 70562 36529
rect 70242 36464 70250 36528
rect 70314 36464 70330 36528
rect 70394 36464 70410 36528
rect 70474 36464 70490 36528
rect 70554 36464 70562 36528
rect 70242 36463 70562 36464
rect 75570 36528 75890 36529
rect 75570 36464 75578 36528
rect 75642 36464 75658 36528
rect 75722 36464 75738 36528
rect 75802 36464 75818 36528
rect 75882 36464 75890 36528
rect 75570 36463 75890 36464
rect 80898 36528 81218 36529
rect 80898 36464 80906 36528
rect 80970 36464 80986 36528
rect 81050 36464 81066 36528
rect 81130 36464 81146 36528
rect 81210 36464 81218 36528
rect 80898 36463 81218 36464
rect 86226 36528 86546 36529
rect 86226 36464 86234 36528
rect 86298 36464 86314 36528
rect 86378 36464 86394 36528
rect 86458 36464 86474 36528
rect 86538 36464 86546 36528
rect 86226 36463 86546 36464
rect 91554 36528 91874 36529
rect 91554 36464 91562 36528
rect 91626 36464 91642 36528
rect 91706 36464 91722 36528
rect 91786 36464 91802 36528
rect 91866 36464 91874 36528
rect 91554 36463 91874 36464
rect 37443 36186 37509 36189
rect 44251 36186 44317 36189
rect 37443 36184 44317 36186
rect 37443 36128 37448 36184
rect 37504 36128 44256 36184
rect 44312 36128 44317 36184
rect 37443 36126 44317 36128
rect 37443 36123 37509 36126
rect 44251 36123 44317 36126
rect 62559 36186 62625 36189
rect 63019 36186 63085 36189
rect 62559 36184 63085 36186
rect 62559 36128 62564 36184
rect 62620 36128 63024 36184
rect 63080 36128 63085 36184
rect 62559 36126 63085 36128
rect 62559 36123 62625 36126
rect 63019 36123 63085 36126
rect 3642 35984 3962 35985
rect 3642 35920 3650 35984
rect 3714 35920 3730 35984
rect 3794 35920 3810 35984
rect 3874 35920 3890 35984
rect 3954 35920 3962 35984
rect 3642 35919 3962 35920
rect 8970 35984 9290 35985
rect 8970 35920 8978 35984
rect 9042 35920 9058 35984
rect 9122 35920 9138 35984
rect 9202 35920 9218 35984
rect 9282 35920 9290 35984
rect 8970 35919 9290 35920
rect 14298 35984 14618 35985
rect 14298 35920 14306 35984
rect 14370 35920 14386 35984
rect 14450 35920 14466 35984
rect 14530 35920 14546 35984
rect 14610 35920 14618 35984
rect 14298 35919 14618 35920
rect 19626 35984 19946 35985
rect 19626 35920 19634 35984
rect 19698 35920 19714 35984
rect 19778 35920 19794 35984
rect 19858 35920 19874 35984
rect 19938 35920 19946 35984
rect 19626 35919 19946 35920
rect 24954 35984 25274 35985
rect 24954 35920 24962 35984
rect 25026 35920 25042 35984
rect 25106 35920 25122 35984
rect 25186 35920 25202 35984
rect 25266 35920 25274 35984
rect 24954 35919 25274 35920
rect 30282 35984 30602 35985
rect 30282 35920 30290 35984
rect 30354 35920 30370 35984
rect 30434 35920 30450 35984
rect 30514 35920 30530 35984
rect 30594 35920 30602 35984
rect 30282 35919 30602 35920
rect 35610 35984 35930 35985
rect 35610 35920 35618 35984
rect 35682 35920 35698 35984
rect 35762 35920 35778 35984
rect 35842 35920 35858 35984
rect 35922 35920 35930 35984
rect 35610 35919 35930 35920
rect 40938 35984 41258 35985
rect 40938 35920 40946 35984
rect 41010 35920 41026 35984
rect 41090 35920 41106 35984
rect 41170 35920 41186 35984
rect 41250 35920 41258 35984
rect 40938 35919 41258 35920
rect 46266 35984 46586 35985
rect 46266 35920 46274 35984
rect 46338 35920 46354 35984
rect 46418 35920 46434 35984
rect 46498 35920 46514 35984
rect 46578 35920 46586 35984
rect 46266 35919 46586 35920
rect 51594 35984 51914 35985
rect 51594 35920 51602 35984
rect 51666 35920 51682 35984
rect 51746 35920 51762 35984
rect 51826 35920 51842 35984
rect 51906 35920 51914 35984
rect 51594 35919 51914 35920
rect 56922 35984 57242 35985
rect 56922 35920 56930 35984
rect 56994 35920 57010 35984
rect 57074 35920 57090 35984
rect 57154 35920 57170 35984
rect 57234 35920 57242 35984
rect 56922 35919 57242 35920
rect 62250 35984 62570 35985
rect 62250 35920 62258 35984
rect 62322 35920 62338 35984
rect 62402 35920 62418 35984
rect 62482 35920 62498 35984
rect 62562 35920 62570 35984
rect 62250 35919 62570 35920
rect 67578 35984 67898 35985
rect 67578 35920 67586 35984
rect 67650 35920 67666 35984
rect 67730 35920 67746 35984
rect 67810 35920 67826 35984
rect 67890 35920 67898 35984
rect 67578 35919 67898 35920
rect 72906 35984 73226 35985
rect 72906 35920 72914 35984
rect 72978 35920 72994 35984
rect 73058 35920 73074 35984
rect 73138 35920 73154 35984
rect 73218 35920 73226 35984
rect 72906 35919 73226 35920
rect 78234 35984 78554 35985
rect 78234 35920 78242 35984
rect 78306 35920 78322 35984
rect 78386 35920 78402 35984
rect 78466 35920 78482 35984
rect 78546 35920 78554 35984
rect 78234 35919 78554 35920
rect 83562 35984 83882 35985
rect 83562 35920 83570 35984
rect 83634 35920 83650 35984
rect 83714 35920 83730 35984
rect 83794 35920 83810 35984
rect 83874 35920 83882 35984
rect 83562 35919 83882 35920
rect 88890 35984 89210 35985
rect 88890 35920 88898 35984
rect 88962 35920 88978 35984
rect 89042 35920 89058 35984
rect 89122 35920 89138 35984
rect 89202 35920 89210 35984
rect 88890 35919 89210 35920
rect 51519 35778 51585 35781
rect 56671 35778 56737 35781
rect 51519 35776 56737 35778
rect 51519 35720 51524 35776
rect 51580 35720 56676 35776
rect 56732 35720 56737 35776
rect 51519 35718 56737 35720
rect 51519 35715 51585 35718
rect 56671 35715 56737 35718
rect 57867 35778 57933 35781
rect 67987 35778 68053 35781
rect 57867 35776 68053 35778
rect 57867 35720 57872 35776
rect 57928 35720 67992 35776
rect 68048 35720 68053 35776
rect 57867 35718 68053 35720
rect 57867 35715 57933 35718
rect 67987 35715 68053 35718
rect 62375 35506 62441 35509
rect 63939 35506 64005 35509
rect 62375 35504 64005 35506
rect 62375 35448 62380 35504
rect 62436 35448 63944 35504
rect 64000 35448 64005 35504
rect 62375 35446 64005 35448
rect 62375 35443 62441 35446
rect 63939 35443 64005 35446
rect 6306 35440 6626 35441
rect 6306 35376 6314 35440
rect 6378 35376 6394 35440
rect 6458 35376 6474 35440
rect 6538 35376 6554 35440
rect 6618 35376 6626 35440
rect 6306 35375 6626 35376
rect 11634 35440 11954 35441
rect 11634 35376 11642 35440
rect 11706 35376 11722 35440
rect 11786 35376 11802 35440
rect 11866 35376 11882 35440
rect 11946 35376 11954 35440
rect 11634 35375 11954 35376
rect 16962 35440 17282 35441
rect 16962 35376 16970 35440
rect 17034 35376 17050 35440
rect 17114 35376 17130 35440
rect 17194 35376 17210 35440
rect 17274 35376 17282 35440
rect 16962 35375 17282 35376
rect 22290 35440 22610 35441
rect 22290 35376 22298 35440
rect 22362 35376 22378 35440
rect 22442 35376 22458 35440
rect 22522 35376 22538 35440
rect 22602 35376 22610 35440
rect 22290 35375 22610 35376
rect 27618 35440 27938 35441
rect 27618 35376 27626 35440
rect 27690 35376 27706 35440
rect 27770 35376 27786 35440
rect 27850 35376 27866 35440
rect 27930 35376 27938 35440
rect 27618 35375 27938 35376
rect 32946 35440 33266 35441
rect 32946 35376 32954 35440
rect 33018 35376 33034 35440
rect 33098 35376 33114 35440
rect 33178 35376 33194 35440
rect 33258 35376 33266 35440
rect 32946 35375 33266 35376
rect 38274 35440 38594 35441
rect 38274 35376 38282 35440
rect 38346 35376 38362 35440
rect 38426 35376 38442 35440
rect 38506 35376 38522 35440
rect 38586 35376 38594 35440
rect 38274 35375 38594 35376
rect 43602 35440 43922 35441
rect 43602 35376 43610 35440
rect 43674 35376 43690 35440
rect 43754 35376 43770 35440
rect 43834 35376 43850 35440
rect 43914 35376 43922 35440
rect 43602 35375 43922 35376
rect 48930 35440 49250 35441
rect 48930 35376 48938 35440
rect 49002 35376 49018 35440
rect 49082 35376 49098 35440
rect 49162 35376 49178 35440
rect 49242 35376 49250 35440
rect 48930 35375 49250 35376
rect 54258 35440 54578 35441
rect 54258 35376 54266 35440
rect 54330 35376 54346 35440
rect 54410 35376 54426 35440
rect 54490 35376 54506 35440
rect 54570 35376 54578 35440
rect 54258 35375 54578 35376
rect 59586 35440 59906 35441
rect 59586 35376 59594 35440
rect 59658 35376 59674 35440
rect 59738 35376 59754 35440
rect 59818 35376 59834 35440
rect 59898 35376 59906 35440
rect 59586 35375 59906 35376
rect 64914 35440 65234 35441
rect 64914 35376 64922 35440
rect 64986 35376 65002 35440
rect 65066 35376 65082 35440
rect 65146 35376 65162 35440
rect 65226 35376 65234 35440
rect 64914 35375 65234 35376
rect 70242 35440 70562 35441
rect 70242 35376 70250 35440
rect 70314 35376 70330 35440
rect 70394 35376 70410 35440
rect 70474 35376 70490 35440
rect 70554 35376 70562 35440
rect 70242 35375 70562 35376
rect 75570 35440 75890 35441
rect 75570 35376 75578 35440
rect 75642 35376 75658 35440
rect 75722 35376 75738 35440
rect 75802 35376 75818 35440
rect 75882 35376 75890 35440
rect 75570 35375 75890 35376
rect 80898 35440 81218 35441
rect 80898 35376 80906 35440
rect 80970 35376 80986 35440
rect 81050 35376 81066 35440
rect 81130 35376 81146 35440
rect 81210 35376 81218 35440
rect 80898 35375 81218 35376
rect 86226 35440 86546 35441
rect 86226 35376 86234 35440
rect 86298 35376 86314 35440
rect 86378 35376 86394 35440
rect 86458 35376 86474 35440
rect 86538 35376 86546 35440
rect 86226 35375 86546 35376
rect 91554 35440 91874 35441
rect 91554 35376 91562 35440
rect 91626 35376 91642 35440
rect 91706 35376 91722 35440
rect 91786 35376 91802 35440
rect 91866 35376 91874 35440
rect 91554 35375 91874 35376
rect 60811 35370 60877 35373
rect 63295 35370 63361 35373
rect 60811 35368 63361 35370
rect 60811 35312 60816 35368
rect 60872 35312 63300 35368
rect 63356 35312 63361 35368
rect 60811 35310 63361 35312
rect 60811 35307 60877 35310
rect 63295 35307 63361 35310
rect 14719 35234 14785 35237
rect 15087 35234 15153 35237
rect 91263 35234 91329 35237
rect 14719 35232 91329 35234
rect 14719 35176 14724 35232
rect 14780 35176 15092 35232
rect 15148 35176 91268 35232
rect 91324 35176 91329 35232
rect 14719 35174 91329 35176
rect 14719 35171 14785 35174
rect 15087 35171 15153 35174
rect 91263 35171 91329 35174
rect 3642 34896 3962 34897
rect 3642 34832 3650 34896
rect 3714 34832 3730 34896
rect 3794 34832 3810 34896
rect 3874 34832 3890 34896
rect 3954 34832 3962 34896
rect 3642 34831 3962 34832
rect 8970 34896 9290 34897
rect 8970 34832 8978 34896
rect 9042 34832 9058 34896
rect 9122 34832 9138 34896
rect 9202 34832 9218 34896
rect 9282 34832 9290 34896
rect 8970 34831 9290 34832
rect 14298 34896 14618 34897
rect 14298 34832 14306 34896
rect 14370 34832 14386 34896
rect 14450 34832 14466 34896
rect 14530 34832 14546 34896
rect 14610 34832 14618 34896
rect 14298 34831 14618 34832
rect 19626 34896 19946 34897
rect 19626 34832 19634 34896
rect 19698 34832 19714 34896
rect 19778 34832 19794 34896
rect 19858 34832 19874 34896
rect 19938 34832 19946 34896
rect 19626 34831 19946 34832
rect 24954 34896 25274 34897
rect 24954 34832 24962 34896
rect 25026 34832 25042 34896
rect 25106 34832 25122 34896
rect 25186 34832 25202 34896
rect 25266 34832 25274 34896
rect 24954 34831 25274 34832
rect 30282 34896 30602 34897
rect 30282 34832 30290 34896
rect 30354 34832 30370 34896
rect 30434 34832 30450 34896
rect 30514 34832 30530 34896
rect 30594 34832 30602 34896
rect 30282 34831 30602 34832
rect 35610 34896 35930 34897
rect 35610 34832 35618 34896
rect 35682 34832 35698 34896
rect 35762 34832 35778 34896
rect 35842 34832 35858 34896
rect 35922 34832 35930 34896
rect 35610 34831 35930 34832
rect 40938 34896 41258 34897
rect 40938 34832 40946 34896
rect 41010 34832 41026 34896
rect 41090 34832 41106 34896
rect 41170 34832 41186 34896
rect 41250 34832 41258 34896
rect 40938 34831 41258 34832
rect 46266 34896 46586 34897
rect 46266 34832 46274 34896
rect 46338 34832 46354 34896
rect 46418 34832 46434 34896
rect 46498 34832 46514 34896
rect 46578 34832 46586 34896
rect 46266 34831 46586 34832
rect 51594 34896 51914 34897
rect 51594 34832 51602 34896
rect 51666 34832 51682 34896
rect 51746 34832 51762 34896
rect 51826 34832 51842 34896
rect 51906 34832 51914 34896
rect 51594 34831 51914 34832
rect 56922 34896 57242 34897
rect 56922 34832 56930 34896
rect 56994 34832 57010 34896
rect 57074 34832 57090 34896
rect 57154 34832 57170 34896
rect 57234 34832 57242 34896
rect 56922 34831 57242 34832
rect 62250 34896 62570 34897
rect 62250 34832 62258 34896
rect 62322 34832 62338 34896
rect 62402 34832 62418 34896
rect 62482 34832 62498 34896
rect 62562 34832 62570 34896
rect 62250 34831 62570 34832
rect 67578 34896 67898 34897
rect 67578 34832 67586 34896
rect 67650 34832 67666 34896
rect 67730 34832 67746 34896
rect 67810 34832 67826 34896
rect 67890 34832 67898 34896
rect 67578 34831 67898 34832
rect 72906 34896 73226 34897
rect 72906 34832 72914 34896
rect 72978 34832 72994 34896
rect 73058 34832 73074 34896
rect 73138 34832 73154 34896
rect 73218 34832 73226 34896
rect 72906 34831 73226 34832
rect 78234 34896 78554 34897
rect 78234 34832 78242 34896
rect 78306 34832 78322 34896
rect 78386 34832 78402 34896
rect 78466 34832 78482 34896
rect 78546 34832 78554 34896
rect 78234 34831 78554 34832
rect 83562 34896 83882 34897
rect 83562 34832 83570 34896
rect 83634 34832 83650 34896
rect 83714 34832 83730 34896
rect 83794 34832 83810 34896
rect 83874 34832 83882 34896
rect 83562 34831 83882 34832
rect 88890 34896 89210 34897
rect 88890 34832 88898 34896
rect 88962 34832 88978 34896
rect 89042 34832 89058 34896
rect 89122 34832 89138 34896
rect 89202 34832 89210 34896
rect 88890 34831 89210 34832
rect 39375 34690 39441 34693
rect 47011 34690 47077 34693
rect 39375 34688 47077 34690
rect 39375 34632 39380 34688
rect 39436 34632 47016 34688
rect 47072 34632 47077 34688
rect 39375 34630 47077 34632
rect 39375 34627 39441 34630
rect 47011 34627 47077 34630
rect 58419 34554 58485 34557
rect 64123 34554 64189 34557
rect 58419 34552 64189 34554
rect 58419 34496 58424 34552
rect 58480 34496 64128 34552
rect 64184 34496 64189 34552
rect 58419 34494 64189 34496
rect 58419 34491 58485 34494
rect 64123 34491 64189 34494
rect 6306 34352 6626 34353
rect 6306 34288 6314 34352
rect 6378 34288 6394 34352
rect 6458 34288 6474 34352
rect 6538 34288 6554 34352
rect 6618 34288 6626 34352
rect 6306 34287 6626 34288
rect 11634 34352 11954 34353
rect 11634 34288 11642 34352
rect 11706 34288 11722 34352
rect 11786 34288 11802 34352
rect 11866 34288 11882 34352
rect 11946 34288 11954 34352
rect 11634 34287 11954 34288
rect 16962 34352 17282 34353
rect 16962 34288 16970 34352
rect 17034 34288 17050 34352
rect 17114 34288 17130 34352
rect 17194 34288 17210 34352
rect 17274 34288 17282 34352
rect 16962 34287 17282 34288
rect 22290 34352 22610 34353
rect 22290 34288 22298 34352
rect 22362 34288 22378 34352
rect 22442 34288 22458 34352
rect 22522 34288 22538 34352
rect 22602 34288 22610 34352
rect 22290 34287 22610 34288
rect 27618 34352 27938 34353
rect 27618 34288 27626 34352
rect 27690 34288 27706 34352
rect 27770 34288 27786 34352
rect 27850 34288 27866 34352
rect 27930 34288 27938 34352
rect 27618 34287 27938 34288
rect 32946 34352 33266 34353
rect 32946 34288 32954 34352
rect 33018 34288 33034 34352
rect 33098 34288 33114 34352
rect 33178 34288 33194 34352
rect 33258 34288 33266 34352
rect 32946 34287 33266 34288
rect 38274 34352 38594 34353
rect 38274 34288 38282 34352
rect 38346 34288 38362 34352
rect 38426 34288 38442 34352
rect 38506 34288 38522 34352
rect 38586 34288 38594 34352
rect 38274 34287 38594 34288
rect 43602 34352 43922 34353
rect 43602 34288 43610 34352
rect 43674 34288 43690 34352
rect 43754 34288 43770 34352
rect 43834 34288 43850 34352
rect 43914 34288 43922 34352
rect 43602 34287 43922 34288
rect 48930 34352 49250 34353
rect 48930 34288 48938 34352
rect 49002 34288 49018 34352
rect 49082 34288 49098 34352
rect 49162 34288 49178 34352
rect 49242 34288 49250 34352
rect 48930 34287 49250 34288
rect 54258 34352 54578 34353
rect 54258 34288 54266 34352
rect 54330 34288 54346 34352
rect 54410 34288 54426 34352
rect 54490 34288 54506 34352
rect 54570 34288 54578 34352
rect 54258 34287 54578 34288
rect 59586 34352 59906 34353
rect 59586 34288 59594 34352
rect 59658 34288 59674 34352
rect 59738 34288 59754 34352
rect 59818 34288 59834 34352
rect 59898 34288 59906 34352
rect 59586 34287 59906 34288
rect 64914 34352 65234 34353
rect 64914 34288 64922 34352
rect 64986 34288 65002 34352
rect 65066 34288 65082 34352
rect 65146 34288 65162 34352
rect 65226 34288 65234 34352
rect 64914 34287 65234 34288
rect 70242 34352 70562 34353
rect 70242 34288 70250 34352
rect 70314 34288 70330 34352
rect 70394 34288 70410 34352
rect 70474 34288 70490 34352
rect 70554 34288 70562 34352
rect 70242 34287 70562 34288
rect 75570 34352 75890 34353
rect 75570 34288 75578 34352
rect 75642 34288 75658 34352
rect 75722 34288 75738 34352
rect 75802 34288 75818 34352
rect 75882 34288 75890 34352
rect 75570 34287 75890 34288
rect 80898 34352 81218 34353
rect 80898 34288 80906 34352
rect 80970 34288 80986 34352
rect 81050 34288 81066 34352
rect 81130 34288 81146 34352
rect 81210 34288 81218 34352
rect 80898 34287 81218 34288
rect 86226 34352 86546 34353
rect 86226 34288 86234 34352
rect 86298 34288 86314 34352
rect 86378 34288 86394 34352
rect 86458 34288 86474 34352
rect 86538 34288 86546 34352
rect 86226 34287 86546 34288
rect 91554 34352 91874 34353
rect 91554 34288 91562 34352
rect 91626 34288 91642 34352
rect 91706 34288 91722 34352
rect 91786 34288 91802 34352
rect 91866 34288 91874 34352
rect 91554 34287 91874 34288
rect 26863 34010 26929 34013
rect 74059 34010 74125 34013
rect 26863 34008 74125 34010
rect 26863 33952 26868 34008
rect 26924 33952 74064 34008
rect 74120 33952 74125 34008
rect 26863 33950 74125 33952
rect 26863 33947 26929 33950
rect 74059 33947 74125 33950
rect 3642 33808 3962 33809
rect 3642 33744 3650 33808
rect 3714 33744 3730 33808
rect 3794 33744 3810 33808
rect 3874 33744 3890 33808
rect 3954 33744 3962 33808
rect 3642 33743 3962 33744
rect 8970 33808 9290 33809
rect 8970 33744 8978 33808
rect 9042 33744 9058 33808
rect 9122 33744 9138 33808
rect 9202 33744 9218 33808
rect 9282 33744 9290 33808
rect 8970 33743 9290 33744
rect 14298 33808 14618 33809
rect 14298 33744 14306 33808
rect 14370 33744 14386 33808
rect 14450 33744 14466 33808
rect 14530 33744 14546 33808
rect 14610 33744 14618 33808
rect 14298 33743 14618 33744
rect 19626 33808 19946 33809
rect 19626 33744 19634 33808
rect 19698 33744 19714 33808
rect 19778 33744 19794 33808
rect 19858 33744 19874 33808
rect 19938 33744 19946 33808
rect 19626 33743 19946 33744
rect 24954 33808 25274 33809
rect 24954 33744 24962 33808
rect 25026 33744 25042 33808
rect 25106 33744 25122 33808
rect 25186 33744 25202 33808
rect 25266 33744 25274 33808
rect 24954 33743 25274 33744
rect 30282 33808 30602 33809
rect 30282 33744 30290 33808
rect 30354 33744 30370 33808
rect 30434 33744 30450 33808
rect 30514 33744 30530 33808
rect 30594 33744 30602 33808
rect 30282 33743 30602 33744
rect 35610 33808 35930 33809
rect 35610 33744 35618 33808
rect 35682 33744 35698 33808
rect 35762 33744 35778 33808
rect 35842 33744 35858 33808
rect 35922 33744 35930 33808
rect 35610 33743 35930 33744
rect 40938 33808 41258 33809
rect 40938 33744 40946 33808
rect 41010 33744 41026 33808
rect 41090 33744 41106 33808
rect 41170 33744 41186 33808
rect 41250 33744 41258 33808
rect 40938 33743 41258 33744
rect 46266 33808 46586 33809
rect 46266 33744 46274 33808
rect 46338 33744 46354 33808
rect 46418 33744 46434 33808
rect 46498 33744 46514 33808
rect 46578 33744 46586 33808
rect 46266 33743 46586 33744
rect 51594 33808 51914 33809
rect 51594 33744 51602 33808
rect 51666 33744 51682 33808
rect 51746 33744 51762 33808
rect 51826 33744 51842 33808
rect 51906 33744 51914 33808
rect 51594 33743 51914 33744
rect 56922 33808 57242 33809
rect 56922 33744 56930 33808
rect 56994 33744 57010 33808
rect 57074 33744 57090 33808
rect 57154 33744 57170 33808
rect 57234 33744 57242 33808
rect 56922 33743 57242 33744
rect 62250 33808 62570 33809
rect 62250 33744 62258 33808
rect 62322 33744 62338 33808
rect 62402 33744 62418 33808
rect 62482 33744 62498 33808
rect 62562 33744 62570 33808
rect 62250 33743 62570 33744
rect 67578 33808 67898 33809
rect 67578 33744 67586 33808
rect 67650 33744 67666 33808
rect 67730 33744 67746 33808
rect 67810 33744 67826 33808
rect 67890 33744 67898 33808
rect 67578 33743 67898 33744
rect 72906 33808 73226 33809
rect 72906 33744 72914 33808
rect 72978 33744 72994 33808
rect 73058 33744 73074 33808
rect 73138 33744 73154 33808
rect 73218 33744 73226 33808
rect 72906 33743 73226 33744
rect 78234 33808 78554 33809
rect 78234 33744 78242 33808
rect 78306 33744 78322 33808
rect 78386 33744 78402 33808
rect 78466 33744 78482 33808
rect 78546 33744 78554 33808
rect 78234 33743 78554 33744
rect 83562 33808 83882 33809
rect 83562 33744 83570 33808
rect 83634 33744 83650 33808
rect 83714 33744 83730 33808
rect 83794 33744 83810 33808
rect 83874 33744 83882 33808
rect 83562 33743 83882 33744
rect 88890 33808 89210 33809
rect 88890 33744 88898 33808
rect 88962 33744 88978 33808
rect 89042 33744 89058 33808
rect 89122 33744 89138 33808
rect 89202 33744 89210 33808
rect 88890 33743 89210 33744
rect 62651 33738 62717 33741
rect 65963 33738 66029 33741
rect 62651 33736 66029 33738
rect 62651 33680 62656 33736
rect 62712 33680 65968 33736
rect 66024 33680 66029 33736
rect 62651 33678 66029 33680
rect 62651 33675 62717 33678
rect 65963 33675 66029 33678
rect 30359 33602 30425 33605
rect 30727 33602 30793 33605
rect 35235 33602 35301 33605
rect 30359 33600 35301 33602
rect 30359 33544 30364 33600
rect 30420 33544 30732 33600
rect 30788 33544 35240 33600
rect 35296 33544 35301 33600
rect 30359 33542 35301 33544
rect 30359 33539 30425 33542
rect 30727 33539 30793 33542
rect 35235 33539 35301 33542
rect 60903 33602 60969 33605
rect 91355 33602 91421 33605
rect 60903 33600 91421 33602
rect 60903 33544 60908 33600
rect 60964 33544 91360 33600
rect 91416 33544 91421 33600
rect 60903 33542 91421 33544
rect 60903 33539 60969 33542
rect 91355 33539 91421 33542
rect 13891 33466 13957 33469
rect 84363 33466 84429 33469
rect 86019 33466 86085 33469
rect 13891 33464 86085 33466
rect 13891 33408 13896 33464
rect 13952 33408 84368 33464
rect 84424 33408 86024 33464
rect 86080 33408 86085 33464
rect 13891 33406 86085 33408
rect 13891 33403 13957 33406
rect 84363 33403 84429 33406
rect 86019 33403 86085 33406
rect 44987 33330 45053 33333
rect 47103 33330 47169 33333
rect 44987 33328 47169 33330
rect 44987 33272 44992 33328
rect 45048 33272 47108 33328
rect 47164 33272 47169 33328
rect 44987 33270 47169 33272
rect 44987 33267 45053 33270
rect 47103 33267 47169 33270
rect 6306 33264 6626 33265
rect 6306 33200 6314 33264
rect 6378 33200 6394 33264
rect 6458 33200 6474 33264
rect 6538 33200 6554 33264
rect 6618 33200 6626 33264
rect 6306 33199 6626 33200
rect 11634 33264 11954 33265
rect 11634 33200 11642 33264
rect 11706 33200 11722 33264
rect 11786 33200 11802 33264
rect 11866 33200 11882 33264
rect 11946 33200 11954 33264
rect 11634 33199 11954 33200
rect 16962 33264 17282 33265
rect 16962 33200 16970 33264
rect 17034 33200 17050 33264
rect 17114 33200 17130 33264
rect 17194 33200 17210 33264
rect 17274 33200 17282 33264
rect 16962 33199 17282 33200
rect 22290 33264 22610 33265
rect 22290 33200 22298 33264
rect 22362 33200 22378 33264
rect 22442 33200 22458 33264
rect 22522 33200 22538 33264
rect 22602 33200 22610 33264
rect 22290 33199 22610 33200
rect 27618 33264 27938 33265
rect 27618 33200 27626 33264
rect 27690 33200 27706 33264
rect 27770 33200 27786 33264
rect 27850 33200 27866 33264
rect 27930 33200 27938 33264
rect 27618 33199 27938 33200
rect 32946 33264 33266 33265
rect 32946 33200 32954 33264
rect 33018 33200 33034 33264
rect 33098 33200 33114 33264
rect 33178 33200 33194 33264
rect 33258 33200 33266 33264
rect 32946 33199 33266 33200
rect 38274 33264 38594 33265
rect 38274 33200 38282 33264
rect 38346 33200 38362 33264
rect 38426 33200 38442 33264
rect 38506 33200 38522 33264
rect 38586 33200 38594 33264
rect 38274 33199 38594 33200
rect 43602 33264 43922 33265
rect 43602 33200 43610 33264
rect 43674 33200 43690 33264
rect 43754 33200 43770 33264
rect 43834 33200 43850 33264
rect 43914 33200 43922 33264
rect 43602 33199 43922 33200
rect 48930 33264 49250 33265
rect 48930 33200 48938 33264
rect 49002 33200 49018 33264
rect 49082 33200 49098 33264
rect 49162 33200 49178 33264
rect 49242 33200 49250 33264
rect 48930 33199 49250 33200
rect 54258 33264 54578 33265
rect 54258 33200 54266 33264
rect 54330 33200 54346 33264
rect 54410 33200 54426 33264
rect 54490 33200 54506 33264
rect 54570 33200 54578 33264
rect 54258 33199 54578 33200
rect 59586 33264 59906 33265
rect 59586 33200 59594 33264
rect 59658 33200 59674 33264
rect 59738 33200 59754 33264
rect 59818 33200 59834 33264
rect 59898 33200 59906 33264
rect 59586 33199 59906 33200
rect 64914 33264 65234 33265
rect 64914 33200 64922 33264
rect 64986 33200 65002 33264
rect 65066 33200 65082 33264
rect 65146 33200 65162 33264
rect 65226 33200 65234 33264
rect 64914 33199 65234 33200
rect 70242 33264 70562 33265
rect 70242 33200 70250 33264
rect 70314 33200 70330 33264
rect 70394 33200 70410 33264
rect 70474 33200 70490 33264
rect 70554 33200 70562 33264
rect 70242 33199 70562 33200
rect 75570 33264 75890 33265
rect 75570 33200 75578 33264
rect 75642 33200 75658 33264
rect 75722 33200 75738 33264
rect 75802 33200 75818 33264
rect 75882 33200 75890 33264
rect 75570 33199 75890 33200
rect 80898 33264 81218 33265
rect 80898 33200 80906 33264
rect 80970 33200 80986 33264
rect 81050 33200 81066 33264
rect 81130 33200 81146 33264
rect 81210 33200 81218 33264
rect 80898 33199 81218 33200
rect 86226 33264 86546 33265
rect 86226 33200 86234 33264
rect 86298 33200 86314 33264
rect 86378 33200 86394 33264
rect 86458 33200 86474 33264
rect 86538 33200 86546 33264
rect 86226 33199 86546 33200
rect 91554 33264 91874 33265
rect 91554 33200 91562 33264
rect 91626 33200 91642 33264
rect 91706 33200 91722 33264
rect 91786 33200 91802 33264
rect 91866 33200 91874 33264
rect 91554 33199 91874 33200
rect 18491 33058 18557 33061
rect 69735 33058 69801 33061
rect 18491 33056 69801 33058
rect 18491 33000 18496 33056
rect 18552 33000 69740 33056
rect 69796 33000 69801 33056
rect 18491 32998 69801 33000
rect 18491 32995 18557 32998
rect 69735 32995 69801 32998
rect 40111 32922 40177 32925
rect 44895 32922 44961 32925
rect 47287 32922 47353 32925
rect 40111 32920 47353 32922
rect 40111 32864 40116 32920
rect 40172 32864 44900 32920
rect 44956 32864 47292 32920
rect 47348 32864 47353 32920
rect 40111 32862 47353 32864
rect 40111 32859 40177 32862
rect 44895 32859 44961 32862
rect 47287 32859 47353 32862
rect 58787 32922 58853 32925
rect 64675 32922 64741 32925
rect 67067 32922 67133 32925
rect 67435 32922 67501 32925
rect 58787 32920 64554 32922
rect 58787 32864 58792 32920
rect 58848 32864 64554 32920
rect 58787 32862 64554 32864
rect 58787 32859 58853 32862
rect 46735 32786 46801 32789
rect 47379 32786 47445 32789
rect 47563 32786 47629 32789
rect 46735 32784 47629 32786
rect 46735 32728 46740 32784
rect 46796 32728 47384 32784
rect 47440 32728 47568 32784
rect 47624 32728 47629 32784
rect 46735 32726 47629 32728
rect 46735 32723 46801 32726
rect 47379 32723 47445 32726
rect 47563 32723 47629 32726
rect 63203 32786 63269 32789
rect 64123 32786 64189 32789
rect 63203 32784 64189 32786
rect 63203 32728 63208 32784
rect 63264 32728 64128 32784
rect 64184 32728 64189 32784
rect 63203 32726 64189 32728
rect 64494 32786 64554 32862
rect 64675 32920 67133 32922
rect 64675 32864 64680 32920
rect 64736 32864 67072 32920
rect 67128 32864 67133 32920
rect 64675 32862 67133 32864
rect 64675 32859 64741 32862
rect 67067 32859 67133 32862
rect 67392 32920 67501 32922
rect 67392 32864 67440 32920
rect 67496 32864 67501 32920
rect 67392 32859 67501 32864
rect 66699 32786 66765 32789
rect 67392 32786 67452 32859
rect 64494 32784 67452 32786
rect 64494 32728 66704 32784
rect 66760 32728 67452 32784
rect 64494 32726 67452 32728
rect 63203 32723 63269 32726
rect 64123 32723 64189 32726
rect 66699 32723 66765 32726
rect 3642 32720 3962 32721
rect 3642 32656 3650 32720
rect 3714 32656 3730 32720
rect 3794 32656 3810 32720
rect 3874 32656 3890 32720
rect 3954 32656 3962 32720
rect 3642 32655 3962 32656
rect 8970 32720 9290 32721
rect 8970 32656 8978 32720
rect 9042 32656 9058 32720
rect 9122 32656 9138 32720
rect 9202 32656 9218 32720
rect 9282 32656 9290 32720
rect 8970 32655 9290 32656
rect 14298 32720 14618 32721
rect 14298 32656 14306 32720
rect 14370 32656 14386 32720
rect 14450 32656 14466 32720
rect 14530 32656 14546 32720
rect 14610 32656 14618 32720
rect 14298 32655 14618 32656
rect 19626 32720 19946 32721
rect 19626 32656 19634 32720
rect 19698 32656 19714 32720
rect 19778 32656 19794 32720
rect 19858 32656 19874 32720
rect 19938 32656 19946 32720
rect 19626 32655 19946 32656
rect 24954 32720 25274 32721
rect 24954 32656 24962 32720
rect 25026 32656 25042 32720
rect 25106 32656 25122 32720
rect 25186 32656 25202 32720
rect 25266 32656 25274 32720
rect 24954 32655 25274 32656
rect 30282 32720 30602 32721
rect 30282 32656 30290 32720
rect 30354 32656 30370 32720
rect 30434 32656 30450 32720
rect 30514 32656 30530 32720
rect 30594 32656 30602 32720
rect 30282 32655 30602 32656
rect 35610 32720 35930 32721
rect 35610 32656 35618 32720
rect 35682 32656 35698 32720
rect 35762 32656 35778 32720
rect 35842 32656 35858 32720
rect 35922 32656 35930 32720
rect 35610 32655 35930 32656
rect 40938 32720 41258 32721
rect 40938 32656 40946 32720
rect 41010 32656 41026 32720
rect 41090 32656 41106 32720
rect 41170 32656 41186 32720
rect 41250 32656 41258 32720
rect 40938 32655 41258 32656
rect 46266 32720 46586 32721
rect 46266 32656 46274 32720
rect 46338 32656 46354 32720
rect 46418 32656 46434 32720
rect 46498 32656 46514 32720
rect 46578 32656 46586 32720
rect 46266 32655 46586 32656
rect 51594 32720 51914 32721
rect 51594 32656 51602 32720
rect 51666 32656 51682 32720
rect 51746 32656 51762 32720
rect 51826 32656 51842 32720
rect 51906 32656 51914 32720
rect 51594 32655 51914 32656
rect 56922 32720 57242 32721
rect 56922 32656 56930 32720
rect 56994 32656 57010 32720
rect 57074 32656 57090 32720
rect 57154 32656 57170 32720
rect 57234 32656 57242 32720
rect 56922 32655 57242 32656
rect 62250 32720 62570 32721
rect 62250 32656 62258 32720
rect 62322 32656 62338 32720
rect 62402 32656 62418 32720
rect 62482 32656 62498 32720
rect 62562 32656 62570 32720
rect 62250 32655 62570 32656
rect 67578 32720 67898 32721
rect 67578 32656 67586 32720
rect 67650 32656 67666 32720
rect 67730 32656 67746 32720
rect 67810 32656 67826 32720
rect 67890 32656 67898 32720
rect 67578 32655 67898 32656
rect 72906 32720 73226 32721
rect 72906 32656 72914 32720
rect 72978 32656 72994 32720
rect 73058 32656 73074 32720
rect 73138 32656 73154 32720
rect 73218 32656 73226 32720
rect 72906 32655 73226 32656
rect 78234 32720 78554 32721
rect 78234 32656 78242 32720
rect 78306 32656 78322 32720
rect 78386 32656 78402 32720
rect 78466 32656 78482 32720
rect 78546 32656 78554 32720
rect 78234 32655 78554 32656
rect 83562 32720 83882 32721
rect 83562 32656 83570 32720
rect 83634 32656 83650 32720
rect 83714 32656 83730 32720
rect 83794 32656 83810 32720
rect 83874 32656 83882 32720
rect 83562 32655 83882 32656
rect 88890 32720 89210 32721
rect 88890 32656 88898 32720
rect 88962 32656 88978 32720
rect 89042 32656 89058 32720
rect 89122 32656 89138 32720
rect 89202 32656 89210 32720
rect 88890 32655 89210 32656
rect 57867 32650 57933 32653
rect 62007 32650 62073 32653
rect 57867 32648 62073 32650
rect 57867 32592 57872 32648
rect 57928 32592 62012 32648
rect 62068 32592 62073 32648
rect 57867 32590 62073 32592
rect 57867 32587 57933 32590
rect 62007 32587 62073 32590
rect 63387 32650 63453 32653
rect 64675 32650 64741 32653
rect 63387 32648 64741 32650
rect 63387 32592 63392 32648
rect 63448 32592 64680 32648
rect 64736 32592 64741 32648
rect 63387 32590 64741 32592
rect 63387 32587 63453 32590
rect 64675 32587 64741 32590
rect 91079 32650 91145 32653
rect 93946 32650 94746 32680
rect 91079 32648 94746 32650
rect 91079 32592 91084 32648
rect 91140 32592 94746 32648
rect 91079 32590 94746 32592
rect 91079 32587 91145 32590
rect 93946 32560 94746 32590
rect 48391 32514 48457 32517
rect 52807 32514 52873 32517
rect 48391 32512 52873 32514
rect 48391 32456 48396 32512
rect 48452 32456 52812 32512
rect 52868 32456 52873 32512
rect 48391 32454 52873 32456
rect 48391 32451 48457 32454
rect 52807 32451 52873 32454
rect 59799 32514 59865 32517
rect 67895 32514 67961 32517
rect 59799 32512 67961 32514
rect 59799 32456 59804 32512
rect 59860 32456 67900 32512
rect 67956 32456 67961 32512
rect 59799 32454 67961 32456
rect 59799 32451 59865 32454
rect 67895 32451 67961 32454
rect 41767 32378 41833 32381
rect 47195 32378 47261 32381
rect 47931 32378 47997 32381
rect 41767 32376 47997 32378
rect 41767 32320 41772 32376
rect 41828 32320 47200 32376
rect 47256 32320 47936 32376
rect 47992 32320 47997 32376
rect 41767 32318 47997 32320
rect 41767 32315 41833 32318
rect 47195 32315 47261 32318
rect 47931 32315 47997 32318
rect 67159 32378 67225 32381
rect 68355 32378 68421 32381
rect 67159 32376 68421 32378
rect 67159 32320 67164 32376
rect 67220 32320 68360 32376
rect 68416 32320 68421 32376
rect 67159 32318 68421 32320
rect 67159 32315 67225 32318
rect 68355 32315 68421 32318
rect 73691 32378 73757 32381
rect 74611 32378 74677 32381
rect 73691 32376 74677 32378
rect 73691 32320 73696 32376
rect 73752 32320 74616 32376
rect 74672 32320 74677 32376
rect 73691 32318 74677 32320
rect 73691 32315 73757 32318
rect 74611 32315 74677 32318
rect 46459 32242 46525 32245
rect 47563 32242 47629 32245
rect 46459 32240 47629 32242
rect 46459 32184 46464 32240
rect 46520 32184 47568 32240
rect 47624 32184 47629 32240
rect 46459 32182 47629 32184
rect 46459 32179 46525 32182
rect 47563 32179 47629 32182
rect 58419 32242 58485 32245
rect 58695 32242 58761 32245
rect 58419 32240 58761 32242
rect 58419 32184 58424 32240
rect 58480 32184 58700 32240
rect 58756 32184 58761 32240
rect 58419 32182 58761 32184
rect 58419 32179 58485 32182
rect 58695 32179 58761 32182
rect 60075 32242 60141 32245
rect 64491 32242 64557 32245
rect 60075 32240 64557 32242
rect 60075 32184 60080 32240
rect 60136 32184 64496 32240
rect 64552 32184 64557 32240
rect 60075 32182 64557 32184
rect 60075 32179 60141 32182
rect 64491 32179 64557 32182
rect 6306 32176 6626 32177
rect 6306 32112 6314 32176
rect 6378 32112 6394 32176
rect 6458 32112 6474 32176
rect 6538 32112 6554 32176
rect 6618 32112 6626 32176
rect 6306 32111 6626 32112
rect 11634 32176 11954 32177
rect 11634 32112 11642 32176
rect 11706 32112 11722 32176
rect 11786 32112 11802 32176
rect 11866 32112 11882 32176
rect 11946 32112 11954 32176
rect 11634 32111 11954 32112
rect 16962 32176 17282 32177
rect 16962 32112 16970 32176
rect 17034 32112 17050 32176
rect 17114 32112 17130 32176
rect 17194 32112 17210 32176
rect 17274 32112 17282 32176
rect 16962 32111 17282 32112
rect 22290 32176 22610 32177
rect 22290 32112 22298 32176
rect 22362 32112 22378 32176
rect 22442 32112 22458 32176
rect 22522 32112 22538 32176
rect 22602 32112 22610 32176
rect 22290 32111 22610 32112
rect 27618 32176 27938 32177
rect 27618 32112 27626 32176
rect 27690 32112 27706 32176
rect 27770 32112 27786 32176
rect 27850 32112 27866 32176
rect 27930 32112 27938 32176
rect 27618 32111 27938 32112
rect 32946 32176 33266 32177
rect 32946 32112 32954 32176
rect 33018 32112 33034 32176
rect 33098 32112 33114 32176
rect 33178 32112 33194 32176
rect 33258 32112 33266 32176
rect 32946 32111 33266 32112
rect 38274 32176 38594 32177
rect 38274 32112 38282 32176
rect 38346 32112 38362 32176
rect 38426 32112 38442 32176
rect 38506 32112 38522 32176
rect 38586 32112 38594 32176
rect 38274 32111 38594 32112
rect 43602 32176 43922 32177
rect 43602 32112 43610 32176
rect 43674 32112 43690 32176
rect 43754 32112 43770 32176
rect 43834 32112 43850 32176
rect 43914 32112 43922 32176
rect 43602 32111 43922 32112
rect 48930 32176 49250 32177
rect 48930 32112 48938 32176
rect 49002 32112 49018 32176
rect 49082 32112 49098 32176
rect 49162 32112 49178 32176
rect 49242 32112 49250 32176
rect 48930 32111 49250 32112
rect 54258 32176 54578 32177
rect 54258 32112 54266 32176
rect 54330 32112 54346 32176
rect 54410 32112 54426 32176
rect 54490 32112 54506 32176
rect 54570 32112 54578 32176
rect 54258 32111 54578 32112
rect 59586 32176 59906 32177
rect 59586 32112 59594 32176
rect 59658 32112 59674 32176
rect 59738 32112 59754 32176
rect 59818 32112 59834 32176
rect 59898 32112 59906 32176
rect 59586 32111 59906 32112
rect 64914 32176 65234 32177
rect 64914 32112 64922 32176
rect 64986 32112 65002 32176
rect 65066 32112 65082 32176
rect 65146 32112 65162 32176
rect 65226 32112 65234 32176
rect 64914 32111 65234 32112
rect 70242 32176 70562 32177
rect 70242 32112 70250 32176
rect 70314 32112 70330 32176
rect 70394 32112 70410 32176
rect 70474 32112 70490 32176
rect 70554 32112 70562 32176
rect 70242 32111 70562 32112
rect 75570 32176 75890 32177
rect 75570 32112 75578 32176
rect 75642 32112 75658 32176
rect 75722 32112 75738 32176
rect 75802 32112 75818 32176
rect 75882 32112 75890 32176
rect 75570 32111 75890 32112
rect 80898 32176 81218 32177
rect 80898 32112 80906 32176
rect 80970 32112 80986 32176
rect 81050 32112 81066 32176
rect 81130 32112 81146 32176
rect 81210 32112 81218 32176
rect 80898 32111 81218 32112
rect 86226 32176 86546 32177
rect 86226 32112 86234 32176
rect 86298 32112 86314 32176
rect 86378 32112 86394 32176
rect 86458 32112 86474 32176
rect 86538 32112 86546 32176
rect 86226 32111 86546 32112
rect 91554 32176 91874 32177
rect 91554 32112 91562 32176
rect 91626 32112 91642 32176
rect 91706 32112 91722 32176
rect 91786 32112 91802 32176
rect 91866 32112 91874 32176
rect 91554 32111 91874 32112
rect 63295 32106 63361 32109
rect 64675 32106 64741 32109
rect 63295 32104 64741 32106
rect 63295 32048 63300 32104
rect 63356 32048 64680 32104
rect 64736 32048 64741 32104
rect 63295 32046 64741 32048
rect 63295 32043 63361 32046
rect 64675 32043 64741 32046
rect 18951 31970 19017 31973
rect 24011 31970 24077 31973
rect 18951 31968 24077 31970
rect 18951 31912 18956 31968
rect 19012 31912 24016 31968
rect 24072 31912 24077 31968
rect 18951 31910 24077 31912
rect 18951 31907 19017 31910
rect 24011 31907 24077 31910
rect 58603 31970 58669 31973
rect 65503 31970 65569 31973
rect 58603 31968 65569 31970
rect 58603 31912 58608 31968
rect 58664 31912 65508 31968
rect 65564 31912 65569 31968
rect 58603 31910 65569 31912
rect 58603 31907 58669 31910
rect 65503 31907 65569 31910
rect 68999 31970 69065 31973
rect 69643 31970 69709 31973
rect 68999 31968 69709 31970
rect 68999 31912 69004 31968
rect 69060 31912 69648 31968
rect 69704 31912 69709 31968
rect 68999 31910 69709 31912
rect 68999 31907 69065 31910
rect 69643 31907 69709 31910
rect 17295 31834 17361 31837
rect 19411 31834 19477 31837
rect 17295 31832 19477 31834
rect 17295 31776 17300 31832
rect 17356 31776 19416 31832
rect 19472 31776 19477 31832
rect 17295 31774 19477 31776
rect 17295 31771 17361 31774
rect 19411 31771 19477 31774
rect 28519 31834 28585 31837
rect 28979 31834 29045 31837
rect 28519 31832 29045 31834
rect 28519 31776 28524 31832
rect 28580 31776 28984 31832
rect 29040 31776 29045 31832
rect 28519 31774 29045 31776
rect 28519 31771 28585 31774
rect 28979 31771 29045 31774
rect 57591 31834 57657 31837
rect 58879 31834 58945 31837
rect 57591 31832 58945 31834
rect 57591 31776 57596 31832
rect 57652 31776 58884 31832
rect 58940 31776 58945 31832
rect 57591 31774 58945 31776
rect 57591 31771 57657 31774
rect 58879 31771 58945 31774
rect 3642 31632 3962 31633
rect 3642 31568 3650 31632
rect 3714 31568 3730 31632
rect 3794 31568 3810 31632
rect 3874 31568 3890 31632
rect 3954 31568 3962 31632
rect 3642 31567 3962 31568
rect 8970 31632 9290 31633
rect 8970 31568 8978 31632
rect 9042 31568 9058 31632
rect 9122 31568 9138 31632
rect 9202 31568 9218 31632
rect 9282 31568 9290 31632
rect 8970 31567 9290 31568
rect 14298 31632 14618 31633
rect 14298 31568 14306 31632
rect 14370 31568 14386 31632
rect 14450 31568 14466 31632
rect 14530 31568 14546 31632
rect 14610 31568 14618 31632
rect 14298 31567 14618 31568
rect 19626 31632 19946 31633
rect 19626 31568 19634 31632
rect 19698 31568 19714 31632
rect 19778 31568 19794 31632
rect 19858 31568 19874 31632
rect 19938 31568 19946 31632
rect 19626 31567 19946 31568
rect 24954 31632 25274 31633
rect 24954 31568 24962 31632
rect 25026 31568 25042 31632
rect 25106 31568 25122 31632
rect 25186 31568 25202 31632
rect 25266 31568 25274 31632
rect 24954 31567 25274 31568
rect 30282 31632 30602 31633
rect 30282 31568 30290 31632
rect 30354 31568 30370 31632
rect 30434 31568 30450 31632
rect 30514 31568 30530 31632
rect 30594 31568 30602 31632
rect 30282 31567 30602 31568
rect 35610 31632 35930 31633
rect 35610 31568 35618 31632
rect 35682 31568 35698 31632
rect 35762 31568 35778 31632
rect 35842 31568 35858 31632
rect 35922 31568 35930 31632
rect 35610 31567 35930 31568
rect 40938 31632 41258 31633
rect 40938 31568 40946 31632
rect 41010 31568 41026 31632
rect 41090 31568 41106 31632
rect 41170 31568 41186 31632
rect 41250 31568 41258 31632
rect 40938 31567 41258 31568
rect 46266 31632 46586 31633
rect 46266 31568 46274 31632
rect 46338 31568 46354 31632
rect 46418 31568 46434 31632
rect 46498 31568 46514 31632
rect 46578 31568 46586 31632
rect 46266 31567 46586 31568
rect 51594 31632 51914 31633
rect 51594 31568 51602 31632
rect 51666 31568 51682 31632
rect 51746 31568 51762 31632
rect 51826 31568 51842 31632
rect 51906 31568 51914 31632
rect 51594 31567 51914 31568
rect 56922 31632 57242 31633
rect 56922 31568 56930 31632
rect 56994 31568 57010 31632
rect 57074 31568 57090 31632
rect 57154 31568 57170 31632
rect 57234 31568 57242 31632
rect 56922 31567 57242 31568
rect 62250 31632 62570 31633
rect 62250 31568 62258 31632
rect 62322 31568 62338 31632
rect 62402 31568 62418 31632
rect 62482 31568 62498 31632
rect 62562 31568 62570 31632
rect 62250 31567 62570 31568
rect 67578 31632 67898 31633
rect 67578 31568 67586 31632
rect 67650 31568 67666 31632
rect 67730 31568 67746 31632
rect 67810 31568 67826 31632
rect 67890 31568 67898 31632
rect 67578 31567 67898 31568
rect 72906 31632 73226 31633
rect 72906 31568 72914 31632
rect 72978 31568 72994 31632
rect 73058 31568 73074 31632
rect 73138 31568 73154 31632
rect 73218 31568 73226 31632
rect 72906 31567 73226 31568
rect 78234 31632 78554 31633
rect 78234 31568 78242 31632
rect 78306 31568 78322 31632
rect 78386 31568 78402 31632
rect 78466 31568 78482 31632
rect 78546 31568 78554 31632
rect 78234 31567 78554 31568
rect 83562 31632 83882 31633
rect 83562 31568 83570 31632
rect 83634 31568 83650 31632
rect 83714 31568 83730 31632
rect 83794 31568 83810 31632
rect 83874 31568 83882 31632
rect 83562 31567 83882 31568
rect 88890 31632 89210 31633
rect 88890 31568 88898 31632
rect 88962 31568 88978 31632
rect 89042 31568 89058 31632
rect 89122 31568 89138 31632
rect 89202 31568 89210 31632
rect 88890 31567 89210 31568
rect 28427 31426 28493 31429
rect 28703 31426 28769 31429
rect 32567 31426 32633 31429
rect 28427 31424 32633 31426
rect 28427 31368 28432 31424
rect 28488 31368 28708 31424
rect 28764 31368 32572 31424
rect 32628 31368 32633 31424
rect 28427 31366 32633 31368
rect 28427 31363 28493 31366
rect 28703 31363 28769 31366
rect 32567 31363 32633 31366
rect 46459 31426 46525 31429
rect 54739 31426 54805 31429
rect 46459 31424 54805 31426
rect 46459 31368 46464 31424
rect 46520 31368 54744 31424
rect 54800 31368 54805 31424
rect 46459 31366 54805 31368
rect 46459 31363 46525 31366
rect 54739 31363 54805 31366
rect 28519 31290 28585 31293
rect 40847 31290 40913 31293
rect 28519 31288 40913 31290
rect 28519 31232 28524 31288
rect 28580 31232 40852 31288
rect 40908 31232 40913 31288
rect 28519 31230 40913 31232
rect 28519 31227 28585 31230
rect 40847 31227 40913 31230
rect 57499 31290 57565 31293
rect 60167 31290 60233 31293
rect 57499 31288 60233 31290
rect 57499 31232 57504 31288
rect 57560 31232 60172 31288
rect 60228 31232 60233 31288
rect 57499 31230 60233 31232
rect 57499 31227 57565 31230
rect 60167 31227 60233 31230
rect 6306 31088 6626 31089
rect 6306 31024 6314 31088
rect 6378 31024 6394 31088
rect 6458 31024 6474 31088
rect 6538 31024 6554 31088
rect 6618 31024 6626 31088
rect 6306 31023 6626 31024
rect 11634 31088 11954 31089
rect 11634 31024 11642 31088
rect 11706 31024 11722 31088
rect 11786 31024 11802 31088
rect 11866 31024 11882 31088
rect 11946 31024 11954 31088
rect 11634 31023 11954 31024
rect 16962 31088 17282 31089
rect 16962 31024 16970 31088
rect 17034 31024 17050 31088
rect 17114 31024 17130 31088
rect 17194 31024 17210 31088
rect 17274 31024 17282 31088
rect 16962 31023 17282 31024
rect 22290 31088 22610 31089
rect 22290 31024 22298 31088
rect 22362 31024 22378 31088
rect 22442 31024 22458 31088
rect 22522 31024 22538 31088
rect 22602 31024 22610 31088
rect 22290 31023 22610 31024
rect 27618 31088 27938 31089
rect 27618 31024 27626 31088
rect 27690 31024 27706 31088
rect 27770 31024 27786 31088
rect 27850 31024 27866 31088
rect 27930 31024 27938 31088
rect 27618 31023 27938 31024
rect 32946 31088 33266 31089
rect 32946 31024 32954 31088
rect 33018 31024 33034 31088
rect 33098 31024 33114 31088
rect 33178 31024 33194 31088
rect 33258 31024 33266 31088
rect 32946 31023 33266 31024
rect 38274 31088 38594 31089
rect 38274 31024 38282 31088
rect 38346 31024 38362 31088
rect 38426 31024 38442 31088
rect 38506 31024 38522 31088
rect 38586 31024 38594 31088
rect 38274 31023 38594 31024
rect 43602 31088 43922 31089
rect 43602 31024 43610 31088
rect 43674 31024 43690 31088
rect 43754 31024 43770 31088
rect 43834 31024 43850 31088
rect 43914 31024 43922 31088
rect 43602 31023 43922 31024
rect 48930 31088 49250 31089
rect 48930 31024 48938 31088
rect 49002 31024 49018 31088
rect 49082 31024 49098 31088
rect 49162 31024 49178 31088
rect 49242 31024 49250 31088
rect 48930 31023 49250 31024
rect 54258 31088 54578 31089
rect 54258 31024 54266 31088
rect 54330 31024 54346 31088
rect 54410 31024 54426 31088
rect 54490 31024 54506 31088
rect 54570 31024 54578 31088
rect 54258 31023 54578 31024
rect 59586 31088 59906 31089
rect 59586 31024 59594 31088
rect 59658 31024 59674 31088
rect 59738 31024 59754 31088
rect 59818 31024 59834 31088
rect 59898 31024 59906 31088
rect 59586 31023 59906 31024
rect 64914 31088 65234 31089
rect 64914 31024 64922 31088
rect 64986 31024 65002 31088
rect 65066 31024 65082 31088
rect 65146 31024 65162 31088
rect 65226 31024 65234 31088
rect 64914 31023 65234 31024
rect 70242 31088 70562 31089
rect 70242 31024 70250 31088
rect 70314 31024 70330 31088
rect 70394 31024 70410 31088
rect 70474 31024 70490 31088
rect 70554 31024 70562 31088
rect 70242 31023 70562 31024
rect 75570 31088 75890 31089
rect 75570 31024 75578 31088
rect 75642 31024 75658 31088
rect 75722 31024 75738 31088
rect 75802 31024 75818 31088
rect 75882 31024 75890 31088
rect 75570 31023 75890 31024
rect 80898 31088 81218 31089
rect 80898 31024 80906 31088
rect 80970 31024 80986 31088
rect 81050 31024 81066 31088
rect 81130 31024 81146 31088
rect 81210 31024 81218 31088
rect 80898 31023 81218 31024
rect 86226 31088 86546 31089
rect 86226 31024 86234 31088
rect 86298 31024 86314 31088
rect 86378 31024 86394 31088
rect 86458 31024 86474 31088
rect 86538 31024 86546 31088
rect 86226 31023 86546 31024
rect 91554 31088 91874 31089
rect 91554 31024 91562 31088
rect 91626 31024 91642 31088
rect 91706 31024 91722 31088
rect 91786 31024 91802 31088
rect 91866 31024 91874 31088
rect 91554 31023 91874 31024
rect 16743 30882 16809 30885
rect 17755 30882 17821 30885
rect 16743 30880 17821 30882
rect 16743 30824 16748 30880
rect 16804 30824 17760 30880
rect 17816 30824 17821 30880
rect 16743 30822 17821 30824
rect 16743 30819 16809 30822
rect 17755 30819 17821 30822
rect 52163 30882 52229 30885
rect 53911 30882 53977 30885
rect 52163 30880 53977 30882
rect 52163 30824 52168 30880
rect 52224 30824 53916 30880
rect 53972 30824 53977 30880
rect 52163 30822 53977 30824
rect 52163 30819 52229 30822
rect 53911 30819 53977 30822
rect 80315 30882 80381 30885
rect 80959 30882 81025 30885
rect 80315 30880 81025 30882
rect 80315 30824 80320 30880
rect 80376 30824 80964 30880
rect 81020 30824 81025 30880
rect 80315 30822 81025 30824
rect 80315 30819 80381 30822
rect 80959 30819 81025 30822
rect 3642 30544 3962 30545
rect 3642 30480 3650 30544
rect 3714 30480 3730 30544
rect 3794 30480 3810 30544
rect 3874 30480 3890 30544
rect 3954 30480 3962 30544
rect 3642 30479 3962 30480
rect 8970 30544 9290 30545
rect 8970 30480 8978 30544
rect 9042 30480 9058 30544
rect 9122 30480 9138 30544
rect 9202 30480 9218 30544
rect 9282 30480 9290 30544
rect 8970 30479 9290 30480
rect 14298 30544 14618 30545
rect 14298 30480 14306 30544
rect 14370 30480 14386 30544
rect 14450 30480 14466 30544
rect 14530 30480 14546 30544
rect 14610 30480 14618 30544
rect 14298 30479 14618 30480
rect 19626 30544 19946 30545
rect 19626 30480 19634 30544
rect 19698 30480 19714 30544
rect 19778 30480 19794 30544
rect 19858 30480 19874 30544
rect 19938 30480 19946 30544
rect 19626 30479 19946 30480
rect 24954 30544 25274 30545
rect 24954 30480 24962 30544
rect 25026 30480 25042 30544
rect 25106 30480 25122 30544
rect 25186 30480 25202 30544
rect 25266 30480 25274 30544
rect 24954 30479 25274 30480
rect 30282 30544 30602 30545
rect 30282 30480 30290 30544
rect 30354 30480 30370 30544
rect 30434 30480 30450 30544
rect 30514 30480 30530 30544
rect 30594 30480 30602 30544
rect 30282 30479 30602 30480
rect 35610 30544 35930 30545
rect 35610 30480 35618 30544
rect 35682 30480 35698 30544
rect 35762 30480 35778 30544
rect 35842 30480 35858 30544
rect 35922 30480 35930 30544
rect 35610 30479 35930 30480
rect 40938 30544 41258 30545
rect 40938 30480 40946 30544
rect 41010 30480 41026 30544
rect 41090 30480 41106 30544
rect 41170 30480 41186 30544
rect 41250 30480 41258 30544
rect 40938 30479 41258 30480
rect 46266 30544 46586 30545
rect 46266 30480 46274 30544
rect 46338 30480 46354 30544
rect 46418 30480 46434 30544
rect 46498 30480 46514 30544
rect 46578 30480 46586 30544
rect 46266 30479 46586 30480
rect 51594 30544 51914 30545
rect 51594 30480 51602 30544
rect 51666 30480 51682 30544
rect 51746 30480 51762 30544
rect 51826 30480 51842 30544
rect 51906 30480 51914 30544
rect 51594 30479 51914 30480
rect 56922 30544 57242 30545
rect 56922 30480 56930 30544
rect 56994 30480 57010 30544
rect 57074 30480 57090 30544
rect 57154 30480 57170 30544
rect 57234 30480 57242 30544
rect 56922 30479 57242 30480
rect 62250 30544 62570 30545
rect 62250 30480 62258 30544
rect 62322 30480 62338 30544
rect 62402 30480 62418 30544
rect 62482 30480 62498 30544
rect 62562 30480 62570 30544
rect 62250 30479 62570 30480
rect 67578 30544 67898 30545
rect 67578 30480 67586 30544
rect 67650 30480 67666 30544
rect 67730 30480 67746 30544
rect 67810 30480 67826 30544
rect 67890 30480 67898 30544
rect 67578 30479 67898 30480
rect 72906 30544 73226 30545
rect 72906 30480 72914 30544
rect 72978 30480 72994 30544
rect 73058 30480 73074 30544
rect 73138 30480 73154 30544
rect 73218 30480 73226 30544
rect 72906 30479 73226 30480
rect 78234 30544 78554 30545
rect 78234 30480 78242 30544
rect 78306 30480 78322 30544
rect 78386 30480 78402 30544
rect 78466 30480 78482 30544
rect 78546 30480 78554 30544
rect 78234 30479 78554 30480
rect 83562 30544 83882 30545
rect 83562 30480 83570 30544
rect 83634 30480 83650 30544
rect 83714 30480 83730 30544
rect 83794 30480 83810 30544
rect 83874 30480 83882 30544
rect 83562 30479 83882 30480
rect 88890 30544 89210 30545
rect 88890 30480 88898 30544
rect 88962 30480 88978 30544
rect 89042 30480 89058 30544
rect 89122 30480 89138 30544
rect 89202 30480 89210 30544
rect 88890 30479 89210 30480
rect 19595 30338 19661 30341
rect 28335 30338 28401 30341
rect 19595 30336 28401 30338
rect 19595 30280 19600 30336
rect 19656 30280 28340 30336
rect 28396 30280 28401 30336
rect 19595 30278 28401 30280
rect 19595 30275 19661 30278
rect 28335 30275 28401 30278
rect 62099 30338 62165 30341
rect 65411 30338 65477 30341
rect 62099 30336 65477 30338
rect 62099 30280 62104 30336
rect 62160 30280 65416 30336
rect 65472 30280 65477 30336
rect 62099 30278 65477 30280
rect 62099 30275 62165 30278
rect 65411 30275 65477 30278
rect 69827 30338 69893 30341
rect 74519 30338 74585 30341
rect 69827 30336 74585 30338
rect 69827 30280 69832 30336
rect 69888 30280 74524 30336
rect 74580 30280 74585 30336
rect 69827 30278 74585 30280
rect 69827 30275 69893 30278
rect 74519 30275 74585 30278
rect 59983 30202 60049 30205
rect 66607 30202 66673 30205
rect 59983 30200 66673 30202
rect 59983 30144 59988 30200
rect 60044 30144 66612 30200
rect 66668 30144 66673 30200
rect 59983 30142 66673 30144
rect 59983 30139 60049 30142
rect 66607 30139 66673 30142
rect 6306 30000 6626 30001
rect 6306 29936 6314 30000
rect 6378 29936 6394 30000
rect 6458 29936 6474 30000
rect 6538 29936 6554 30000
rect 6618 29936 6626 30000
rect 6306 29935 6626 29936
rect 11634 30000 11954 30001
rect 11634 29936 11642 30000
rect 11706 29936 11722 30000
rect 11786 29936 11802 30000
rect 11866 29936 11882 30000
rect 11946 29936 11954 30000
rect 11634 29935 11954 29936
rect 16962 30000 17282 30001
rect 16962 29936 16970 30000
rect 17034 29936 17050 30000
rect 17114 29936 17130 30000
rect 17194 29936 17210 30000
rect 17274 29936 17282 30000
rect 16962 29935 17282 29936
rect 22290 30000 22610 30001
rect 22290 29936 22298 30000
rect 22362 29936 22378 30000
rect 22442 29936 22458 30000
rect 22522 29936 22538 30000
rect 22602 29936 22610 30000
rect 22290 29935 22610 29936
rect 27618 30000 27938 30001
rect 27618 29936 27626 30000
rect 27690 29936 27706 30000
rect 27770 29936 27786 30000
rect 27850 29936 27866 30000
rect 27930 29936 27938 30000
rect 27618 29935 27938 29936
rect 32946 30000 33266 30001
rect 32946 29936 32954 30000
rect 33018 29936 33034 30000
rect 33098 29936 33114 30000
rect 33178 29936 33194 30000
rect 33258 29936 33266 30000
rect 32946 29935 33266 29936
rect 38274 30000 38594 30001
rect 38274 29936 38282 30000
rect 38346 29936 38362 30000
rect 38426 29936 38442 30000
rect 38506 29936 38522 30000
rect 38586 29936 38594 30000
rect 38274 29935 38594 29936
rect 43602 30000 43922 30001
rect 43602 29936 43610 30000
rect 43674 29936 43690 30000
rect 43754 29936 43770 30000
rect 43834 29936 43850 30000
rect 43914 29936 43922 30000
rect 43602 29935 43922 29936
rect 48930 30000 49250 30001
rect 48930 29936 48938 30000
rect 49002 29936 49018 30000
rect 49082 29936 49098 30000
rect 49162 29936 49178 30000
rect 49242 29936 49250 30000
rect 48930 29935 49250 29936
rect 54258 30000 54578 30001
rect 54258 29936 54266 30000
rect 54330 29936 54346 30000
rect 54410 29936 54426 30000
rect 54490 29936 54506 30000
rect 54570 29936 54578 30000
rect 54258 29935 54578 29936
rect 59586 30000 59906 30001
rect 59586 29936 59594 30000
rect 59658 29936 59674 30000
rect 59738 29936 59754 30000
rect 59818 29936 59834 30000
rect 59898 29936 59906 30000
rect 59586 29935 59906 29936
rect 64914 30000 65234 30001
rect 64914 29936 64922 30000
rect 64986 29936 65002 30000
rect 65066 29936 65082 30000
rect 65146 29936 65162 30000
rect 65226 29936 65234 30000
rect 64914 29935 65234 29936
rect 70242 30000 70562 30001
rect 70242 29936 70250 30000
rect 70314 29936 70330 30000
rect 70394 29936 70410 30000
rect 70474 29936 70490 30000
rect 70554 29936 70562 30000
rect 70242 29935 70562 29936
rect 75570 30000 75890 30001
rect 75570 29936 75578 30000
rect 75642 29936 75658 30000
rect 75722 29936 75738 30000
rect 75802 29936 75818 30000
rect 75882 29936 75890 30000
rect 75570 29935 75890 29936
rect 80898 30000 81218 30001
rect 80898 29936 80906 30000
rect 80970 29936 80986 30000
rect 81050 29936 81066 30000
rect 81130 29936 81146 30000
rect 81210 29936 81218 30000
rect 80898 29935 81218 29936
rect 86226 30000 86546 30001
rect 86226 29936 86234 30000
rect 86298 29936 86314 30000
rect 86378 29936 86394 30000
rect 86458 29936 86474 30000
rect 86538 29936 86546 30000
rect 86226 29935 86546 29936
rect 91554 30000 91874 30001
rect 91554 29936 91562 30000
rect 91626 29936 91642 30000
rect 91706 29936 91722 30000
rect 91786 29936 91802 30000
rect 91866 29936 91874 30000
rect 91554 29935 91874 29936
rect 22723 29930 22789 29933
rect 27415 29930 27481 29933
rect 22723 29928 27481 29930
rect 22723 29872 22728 29928
rect 22784 29872 27420 29928
rect 27476 29872 27481 29928
rect 22723 29870 27481 29872
rect 22723 29867 22789 29870
rect 27415 29867 27481 29870
rect 74979 29794 75045 29797
rect 76635 29794 76701 29797
rect 74979 29792 76701 29794
rect 74979 29736 74984 29792
rect 75040 29736 76640 29792
rect 76696 29736 76701 29792
rect 74979 29734 76701 29736
rect 74979 29731 75045 29734
rect 76635 29731 76701 29734
rect 52255 29658 52321 29661
rect 54463 29658 54529 29661
rect 52255 29656 54529 29658
rect 52255 29600 52260 29656
rect 52316 29600 54468 29656
rect 54524 29600 54529 29656
rect 52255 29598 54529 29600
rect 52255 29595 52321 29598
rect 54463 29595 54529 29598
rect 3642 29456 3962 29457
rect 3642 29392 3650 29456
rect 3714 29392 3730 29456
rect 3794 29392 3810 29456
rect 3874 29392 3890 29456
rect 3954 29392 3962 29456
rect 3642 29391 3962 29392
rect 8970 29456 9290 29457
rect 8970 29392 8978 29456
rect 9042 29392 9058 29456
rect 9122 29392 9138 29456
rect 9202 29392 9218 29456
rect 9282 29392 9290 29456
rect 8970 29391 9290 29392
rect 14298 29456 14618 29457
rect 14298 29392 14306 29456
rect 14370 29392 14386 29456
rect 14450 29392 14466 29456
rect 14530 29392 14546 29456
rect 14610 29392 14618 29456
rect 14298 29391 14618 29392
rect 19626 29456 19946 29457
rect 19626 29392 19634 29456
rect 19698 29392 19714 29456
rect 19778 29392 19794 29456
rect 19858 29392 19874 29456
rect 19938 29392 19946 29456
rect 19626 29391 19946 29392
rect 24954 29456 25274 29457
rect 24954 29392 24962 29456
rect 25026 29392 25042 29456
rect 25106 29392 25122 29456
rect 25186 29392 25202 29456
rect 25266 29392 25274 29456
rect 24954 29391 25274 29392
rect 30282 29456 30602 29457
rect 30282 29392 30290 29456
rect 30354 29392 30370 29456
rect 30434 29392 30450 29456
rect 30514 29392 30530 29456
rect 30594 29392 30602 29456
rect 30282 29391 30602 29392
rect 35610 29456 35930 29457
rect 35610 29392 35618 29456
rect 35682 29392 35698 29456
rect 35762 29392 35778 29456
rect 35842 29392 35858 29456
rect 35922 29392 35930 29456
rect 35610 29391 35930 29392
rect 40938 29456 41258 29457
rect 40938 29392 40946 29456
rect 41010 29392 41026 29456
rect 41090 29392 41106 29456
rect 41170 29392 41186 29456
rect 41250 29392 41258 29456
rect 40938 29391 41258 29392
rect 46266 29456 46586 29457
rect 46266 29392 46274 29456
rect 46338 29392 46354 29456
rect 46418 29392 46434 29456
rect 46498 29392 46514 29456
rect 46578 29392 46586 29456
rect 46266 29391 46586 29392
rect 51594 29456 51914 29457
rect 51594 29392 51602 29456
rect 51666 29392 51682 29456
rect 51746 29392 51762 29456
rect 51826 29392 51842 29456
rect 51906 29392 51914 29456
rect 51594 29391 51914 29392
rect 56922 29456 57242 29457
rect 56922 29392 56930 29456
rect 56994 29392 57010 29456
rect 57074 29392 57090 29456
rect 57154 29392 57170 29456
rect 57234 29392 57242 29456
rect 56922 29391 57242 29392
rect 62250 29456 62570 29457
rect 62250 29392 62258 29456
rect 62322 29392 62338 29456
rect 62402 29392 62418 29456
rect 62482 29392 62498 29456
rect 62562 29392 62570 29456
rect 62250 29391 62570 29392
rect 67578 29456 67898 29457
rect 67578 29392 67586 29456
rect 67650 29392 67666 29456
rect 67730 29392 67746 29456
rect 67810 29392 67826 29456
rect 67890 29392 67898 29456
rect 67578 29391 67898 29392
rect 72906 29456 73226 29457
rect 72906 29392 72914 29456
rect 72978 29392 72994 29456
rect 73058 29392 73074 29456
rect 73138 29392 73154 29456
rect 73218 29392 73226 29456
rect 72906 29391 73226 29392
rect 78234 29456 78554 29457
rect 78234 29392 78242 29456
rect 78306 29392 78322 29456
rect 78386 29392 78402 29456
rect 78466 29392 78482 29456
rect 78546 29392 78554 29456
rect 78234 29391 78554 29392
rect 83562 29456 83882 29457
rect 83562 29392 83570 29456
rect 83634 29392 83650 29456
rect 83714 29392 83730 29456
rect 83794 29392 83810 29456
rect 83874 29392 83882 29456
rect 83562 29391 83882 29392
rect 88890 29456 89210 29457
rect 88890 29392 88898 29456
rect 88962 29392 88978 29456
rect 89042 29392 89058 29456
rect 89122 29392 89138 29456
rect 89202 29392 89210 29456
rect 88890 29391 89210 29392
rect 60351 29250 60417 29253
rect 64491 29250 64557 29253
rect 60351 29248 64557 29250
rect 60351 29192 60356 29248
rect 60412 29192 64496 29248
rect 64552 29192 64557 29248
rect 60351 29190 64557 29192
rect 60351 29187 60417 29190
rect 64491 29187 64557 29190
rect 33211 29114 33277 29117
rect 37811 29114 37877 29117
rect 33211 29112 37877 29114
rect 33211 29056 33216 29112
rect 33272 29056 37816 29112
rect 37872 29056 37877 29112
rect 33211 29054 37877 29056
rect 33211 29051 33277 29054
rect 37811 29051 37877 29054
rect 38271 29114 38337 29117
rect 45999 29114 46065 29117
rect 38271 29112 46065 29114
rect 38271 29056 38276 29112
rect 38332 29056 46004 29112
rect 46060 29056 46065 29112
rect 38271 29054 46065 29056
rect 38271 29051 38337 29054
rect 45999 29051 46065 29054
rect 52623 29114 52689 29117
rect 56579 29114 56645 29117
rect 52623 29112 56645 29114
rect 52623 29056 52628 29112
rect 52684 29056 56584 29112
rect 56640 29056 56645 29112
rect 52623 29054 56645 29056
rect 52623 29051 52689 29054
rect 56579 29051 56645 29054
rect 6306 28912 6626 28913
rect 6306 28848 6314 28912
rect 6378 28848 6394 28912
rect 6458 28848 6474 28912
rect 6538 28848 6554 28912
rect 6618 28848 6626 28912
rect 6306 28847 6626 28848
rect 11634 28912 11954 28913
rect 11634 28848 11642 28912
rect 11706 28848 11722 28912
rect 11786 28848 11802 28912
rect 11866 28848 11882 28912
rect 11946 28848 11954 28912
rect 11634 28847 11954 28848
rect 16962 28912 17282 28913
rect 16962 28848 16970 28912
rect 17034 28848 17050 28912
rect 17114 28848 17130 28912
rect 17194 28848 17210 28912
rect 17274 28848 17282 28912
rect 16962 28847 17282 28848
rect 22290 28912 22610 28913
rect 22290 28848 22298 28912
rect 22362 28848 22378 28912
rect 22442 28848 22458 28912
rect 22522 28848 22538 28912
rect 22602 28848 22610 28912
rect 22290 28847 22610 28848
rect 27618 28912 27938 28913
rect 27618 28848 27626 28912
rect 27690 28848 27706 28912
rect 27770 28848 27786 28912
rect 27850 28848 27866 28912
rect 27930 28848 27938 28912
rect 27618 28847 27938 28848
rect 32946 28912 33266 28913
rect 32946 28848 32954 28912
rect 33018 28848 33034 28912
rect 33098 28848 33114 28912
rect 33178 28848 33194 28912
rect 33258 28848 33266 28912
rect 32946 28847 33266 28848
rect 38274 28912 38594 28913
rect 38274 28848 38282 28912
rect 38346 28848 38362 28912
rect 38426 28848 38442 28912
rect 38506 28848 38522 28912
rect 38586 28848 38594 28912
rect 38274 28847 38594 28848
rect 43602 28912 43922 28913
rect 43602 28848 43610 28912
rect 43674 28848 43690 28912
rect 43754 28848 43770 28912
rect 43834 28848 43850 28912
rect 43914 28848 43922 28912
rect 43602 28847 43922 28848
rect 48930 28912 49250 28913
rect 48930 28848 48938 28912
rect 49002 28848 49018 28912
rect 49082 28848 49098 28912
rect 49162 28848 49178 28912
rect 49242 28848 49250 28912
rect 48930 28847 49250 28848
rect 54258 28912 54578 28913
rect 54258 28848 54266 28912
rect 54330 28848 54346 28912
rect 54410 28848 54426 28912
rect 54490 28848 54506 28912
rect 54570 28848 54578 28912
rect 54258 28847 54578 28848
rect 59586 28912 59906 28913
rect 59586 28848 59594 28912
rect 59658 28848 59674 28912
rect 59738 28848 59754 28912
rect 59818 28848 59834 28912
rect 59898 28848 59906 28912
rect 59586 28847 59906 28848
rect 64914 28912 65234 28913
rect 64914 28848 64922 28912
rect 64986 28848 65002 28912
rect 65066 28848 65082 28912
rect 65146 28848 65162 28912
rect 65226 28848 65234 28912
rect 64914 28847 65234 28848
rect 70242 28912 70562 28913
rect 70242 28848 70250 28912
rect 70314 28848 70330 28912
rect 70394 28848 70410 28912
rect 70474 28848 70490 28912
rect 70554 28848 70562 28912
rect 70242 28847 70562 28848
rect 75570 28912 75890 28913
rect 75570 28848 75578 28912
rect 75642 28848 75658 28912
rect 75722 28848 75738 28912
rect 75802 28848 75818 28912
rect 75882 28848 75890 28912
rect 75570 28847 75890 28848
rect 80898 28912 81218 28913
rect 80898 28848 80906 28912
rect 80970 28848 80986 28912
rect 81050 28848 81066 28912
rect 81130 28848 81146 28912
rect 81210 28848 81218 28912
rect 80898 28847 81218 28848
rect 86226 28912 86546 28913
rect 86226 28848 86234 28912
rect 86298 28848 86314 28912
rect 86378 28848 86394 28912
rect 86458 28848 86474 28912
rect 86538 28848 86546 28912
rect 86226 28847 86546 28848
rect 91554 28912 91874 28913
rect 91554 28848 91562 28912
rect 91626 28848 91642 28912
rect 91706 28848 91722 28912
rect 91786 28848 91802 28912
rect 91866 28848 91874 28912
rect 91554 28847 91874 28848
rect 23827 28706 23893 28709
rect 24839 28706 24905 28709
rect 23827 28704 24905 28706
rect 23827 28648 23832 28704
rect 23888 28648 24844 28704
rect 24900 28648 24905 28704
rect 23827 28646 24905 28648
rect 23827 28643 23893 28646
rect 24839 28643 24905 28646
rect 25759 28706 25825 28709
rect 27967 28706 28033 28709
rect 25759 28704 28033 28706
rect 25759 28648 25764 28704
rect 25820 28648 27972 28704
rect 28028 28648 28033 28704
rect 25759 28646 28033 28648
rect 25759 28643 25825 28646
rect 27967 28643 28033 28646
rect 52071 28706 52137 28709
rect 52991 28706 53057 28709
rect 52071 28704 53057 28706
rect 52071 28648 52076 28704
rect 52132 28648 52996 28704
rect 53052 28648 53057 28704
rect 52071 28646 53057 28648
rect 52071 28643 52137 28646
rect 52991 28643 53057 28646
rect 22815 28570 22881 28573
rect 28519 28570 28585 28573
rect 22815 28568 28585 28570
rect 22815 28512 22820 28568
rect 22876 28512 28524 28568
rect 28580 28512 28585 28568
rect 22815 28510 28585 28512
rect 22815 28507 22881 28510
rect 28519 28507 28585 28510
rect 3642 28368 3962 28369
rect 3642 28304 3650 28368
rect 3714 28304 3730 28368
rect 3794 28304 3810 28368
rect 3874 28304 3890 28368
rect 3954 28304 3962 28368
rect 3642 28303 3962 28304
rect 8970 28368 9290 28369
rect 8970 28304 8978 28368
rect 9042 28304 9058 28368
rect 9122 28304 9138 28368
rect 9202 28304 9218 28368
rect 9282 28304 9290 28368
rect 8970 28303 9290 28304
rect 14298 28368 14618 28369
rect 14298 28304 14306 28368
rect 14370 28304 14386 28368
rect 14450 28304 14466 28368
rect 14530 28304 14546 28368
rect 14610 28304 14618 28368
rect 14298 28303 14618 28304
rect 19626 28368 19946 28369
rect 19626 28304 19634 28368
rect 19698 28304 19714 28368
rect 19778 28304 19794 28368
rect 19858 28304 19874 28368
rect 19938 28304 19946 28368
rect 19626 28303 19946 28304
rect 24954 28368 25274 28369
rect 24954 28304 24962 28368
rect 25026 28304 25042 28368
rect 25106 28304 25122 28368
rect 25186 28304 25202 28368
rect 25266 28304 25274 28368
rect 24954 28303 25274 28304
rect 30282 28368 30602 28369
rect 30282 28304 30290 28368
rect 30354 28304 30370 28368
rect 30434 28304 30450 28368
rect 30514 28304 30530 28368
rect 30594 28304 30602 28368
rect 30282 28303 30602 28304
rect 35610 28368 35930 28369
rect 35610 28304 35618 28368
rect 35682 28304 35698 28368
rect 35762 28304 35778 28368
rect 35842 28304 35858 28368
rect 35922 28304 35930 28368
rect 35610 28303 35930 28304
rect 40938 28368 41258 28369
rect 40938 28304 40946 28368
rect 41010 28304 41026 28368
rect 41090 28304 41106 28368
rect 41170 28304 41186 28368
rect 41250 28304 41258 28368
rect 40938 28303 41258 28304
rect 46266 28368 46586 28369
rect 46266 28304 46274 28368
rect 46338 28304 46354 28368
rect 46418 28304 46434 28368
rect 46498 28304 46514 28368
rect 46578 28304 46586 28368
rect 46266 28303 46586 28304
rect 51594 28368 51914 28369
rect 51594 28304 51602 28368
rect 51666 28304 51682 28368
rect 51746 28304 51762 28368
rect 51826 28304 51842 28368
rect 51906 28304 51914 28368
rect 51594 28303 51914 28304
rect 56922 28368 57242 28369
rect 56922 28304 56930 28368
rect 56994 28304 57010 28368
rect 57074 28304 57090 28368
rect 57154 28304 57170 28368
rect 57234 28304 57242 28368
rect 56922 28303 57242 28304
rect 62250 28368 62570 28369
rect 62250 28304 62258 28368
rect 62322 28304 62338 28368
rect 62402 28304 62418 28368
rect 62482 28304 62498 28368
rect 62562 28304 62570 28368
rect 62250 28303 62570 28304
rect 67578 28368 67898 28369
rect 67578 28304 67586 28368
rect 67650 28304 67666 28368
rect 67730 28304 67746 28368
rect 67810 28304 67826 28368
rect 67890 28304 67898 28368
rect 67578 28303 67898 28304
rect 72906 28368 73226 28369
rect 72906 28304 72914 28368
rect 72978 28304 72994 28368
rect 73058 28304 73074 28368
rect 73138 28304 73154 28368
rect 73218 28304 73226 28368
rect 72906 28303 73226 28304
rect 78234 28368 78554 28369
rect 78234 28304 78242 28368
rect 78306 28304 78322 28368
rect 78386 28304 78402 28368
rect 78466 28304 78482 28368
rect 78546 28304 78554 28368
rect 78234 28303 78554 28304
rect 83562 28368 83882 28369
rect 83562 28304 83570 28368
rect 83634 28304 83650 28368
rect 83714 28304 83730 28368
rect 83794 28304 83810 28368
rect 83874 28304 83882 28368
rect 83562 28303 83882 28304
rect 88890 28368 89210 28369
rect 88890 28304 88898 28368
rect 88962 28304 88978 28368
rect 89042 28304 89058 28368
rect 89122 28304 89138 28368
rect 89202 28304 89210 28368
rect 88890 28303 89210 28304
rect 12695 28162 12761 28165
rect 68171 28162 68237 28165
rect 12695 28160 68237 28162
rect 12695 28104 12700 28160
rect 12756 28104 68176 28160
rect 68232 28104 68237 28160
rect 12695 28102 68237 28104
rect 12695 28099 12761 28102
rect 68171 28099 68237 28102
rect 18859 28026 18925 28029
rect 24379 28026 24445 28029
rect 18859 28024 24445 28026
rect 18859 27968 18864 28024
rect 18920 27968 24384 28024
rect 24440 27968 24445 28024
rect 18859 27966 24445 27968
rect 18859 27963 18925 27966
rect 24379 27963 24445 27966
rect 30359 28026 30425 28029
rect 31371 28026 31437 28029
rect 36707 28026 36773 28029
rect 30359 28024 31437 28026
rect 30359 27968 30364 28024
rect 30420 27968 31376 28024
rect 31432 27968 31437 28024
rect 30359 27966 31437 27968
rect 30359 27963 30425 27966
rect 31371 27963 31437 27966
rect 31512 28024 36773 28026
rect 31512 27968 36712 28024
rect 36768 27968 36773 28024
rect 31512 27966 36773 27968
rect 31279 27890 31345 27893
rect 31512 27890 31572 27966
rect 36707 27963 36773 27966
rect 48207 28026 48273 28029
rect 51519 28026 51585 28029
rect 48207 28024 51585 28026
rect 48207 27968 48212 28024
rect 48268 27968 51524 28024
rect 51580 27968 51585 28024
rect 48207 27966 51585 27968
rect 48207 27963 48273 27966
rect 51519 27963 51585 27966
rect 31279 27888 31572 27890
rect 31279 27832 31284 27888
rect 31340 27832 31572 27888
rect 31279 27830 31572 27832
rect 50415 27890 50481 27893
rect 51151 27890 51217 27893
rect 54003 27890 54069 27893
rect 50415 27888 54069 27890
rect 50415 27832 50420 27888
rect 50476 27832 51156 27888
rect 51212 27832 54008 27888
rect 54064 27832 54069 27888
rect 50415 27830 54069 27832
rect 31279 27827 31345 27830
rect 50415 27827 50481 27830
rect 51151 27827 51217 27830
rect 54003 27827 54069 27830
rect 6306 27824 6626 27825
rect 6306 27760 6314 27824
rect 6378 27760 6394 27824
rect 6458 27760 6474 27824
rect 6538 27760 6554 27824
rect 6618 27760 6626 27824
rect 6306 27759 6626 27760
rect 11634 27824 11954 27825
rect 11634 27760 11642 27824
rect 11706 27760 11722 27824
rect 11786 27760 11802 27824
rect 11866 27760 11882 27824
rect 11946 27760 11954 27824
rect 11634 27759 11954 27760
rect 16962 27824 17282 27825
rect 16962 27760 16970 27824
rect 17034 27760 17050 27824
rect 17114 27760 17130 27824
rect 17194 27760 17210 27824
rect 17274 27760 17282 27824
rect 16962 27759 17282 27760
rect 22290 27824 22610 27825
rect 22290 27760 22298 27824
rect 22362 27760 22378 27824
rect 22442 27760 22458 27824
rect 22522 27760 22538 27824
rect 22602 27760 22610 27824
rect 22290 27759 22610 27760
rect 27618 27824 27938 27825
rect 27618 27760 27626 27824
rect 27690 27760 27706 27824
rect 27770 27760 27786 27824
rect 27850 27760 27866 27824
rect 27930 27760 27938 27824
rect 27618 27759 27938 27760
rect 32946 27824 33266 27825
rect 32946 27760 32954 27824
rect 33018 27760 33034 27824
rect 33098 27760 33114 27824
rect 33178 27760 33194 27824
rect 33258 27760 33266 27824
rect 32946 27759 33266 27760
rect 38274 27824 38594 27825
rect 38274 27760 38282 27824
rect 38346 27760 38362 27824
rect 38426 27760 38442 27824
rect 38506 27760 38522 27824
rect 38586 27760 38594 27824
rect 38274 27759 38594 27760
rect 43602 27824 43922 27825
rect 43602 27760 43610 27824
rect 43674 27760 43690 27824
rect 43754 27760 43770 27824
rect 43834 27760 43850 27824
rect 43914 27760 43922 27824
rect 43602 27759 43922 27760
rect 48930 27824 49250 27825
rect 48930 27760 48938 27824
rect 49002 27760 49018 27824
rect 49082 27760 49098 27824
rect 49162 27760 49178 27824
rect 49242 27760 49250 27824
rect 48930 27759 49250 27760
rect 54258 27824 54578 27825
rect 54258 27760 54266 27824
rect 54330 27760 54346 27824
rect 54410 27760 54426 27824
rect 54490 27760 54506 27824
rect 54570 27760 54578 27824
rect 54258 27759 54578 27760
rect 59586 27824 59906 27825
rect 59586 27760 59594 27824
rect 59658 27760 59674 27824
rect 59738 27760 59754 27824
rect 59818 27760 59834 27824
rect 59898 27760 59906 27824
rect 59586 27759 59906 27760
rect 64914 27824 65234 27825
rect 64914 27760 64922 27824
rect 64986 27760 65002 27824
rect 65066 27760 65082 27824
rect 65146 27760 65162 27824
rect 65226 27760 65234 27824
rect 64914 27759 65234 27760
rect 70242 27824 70562 27825
rect 70242 27760 70250 27824
rect 70314 27760 70330 27824
rect 70394 27760 70410 27824
rect 70474 27760 70490 27824
rect 70554 27760 70562 27824
rect 70242 27759 70562 27760
rect 75570 27824 75890 27825
rect 75570 27760 75578 27824
rect 75642 27760 75658 27824
rect 75722 27760 75738 27824
rect 75802 27760 75818 27824
rect 75882 27760 75890 27824
rect 75570 27759 75890 27760
rect 80898 27824 81218 27825
rect 80898 27760 80906 27824
rect 80970 27760 80986 27824
rect 81050 27760 81066 27824
rect 81130 27760 81146 27824
rect 81210 27760 81218 27824
rect 80898 27759 81218 27760
rect 86226 27824 86546 27825
rect 86226 27760 86234 27824
rect 86298 27760 86314 27824
rect 86378 27760 86394 27824
rect 86458 27760 86474 27824
rect 86538 27760 86546 27824
rect 86226 27759 86546 27760
rect 91554 27824 91874 27825
rect 91554 27760 91562 27824
rect 91626 27760 91642 27824
rect 91706 27760 91722 27824
rect 91786 27760 91802 27824
rect 91866 27760 91874 27824
rect 91554 27759 91874 27760
rect 29899 27754 29965 27757
rect 31463 27754 31529 27757
rect 29899 27752 31529 27754
rect 29899 27696 29904 27752
rect 29960 27696 31468 27752
rect 31524 27696 31529 27752
rect 29899 27694 31529 27696
rect 29899 27691 29965 27694
rect 31463 27691 31529 27694
rect 12603 27618 12669 27621
rect 17111 27618 17177 27621
rect 12603 27616 17177 27618
rect 12603 27560 12608 27616
rect 12664 27560 17116 27616
rect 17172 27560 17177 27616
rect 12603 27558 17177 27560
rect 12603 27555 12669 27558
rect 17111 27555 17177 27558
rect 29807 27618 29873 27621
rect 31187 27618 31253 27621
rect 29807 27616 31253 27618
rect 29807 27560 29812 27616
rect 29868 27560 31192 27616
rect 31248 27560 31253 27616
rect 29807 27558 31253 27560
rect 29807 27555 29873 27558
rect 31187 27555 31253 27558
rect 10119 27482 10185 27485
rect 16559 27482 16625 27485
rect 10119 27480 16625 27482
rect 10119 27424 10124 27480
rect 10180 27424 16564 27480
rect 16620 27424 16625 27480
rect 10119 27422 16625 27424
rect 10119 27419 10185 27422
rect 16559 27419 16625 27422
rect 23735 27482 23801 27485
rect 25207 27482 25273 27485
rect 23735 27480 25273 27482
rect 23735 27424 23740 27480
rect 23796 27424 25212 27480
rect 25268 27424 25273 27480
rect 23735 27422 25273 27424
rect 23735 27419 23801 27422
rect 25207 27419 25273 27422
rect 30175 27482 30241 27485
rect 31739 27482 31805 27485
rect 30175 27480 31805 27482
rect 30175 27424 30180 27480
rect 30236 27424 31744 27480
rect 31800 27424 31805 27480
rect 30175 27422 31805 27424
rect 30175 27419 30241 27422
rect 31739 27419 31805 27422
rect 48391 27482 48457 27485
rect 52899 27482 52965 27485
rect 48391 27480 52965 27482
rect 48391 27424 48396 27480
rect 48452 27424 52904 27480
rect 52960 27424 52965 27480
rect 48391 27422 52965 27424
rect 48391 27419 48457 27422
rect 52899 27419 52965 27422
rect 3642 27280 3962 27281
rect 3642 27216 3650 27280
rect 3714 27216 3730 27280
rect 3794 27216 3810 27280
rect 3874 27216 3890 27280
rect 3954 27216 3962 27280
rect 3642 27215 3962 27216
rect 8970 27280 9290 27281
rect 8970 27216 8978 27280
rect 9042 27216 9058 27280
rect 9122 27216 9138 27280
rect 9202 27216 9218 27280
rect 9282 27216 9290 27280
rect 8970 27215 9290 27216
rect 14298 27280 14618 27281
rect 14298 27216 14306 27280
rect 14370 27216 14386 27280
rect 14450 27216 14466 27280
rect 14530 27216 14546 27280
rect 14610 27216 14618 27280
rect 14298 27215 14618 27216
rect 19626 27280 19946 27281
rect 19626 27216 19634 27280
rect 19698 27216 19714 27280
rect 19778 27216 19794 27280
rect 19858 27216 19874 27280
rect 19938 27216 19946 27280
rect 19626 27215 19946 27216
rect 24954 27280 25274 27281
rect 24954 27216 24962 27280
rect 25026 27216 25042 27280
rect 25106 27216 25122 27280
rect 25186 27216 25202 27280
rect 25266 27216 25274 27280
rect 24954 27215 25274 27216
rect 30282 27280 30602 27281
rect 30282 27216 30290 27280
rect 30354 27216 30370 27280
rect 30434 27216 30450 27280
rect 30514 27216 30530 27280
rect 30594 27216 30602 27280
rect 30282 27215 30602 27216
rect 35610 27280 35930 27281
rect 35610 27216 35618 27280
rect 35682 27216 35698 27280
rect 35762 27216 35778 27280
rect 35842 27216 35858 27280
rect 35922 27216 35930 27280
rect 35610 27215 35930 27216
rect 40938 27280 41258 27281
rect 40938 27216 40946 27280
rect 41010 27216 41026 27280
rect 41090 27216 41106 27280
rect 41170 27216 41186 27280
rect 41250 27216 41258 27280
rect 40938 27215 41258 27216
rect 46266 27280 46586 27281
rect 46266 27216 46274 27280
rect 46338 27216 46354 27280
rect 46418 27216 46434 27280
rect 46498 27216 46514 27280
rect 46578 27216 46586 27280
rect 46266 27215 46586 27216
rect 51594 27280 51914 27281
rect 51594 27216 51602 27280
rect 51666 27216 51682 27280
rect 51746 27216 51762 27280
rect 51826 27216 51842 27280
rect 51906 27216 51914 27280
rect 51594 27215 51914 27216
rect 56922 27280 57242 27281
rect 56922 27216 56930 27280
rect 56994 27216 57010 27280
rect 57074 27216 57090 27280
rect 57154 27216 57170 27280
rect 57234 27216 57242 27280
rect 56922 27215 57242 27216
rect 62250 27280 62570 27281
rect 62250 27216 62258 27280
rect 62322 27216 62338 27280
rect 62402 27216 62418 27280
rect 62482 27216 62498 27280
rect 62562 27216 62570 27280
rect 62250 27215 62570 27216
rect 67578 27280 67898 27281
rect 67578 27216 67586 27280
rect 67650 27216 67666 27280
rect 67730 27216 67746 27280
rect 67810 27216 67826 27280
rect 67890 27216 67898 27280
rect 67578 27215 67898 27216
rect 72906 27280 73226 27281
rect 72906 27216 72914 27280
rect 72978 27216 72994 27280
rect 73058 27216 73074 27280
rect 73138 27216 73154 27280
rect 73218 27216 73226 27280
rect 72906 27215 73226 27216
rect 78234 27280 78554 27281
rect 78234 27216 78242 27280
rect 78306 27216 78322 27280
rect 78386 27216 78402 27280
rect 78466 27216 78482 27280
rect 78546 27216 78554 27280
rect 78234 27215 78554 27216
rect 83562 27280 83882 27281
rect 83562 27216 83570 27280
rect 83634 27216 83650 27280
rect 83714 27216 83730 27280
rect 83794 27216 83810 27280
rect 83874 27216 83882 27280
rect 83562 27215 83882 27216
rect 88890 27280 89210 27281
rect 88890 27216 88898 27280
rect 88962 27216 88978 27280
rect 89042 27216 89058 27280
rect 89122 27216 89138 27280
rect 89202 27216 89210 27280
rect 88890 27215 89210 27216
rect 29715 27074 29781 27077
rect 31647 27074 31713 27077
rect 29715 27072 31713 27074
rect 29715 27016 29720 27072
rect 29776 27016 31652 27072
rect 31708 27016 31713 27072
rect 29715 27014 31713 27016
rect 29715 27011 29781 27014
rect 31647 27011 31713 27014
rect 51059 27074 51125 27077
rect 52899 27074 52965 27077
rect 51059 27072 52965 27074
rect 51059 27016 51064 27072
rect 51120 27016 52904 27072
rect 52960 27016 52965 27072
rect 51059 27014 52965 27016
rect 51059 27011 51125 27014
rect 52899 27011 52965 27014
rect 29347 26938 29413 26941
rect 30359 26938 30425 26941
rect 29347 26936 30425 26938
rect 29347 26880 29352 26936
rect 29408 26880 30364 26936
rect 30420 26880 30425 26936
rect 29347 26878 30425 26880
rect 29347 26875 29413 26878
rect 30359 26875 30425 26878
rect 30727 26938 30793 26941
rect 31371 26938 31437 26941
rect 30727 26936 31437 26938
rect 30727 26880 30732 26936
rect 30788 26880 31376 26936
rect 31432 26880 31437 26936
rect 30727 26878 31437 26880
rect 30727 26875 30793 26878
rect 31371 26875 31437 26878
rect 6306 26736 6626 26737
rect 6306 26672 6314 26736
rect 6378 26672 6394 26736
rect 6458 26672 6474 26736
rect 6538 26672 6554 26736
rect 6618 26672 6626 26736
rect 6306 26671 6626 26672
rect 11634 26736 11954 26737
rect 11634 26672 11642 26736
rect 11706 26672 11722 26736
rect 11786 26672 11802 26736
rect 11866 26672 11882 26736
rect 11946 26672 11954 26736
rect 11634 26671 11954 26672
rect 16962 26736 17282 26737
rect 16962 26672 16970 26736
rect 17034 26672 17050 26736
rect 17114 26672 17130 26736
rect 17194 26672 17210 26736
rect 17274 26672 17282 26736
rect 16962 26671 17282 26672
rect 22290 26736 22610 26737
rect 22290 26672 22298 26736
rect 22362 26672 22378 26736
rect 22442 26672 22458 26736
rect 22522 26672 22538 26736
rect 22602 26672 22610 26736
rect 22290 26671 22610 26672
rect 27618 26736 27938 26737
rect 27618 26672 27626 26736
rect 27690 26672 27706 26736
rect 27770 26672 27786 26736
rect 27850 26672 27866 26736
rect 27930 26672 27938 26736
rect 27618 26671 27938 26672
rect 32946 26736 33266 26737
rect 32946 26672 32954 26736
rect 33018 26672 33034 26736
rect 33098 26672 33114 26736
rect 33178 26672 33194 26736
rect 33258 26672 33266 26736
rect 32946 26671 33266 26672
rect 38274 26736 38594 26737
rect 38274 26672 38282 26736
rect 38346 26672 38362 26736
rect 38426 26672 38442 26736
rect 38506 26672 38522 26736
rect 38586 26672 38594 26736
rect 38274 26671 38594 26672
rect 43602 26736 43922 26737
rect 43602 26672 43610 26736
rect 43674 26672 43690 26736
rect 43754 26672 43770 26736
rect 43834 26672 43850 26736
rect 43914 26672 43922 26736
rect 43602 26671 43922 26672
rect 48930 26736 49250 26737
rect 48930 26672 48938 26736
rect 49002 26672 49018 26736
rect 49082 26672 49098 26736
rect 49162 26672 49178 26736
rect 49242 26672 49250 26736
rect 48930 26671 49250 26672
rect 54258 26736 54578 26737
rect 54258 26672 54266 26736
rect 54330 26672 54346 26736
rect 54410 26672 54426 26736
rect 54490 26672 54506 26736
rect 54570 26672 54578 26736
rect 54258 26671 54578 26672
rect 59586 26736 59906 26737
rect 59586 26672 59594 26736
rect 59658 26672 59674 26736
rect 59738 26672 59754 26736
rect 59818 26672 59834 26736
rect 59898 26672 59906 26736
rect 59586 26671 59906 26672
rect 64914 26736 65234 26737
rect 64914 26672 64922 26736
rect 64986 26672 65002 26736
rect 65066 26672 65082 26736
rect 65146 26672 65162 26736
rect 65226 26672 65234 26736
rect 64914 26671 65234 26672
rect 70242 26736 70562 26737
rect 70242 26672 70250 26736
rect 70314 26672 70330 26736
rect 70394 26672 70410 26736
rect 70474 26672 70490 26736
rect 70554 26672 70562 26736
rect 70242 26671 70562 26672
rect 75570 26736 75890 26737
rect 75570 26672 75578 26736
rect 75642 26672 75658 26736
rect 75722 26672 75738 26736
rect 75802 26672 75818 26736
rect 75882 26672 75890 26736
rect 75570 26671 75890 26672
rect 80898 26736 81218 26737
rect 80898 26672 80906 26736
rect 80970 26672 80986 26736
rect 81050 26672 81066 26736
rect 81130 26672 81146 26736
rect 81210 26672 81218 26736
rect 80898 26671 81218 26672
rect 86226 26736 86546 26737
rect 86226 26672 86234 26736
rect 86298 26672 86314 26736
rect 86378 26672 86394 26736
rect 86458 26672 86474 26736
rect 86538 26672 86546 26736
rect 86226 26671 86546 26672
rect 91554 26736 91874 26737
rect 91554 26672 91562 26736
rect 91626 26672 91642 26736
rect 91706 26672 91722 26736
rect 91786 26672 91802 26736
rect 91866 26672 91874 26736
rect 91554 26671 91874 26672
rect 3642 26192 3962 26193
rect 3642 26128 3650 26192
rect 3714 26128 3730 26192
rect 3794 26128 3810 26192
rect 3874 26128 3890 26192
rect 3954 26128 3962 26192
rect 3642 26127 3962 26128
rect 35610 26192 35930 26193
rect 35610 26128 35618 26192
rect 35682 26128 35698 26192
rect 35762 26128 35778 26192
rect 35842 26128 35858 26192
rect 35922 26128 35930 26192
rect 35610 26127 35930 26128
rect 40938 26192 41258 26193
rect 40938 26128 40946 26192
rect 41010 26128 41026 26192
rect 41090 26128 41106 26192
rect 41170 26128 41186 26192
rect 41250 26128 41258 26192
rect 40938 26127 41258 26128
rect 6306 25648 6626 25649
rect 6306 25584 6314 25648
rect 6378 25584 6394 25648
rect 6458 25584 6474 25648
rect 6538 25584 6554 25648
rect 6618 25584 6626 25648
rect 6306 25583 6626 25584
rect 38274 25648 38594 25649
rect 38274 25584 38282 25648
rect 38346 25584 38362 25648
rect 38426 25584 38442 25648
rect 38506 25584 38522 25648
rect 38586 25584 38594 25648
rect 38274 25583 38594 25584
rect 3642 25104 3962 25105
rect 3642 25040 3650 25104
rect 3714 25040 3730 25104
rect 3794 25040 3810 25104
rect 3874 25040 3890 25104
rect 3954 25040 3962 25104
rect 3642 25039 3962 25040
rect 35610 25104 35930 25105
rect 35610 25040 35618 25104
rect 35682 25040 35698 25104
rect 35762 25040 35778 25104
rect 35842 25040 35858 25104
rect 35922 25040 35930 25104
rect 35610 25039 35930 25040
rect 40938 25104 41258 25105
rect 40938 25040 40946 25104
rect 41010 25040 41026 25104
rect 41090 25040 41106 25104
rect 41170 25040 41186 25104
rect 41250 25040 41258 25104
rect 40938 25039 41258 25040
rect 6306 24560 6626 24561
rect 6306 24496 6314 24560
rect 6378 24496 6394 24560
rect 6458 24496 6474 24560
rect 6538 24496 6554 24560
rect 6618 24496 6626 24560
rect 6306 24495 6626 24496
rect 38274 24560 38594 24561
rect 38274 24496 38282 24560
rect 38346 24496 38362 24560
rect 38426 24496 38442 24560
rect 38506 24496 38522 24560
rect 38586 24496 38594 24560
rect 38274 24495 38594 24496
rect 3642 24016 3962 24017
rect 3642 23952 3650 24016
rect 3714 23952 3730 24016
rect 3794 23952 3810 24016
rect 3874 23952 3890 24016
rect 3954 23952 3962 24016
rect 3642 23951 3962 23952
rect 35610 24016 35930 24017
rect 35610 23952 35618 24016
rect 35682 23952 35698 24016
rect 35762 23952 35778 24016
rect 35842 23952 35858 24016
rect 35922 23952 35930 24016
rect 35610 23951 35930 23952
rect 40938 24016 41258 24017
rect 40938 23952 40946 24016
rect 41010 23952 41026 24016
rect 41090 23952 41106 24016
rect 41170 23952 41186 24016
rect 41250 23952 41258 24016
rect 40938 23951 41258 23952
rect 46091 23606 46157 23609
rect 46091 23604 46262 23606
rect 46091 23548 46096 23604
rect 46152 23548 46262 23604
rect 46091 23546 46262 23548
rect 46091 23543 46157 23546
rect 34315 23538 34381 23541
rect 31174 23536 34381 23538
rect 31174 23480 34320 23536
rect 34376 23480 34381 23536
rect 31174 23478 34381 23480
rect 34315 23475 34381 23478
rect 68355 23538 68421 23541
rect 68355 23536 70734 23538
rect 68355 23480 68360 23536
rect 68416 23480 70734 23536
rect 68355 23478 70734 23480
rect 68355 23475 68421 23478
rect 6306 23472 6626 23473
rect 6306 23408 6314 23472
rect 6378 23408 6394 23472
rect 6458 23408 6474 23472
rect 6538 23408 6554 23472
rect 6618 23408 6626 23472
rect 6306 23407 6626 23408
rect 38274 23472 38594 23473
rect 38274 23408 38282 23472
rect 38346 23408 38362 23472
rect 38426 23408 38442 23472
rect 38506 23408 38522 23472
rect 38586 23408 38594 23472
rect 38274 23407 38594 23408
rect 31371 23062 31437 23065
rect 31174 23060 31437 23062
rect 31174 23004 31376 23060
rect 31432 23004 31437 23060
rect 31174 23002 31437 23004
rect 31371 22999 31437 23002
rect 43515 22994 43581 22997
rect 45680 22994 46262 23006
rect 43515 22992 46262 22994
rect 43515 22936 43520 22992
rect 43576 22946 46262 22992
rect 70011 22994 70077 22997
rect 70011 22992 70734 22994
rect 43576 22936 45740 22946
rect 43515 22934 45740 22936
rect 70011 22936 70016 22992
rect 70072 22936 70734 22992
rect 70011 22934 70734 22936
rect 43515 22931 43581 22934
rect 70011 22931 70077 22934
rect 3642 22928 3962 22929
rect 3642 22864 3650 22928
rect 3714 22864 3730 22928
rect 3794 22864 3810 22928
rect 3874 22864 3890 22928
rect 3954 22864 3962 22928
rect 3642 22863 3962 22864
rect 35610 22928 35930 22929
rect 35610 22864 35618 22928
rect 35682 22864 35698 22928
rect 35762 22864 35778 22928
rect 35842 22864 35858 22928
rect 35922 22864 35930 22928
rect 35610 22863 35930 22864
rect 40938 22928 41258 22929
rect 40938 22864 40946 22928
rect 41010 22864 41026 22928
rect 41090 22864 41106 22928
rect 41170 22864 41186 22928
rect 41250 22864 41258 22928
rect 40938 22863 41258 22864
rect 3352 22660 3358 22724
rect 3422 22722 3428 22724
rect 3495 22722 3561 22725
rect 3422 22720 3561 22722
rect 3422 22664 3500 22720
rect 3556 22664 3561 22720
rect 3422 22662 3561 22664
rect 3422 22660 3428 22662
rect 3495 22659 3561 22662
rect 70195 22518 70261 22521
rect 70195 22516 70734 22518
rect 31504 22450 31510 22452
rect 31174 22390 31510 22450
rect 31504 22388 31510 22390
rect 31574 22450 31580 22452
rect 34775 22450 34841 22453
rect 31574 22448 34841 22450
rect 31574 22392 34780 22448
rect 34836 22392 34841 22448
rect 31574 22390 34841 22392
rect 31574 22388 31580 22390
rect 34775 22387 34841 22390
rect 43055 22450 43121 22453
rect 45680 22450 46262 22462
rect 70195 22460 70200 22516
rect 70256 22460 70734 22516
rect 70195 22458 70734 22460
rect 70195 22455 70261 22458
rect 43055 22448 46262 22450
rect 43055 22392 43060 22448
rect 43116 22402 46262 22448
rect 43116 22392 45740 22402
rect 43055 22390 45740 22392
rect 43055 22387 43121 22390
rect 6306 22384 6626 22385
rect 6306 22320 6314 22384
rect 6378 22320 6394 22384
rect 6458 22320 6474 22384
rect 6538 22320 6554 22384
rect 6618 22320 6626 22384
rect 6306 22319 6626 22320
rect 38274 22384 38594 22385
rect 38274 22320 38282 22384
rect 38346 22320 38362 22384
rect 38426 22320 38442 22384
rect 38506 22320 38522 22384
rect 38586 22320 38594 22384
rect 38274 22319 38594 22320
rect 3642 21840 3962 21841
rect 3642 21776 3650 21840
rect 3714 21776 3730 21840
rect 3794 21776 3810 21840
rect 3874 21776 3890 21840
rect 3954 21776 3962 21840
rect 3642 21775 3962 21776
rect 35610 21840 35930 21841
rect 35610 21776 35618 21840
rect 35682 21776 35698 21840
rect 35762 21776 35778 21840
rect 35842 21776 35858 21840
rect 35922 21776 35930 21840
rect 35610 21775 35930 21776
rect 40938 21840 41258 21841
rect 40938 21776 40946 21840
rect 41010 21776 41026 21840
rect 41090 21776 41106 21840
rect 41170 21776 41186 21840
rect 41250 21776 41258 21840
rect 40938 21775 41258 21776
rect 36983 21498 37049 21501
rect 37944 21498 37950 21500
rect 36983 21496 37950 21498
rect 36983 21440 36988 21496
rect 37044 21440 37950 21496
rect 36983 21438 37950 21440
rect 36983 21435 37049 21438
rect 37944 21436 37950 21438
rect 38014 21436 38020 21500
rect 33947 21362 34013 21365
rect 34775 21362 34841 21365
rect 31174 21360 34841 21362
rect 31174 21304 33952 21360
rect 34008 21304 34780 21360
rect 34836 21304 34841 21360
rect 31174 21302 34841 21304
rect 33947 21299 34013 21302
rect 34775 21299 34841 21302
rect 43055 21362 43121 21365
rect 45680 21362 46262 21374
rect 43055 21360 46262 21362
rect 43055 21304 43060 21360
rect 43116 21314 46262 21360
rect 67159 21362 67225 21365
rect 67159 21360 70734 21362
rect 43116 21304 45740 21314
rect 43055 21302 45740 21304
rect 67159 21304 67164 21360
rect 67220 21304 70734 21360
rect 67159 21302 70734 21304
rect 43055 21299 43121 21302
rect 67159 21299 67225 21302
rect 6306 21296 6626 21297
rect 6306 21232 6314 21296
rect 6378 21232 6394 21296
rect 6458 21232 6474 21296
rect 6538 21232 6554 21296
rect 6618 21232 6626 21296
rect 6306 21231 6626 21232
rect 38274 21296 38594 21297
rect 38274 21232 38282 21296
rect 38346 21232 38362 21296
rect 38426 21232 38442 21296
rect 38506 21232 38522 21296
rect 38586 21232 38594 21296
rect 38274 21231 38594 21232
rect 3642 20752 3962 20753
rect 3642 20688 3650 20752
rect 3714 20688 3730 20752
rect 3794 20688 3810 20752
rect 3874 20688 3890 20752
rect 3954 20688 3962 20752
rect 3642 20687 3962 20688
rect 35610 20752 35930 20753
rect 35610 20688 35618 20752
rect 35682 20688 35698 20752
rect 35762 20688 35778 20752
rect 35842 20688 35858 20752
rect 35922 20688 35930 20752
rect 35610 20687 35930 20688
rect 40938 20752 41258 20753
rect 40938 20688 40946 20752
rect 41010 20688 41026 20752
rect 41090 20688 41106 20752
rect 41170 20688 41186 20752
rect 41250 20688 41258 20752
rect 40938 20687 41258 20688
rect 66832 20620 66838 20684
rect 66902 20682 66908 20684
rect 67067 20682 67133 20685
rect 66902 20680 67133 20682
rect 66902 20624 67072 20680
rect 67128 20624 67133 20680
rect 66902 20622 67133 20624
rect 66902 20620 66908 20622
rect 67067 20619 67133 20622
rect 31504 20274 31510 20276
rect 31174 20214 31510 20274
rect 31504 20212 31510 20214
rect 31574 20274 31580 20276
rect 34407 20274 34473 20277
rect 31574 20272 34473 20274
rect 31574 20216 34412 20272
rect 34468 20216 34473 20272
rect 31574 20214 34473 20216
rect 31574 20212 31580 20214
rect 34407 20211 34473 20214
rect 43055 20274 43121 20277
rect 45680 20274 46262 20286
rect 43055 20272 46262 20274
rect 43055 20216 43060 20272
rect 43116 20226 46262 20272
rect 68171 20274 68237 20277
rect 68171 20272 70734 20274
rect 43116 20216 45740 20226
rect 43055 20214 45740 20216
rect 68171 20216 68176 20272
rect 68232 20216 70734 20272
rect 68171 20214 70734 20216
rect 43055 20211 43121 20214
rect 68171 20211 68237 20214
rect 6306 20208 6626 20209
rect 6306 20144 6314 20208
rect 6378 20144 6394 20208
rect 6458 20144 6474 20208
rect 6538 20144 6554 20208
rect 6618 20144 6626 20208
rect 6306 20143 6626 20144
rect 38274 20208 38594 20209
rect 38274 20144 38282 20208
rect 38346 20144 38362 20208
rect 38426 20144 38442 20208
rect 38506 20144 38522 20208
rect 38586 20144 38594 20208
rect 38274 20143 38594 20144
rect 6807 20004 6873 20005
rect 6807 20002 6854 20004
rect 6762 20000 6854 20002
rect 6762 19944 6812 20000
rect 6762 19942 6854 19944
rect 6807 19940 6854 19942
rect 6918 19940 6924 20004
rect 41491 20002 41557 20005
rect 41624 20002 41630 20004
rect 41491 20000 41630 20002
rect 41491 19944 41496 20000
rect 41552 19944 41630 20000
rect 41491 19942 41630 19944
rect 6807 19939 6873 19940
rect 41491 19939 41557 19942
rect 41624 19940 41630 19942
rect 41694 19940 41700 20004
rect 67016 19940 67022 20004
rect 67086 20002 67092 20004
rect 67159 20002 67225 20005
rect 67086 20000 67225 20002
rect 67086 19944 67164 20000
rect 67220 19944 67225 20000
rect 67086 19942 67225 19944
rect 67086 19940 67092 19942
rect 67159 19939 67225 19942
rect 3642 19664 3962 19665
rect 3642 19600 3650 19664
rect 3714 19600 3730 19664
rect 3794 19600 3810 19664
rect 3874 19600 3890 19664
rect 3954 19600 3962 19664
rect 3642 19599 3962 19600
rect 35610 19664 35930 19665
rect 35610 19600 35618 19664
rect 35682 19600 35698 19664
rect 35762 19600 35778 19664
rect 35842 19600 35858 19664
rect 35922 19600 35930 19664
rect 35610 19599 35930 19600
rect 40938 19664 41258 19665
rect 40938 19600 40946 19664
rect 41010 19600 41026 19664
rect 41090 19600 41106 19664
rect 41170 19600 41186 19664
rect 41250 19600 41258 19664
rect 40938 19599 41258 19600
rect 4139 19322 4205 19325
rect 4272 19322 4278 19324
rect 4139 19320 4278 19322
rect 4139 19264 4144 19320
rect 4200 19264 4278 19320
rect 4139 19262 4278 19264
rect 4139 19259 4205 19262
rect 4272 19260 4278 19262
rect 4342 19260 4348 19324
rect 31504 19186 31510 19188
rect 31174 19126 31510 19186
rect 31504 19124 31510 19126
rect 31574 19186 31580 19188
rect 34407 19186 34473 19189
rect 31574 19184 34473 19186
rect 31574 19128 34412 19184
rect 34468 19128 34473 19184
rect 31574 19126 34473 19128
rect 31574 19124 31580 19126
rect 34407 19123 34473 19126
rect 42319 19186 42385 19189
rect 45680 19186 46262 19198
rect 42319 19184 46262 19186
rect 42319 19128 42324 19184
rect 42380 19138 46262 19184
rect 68263 19186 68329 19189
rect 68263 19184 70734 19186
rect 42380 19128 45740 19138
rect 42319 19126 45740 19128
rect 68263 19128 68268 19184
rect 68324 19128 70734 19184
rect 68263 19126 70734 19128
rect 42319 19123 42385 19126
rect 68263 19123 68329 19126
rect 6306 19120 6626 19121
rect 6306 19056 6314 19120
rect 6378 19056 6394 19120
rect 6458 19056 6474 19120
rect 6538 19056 6554 19120
rect 6618 19056 6626 19120
rect 6306 19055 6626 19056
rect 38274 19120 38594 19121
rect 38274 19056 38282 19120
rect 38346 19056 38362 19120
rect 38426 19056 38442 19120
rect 38506 19056 38522 19120
rect 38586 19056 38594 19120
rect 38274 19055 38594 19056
rect 3642 18576 3962 18577
rect 3642 18512 3650 18576
rect 3714 18512 3730 18576
rect 3794 18512 3810 18576
rect 3874 18512 3890 18576
rect 3954 18512 3962 18576
rect 3642 18511 3962 18512
rect 35610 18576 35930 18577
rect 35610 18512 35618 18576
rect 35682 18512 35698 18576
rect 35762 18512 35778 18576
rect 35842 18512 35858 18576
rect 35922 18512 35930 18576
rect 35610 18511 35930 18512
rect 40938 18576 41258 18577
rect 40938 18512 40946 18576
rect 41010 18512 41026 18576
rect 41090 18512 41106 18576
rect 41170 18512 41186 18576
rect 41250 18512 41258 18576
rect 40938 18511 41258 18512
rect 68263 18506 68329 18509
rect 70379 18506 70445 18509
rect 68263 18504 70445 18506
rect 68263 18448 68268 18504
rect 68324 18448 70384 18504
rect 70440 18448 70445 18504
rect 68263 18446 70445 18448
rect 68263 18443 68329 18446
rect 70379 18443 70445 18446
rect 31504 18098 31510 18100
rect 31174 18038 31510 18098
rect 31504 18036 31510 18038
rect 31574 18098 31580 18100
rect 34407 18098 34473 18101
rect 31574 18096 34473 18098
rect 31574 18040 34412 18096
rect 34468 18040 34473 18096
rect 31574 18038 34473 18040
rect 31574 18036 31580 18038
rect 34407 18035 34473 18038
rect 43515 18098 43581 18101
rect 45680 18098 46262 18110
rect 43515 18096 46262 18098
rect 43515 18040 43520 18096
rect 43576 18050 46262 18096
rect 67067 18098 67133 18101
rect 67067 18096 70734 18098
rect 43576 18040 45740 18050
rect 43515 18038 45740 18040
rect 67067 18040 67072 18096
rect 67128 18040 70734 18096
rect 67067 18038 70734 18040
rect 43515 18035 43581 18038
rect 67067 18035 67133 18038
rect 6306 18032 6626 18033
rect 6306 17968 6314 18032
rect 6378 17968 6394 18032
rect 6458 17968 6474 18032
rect 6538 17968 6554 18032
rect 6618 17968 6626 18032
rect 6306 17967 6626 17968
rect 38274 18032 38594 18033
rect 38274 17968 38282 18032
rect 38346 17968 38362 18032
rect 38426 17968 38442 18032
rect 38506 17968 38522 18032
rect 38586 17968 38594 18032
rect 38274 17967 38594 17968
rect 42043 17964 42109 17965
rect 41992 17900 41998 17964
rect 42062 17962 42109 17964
rect 42062 17960 42154 17962
rect 42104 17904 42154 17960
rect 42062 17902 42154 17904
rect 42062 17900 42109 17902
rect 67752 17900 67758 17964
rect 67822 17962 67828 17964
rect 68263 17962 68329 17965
rect 67822 17960 68329 17962
rect 67822 17904 68268 17960
rect 68324 17904 68329 17960
rect 67822 17902 68329 17904
rect 67822 17900 67828 17902
rect 42043 17899 42109 17900
rect 68263 17899 68329 17902
rect 7267 17554 7333 17557
rect 7400 17554 7406 17556
rect 7267 17552 7406 17554
rect 7267 17496 7272 17552
rect 7328 17496 7406 17552
rect 7267 17494 7406 17496
rect 7267 17491 7333 17494
rect 7400 17492 7406 17494
rect 7470 17492 7476 17556
rect 3642 17488 3962 17489
rect 3642 17424 3650 17488
rect 3714 17424 3730 17488
rect 3794 17424 3810 17488
rect 3874 17424 3890 17488
rect 3954 17424 3962 17488
rect 3642 17423 3962 17424
rect 35610 17488 35930 17489
rect 35610 17424 35618 17488
rect 35682 17424 35698 17488
rect 35762 17424 35778 17488
rect 35842 17424 35858 17488
rect 35922 17424 35930 17488
rect 35610 17423 35930 17424
rect 40938 17488 41258 17489
rect 40938 17424 40946 17488
rect 41010 17424 41026 17488
rect 41090 17424 41106 17488
rect 41170 17424 41186 17488
rect 41250 17424 41258 17488
rect 40938 17423 41258 17424
rect 5059 17282 5125 17285
rect 5192 17282 5198 17284
rect 5059 17280 5198 17282
rect 5059 17224 5064 17280
rect 5120 17224 5198 17280
rect 5059 17222 5198 17224
rect 5059 17219 5125 17222
rect 5192 17220 5198 17222
rect 5262 17220 5268 17284
rect 38823 17146 38889 17149
rect 40755 17146 40821 17149
rect 38823 17144 40821 17146
rect 38823 17088 38828 17144
rect 38884 17088 40760 17144
rect 40816 17088 40821 17144
rect 38823 17086 40821 17088
rect 38823 17083 38889 17086
rect 40755 17083 40821 17086
rect 70471 17078 70537 17081
rect 70471 17076 70734 17078
rect 31504 17010 31510 17012
rect 31174 16950 31510 17010
rect 31504 16948 31510 16950
rect 31574 17010 31580 17012
rect 34407 17010 34473 17013
rect 31574 17008 34473 17010
rect 31574 16952 34412 17008
rect 34468 16952 34473 17008
rect 31574 16950 34473 16952
rect 31574 16948 31580 16950
rect 34407 16947 34473 16950
rect 43331 17010 43397 17013
rect 45680 17010 46262 17022
rect 70471 17020 70476 17076
rect 70532 17020 70734 17076
rect 70471 17018 70734 17020
rect 70471 17015 70537 17018
rect 43331 17008 46262 17010
rect 43331 16952 43336 17008
rect 43392 16962 46262 17008
rect 43392 16952 45740 16962
rect 43331 16950 45740 16952
rect 43331 16947 43397 16950
rect 6306 16944 6626 16945
rect 6306 16880 6314 16944
rect 6378 16880 6394 16944
rect 6458 16880 6474 16944
rect 6538 16880 6554 16944
rect 6618 16880 6626 16944
rect 6306 16879 6626 16880
rect 38274 16944 38594 16945
rect 38274 16880 38282 16944
rect 38346 16880 38362 16944
rect 38426 16880 38442 16944
rect 38506 16880 38522 16944
rect 38586 16880 38594 16944
rect 38274 16879 38594 16880
rect 5703 16604 5769 16605
rect 36339 16604 36405 16605
rect 5703 16602 5750 16604
rect 5658 16600 5750 16602
rect 5658 16544 5708 16600
rect 5658 16542 5750 16544
rect 5703 16540 5750 16542
rect 5814 16540 5820 16604
rect 36288 16540 36294 16604
rect 36358 16602 36405 16604
rect 41675 16602 41741 16605
rect 68355 16604 68421 16605
rect 41808 16602 41814 16604
rect 36358 16600 36450 16602
rect 36400 16544 36450 16600
rect 36358 16542 36450 16544
rect 41675 16600 41814 16602
rect 41675 16544 41680 16600
rect 41736 16544 41814 16600
rect 41675 16542 41814 16544
rect 36358 16540 36405 16542
rect 5703 16539 5769 16540
rect 36339 16539 36405 16540
rect 41675 16539 41741 16542
rect 41808 16540 41814 16542
rect 41878 16540 41884 16604
rect 68304 16602 68310 16604
rect 68264 16542 68310 16602
rect 68374 16600 68421 16604
rect 68416 16544 68421 16600
rect 68304 16540 68310 16542
rect 68374 16540 68421 16544
rect 68355 16539 68421 16540
rect 3642 16400 3962 16401
rect 3642 16336 3650 16400
rect 3714 16336 3730 16400
rect 3794 16336 3810 16400
rect 3874 16336 3890 16400
rect 3954 16336 3962 16400
rect 3642 16335 3962 16336
rect 35610 16400 35930 16401
rect 35610 16336 35618 16400
rect 35682 16336 35698 16400
rect 35762 16336 35778 16400
rect 35842 16336 35858 16400
rect 35922 16336 35930 16400
rect 35610 16335 35930 16336
rect 40938 16400 41258 16401
rect 40938 16336 40946 16400
rect 41010 16336 41026 16400
rect 41090 16336 41106 16400
rect 41170 16336 41186 16400
rect 41250 16336 41258 16400
rect 40938 16335 41258 16336
rect 6306 15856 6626 15857
rect 6306 15792 6314 15856
rect 6378 15792 6394 15856
rect 6458 15792 6474 15856
rect 6538 15792 6554 15856
rect 6618 15792 6626 15856
rect 6306 15791 6626 15792
rect 38274 15856 38594 15857
rect 38274 15792 38282 15856
rect 38346 15792 38362 15856
rect 38426 15792 38442 15856
rect 38506 15792 38522 15856
rect 38586 15792 38594 15856
rect 38274 15791 38594 15792
rect 3642 15312 3962 15313
rect 3642 15248 3650 15312
rect 3714 15248 3730 15312
rect 3794 15248 3810 15312
rect 3874 15248 3890 15312
rect 3954 15248 3962 15312
rect 3642 15247 3962 15248
rect 35610 15312 35930 15313
rect 35610 15248 35618 15312
rect 35682 15248 35698 15312
rect 35762 15248 35778 15312
rect 35842 15248 35858 15312
rect 35922 15248 35930 15312
rect 35610 15247 35930 15248
rect 40938 15312 41258 15313
rect 40938 15248 40946 15312
rect 41010 15248 41026 15312
rect 41090 15248 41106 15312
rect 41170 15248 41186 15312
rect 41250 15248 41258 15312
rect 40938 15247 41258 15248
rect 6991 15242 7057 15245
rect 7216 15242 7222 15244
rect 6991 15240 7222 15242
rect 6991 15184 6996 15240
rect 7052 15184 7222 15240
rect 6991 15182 7222 15184
rect 6991 15179 7057 15182
rect 7216 15180 7222 15182
rect 7286 15180 7292 15244
rect 70471 14902 70537 14905
rect 70471 14900 70734 14902
rect 31504 14834 31510 14836
rect 31174 14774 31510 14834
rect 31504 14772 31510 14774
rect 31574 14834 31580 14836
rect 34407 14834 34473 14837
rect 31574 14832 34473 14834
rect 31574 14776 34412 14832
rect 34468 14776 34473 14832
rect 31574 14774 34473 14776
rect 31574 14772 31580 14774
rect 34407 14771 34473 14774
rect 43515 14834 43581 14837
rect 45680 14834 46262 14846
rect 70471 14844 70476 14900
rect 70532 14844 70734 14900
rect 70471 14842 70734 14844
rect 70471 14839 70537 14842
rect 43515 14832 46262 14834
rect 43515 14776 43520 14832
rect 43576 14786 46262 14832
rect 43576 14776 45740 14786
rect 43515 14774 45740 14776
rect 43515 14771 43581 14774
rect 6306 14768 6626 14769
rect 6306 14704 6314 14768
rect 6378 14704 6394 14768
rect 6458 14704 6474 14768
rect 6538 14704 6554 14768
rect 6618 14704 6626 14768
rect 6306 14703 6626 14704
rect 38274 14768 38594 14769
rect 38274 14704 38282 14768
rect 38346 14704 38362 14768
rect 38426 14704 38442 14768
rect 38506 14704 38522 14768
rect 38586 14704 38594 14768
rect 38274 14703 38594 14704
rect 7359 14564 7425 14565
rect 7359 14562 7406 14564
rect 7314 14560 7406 14562
rect 7314 14504 7364 14560
rect 7314 14502 7406 14504
rect 7359 14500 7406 14502
rect 7470 14500 7476 14564
rect 7359 14499 7425 14500
rect 3642 14224 3962 14225
rect 3642 14160 3650 14224
rect 3714 14160 3730 14224
rect 3794 14160 3810 14224
rect 3874 14160 3890 14224
rect 3954 14160 3962 14224
rect 3642 14159 3962 14160
rect 35610 14224 35930 14225
rect 35610 14160 35618 14224
rect 35682 14160 35698 14224
rect 35762 14160 35778 14224
rect 35842 14160 35858 14224
rect 35922 14160 35930 14224
rect 35610 14159 35930 14160
rect 40938 14224 41258 14225
rect 40938 14160 40946 14224
rect 41010 14160 41026 14224
rect 41090 14160 41106 14224
rect 41170 14160 41186 14224
rect 41250 14160 41258 14224
rect 40938 14159 41258 14160
rect 6306 13680 6626 13681
rect 6306 13616 6314 13680
rect 6378 13616 6394 13680
rect 6458 13616 6474 13680
rect 6538 13616 6554 13680
rect 6618 13616 6626 13680
rect 6306 13615 6626 13616
rect 38274 13680 38594 13681
rect 38274 13616 38282 13680
rect 38346 13616 38362 13680
rect 38426 13616 38442 13680
rect 38506 13616 38522 13680
rect 38586 13616 38594 13680
rect 38274 13615 38594 13616
rect 3642 13136 3962 13137
rect 3642 13072 3650 13136
rect 3714 13072 3730 13136
rect 3794 13072 3810 13136
rect 3874 13072 3890 13136
rect 3954 13072 3962 13136
rect 3642 13071 3962 13072
rect 35610 13136 35930 13137
rect 35610 13072 35618 13136
rect 35682 13072 35698 13136
rect 35762 13072 35778 13136
rect 35842 13072 35858 13136
rect 35922 13072 35930 13136
rect 35610 13071 35930 13072
rect 40938 13136 41258 13137
rect 40938 13072 40946 13136
rect 41010 13072 41026 13136
rect 41090 13072 41106 13136
rect 41170 13072 41186 13136
rect 41250 13072 41258 13136
rect 40938 13071 41258 13072
rect 6306 12592 6626 12593
rect 6306 12528 6314 12592
rect 6378 12528 6394 12592
rect 6458 12528 6474 12592
rect 6538 12528 6554 12592
rect 6618 12528 6626 12592
rect 6306 12527 6626 12528
rect 38274 12592 38594 12593
rect 38274 12528 38282 12592
rect 38346 12528 38362 12592
rect 38426 12528 38442 12592
rect 38506 12528 38522 12592
rect 38586 12528 38594 12592
rect 38274 12527 38594 12528
rect 3642 12048 3962 12049
rect 3642 11984 3650 12048
rect 3714 11984 3730 12048
rect 3794 11984 3810 12048
rect 3874 11984 3890 12048
rect 3954 11984 3962 12048
rect 3642 11983 3962 11984
rect 35610 12048 35930 12049
rect 35610 11984 35618 12048
rect 35682 11984 35698 12048
rect 35762 11984 35778 12048
rect 35842 11984 35858 12048
rect 35922 11984 35930 12048
rect 35610 11983 35930 11984
rect 40938 12048 41258 12049
rect 40938 11984 40946 12048
rect 41010 11984 41026 12048
rect 41090 11984 41106 12048
rect 41170 11984 41186 12048
rect 41250 11984 41258 12048
rect 40938 11983 41258 11984
rect 6306 11504 6626 11505
rect 6306 11440 6314 11504
rect 6378 11440 6394 11504
rect 6458 11440 6474 11504
rect 6538 11440 6554 11504
rect 6618 11440 6626 11504
rect 6306 11439 6626 11440
rect 38274 11504 38594 11505
rect 38274 11440 38282 11504
rect 38346 11440 38362 11504
rect 38426 11440 38442 11504
rect 38506 11440 38522 11504
rect 38586 11440 38594 11504
rect 38274 11439 38594 11440
rect 3642 10960 3962 10961
rect 3642 10896 3650 10960
rect 3714 10896 3730 10960
rect 3794 10896 3810 10960
rect 3874 10896 3890 10960
rect 3954 10896 3962 10960
rect 3642 10895 3962 10896
rect 35610 10960 35930 10961
rect 35610 10896 35618 10960
rect 35682 10896 35698 10960
rect 35762 10896 35778 10960
rect 35842 10896 35858 10960
rect 35922 10896 35930 10960
rect 35610 10895 35930 10896
rect 40938 10960 41258 10961
rect 40938 10896 40946 10960
rect 41010 10896 41026 10960
rect 41090 10896 41106 10960
rect 41170 10896 41186 10960
rect 41250 10896 41258 10960
rect 40938 10895 41258 10896
rect 31504 10482 31510 10484
rect 31174 10422 31510 10482
rect 31504 10420 31510 10422
rect 31574 10482 31580 10484
rect 34407 10482 34473 10485
rect 31574 10480 34473 10482
rect 31574 10424 34412 10480
rect 34468 10424 34473 10480
rect 31574 10422 34473 10424
rect 31574 10420 31580 10422
rect 34407 10419 34473 10422
rect 43515 10482 43581 10485
rect 45680 10482 46262 10494
rect 43515 10480 46262 10482
rect 43515 10424 43520 10480
rect 43576 10434 46262 10480
rect 68263 10482 68329 10485
rect 68263 10480 70734 10482
rect 43576 10424 45740 10434
rect 43515 10422 45740 10424
rect 68263 10424 68268 10480
rect 68324 10424 70734 10480
rect 68263 10422 70734 10424
rect 43515 10419 43581 10422
rect 68263 10419 68329 10422
rect 6306 10416 6626 10417
rect 6306 10352 6314 10416
rect 6378 10352 6394 10416
rect 6458 10352 6474 10416
rect 6538 10352 6554 10416
rect 6618 10352 6626 10416
rect 6306 10351 6626 10352
rect 38274 10416 38594 10417
rect 38274 10352 38282 10416
rect 38346 10352 38362 10416
rect 38426 10352 38442 10416
rect 38506 10352 38522 10416
rect 38586 10352 38594 10416
rect 38274 10351 38594 10352
rect 3642 9872 3962 9873
rect 3642 9808 3650 9872
rect 3714 9808 3730 9872
rect 3794 9808 3810 9872
rect 3874 9808 3890 9872
rect 3954 9808 3962 9872
rect 3642 9807 3962 9808
rect 35610 9872 35930 9873
rect 35610 9808 35618 9872
rect 35682 9808 35698 9872
rect 35762 9808 35778 9872
rect 35842 9808 35858 9872
rect 35922 9808 35930 9872
rect 35610 9807 35930 9808
rect 40938 9872 41258 9873
rect 40938 9808 40946 9872
rect 41010 9808 41026 9872
rect 41090 9808 41106 9872
rect 41170 9808 41186 9872
rect 41250 9808 41258 9872
rect 40938 9807 41258 9808
rect 91171 9530 91237 9533
rect 93946 9530 94746 9560
rect 91171 9528 94746 9530
rect 91171 9472 91176 9528
rect 91232 9472 94746 9528
rect 91171 9470 94746 9472
rect 91171 9467 91237 9470
rect 93946 9440 94746 9470
rect 6306 9328 6626 9329
rect 6306 9264 6314 9328
rect 6378 9264 6394 9328
rect 6458 9264 6474 9328
rect 6538 9264 6554 9328
rect 6618 9264 6626 9328
rect 6306 9263 6626 9264
rect 38274 9328 38594 9329
rect 38274 9264 38282 9328
rect 38346 9264 38362 9328
rect 38426 9264 38442 9328
rect 38506 9264 38522 9328
rect 38586 9264 38594 9328
rect 38274 9263 38594 9264
rect 3642 8784 3962 8785
rect 3642 8720 3650 8784
rect 3714 8720 3730 8784
rect 3794 8720 3810 8784
rect 3874 8720 3890 8784
rect 3954 8720 3962 8784
rect 3642 8719 3962 8720
rect 35610 8784 35930 8785
rect 35610 8720 35618 8784
rect 35682 8720 35698 8784
rect 35762 8720 35778 8784
rect 35842 8720 35858 8784
rect 35922 8720 35930 8784
rect 35610 8719 35930 8720
rect 40938 8784 41258 8785
rect 40938 8720 40946 8784
rect 41010 8720 41026 8784
rect 41090 8720 41106 8784
rect 41170 8720 41186 8784
rect 41250 8720 41258 8784
rect 40938 8719 41258 8720
rect 6306 8240 6626 8241
rect 6306 8176 6314 8240
rect 6378 8176 6394 8240
rect 6458 8176 6474 8240
rect 6538 8176 6554 8240
rect 6618 8176 6626 8240
rect 6306 8175 6626 8176
rect 38274 8240 38594 8241
rect 38274 8176 38282 8240
rect 38346 8176 38362 8240
rect 38426 8176 38442 8240
rect 38506 8176 38522 8240
rect 38586 8176 38594 8240
rect 38274 8175 38594 8176
rect 3642 7696 3962 7697
rect 3642 7632 3650 7696
rect 3714 7632 3730 7696
rect 3794 7632 3810 7696
rect 3874 7632 3890 7696
rect 3954 7632 3962 7696
rect 3642 7631 3962 7632
rect 35610 7696 35930 7697
rect 35610 7632 35618 7696
rect 35682 7632 35698 7696
rect 35762 7632 35778 7696
rect 35842 7632 35858 7696
rect 35922 7632 35930 7696
rect 35610 7631 35930 7632
rect 40938 7696 41258 7697
rect 40938 7632 40946 7696
rect 41010 7632 41026 7696
rect 41090 7632 41106 7696
rect 41170 7632 41186 7696
rect 41250 7632 41258 7696
rect 40938 7631 41258 7632
rect 6306 7152 6626 7153
rect 6306 7088 6314 7152
rect 6378 7088 6394 7152
rect 6458 7088 6474 7152
rect 6538 7088 6554 7152
rect 6618 7088 6626 7152
rect 6306 7087 6626 7088
rect 38274 7152 38594 7153
rect 38274 7088 38282 7152
rect 38346 7088 38362 7152
rect 38426 7088 38442 7152
rect 38506 7088 38522 7152
rect 38586 7088 38594 7152
rect 38274 7087 38594 7088
rect 3642 6608 3962 6609
rect 3642 6544 3650 6608
rect 3714 6544 3730 6608
rect 3794 6544 3810 6608
rect 3874 6544 3890 6608
rect 3954 6544 3962 6608
rect 3642 6543 3962 6544
rect 35610 6608 35930 6609
rect 35610 6544 35618 6608
rect 35682 6544 35698 6608
rect 35762 6544 35778 6608
rect 35842 6544 35858 6608
rect 35922 6544 35930 6608
rect 35610 6543 35930 6544
rect 40938 6608 41258 6609
rect 40938 6544 40946 6608
rect 41010 6544 41026 6608
rect 41090 6544 41106 6608
rect 41170 6544 41186 6608
rect 41250 6544 41258 6608
rect 40938 6543 41258 6544
rect 6306 6064 6626 6065
rect 6306 6000 6314 6064
rect 6378 6000 6394 6064
rect 6458 6000 6474 6064
rect 6538 6000 6554 6064
rect 6618 6000 6626 6064
rect 6306 5999 6626 6000
rect 38274 6064 38594 6065
rect 38274 6000 38282 6064
rect 38346 6000 38362 6064
rect 38426 6000 38442 6064
rect 38506 6000 38522 6064
rect 38586 6000 38594 6064
rect 38274 5999 38594 6000
rect 3642 5520 3962 5521
rect 3642 5456 3650 5520
rect 3714 5456 3730 5520
rect 3794 5456 3810 5520
rect 3874 5456 3890 5520
rect 3954 5456 3962 5520
rect 3642 5455 3962 5456
rect 35610 5520 35930 5521
rect 35610 5456 35618 5520
rect 35682 5456 35698 5520
rect 35762 5456 35778 5520
rect 35842 5456 35858 5520
rect 35922 5456 35930 5520
rect 35610 5455 35930 5456
rect 40938 5520 41258 5521
rect 40938 5456 40946 5520
rect 41010 5456 41026 5520
rect 41090 5456 41106 5520
rect 41170 5456 41186 5520
rect 41250 5456 41258 5520
rect 40938 5455 41258 5456
rect 6306 4976 6626 4977
rect 6306 4912 6314 4976
rect 6378 4912 6394 4976
rect 6458 4912 6474 4976
rect 6538 4912 6554 4976
rect 6618 4912 6626 4976
rect 6306 4911 6626 4912
rect 38274 4976 38594 4977
rect 38274 4912 38282 4976
rect 38346 4912 38362 4976
rect 38426 4912 38442 4976
rect 38506 4912 38522 4976
rect 38586 4912 38594 4976
rect 38274 4911 38594 4912
rect 3642 4432 3962 4433
rect 3642 4368 3650 4432
rect 3714 4368 3730 4432
rect 3794 4368 3810 4432
rect 3874 4368 3890 4432
rect 3954 4368 3962 4432
rect 3642 4367 3962 4368
rect 35610 4432 35930 4433
rect 35610 4368 35618 4432
rect 35682 4368 35698 4432
rect 35762 4368 35778 4432
rect 35842 4368 35858 4432
rect 35922 4368 35930 4432
rect 35610 4367 35930 4368
rect 40938 4432 41258 4433
rect 40938 4368 40946 4432
rect 41010 4368 41026 4432
rect 41090 4368 41106 4432
rect 41170 4368 41186 4432
rect 41250 4368 41258 4432
rect 40938 4367 41258 4368
rect 6306 3888 6626 3889
rect 6306 3824 6314 3888
rect 6378 3824 6394 3888
rect 6458 3824 6474 3888
rect 6538 3824 6554 3888
rect 6618 3824 6626 3888
rect 6306 3823 6626 3824
rect 38274 3888 38594 3889
rect 38274 3824 38282 3888
rect 38346 3824 38362 3888
rect 38426 3824 38442 3888
rect 38506 3824 38522 3888
rect 38586 3824 38594 3888
rect 38274 3823 38594 3824
rect 3642 3344 3962 3345
rect 3642 3280 3650 3344
rect 3714 3280 3730 3344
rect 3794 3280 3810 3344
rect 3874 3280 3890 3344
rect 3954 3280 3962 3344
rect 3642 3279 3962 3280
rect 35610 3344 35930 3345
rect 35610 3280 35618 3344
rect 35682 3280 35698 3344
rect 35762 3280 35778 3344
rect 35842 3280 35858 3344
rect 35922 3280 35930 3344
rect 35610 3279 35930 3280
rect 40938 3344 41258 3345
rect 40938 3280 40946 3344
rect 41010 3280 41026 3344
rect 41090 3280 41106 3344
rect 41170 3280 41186 3344
rect 41250 3280 41258 3344
rect 40938 3279 41258 3280
rect 6306 2800 6626 2801
rect 6306 2736 6314 2800
rect 6378 2736 6394 2800
rect 6458 2736 6474 2800
rect 6538 2736 6554 2800
rect 6618 2736 6626 2800
rect 6306 2735 6626 2736
rect 38274 2800 38594 2801
rect 38274 2736 38282 2800
rect 38346 2736 38362 2800
rect 38426 2736 38442 2800
rect 38506 2736 38522 2800
rect 38586 2736 38594 2800
rect 38274 2735 38594 2736
rect 31371 2322 31437 2325
rect 31174 2320 31437 2322
rect 31174 2264 31376 2320
rect 31432 2264 31437 2320
rect 31174 2262 31437 2264
rect 31371 2259 31437 2262
rect 43239 2322 43305 2325
rect 45680 2322 46262 2362
rect 43239 2320 46262 2322
rect 43239 2264 43244 2320
rect 43300 2302 46262 2320
rect 69735 2322 69801 2325
rect 69735 2320 70734 2322
rect 43300 2264 45740 2302
rect 43239 2262 45740 2264
rect 69735 2264 69740 2320
rect 69796 2264 70734 2320
rect 69735 2262 70734 2264
rect 43239 2259 43305 2262
rect 69735 2259 69801 2262
rect 3642 2256 3962 2257
rect 3642 2192 3650 2256
rect 3714 2192 3730 2256
rect 3794 2192 3810 2256
rect 3874 2192 3890 2256
rect 3954 2192 3962 2256
rect 3642 2191 3962 2192
rect 35610 2256 35930 2257
rect 35610 2192 35618 2256
rect 35682 2192 35698 2256
rect 35762 2192 35778 2256
rect 35842 2192 35858 2256
rect 35922 2192 35930 2256
rect 35610 2191 35930 2192
rect 40938 2256 41258 2257
rect 40938 2192 40946 2256
rect 41010 2192 41026 2256
rect 41090 2192 41106 2256
rect 41170 2192 41186 2256
rect 41250 2192 41258 2256
rect 40938 2191 41258 2192
rect 6306 1712 6626 1713
rect 6306 1648 6314 1712
rect 6378 1648 6394 1712
rect 6458 1648 6474 1712
rect 6538 1648 6554 1712
rect 6618 1648 6626 1712
rect 6306 1647 6626 1648
rect 38274 1712 38594 1713
rect 38274 1648 38282 1712
rect 38346 1648 38362 1712
rect 38426 1648 38442 1712
rect 38506 1648 38522 1712
rect 38586 1648 38594 1712
rect 38274 1647 38594 1648
rect 3642 1168 3962 1169
rect 3642 1104 3650 1168
rect 3714 1104 3730 1168
rect 3794 1104 3810 1168
rect 3874 1104 3890 1168
rect 3954 1104 3962 1168
rect 3642 1103 3962 1104
rect 35610 1168 35930 1169
rect 35610 1104 35618 1168
rect 35682 1104 35698 1168
rect 35762 1104 35778 1168
rect 35842 1104 35858 1168
rect 35922 1104 35930 1168
rect 35610 1103 35930 1104
rect 40938 1168 41258 1169
rect 40938 1104 40946 1168
rect 41010 1104 41026 1168
rect 41090 1104 41106 1168
rect 41170 1104 41186 1168
rect 41250 1104 41258 1168
rect 40938 1103 41258 1104
rect 6306 624 6626 625
rect 6306 560 6314 624
rect 6378 560 6394 624
rect 6458 560 6474 624
rect 6538 560 6554 624
rect 6618 560 6626 624
rect 6306 559 6626 560
rect 38274 624 38594 625
rect 38274 560 38282 624
rect 38346 560 38362 624
rect 38426 560 38442 624
rect 38506 560 38522 624
rect 38586 560 38594 624
rect 38274 559 38594 560
rect 3642 80 3962 81
rect 3642 16 3650 80
rect 3714 16 3730 80
rect 3794 16 3810 80
rect 3874 16 3890 80
rect 3954 16 3962 80
rect 3642 15 3962 16
rect 35610 80 35930 81
rect 35610 16 35618 80
rect 35682 16 35698 80
rect 35762 16 35778 80
rect 35842 16 35858 80
rect 35922 16 35930 80
rect 35610 15 35930 16
rect 40938 80 41258 81
rect 40938 16 40946 80
rect 41010 16 41026 80
rect 41090 16 41106 80
rect 41170 16 41186 80
rect 41250 16 41258 80
rect 40938 15 41258 16
<< via3 >>
rect 6314 41964 6378 41968
rect 6314 41908 6318 41964
rect 6318 41908 6374 41964
rect 6374 41908 6378 41964
rect 6314 41904 6378 41908
rect 6394 41964 6458 41968
rect 6394 41908 6398 41964
rect 6398 41908 6454 41964
rect 6454 41908 6458 41964
rect 6394 41904 6458 41908
rect 6474 41964 6538 41968
rect 6474 41908 6478 41964
rect 6478 41908 6534 41964
rect 6534 41908 6538 41964
rect 6474 41904 6538 41908
rect 6554 41964 6618 41968
rect 6554 41908 6558 41964
rect 6558 41908 6614 41964
rect 6614 41908 6618 41964
rect 6554 41904 6618 41908
rect 11642 41964 11706 41968
rect 11642 41908 11646 41964
rect 11646 41908 11702 41964
rect 11702 41908 11706 41964
rect 11642 41904 11706 41908
rect 11722 41964 11786 41968
rect 11722 41908 11726 41964
rect 11726 41908 11782 41964
rect 11782 41908 11786 41964
rect 11722 41904 11786 41908
rect 11802 41964 11866 41968
rect 11802 41908 11806 41964
rect 11806 41908 11862 41964
rect 11862 41908 11866 41964
rect 11802 41904 11866 41908
rect 11882 41964 11946 41968
rect 11882 41908 11886 41964
rect 11886 41908 11942 41964
rect 11942 41908 11946 41964
rect 11882 41904 11946 41908
rect 16970 41964 17034 41968
rect 16970 41908 16974 41964
rect 16974 41908 17030 41964
rect 17030 41908 17034 41964
rect 16970 41904 17034 41908
rect 17050 41964 17114 41968
rect 17050 41908 17054 41964
rect 17054 41908 17110 41964
rect 17110 41908 17114 41964
rect 17050 41904 17114 41908
rect 17130 41964 17194 41968
rect 17130 41908 17134 41964
rect 17134 41908 17190 41964
rect 17190 41908 17194 41964
rect 17130 41904 17194 41908
rect 17210 41964 17274 41968
rect 17210 41908 17214 41964
rect 17214 41908 17270 41964
rect 17270 41908 17274 41964
rect 17210 41904 17274 41908
rect 22298 41964 22362 41968
rect 22298 41908 22302 41964
rect 22302 41908 22358 41964
rect 22358 41908 22362 41964
rect 22298 41904 22362 41908
rect 22378 41964 22442 41968
rect 22378 41908 22382 41964
rect 22382 41908 22438 41964
rect 22438 41908 22442 41964
rect 22378 41904 22442 41908
rect 22458 41964 22522 41968
rect 22458 41908 22462 41964
rect 22462 41908 22518 41964
rect 22518 41908 22522 41964
rect 22458 41904 22522 41908
rect 22538 41964 22602 41968
rect 22538 41908 22542 41964
rect 22542 41908 22598 41964
rect 22598 41908 22602 41964
rect 22538 41904 22602 41908
rect 27626 41964 27690 41968
rect 27626 41908 27630 41964
rect 27630 41908 27686 41964
rect 27686 41908 27690 41964
rect 27626 41904 27690 41908
rect 27706 41964 27770 41968
rect 27706 41908 27710 41964
rect 27710 41908 27766 41964
rect 27766 41908 27770 41964
rect 27706 41904 27770 41908
rect 27786 41964 27850 41968
rect 27786 41908 27790 41964
rect 27790 41908 27846 41964
rect 27846 41908 27850 41964
rect 27786 41904 27850 41908
rect 27866 41964 27930 41968
rect 27866 41908 27870 41964
rect 27870 41908 27926 41964
rect 27926 41908 27930 41964
rect 27866 41904 27930 41908
rect 32954 41964 33018 41968
rect 32954 41908 32958 41964
rect 32958 41908 33014 41964
rect 33014 41908 33018 41964
rect 32954 41904 33018 41908
rect 33034 41964 33098 41968
rect 33034 41908 33038 41964
rect 33038 41908 33094 41964
rect 33094 41908 33098 41964
rect 33034 41904 33098 41908
rect 33114 41964 33178 41968
rect 33114 41908 33118 41964
rect 33118 41908 33174 41964
rect 33174 41908 33178 41964
rect 33114 41904 33178 41908
rect 33194 41964 33258 41968
rect 33194 41908 33198 41964
rect 33198 41908 33254 41964
rect 33254 41908 33258 41964
rect 33194 41904 33258 41908
rect 38282 41964 38346 41968
rect 38282 41908 38286 41964
rect 38286 41908 38342 41964
rect 38342 41908 38346 41964
rect 38282 41904 38346 41908
rect 38362 41964 38426 41968
rect 38362 41908 38366 41964
rect 38366 41908 38422 41964
rect 38422 41908 38426 41964
rect 38362 41904 38426 41908
rect 38442 41964 38506 41968
rect 38442 41908 38446 41964
rect 38446 41908 38502 41964
rect 38502 41908 38506 41964
rect 38442 41904 38506 41908
rect 38522 41964 38586 41968
rect 38522 41908 38526 41964
rect 38526 41908 38582 41964
rect 38582 41908 38586 41964
rect 38522 41904 38586 41908
rect 43610 41964 43674 41968
rect 43610 41908 43614 41964
rect 43614 41908 43670 41964
rect 43670 41908 43674 41964
rect 43610 41904 43674 41908
rect 43690 41964 43754 41968
rect 43690 41908 43694 41964
rect 43694 41908 43750 41964
rect 43750 41908 43754 41964
rect 43690 41904 43754 41908
rect 43770 41964 43834 41968
rect 43770 41908 43774 41964
rect 43774 41908 43830 41964
rect 43830 41908 43834 41964
rect 43770 41904 43834 41908
rect 43850 41964 43914 41968
rect 43850 41908 43854 41964
rect 43854 41908 43910 41964
rect 43910 41908 43914 41964
rect 43850 41904 43914 41908
rect 48938 41964 49002 41968
rect 48938 41908 48942 41964
rect 48942 41908 48998 41964
rect 48998 41908 49002 41964
rect 48938 41904 49002 41908
rect 49018 41964 49082 41968
rect 49018 41908 49022 41964
rect 49022 41908 49078 41964
rect 49078 41908 49082 41964
rect 49018 41904 49082 41908
rect 49098 41964 49162 41968
rect 49098 41908 49102 41964
rect 49102 41908 49158 41964
rect 49158 41908 49162 41964
rect 49098 41904 49162 41908
rect 49178 41964 49242 41968
rect 49178 41908 49182 41964
rect 49182 41908 49238 41964
rect 49238 41908 49242 41964
rect 49178 41904 49242 41908
rect 54266 41964 54330 41968
rect 54266 41908 54270 41964
rect 54270 41908 54326 41964
rect 54326 41908 54330 41964
rect 54266 41904 54330 41908
rect 54346 41964 54410 41968
rect 54346 41908 54350 41964
rect 54350 41908 54406 41964
rect 54406 41908 54410 41964
rect 54346 41904 54410 41908
rect 54426 41964 54490 41968
rect 54426 41908 54430 41964
rect 54430 41908 54486 41964
rect 54486 41908 54490 41964
rect 54426 41904 54490 41908
rect 54506 41964 54570 41968
rect 54506 41908 54510 41964
rect 54510 41908 54566 41964
rect 54566 41908 54570 41964
rect 54506 41904 54570 41908
rect 59594 41964 59658 41968
rect 59594 41908 59598 41964
rect 59598 41908 59654 41964
rect 59654 41908 59658 41964
rect 59594 41904 59658 41908
rect 59674 41964 59738 41968
rect 59674 41908 59678 41964
rect 59678 41908 59734 41964
rect 59734 41908 59738 41964
rect 59674 41904 59738 41908
rect 59754 41964 59818 41968
rect 59754 41908 59758 41964
rect 59758 41908 59814 41964
rect 59814 41908 59818 41964
rect 59754 41904 59818 41908
rect 59834 41964 59898 41968
rect 59834 41908 59838 41964
rect 59838 41908 59894 41964
rect 59894 41908 59898 41964
rect 59834 41904 59898 41908
rect 64922 41964 64986 41968
rect 64922 41908 64926 41964
rect 64926 41908 64982 41964
rect 64982 41908 64986 41964
rect 64922 41904 64986 41908
rect 65002 41964 65066 41968
rect 65002 41908 65006 41964
rect 65006 41908 65062 41964
rect 65062 41908 65066 41964
rect 65002 41904 65066 41908
rect 65082 41964 65146 41968
rect 65082 41908 65086 41964
rect 65086 41908 65142 41964
rect 65142 41908 65146 41964
rect 65082 41904 65146 41908
rect 65162 41964 65226 41968
rect 65162 41908 65166 41964
rect 65166 41908 65222 41964
rect 65222 41908 65226 41964
rect 65162 41904 65226 41908
rect 70250 41964 70314 41968
rect 70250 41908 70254 41964
rect 70254 41908 70310 41964
rect 70310 41908 70314 41964
rect 70250 41904 70314 41908
rect 70330 41964 70394 41968
rect 70330 41908 70334 41964
rect 70334 41908 70390 41964
rect 70390 41908 70394 41964
rect 70330 41904 70394 41908
rect 70410 41964 70474 41968
rect 70410 41908 70414 41964
rect 70414 41908 70470 41964
rect 70470 41908 70474 41964
rect 70410 41904 70474 41908
rect 70490 41964 70554 41968
rect 70490 41908 70494 41964
rect 70494 41908 70550 41964
rect 70550 41908 70554 41964
rect 70490 41904 70554 41908
rect 75578 41964 75642 41968
rect 75578 41908 75582 41964
rect 75582 41908 75638 41964
rect 75638 41908 75642 41964
rect 75578 41904 75642 41908
rect 75658 41964 75722 41968
rect 75658 41908 75662 41964
rect 75662 41908 75718 41964
rect 75718 41908 75722 41964
rect 75658 41904 75722 41908
rect 75738 41964 75802 41968
rect 75738 41908 75742 41964
rect 75742 41908 75798 41964
rect 75798 41908 75802 41964
rect 75738 41904 75802 41908
rect 75818 41964 75882 41968
rect 75818 41908 75822 41964
rect 75822 41908 75878 41964
rect 75878 41908 75882 41964
rect 75818 41904 75882 41908
rect 80906 41964 80970 41968
rect 80906 41908 80910 41964
rect 80910 41908 80966 41964
rect 80966 41908 80970 41964
rect 80906 41904 80970 41908
rect 80986 41964 81050 41968
rect 80986 41908 80990 41964
rect 80990 41908 81046 41964
rect 81046 41908 81050 41964
rect 80986 41904 81050 41908
rect 81066 41964 81130 41968
rect 81066 41908 81070 41964
rect 81070 41908 81126 41964
rect 81126 41908 81130 41964
rect 81066 41904 81130 41908
rect 81146 41964 81210 41968
rect 81146 41908 81150 41964
rect 81150 41908 81206 41964
rect 81206 41908 81210 41964
rect 81146 41904 81210 41908
rect 86234 41964 86298 41968
rect 86234 41908 86238 41964
rect 86238 41908 86294 41964
rect 86294 41908 86298 41964
rect 86234 41904 86298 41908
rect 86314 41964 86378 41968
rect 86314 41908 86318 41964
rect 86318 41908 86374 41964
rect 86374 41908 86378 41964
rect 86314 41904 86378 41908
rect 86394 41964 86458 41968
rect 86394 41908 86398 41964
rect 86398 41908 86454 41964
rect 86454 41908 86458 41964
rect 86394 41904 86458 41908
rect 86474 41964 86538 41968
rect 86474 41908 86478 41964
rect 86478 41908 86534 41964
rect 86534 41908 86538 41964
rect 86474 41904 86538 41908
rect 91562 41964 91626 41968
rect 91562 41908 91566 41964
rect 91566 41908 91622 41964
rect 91622 41908 91626 41964
rect 91562 41904 91626 41908
rect 91642 41964 91706 41968
rect 91642 41908 91646 41964
rect 91646 41908 91702 41964
rect 91702 41908 91706 41964
rect 91642 41904 91706 41908
rect 91722 41964 91786 41968
rect 91722 41908 91726 41964
rect 91726 41908 91782 41964
rect 91782 41908 91786 41964
rect 91722 41904 91786 41908
rect 91802 41964 91866 41968
rect 91802 41908 91806 41964
rect 91806 41908 91862 41964
rect 91862 41908 91866 41964
rect 91802 41904 91866 41908
rect 3650 41420 3714 41424
rect 3650 41364 3654 41420
rect 3654 41364 3710 41420
rect 3710 41364 3714 41420
rect 3650 41360 3714 41364
rect 3730 41420 3794 41424
rect 3730 41364 3734 41420
rect 3734 41364 3790 41420
rect 3790 41364 3794 41420
rect 3730 41360 3794 41364
rect 3810 41420 3874 41424
rect 3810 41364 3814 41420
rect 3814 41364 3870 41420
rect 3870 41364 3874 41420
rect 3810 41360 3874 41364
rect 3890 41420 3954 41424
rect 3890 41364 3894 41420
rect 3894 41364 3950 41420
rect 3950 41364 3954 41420
rect 3890 41360 3954 41364
rect 8978 41420 9042 41424
rect 8978 41364 8982 41420
rect 8982 41364 9038 41420
rect 9038 41364 9042 41420
rect 8978 41360 9042 41364
rect 9058 41420 9122 41424
rect 9058 41364 9062 41420
rect 9062 41364 9118 41420
rect 9118 41364 9122 41420
rect 9058 41360 9122 41364
rect 9138 41420 9202 41424
rect 9138 41364 9142 41420
rect 9142 41364 9198 41420
rect 9198 41364 9202 41420
rect 9138 41360 9202 41364
rect 9218 41420 9282 41424
rect 9218 41364 9222 41420
rect 9222 41364 9278 41420
rect 9278 41364 9282 41420
rect 9218 41360 9282 41364
rect 14306 41420 14370 41424
rect 14306 41364 14310 41420
rect 14310 41364 14366 41420
rect 14366 41364 14370 41420
rect 14306 41360 14370 41364
rect 14386 41420 14450 41424
rect 14386 41364 14390 41420
rect 14390 41364 14446 41420
rect 14446 41364 14450 41420
rect 14386 41360 14450 41364
rect 14466 41420 14530 41424
rect 14466 41364 14470 41420
rect 14470 41364 14526 41420
rect 14526 41364 14530 41420
rect 14466 41360 14530 41364
rect 14546 41420 14610 41424
rect 14546 41364 14550 41420
rect 14550 41364 14606 41420
rect 14606 41364 14610 41420
rect 14546 41360 14610 41364
rect 19634 41420 19698 41424
rect 19634 41364 19638 41420
rect 19638 41364 19694 41420
rect 19694 41364 19698 41420
rect 19634 41360 19698 41364
rect 19714 41420 19778 41424
rect 19714 41364 19718 41420
rect 19718 41364 19774 41420
rect 19774 41364 19778 41420
rect 19714 41360 19778 41364
rect 19794 41420 19858 41424
rect 19794 41364 19798 41420
rect 19798 41364 19854 41420
rect 19854 41364 19858 41420
rect 19794 41360 19858 41364
rect 19874 41420 19938 41424
rect 19874 41364 19878 41420
rect 19878 41364 19934 41420
rect 19934 41364 19938 41420
rect 19874 41360 19938 41364
rect 24962 41420 25026 41424
rect 24962 41364 24966 41420
rect 24966 41364 25022 41420
rect 25022 41364 25026 41420
rect 24962 41360 25026 41364
rect 25042 41420 25106 41424
rect 25042 41364 25046 41420
rect 25046 41364 25102 41420
rect 25102 41364 25106 41420
rect 25042 41360 25106 41364
rect 25122 41420 25186 41424
rect 25122 41364 25126 41420
rect 25126 41364 25182 41420
rect 25182 41364 25186 41420
rect 25122 41360 25186 41364
rect 25202 41420 25266 41424
rect 25202 41364 25206 41420
rect 25206 41364 25262 41420
rect 25262 41364 25266 41420
rect 25202 41360 25266 41364
rect 30290 41420 30354 41424
rect 30290 41364 30294 41420
rect 30294 41364 30350 41420
rect 30350 41364 30354 41420
rect 30290 41360 30354 41364
rect 30370 41420 30434 41424
rect 30370 41364 30374 41420
rect 30374 41364 30430 41420
rect 30430 41364 30434 41420
rect 30370 41360 30434 41364
rect 30450 41420 30514 41424
rect 30450 41364 30454 41420
rect 30454 41364 30510 41420
rect 30510 41364 30514 41420
rect 30450 41360 30514 41364
rect 30530 41420 30594 41424
rect 30530 41364 30534 41420
rect 30534 41364 30590 41420
rect 30590 41364 30594 41420
rect 30530 41360 30594 41364
rect 35618 41420 35682 41424
rect 35618 41364 35622 41420
rect 35622 41364 35678 41420
rect 35678 41364 35682 41420
rect 35618 41360 35682 41364
rect 35698 41420 35762 41424
rect 35698 41364 35702 41420
rect 35702 41364 35758 41420
rect 35758 41364 35762 41420
rect 35698 41360 35762 41364
rect 35778 41420 35842 41424
rect 35778 41364 35782 41420
rect 35782 41364 35838 41420
rect 35838 41364 35842 41420
rect 35778 41360 35842 41364
rect 35858 41420 35922 41424
rect 35858 41364 35862 41420
rect 35862 41364 35918 41420
rect 35918 41364 35922 41420
rect 35858 41360 35922 41364
rect 40946 41420 41010 41424
rect 40946 41364 40950 41420
rect 40950 41364 41006 41420
rect 41006 41364 41010 41420
rect 40946 41360 41010 41364
rect 41026 41420 41090 41424
rect 41026 41364 41030 41420
rect 41030 41364 41086 41420
rect 41086 41364 41090 41420
rect 41026 41360 41090 41364
rect 41106 41420 41170 41424
rect 41106 41364 41110 41420
rect 41110 41364 41166 41420
rect 41166 41364 41170 41420
rect 41106 41360 41170 41364
rect 41186 41420 41250 41424
rect 41186 41364 41190 41420
rect 41190 41364 41246 41420
rect 41246 41364 41250 41420
rect 41186 41360 41250 41364
rect 46274 41420 46338 41424
rect 46274 41364 46278 41420
rect 46278 41364 46334 41420
rect 46334 41364 46338 41420
rect 46274 41360 46338 41364
rect 46354 41420 46418 41424
rect 46354 41364 46358 41420
rect 46358 41364 46414 41420
rect 46414 41364 46418 41420
rect 46354 41360 46418 41364
rect 46434 41420 46498 41424
rect 46434 41364 46438 41420
rect 46438 41364 46494 41420
rect 46494 41364 46498 41420
rect 46434 41360 46498 41364
rect 46514 41420 46578 41424
rect 46514 41364 46518 41420
rect 46518 41364 46574 41420
rect 46574 41364 46578 41420
rect 46514 41360 46578 41364
rect 51602 41420 51666 41424
rect 51602 41364 51606 41420
rect 51606 41364 51662 41420
rect 51662 41364 51666 41420
rect 51602 41360 51666 41364
rect 51682 41420 51746 41424
rect 51682 41364 51686 41420
rect 51686 41364 51742 41420
rect 51742 41364 51746 41420
rect 51682 41360 51746 41364
rect 51762 41420 51826 41424
rect 51762 41364 51766 41420
rect 51766 41364 51822 41420
rect 51822 41364 51826 41420
rect 51762 41360 51826 41364
rect 51842 41420 51906 41424
rect 51842 41364 51846 41420
rect 51846 41364 51902 41420
rect 51902 41364 51906 41420
rect 51842 41360 51906 41364
rect 56930 41420 56994 41424
rect 56930 41364 56934 41420
rect 56934 41364 56990 41420
rect 56990 41364 56994 41420
rect 56930 41360 56994 41364
rect 57010 41420 57074 41424
rect 57010 41364 57014 41420
rect 57014 41364 57070 41420
rect 57070 41364 57074 41420
rect 57010 41360 57074 41364
rect 57090 41420 57154 41424
rect 57090 41364 57094 41420
rect 57094 41364 57150 41420
rect 57150 41364 57154 41420
rect 57090 41360 57154 41364
rect 57170 41420 57234 41424
rect 57170 41364 57174 41420
rect 57174 41364 57230 41420
rect 57230 41364 57234 41420
rect 57170 41360 57234 41364
rect 62258 41420 62322 41424
rect 62258 41364 62262 41420
rect 62262 41364 62318 41420
rect 62318 41364 62322 41420
rect 62258 41360 62322 41364
rect 62338 41420 62402 41424
rect 62338 41364 62342 41420
rect 62342 41364 62398 41420
rect 62398 41364 62402 41420
rect 62338 41360 62402 41364
rect 62418 41420 62482 41424
rect 62418 41364 62422 41420
rect 62422 41364 62478 41420
rect 62478 41364 62482 41420
rect 62418 41360 62482 41364
rect 62498 41420 62562 41424
rect 62498 41364 62502 41420
rect 62502 41364 62558 41420
rect 62558 41364 62562 41420
rect 62498 41360 62562 41364
rect 67586 41420 67650 41424
rect 67586 41364 67590 41420
rect 67590 41364 67646 41420
rect 67646 41364 67650 41420
rect 67586 41360 67650 41364
rect 67666 41420 67730 41424
rect 67666 41364 67670 41420
rect 67670 41364 67726 41420
rect 67726 41364 67730 41420
rect 67666 41360 67730 41364
rect 67746 41420 67810 41424
rect 67746 41364 67750 41420
rect 67750 41364 67806 41420
rect 67806 41364 67810 41420
rect 67746 41360 67810 41364
rect 67826 41420 67890 41424
rect 67826 41364 67830 41420
rect 67830 41364 67886 41420
rect 67886 41364 67890 41420
rect 67826 41360 67890 41364
rect 72914 41420 72978 41424
rect 72914 41364 72918 41420
rect 72918 41364 72974 41420
rect 72974 41364 72978 41420
rect 72914 41360 72978 41364
rect 72994 41420 73058 41424
rect 72994 41364 72998 41420
rect 72998 41364 73054 41420
rect 73054 41364 73058 41420
rect 72994 41360 73058 41364
rect 73074 41420 73138 41424
rect 73074 41364 73078 41420
rect 73078 41364 73134 41420
rect 73134 41364 73138 41420
rect 73074 41360 73138 41364
rect 73154 41420 73218 41424
rect 73154 41364 73158 41420
rect 73158 41364 73214 41420
rect 73214 41364 73218 41420
rect 73154 41360 73218 41364
rect 78242 41420 78306 41424
rect 78242 41364 78246 41420
rect 78246 41364 78302 41420
rect 78302 41364 78306 41420
rect 78242 41360 78306 41364
rect 78322 41420 78386 41424
rect 78322 41364 78326 41420
rect 78326 41364 78382 41420
rect 78382 41364 78386 41420
rect 78322 41360 78386 41364
rect 78402 41420 78466 41424
rect 78402 41364 78406 41420
rect 78406 41364 78462 41420
rect 78462 41364 78466 41420
rect 78402 41360 78466 41364
rect 78482 41420 78546 41424
rect 78482 41364 78486 41420
rect 78486 41364 78542 41420
rect 78542 41364 78546 41420
rect 78482 41360 78546 41364
rect 83570 41420 83634 41424
rect 83570 41364 83574 41420
rect 83574 41364 83630 41420
rect 83630 41364 83634 41420
rect 83570 41360 83634 41364
rect 83650 41420 83714 41424
rect 83650 41364 83654 41420
rect 83654 41364 83710 41420
rect 83710 41364 83714 41420
rect 83650 41360 83714 41364
rect 83730 41420 83794 41424
rect 83730 41364 83734 41420
rect 83734 41364 83790 41420
rect 83790 41364 83794 41420
rect 83730 41360 83794 41364
rect 83810 41420 83874 41424
rect 83810 41364 83814 41420
rect 83814 41364 83870 41420
rect 83870 41364 83874 41420
rect 83810 41360 83874 41364
rect 88898 41420 88962 41424
rect 88898 41364 88902 41420
rect 88902 41364 88958 41420
rect 88958 41364 88962 41420
rect 88898 41360 88962 41364
rect 88978 41420 89042 41424
rect 88978 41364 88982 41420
rect 88982 41364 89038 41420
rect 89038 41364 89042 41420
rect 88978 41360 89042 41364
rect 89058 41420 89122 41424
rect 89058 41364 89062 41420
rect 89062 41364 89118 41420
rect 89118 41364 89122 41420
rect 89058 41360 89122 41364
rect 89138 41420 89202 41424
rect 89138 41364 89142 41420
rect 89142 41364 89198 41420
rect 89198 41364 89202 41420
rect 89138 41360 89202 41364
rect 6314 40876 6378 40880
rect 6314 40820 6318 40876
rect 6318 40820 6374 40876
rect 6374 40820 6378 40876
rect 6314 40816 6378 40820
rect 6394 40876 6458 40880
rect 6394 40820 6398 40876
rect 6398 40820 6454 40876
rect 6454 40820 6458 40876
rect 6394 40816 6458 40820
rect 6474 40876 6538 40880
rect 6474 40820 6478 40876
rect 6478 40820 6534 40876
rect 6534 40820 6538 40876
rect 6474 40816 6538 40820
rect 6554 40876 6618 40880
rect 6554 40820 6558 40876
rect 6558 40820 6614 40876
rect 6614 40820 6618 40876
rect 6554 40816 6618 40820
rect 11642 40876 11706 40880
rect 11642 40820 11646 40876
rect 11646 40820 11702 40876
rect 11702 40820 11706 40876
rect 11642 40816 11706 40820
rect 11722 40876 11786 40880
rect 11722 40820 11726 40876
rect 11726 40820 11782 40876
rect 11782 40820 11786 40876
rect 11722 40816 11786 40820
rect 11802 40876 11866 40880
rect 11802 40820 11806 40876
rect 11806 40820 11862 40876
rect 11862 40820 11866 40876
rect 11802 40816 11866 40820
rect 11882 40876 11946 40880
rect 11882 40820 11886 40876
rect 11886 40820 11942 40876
rect 11942 40820 11946 40876
rect 11882 40816 11946 40820
rect 16970 40876 17034 40880
rect 16970 40820 16974 40876
rect 16974 40820 17030 40876
rect 17030 40820 17034 40876
rect 16970 40816 17034 40820
rect 17050 40876 17114 40880
rect 17050 40820 17054 40876
rect 17054 40820 17110 40876
rect 17110 40820 17114 40876
rect 17050 40816 17114 40820
rect 17130 40876 17194 40880
rect 17130 40820 17134 40876
rect 17134 40820 17190 40876
rect 17190 40820 17194 40876
rect 17130 40816 17194 40820
rect 17210 40876 17274 40880
rect 17210 40820 17214 40876
rect 17214 40820 17270 40876
rect 17270 40820 17274 40876
rect 17210 40816 17274 40820
rect 22298 40876 22362 40880
rect 22298 40820 22302 40876
rect 22302 40820 22358 40876
rect 22358 40820 22362 40876
rect 22298 40816 22362 40820
rect 22378 40876 22442 40880
rect 22378 40820 22382 40876
rect 22382 40820 22438 40876
rect 22438 40820 22442 40876
rect 22378 40816 22442 40820
rect 22458 40876 22522 40880
rect 22458 40820 22462 40876
rect 22462 40820 22518 40876
rect 22518 40820 22522 40876
rect 22458 40816 22522 40820
rect 22538 40876 22602 40880
rect 22538 40820 22542 40876
rect 22542 40820 22598 40876
rect 22598 40820 22602 40876
rect 22538 40816 22602 40820
rect 27626 40876 27690 40880
rect 27626 40820 27630 40876
rect 27630 40820 27686 40876
rect 27686 40820 27690 40876
rect 27626 40816 27690 40820
rect 27706 40876 27770 40880
rect 27706 40820 27710 40876
rect 27710 40820 27766 40876
rect 27766 40820 27770 40876
rect 27706 40816 27770 40820
rect 27786 40876 27850 40880
rect 27786 40820 27790 40876
rect 27790 40820 27846 40876
rect 27846 40820 27850 40876
rect 27786 40816 27850 40820
rect 27866 40876 27930 40880
rect 27866 40820 27870 40876
rect 27870 40820 27926 40876
rect 27926 40820 27930 40876
rect 27866 40816 27930 40820
rect 32954 40876 33018 40880
rect 32954 40820 32958 40876
rect 32958 40820 33014 40876
rect 33014 40820 33018 40876
rect 32954 40816 33018 40820
rect 33034 40876 33098 40880
rect 33034 40820 33038 40876
rect 33038 40820 33094 40876
rect 33094 40820 33098 40876
rect 33034 40816 33098 40820
rect 33114 40876 33178 40880
rect 33114 40820 33118 40876
rect 33118 40820 33174 40876
rect 33174 40820 33178 40876
rect 33114 40816 33178 40820
rect 33194 40876 33258 40880
rect 33194 40820 33198 40876
rect 33198 40820 33254 40876
rect 33254 40820 33258 40876
rect 33194 40816 33258 40820
rect 38282 40876 38346 40880
rect 38282 40820 38286 40876
rect 38286 40820 38342 40876
rect 38342 40820 38346 40876
rect 38282 40816 38346 40820
rect 38362 40876 38426 40880
rect 38362 40820 38366 40876
rect 38366 40820 38422 40876
rect 38422 40820 38426 40876
rect 38362 40816 38426 40820
rect 38442 40876 38506 40880
rect 38442 40820 38446 40876
rect 38446 40820 38502 40876
rect 38502 40820 38506 40876
rect 38442 40816 38506 40820
rect 38522 40876 38586 40880
rect 38522 40820 38526 40876
rect 38526 40820 38582 40876
rect 38582 40820 38586 40876
rect 38522 40816 38586 40820
rect 43610 40876 43674 40880
rect 43610 40820 43614 40876
rect 43614 40820 43670 40876
rect 43670 40820 43674 40876
rect 43610 40816 43674 40820
rect 43690 40876 43754 40880
rect 43690 40820 43694 40876
rect 43694 40820 43750 40876
rect 43750 40820 43754 40876
rect 43690 40816 43754 40820
rect 43770 40876 43834 40880
rect 43770 40820 43774 40876
rect 43774 40820 43830 40876
rect 43830 40820 43834 40876
rect 43770 40816 43834 40820
rect 43850 40876 43914 40880
rect 43850 40820 43854 40876
rect 43854 40820 43910 40876
rect 43910 40820 43914 40876
rect 43850 40816 43914 40820
rect 48938 40876 49002 40880
rect 48938 40820 48942 40876
rect 48942 40820 48998 40876
rect 48998 40820 49002 40876
rect 48938 40816 49002 40820
rect 49018 40876 49082 40880
rect 49018 40820 49022 40876
rect 49022 40820 49078 40876
rect 49078 40820 49082 40876
rect 49018 40816 49082 40820
rect 49098 40876 49162 40880
rect 49098 40820 49102 40876
rect 49102 40820 49158 40876
rect 49158 40820 49162 40876
rect 49098 40816 49162 40820
rect 49178 40876 49242 40880
rect 49178 40820 49182 40876
rect 49182 40820 49238 40876
rect 49238 40820 49242 40876
rect 49178 40816 49242 40820
rect 54266 40876 54330 40880
rect 54266 40820 54270 40876
rect 54270 40820 54326 40876
rect 54326 40820 54330 40876
rect 54266 40816 54330 40820
rect 54346 40876 54410 40880
rect 54346 40820 54350 40876
rect 54350 40820 54406 40876
rect 54406 40820 54410 40876
rect 54346 40816 54410 40820
rect 54426 40876 54490 40880
rect 54426 40820 54430 40876
rect 54430 40820 54486 40876
rect 54486 40820 54490 40876
rect 54426 40816 54490 40820
rect 54506 40876 54570 40880
rect 54506 40820 54510 40876
rect 54510 40820 54566 40876
rect 54566 40820 54570 40876
rect 54506 40816 54570 40820
rect 59594 40876 59658 40880
rect 59594 40820 59598 40876
rect 59598 40820 59654 40876
rect 59654 40820 59658 40876
rect 59594 40816 59658 40820
rect 59674 40876 59738 40880
rect 59674 40820 59678 40876
rect 59678 40820 59734 40876
rect 59734 40820 59738 40876
rect 59674 40816 59738 40820
rect 59754 40876 59818 40880
rect 59754 40820 59758 40876
rect 59758 40820 59814 40876
rect 59814 40820 59818 40876
rect 59754 40816 59818 40820
rect 59834 40876 59898 40880
rect 59834 40820 59838 40876
rect 59838 40820 59894 40876
rect 59894 40820 59898 40876
rect 59834 40816 59898 40820
rect 64922 40876 64986 40880
rect 64922 40820 64926 40876
rect 64926 40820 64982 40876
rect 64982 40820 64986 40876
rect 64922 40816 64986 40820
rect 65002 40876 65066 40880
rect 65002 40820 65006 40876
rect 65006 40820 65062 40876
rect 65062 40820 65066 40876
rect 65002 40816 65066 40820
rect 65082 40876 65146 40880
rect 65082 40820 65086 40876
rect 65086 40820 65142 40876
rect 65142 40820 65146 40876
rect 65082 40816 65146 40820
rect 65162 40876 65226 40880
rect 65162 40820 65166 40876
rect 65166 40820 65222 40876
rect 65222 40820 65226 40876
rect 65162 40816 65226 40820
rect 70250 40876 70314 40880
rect 70250 40820 70254 40876
rect 70254 40820 70310 40876
rect 70310 40820 70314 40876
rect 70250 40816 70314 40820
rect 70330 40876 70394 40880
rect 70330 40820 70334 40876
rect 70334 40820 70390 40876
rect 70390 40820 70394 40876
rect 70330 40816 70394 40820
rect 70410 40876 70474 40880
rect 70410 40820 70414 40876
rect 70414 40820 70470 40876
rect 70470 40820 70474 40876
rect 70410 40816 70474 40820
rect 70490 40876 70554 40880
rect 70490 40820 70494 40876
rect 70494 40820 70550 40876
rect 70550 40820 70554 40876
rect 70490 40816 70554 40820
rect 75578 40876 75642 40880
rect 75578 40820 75582 40876
rect 75582 40820 75638 40876
rect 75638 40820 75642 40876
rect 75578 40816 75642 40820
rect 75658 40876 75722 40880
rect 75658 40820 75662 40876
rect 75662 40820 75718 40876
rect 75718 40820 75722 40876
rect 75658 40816 75722 40820
rect 75738 40876 75802 40880
rect 75738 40820 75742 40876
rect 75742 40820 75798 40876
rect 75798 40820 75802 40876
rect 75738 40816 75802 40820
rect 75818 40876 75882 40880
rect 75818 40820 75822 40876
rect 75822 40820 75878 40876
rect 75878 40820 75882 40876
rect 75818 40816 75882 40820
rect 80906 40876 80970 40880
rect 80906 40820 80910 40876
rect 80910 40820 80966 40876
rect 80966 40820 80970 40876
rect 80906 40816 80970 40820
rect 80986 40876 81050 40880
rect 80986 40820 80990 40876
rect 80990 40820 81046 40876
rect 81046 40820 81050 40876
rect 80986 40816 81050 40820
rect 81066 40876 81130 40880
rect 81066 40820 81070 40876
rect 81070 40820 81126 40876
rect 81126 40820 81130 40876
rect 81066 40816 81130 40820
rect 81146 40876 81210 40880
rect 81146 40820 81150 40876
rect 81150 40820 81206 40876
rect 81206 40820 81210 40876
rect 81146 40816 81210 40820
rect 86234 40876 86298 40880
rect 86234 40820 86238 40876
rect 86238 40820 86294 40876
rect 86294 40820 86298 40876
rect 86234 40816 86298 40820
rect 86314 40876 86378 40880
rect 86314 40820 86318 40876
rect 86318 40820 86374 40876
rect 86374 40820 86378 40876
rect 86314 40816 86378 40820
rect 86394 40876 86458 40880
rect 86394 40820 86398 40876
rect 86398 40820 86454 40876
rect 86454 40820 86458 40876
rect 86394 40816 86458 40820
rect 86474 40876 86538 40880
rect 86474 40820 86478 40876
rect 86478 40820 86534 40876
rect 86534 40820 86538 40876
rect 86474 40816 86538 40820
rect 91562 40876 91626 40880
rect 91562 40820 91566 40876
rect 91566 40820 91622 40876
rect 91622 40820 91626 40876
rect 91562 40816 91626 40820
rect 91642 40876 91706 40880
rect 91642 40820 91646 40876
rect 91646 40820 91702 40876
rect 91702 40820 91706 40876
rect 91642 40816 91706 40820
rect 91722 40876 91786 40880
rect 91722 40820 91726 40876
rect 91726 40820 91782 40876
rect 91782 40820 91786 40876
rect 91722 40816 91786 40820
rect 91802 40876 91866 40880
rect 91802 40820 91806 40876
rect 91806 40820 91862 40876
rect 91862 40820 91866 40876
rect 91802 40816 91866 40820
rect 3650 40332 3714 40336
rect 3650 40276 3654 40332
rect 3654 40276 3710 40332
rect 3710 40276 3714 40332
rect 3650 40272 3714 40276
rect 3730 40332 3794 40336
rect 3730 40276 3734 40332
rect 3734 40276 3790 40332
rect 3790 40276 3794 40332
rect 3730 40272 3794 40276
rect 3810 40332 3874 40336
rect 3810 40276 3814 40332
rect 3814 40276 3870 40332
rect 3870 40276 3874 40332
rect 3810 40272 3874 40276
rect 3890 40332 3954 40336
rect 3890 40276 3894 40332
rect 3894 40276 3950 40332
rect 3950 40276 3954 40332
rect 3890 40272 3954 40276
rect 8978 40332 9042 40336
rect 8978 40276 8982 40332
rect 8982 40276 9038 40332
rect 9038 40276 9042 40332
rect 8978 40272 9042 40276
rect 9058 40332 9122 40336
rect 9058 40276 9062 40332
rect 9062 40276 9118 40332
rect 9118 40276 9122 40332
rect 9058 40272 9122 40276
rect 9138 40332 9202 40336
rect 9138 40276 9142 40332
rect 9142 40276 9198 40332
rect 9198 40276 9202 40332
rect 9138 40272 9202 40276
rect 9218 40332 9282 40336
rect 9218 40276 9222 40332
rect 9222 40276 9278 40332
rect 9278 40276 9282 40332
rect 9218 40272 9282 40276
rect 14306 40332 14370 40336
rect 14306 40276 14310 40332
rect 14310 40276 14366 40332
rect 14366 40276 14370 40332
rect 14306 40272 14370 40276
rect 14386 40332 14450 40336
rect 14386 40276 14390 40332
rect 14390 40276 14446 40332
rect 14446 40276 14450 40332
rect 14386 40272 14450 40276
rect 14466 40332 14530 40336
rect 14466 40276 14470 40332
rect 14470 40276 14526 40332
rect 14526 40276 14530 40332
rect 14466 40272 14530 40276
rect 14546 40332 14610 40336
rect 14546 40276 14550 40332
rect 14550 40276 14606 40332
rect 14606 40276 14610 40332
rect 14546 40272 14610 40276
rect 19634 40332 19698 40336
rect 19634 40276 19638 40332
rect 19638 40276 19694 40332
rect 19694 40276 19698 40332
rect 19634 40272 19698 40276
rect 19714 40332 19778 40336
rect 19714 40276 19718 40332
rect 19718 40276 19774 40332
rect 19774 40276 19778 40332
rect 19714 40272 19778 40276
rect 19794 40332 19858 40336
rect 19794 40276 19798 40332
rect 19798 40276 19854 40332
rect 19854 40276 19858 40332
rect 19794 40272 19858 40276
rect 19874 40332 19938 40336
rect 19874 40276 19878 40332
rect 19878 40276 19934 40332
rect 19934 40276 19938 40332
rect 19874 40272 19938 40276
rect 24962 40332 25026 40336
rect 24962 40276 24966 40332
rect 24966 40276 25022 40332
rect 25022 40276 25026 40332
rect 24962 40272 25026 40276
rect 25042 40332 25106 40336
rect 25042 40276 25046 40332
rect 25046 40276 25102 40332
rect 25102 40276 25106 40332
rect 25042 40272 25106 40276
rect 25122 40332 25186 40336
rect 25122 40276 25126 40332
rect 25126 40276 25182 40332
rect 25182 40276 25186 40332
rect 25122 40272 25186 40276
rect 25202 40332 25266 40336
rect 25202 40276 25206 40332
rect 25206 40276 25262 40332
rect 25262 40276 25266 40332
rect 25202 40272 25266 40276
rect 30290 40332 30354 40336
rect 30290 40276 30294 40332
rect 30294 40276 30350 40332
rect 30350 40276 30354 40332
rect 30290 40272 30354 40276
rect 30370 40332 30434 40336
rect 30370 40276 30374 40332
rect 30374 40276 30430 40332
rect 30430 40276 30434 40332
rect 30370 40272 30434 40276
rect 30450 40332 30514 40336
rect 30450 40276 30454 40332
rect 30454 40276 30510 40332
rect 30510 40276 30514 40332
rect 30450 40272 30514 40276
rect 30530 40332 30594 40336
rect 30530 40276 30534 40332
rect 30534 40276 30590 40332
rect 30590 40276 30594 40332
rect 30530 40272 30594 40276
rect 35618 40332 35682 40336
rect 35618 40276 35622 40332
rect 35622 40276 35678 40332
rect 35678 40276 35682 40332
rect 35618 40272 35682 40276
rect 35698 40332 35762 40336
rect 35698 40276 35702 40332
rect 35702 40276 35758 40332
rect 35758 40276 35762 40332
rect 35698 40272 35762 40276
rect 35778 40332 35842 40336
rect 35778 40276 35782 40332
rect 35782 40276 35838 40332
rect 35838 40276 35842 40332
rect 35778 40272 35842 40276
rect 35858 40332 35922 40336
rect 35858 40276 35862 40332
rect 35862 40276 35918 40332
rect 35918 40276 35922 40332
rect 35858 40272 35922 40276
rect 40946 40332 41010 40336
rect 40946 40276 40950 40332
rect 40950 40276 41006 40332
rect 41006 40276 41010 40332
rect 40946 40272 41010 40276
rect 41026 40332 41090 40336
rect 41026 40276 41030 40332
rect 41030 40276 41086 40332
rect 41086 40276 41090 40332
rect 41026 40272 41090 40276
rect 41106 40332 41170 40336
rect 41106 40276 41110 40332
rect 41110 40276 41166 40332
rect 41166 40276 41170 40332
rect 41106 40272 41170 40276
rect 41186 40332 41250 40336
rect 41186 40276 41190 40332
rect 41190 40276 41246 40332
rect 41246 40276 41250 40332
rect 41186 40272 41250 40276
rect 46274 40332 46338 40336
rect 46274 40276 46278 40332
rect 46278 40276 46334 40332
rect 46334 40276 46338 40332
rect 46274 40272 46338 40276
rect 46354 40332 46418 40336
rect 46354 40276 46358 40332
rect 46358 40276 46414 40332
rect 46414 40276 46418 40332
rect 46354 40272 46418 40276
rect 46434 40332 46498 40336
rect 46434 40276 46438 40332
rect 46438 40276 46494 40332
rect 46494 40276 46498 40332
rect 46434 40272 46498 40276
rect 46514 40332 46578 40336
rect 46514 40276 46518 40332
rect 46518 40276 46574 40332
rect 46574 40276 46578 40332
rect 46514 40272 46578 40276
rect 51602 40332 51666 40336
rect 51602 40276 51606 40332
rect 51606 40276 51662 40332
rect 51662 40276 51666 40332
rect 51602 40272 51666 40276
rect 51682 40332 51746 40336
rect 51682 40276 51686 40332
rect 51686 40276 51742 40332
rect 51742 40276 51746 40332
rect 51682 40272 51746 40276
rect 51762 40332 51826 40336
rect 51762 40276 51766 40332
rect 51766 40276 51822 40332
rect 51822 40276 51826 40332
rect 51762 40272 51826 40276
rect 51842 40332 51906 40336
rect 51842 40276 51846 40332
rect 51846 40276 51902 40332
rect 51902 40276 51906 40332
rect 51842 40272 51906 40276
rect 56930 40332 56994 40336
rect 56930 40276 56934 40332
rect 56934 40276 56990 40332
rect 56990 40276 56994 40332
rect 56930 40272 56994 40276
rect 57010 40332 57074 40336
rect 57010 40276 57014 40332
rect 57014 40276 57070 40332
rect 57070 40276 57074 40332
rect 57010 40272 57074 40276
rect 57090 40332 57154 40336
rect 57090 40276 57094 40332
rect 57094 40276 57150 40332
rect 57150 40276 57154 40332
rect 57090 40272 57154 40276
rect 57170 40332 57234 40336
rect 57170 40276 57174 40332
rect 57174 40276 57230 40332
rect 57230 40276 57234 40332
rect 57170 40272 57234 40276
rect 62258 40332 62322 40336
rect 62258 40276 62262 40332
rect 62262 40276 62318 40332
rect 62318 40276 62322 40332
rect 62258 40272 62322 40276
rect 62338 40332 62402 40336
rect 62338 40276 62342 40332
rect 62342 40276 62398 40332
rect 62398 40276 62402 40332
rect 62338 40272 62402 40276
rect 62418 40332 62482 40336
rect 62418 40276 62422 40332
rect 62422 40276 62478 40332
rect 62478 40276 62482 40332
rect 62418 40272 62482 40276
rect 62498 40332 62562 40336
rect 62498 40276 62502 40332
rect 62502 40276 62558 40332
rect 62558 40276 62562 40332
rect 62498 40272 62562 40276
rect 67586 40332 67650 40336
rect 67586 40276 67590 40332
rect 67590 40276 67646 40332
rect 67646 40276 67650 40332
rect 67586 40272 67650 40276
rect 67666 40332 67730 40336
rect 67666 40276 67670 40332
rect 67670 40276 67726 40332
rect 67726 40276 67730 40332
rect 67666 40272 67730 40276
rect 67746 40332 67810 40336
rect 67746 40276 67750 40332
rect 67750 40276 67806 40332
rect 67806 40276 67810 40332
rect 67746 40272 67810 40276
rect 67826 40332 67890 40336
rect 67826 40276 67830 40332
rect 67830 40276 67886 40332
rect 67886 40276 67890 40332
rect 67826 40272 67890 40276
rect 72914 40332 72978 40336
rect 72914 40276 72918 40332
rect 72918 40276 72974 40332
rect 72974 40276 72978 40332
rect 72914 40272 72978 40276
rect 72994 40332 73058 40336
rect 72994 40276 72998 40332
rect 72998 40276 73054 40332
rect 73054 40276 73058 40332
rect 72994 40272 73058 40276
rect 73074 40332 73138 40336
rect 73074 40276 73078 40332
rect 73078 40276 73134 40332
rect 73134 40276 73138 40332
rect 73074 40272 73138 40276
rect 73154 40332 73218 40336
rect 73154 40276 73158 40332
rect 73158 40276 73214 40332
rect 73214 40276 73218 40332
rect 73154 40272 73218 40276
rect 78242 40332 78306 40336
rect 78242 40276 78246 40332
rect 78246 40276 78302 40332
rect 78302 40276 78306 40332
rect 78242 40272 78306 40276
rect 78322 40332 78386 40336
rect 78322 40276 78326 40332
rect 78326 40276 78382 40332
rect 78382 40276 78386 40332
rect 78322 40272 78386 40276
rect 78402 40332 78466 40336
rect 78402 40276 78406 40332
rect 78406 40276 78462 40332
rect 78462 40276 78466 40332
rect 78402 40272 78466 40276
rect 78482 40332 78546 40336
rect 78482 40276 78486 40332
rect 78486 40276 78542 40332
rect 78542 40276 78546 40332
rect 78482 40272 78546 40276
rect 83570 40332 83634 40336
rect 83570 40276 83574 40332
rect 83574 40276 83630 40332
rect 83630 40276 83634 40332
rect 83570 40272 83634 40276
rect 83650 40332 83714 40336
rect 83650 40276 83654 40332
rect 83654 40276 83710 40332
rect 83710 40276 83714 40332
rect 83650 40272 83714 40276
rect 83730 40332 83794 40336
rect 83730 40276 83734 40332
rect 83734 40276 83790 40332
rect 83790 40276 83794 40332
rect 83730 40272 83794 40276
rect 83810 40332 83874 40336
rect 83810 40276 83814 40332
rect 83814 40276 83870 40332
rect 83870 40276 83874 40332
rect 83810 40272 83874 40276
rect 88898 40332 88962 40336
rect 88898 40276 88902 40332
rect 88902 40276 88958 40332
rect 88958 40276 88962 40332
rect 88898 40272 88962 40276
rect 88978 40332 89042 40336
rect 88978 40276 88982 40332
rect 88982 40276 89038 40332
rect 89038 40276 89042 40332
rect 88978 40272 89042 40276
rect 89058 40332 89122 40336
rect 89058 40276 89062 40332
rect 89062 40276 89118 40332
rect 89118 40276 89122 40332
rect 89058 40272 89122 40276
rect 89138 40332 89202 40336
rect 89138 40276 89142 40332
rect 89142 40276 89198 40332
rect 89198 40276 89202 40332
rect 89138 40272 89202 40276
rect 6314 39788 6378 39792
rect 6314 39732 6318 39788
rect 6318 39732 6374 39788
rect 6374 39732 6378 39788
rect 6314 39728 6378 39732
rect 6394 39788 6458 39792
rect 6394 39732 6398 39788
rect 6398 39732 6454 39788
rect 6454 39732 6458 39788
rect 6394 39728 6458 39732
rect 6474 39788 6538 39792
rect 6474 39732 6478 39788
rect 6478 39732 6534 39788
rect 6534 39732 6538 39788
rect 6474 39728 6538 39732
rect 6554 39788 6618 39792
rect 6554 39732 6558 39788
rect 6558 39732 6614 39788
rect 6614 39732 6618 39788
rect 6554 39728 6618 39732
rect 11642 39788 11706 39792
rect 11642 39732 11646 39788
rect 11646 39732 11702 39788
rect 11702 39732 11706 39788
rect 11642 39728 11706 39732
rect 11722 39788 11786 39792
rect 11722 39732 11726 39788
rect 11726 39732 11782 39788
rect 11782 39732 11786 39788
rect 11722 39728 11786 39732
rect 11802 39788 11866 39792
rect 11802 39732 11806 39788
rect 11806 39732 11862 39788
rect 11862 39732 11866 39788
rect 11802 39728 11866 39732
rect 11882 39788 11946 39792
rect 11882 39732 11886 39788
rect 11886 39732 11942 39788
rect 11942 39732 11946 39788
rect 11882 39728 11946 39732
rect 16970 39788 17034 39792
rect 16970 39732 16974 39788
rect 16974 39732 17030 39788
rect 17030 39732 17034 39788
rect 16970 39728 17034 39732
rect 17050 39788 17114 39792
rect 17050 39732 17054 39788
rect 17054 39732 17110 39788
rect 17110 39732 17114 39788
rect 17050 39728 17114 39732
rect 17130 39788 17194 39792
rect 17130 39732 17134 39788
rect 17134 39732 17190 39788
rect 17190 39732 17194 39788
rect 17130 39728 17194 39732
rect 17210 39788 17274 39792
rect 17210 39732 17214 39788
rect 17214 39732 17270 39788
rect 17270 39732 17274 39788
rect 17210 39728 17274 39732
rect 22298 39788 22362 39792
rect 22298 39732 22302 39788
rect 22302 39732 22358 39788
rect 22358 39732 22362 39788
rect 22298 39728 22362 39732
rect 22378 39788 22442 39792
rect 22378 39732 22382 39788
rect 22382 39732 22438 39788
rect 22438 39732 22442 39788
rect 22378 39728 22442 39732
rect 22458 39788 22522 39792
rect 22458 39732 22462 39788
rect 22462 39732 22518 39788
rect 22518 39732 22522 39788
rect 22458 39728 22522 39732
rect 22538 39788 22602 39792
rect 22538 39732 22542 39788
rect 22542 39732 22598 39788
rect 22598 39732 22602 39788
rect 22538 39728 22602 39732
rect 27626 39788 27690 39792
rect 27626 39732 27630 39788
rect 27630 39732 27686 39788
rect 27686 39732 27690 39788
rect 27626 39728 27690 39732
rect 27706 39788 27770 39792
rect 27706 39732 27710 39788
rect 27710 39732 27766 39788
rect 27766 39732 27770 39788
rect 27706 39728 27770 39732
rect 27786 39788 27850 39792
rect 27786 39732 27790 39788
rect 27790 39732 27846 39788
rect 27846 39732 27850 39788
rect 27786 39728 27850 39732
rect 27866 39788 27930 39792
rect 27866 39732 27870 39788
rect 27870 39732 27926 39788
rect 27926 39732 27930 39788
rect 27866 39728 27930 39732
rect 32954 39788 33018 39792
rect 32954 39732 32958 39788
rect 32958 39732 33014 39788
rect 33014 39732 33018 39788
rect 32954 39728 33018 39732
rect 33034 39788 33098 39792
rect 33034 39732 33038 39788
rect 33038 39732 33094 39788
rect 33094 39732 33098 39788
rect 33034 39728 33098 39732
rect 33114 39788 33178 39792
rect 33114 39732 33118 39788
rect 33118 39732 33174 39788
rect 33174 39732 33178 39788
rect 33114 39728 33178 39732
rect 33194 39788 33258 39792
rect 33194 39732 33198 39788
rect 33198 39732 33254 39788
rect 33254 39732 33258 39788
rect 33194 39728 33258 39732
rect 38282 39788 38346 39792
rect 38282 39732 38286 39788
rect 38286 39732 38342 39788
rect 38342 39732 38346 39788
rect 38282 39728 38346 39732
rect 38362 39788 38426 39792
rect 38362 39732 38366 39788
rect 38366 39732 38422 39788
rect 38422 39732 38426 39788
rect 38362 39728 38426 39732
rect 38442 39788 38506 39792
rect 38442 39732 38446 39788
rect 38446 39732 38502 39788
rect 38502 39732 38506 39788
rect 38442 39728 38506 39732
rect 38522 39788 38586 39792
rect 38522 39732 38526 39788
rect 38526 39732 38582 39788
rect 38582 39732 38586 39788
rect 38522 39728 38586 39732
rect 43610 39788 43674 39792
rect 43610 39732 43614 39788
rect 43614 39732 43670 39788
rect 43670 39732 43674 39788
rect 43610 39728 43674 39732
rect 43690 39788 43754 39792
rect 43690 39732 43694 39788
rect 43694 39732 43750 39788
rect 43750 39732 43754 39788
rect 43690 39728 43754 39732
rect 43770 39788 43834 39792
rect 43770 39732 43774 39788
rect 43774 39732 43830 39788
rect 43830 39732 43834 39788
rect 43770 39728 43834 39732
rect 43850 39788 43914 39792
rect 43850 39732 43854 39788
rect 43854 39732 43910 39788
rect 43910 39732 43914 39788
rect 43850 39728 43914 39732
rect 48938 39788 49002 39792
rect 48938 39732 48942 39788
rect 48942 39732 48998 39788
rect 48998 39732 49002 39788
rect 48938 39728 49002 39732
rect 49018 39788 49082 39792
rect 49018 39732 49022 39788
rect 49022 39732 49078 39788
rect 49078 39732 49082 39788
rect 49018 39728 49082 39732
rect 49098 39788 49162 39792
rect 49098 39732 49102 39788
rect 49102 39732 49158 39788
rect 49158 39732 49162 39788
rect 49098 39728 49162 39732
rect 49178 39788 49242 39792
rect 49178 39732 49182 39788
rect 49182 39732 49238 39788
rect 49238 39732 49242 39788
rect 49178 39728 49242 39732
rect 54266 39788 54330 39792
rect 54266 39732 54270 39788
rect 54270 39732 54326 39788
rect 54326 39732 54330 39788
rect 54266 39728 54330 39732
rect 54346 39788 54410 39792
rect 54346 39732 54350 39788
rect 54350 39732 54406 39788
rect 54406 39732 54410 39788
rect 54346 39728 54410 39732
rect 54426 39788 54490 39792
rect 54426 39732 54430 39788
rect 54430 39732 54486 39788
rect 54486 39732 54490 39788
rect 54426 39728 54490 39732
rect 54506 39788 54570 39792
rect 54506 39732 54510 39788
rect 54510 39732 54566 39788
rect 54566 39732 54570 39788
rect 54506 39728 54570 39732
rect 59594 39788 59658 39792
rect 59594 39732 59598 39788
rect 59598 39732 59654 39788
rect 59654 39732 59658 39788
rect 59594 39728 59658 39732
rect 59674 39788 59738 39792
rect 59674 39732 59678 39788
rect 59678 39732 59734 39788
rect 59734 39732 59738 39788
rect 59674 39728 59738 39732
rect 59754 39788 59818 39792
rect 59754 39732 59758 39788
rect 59758 39732 59814 39788
rect 59814 39732 59818 39788
rect 59754 39728 59818 39732
rect 59834 39788 59898 39792
rect 59834 39732 59838 39788
rect 59838 39732 59894 39788
rect 59894 39732 59898 39788
rect 59834 39728 59898 39732
rect 64922 39788 64986 39792
rect 64922 39732 64926 39788
rect 64926 39732 64982 39788
rect 64982 39732 64986 39788
rect 64922 39728 64986 39732
rect 65002 39788 65066 39792
rect 65002 39732 65006 39788
rect 65006 39732 65062 39788
rect 65062 39732 65066 39788
rect 65002 39728 65066 39732
rect 65082 39788 65146 39792
rect 65082 39732 65086 39788
rect 65086 39732 65142 39788
rect 65142 39732 65146 39788
rect 65082 39728 65146 39732
rect 65162 39788 65226 39792
rect 65162 39732 65166 39788
rect 65166 39732 65222 39788
rect 65222 39732 65226 39788
rect 65162 39728 65226 39732
rect 70250 39788 70314 39792
rect 70250 39732 70254 39788
rect 70254 39732 70310 39788
rect 70310 39732 70314 39788
rect 70250 39728 70314 39732
rect 70330 39788 70394 39792
rect 70330 39732 70334 39788
rect 70334 39732 70390 39788
rect 70390 39732 70394 39788
rect 70330 39728 70394 39732
rect 70410 39788 70474 39792
rect 70410 39732 70414 39788
rect 70414 39732 70470 39788
rect 70470 39732 70474 39788
rect 70410 39728 70474 39732
rect 70490 39788 70554 39792
rect 70490 39732 70494 39788
rect 70494 39732 70550 39788
rect 70550 39732 70554 39788
rect 70490 39728 70554 39732
rect 75578 39788 75642 39792
rect 75578 39732 75582 39788
rect 75582 39732 75638 39788
rect 75638 39732 75642 39788
rect 75578 39728 75642 39732
rect 75658 39788 75722 39792
rect 75658 39732 75662 39788
rect 75662 39732 75718 39788
rect 75718 39732 75722 39788
rect 75658 39728 75722 39732
rect 75738 39788 75802 39792
rect 75738 39732 75742 39788
rect 75742 39732 75798 39788
rect 75798 39732 75802 39788
rect 75738 39728 75802 39732
rect 75818 39788 75882 39792
rect 75818 39732 75822 39788
rect 75822 39732 75878 39788
rect 75878 39732 75882 39788
rect 75818 39728 75882 39732
rect 80906 39788 80970 39792
rect 80906 39732 80910 39788
rect 80910 39732 80966 39788
rect 80966 39732 80970 39788
rect 80906 39728 80970 39732
rect 80986 39788 81050 39792
rect 80986 39732 80990 39788
rect 80990 39732 81046 39788
rect 81046 39732 81050 39788
rect 80986 39728 81050 39732
rect 81066 39788 81130 39792
rect 81066 39732 81070 39788
rect 81070 39732 81126 39788
rect 81126 39732 81130 39788
rect 81066 39728 81130 39732
rect 81146 39788 81210 39792
rect 81146 39732 81150 39788
rect 81150 39732 81206 39788
rect 81206 39732 81210 39788
rect 81146 39728 81210 39732
rect 86234 39788 86298 39792
rect 86234 39732 86238 39788
rect 86238 39732 86294 39788
rect 86294 39732 86298 39788
rect 86234 39728 86298 39732
rect 86314 39788 86378 39792
rect 86314 39732 86318 39788
rect 86318 39732 86374 39788
rect 86374 39732 86378 39788
rect 86314 39728 86378 39732
rect 86394 39788 86458 39792
rect 86394 39732 86398 39788
rect 86398 39732 86454 39788
rect 86454 39732 86458 39788
rect 86394 39728 86458 39732
rect 86474 39788 86538 39792
rect 86474 39732 86478 39788
rect 86478 39732 86534 39788
rect 86534 39732 86538 39788
rect 86474 39728 86538 39732
rect 91562 39788 91626 39792
rect 91562 39732 91566 39788
rect 91566 39732 91622 39788
rect 91622 39732 91626 39788
rect 91562 39728 91626 39732
rect 91642 39788 91706 39792
rect 91642 39732 91646 39788
rect 91646 39732 91702 39788
rect 91702 39732 91706 39788
rect 91642 39728 91706 39732
rect 91722 39788 91786 39792
rect 91722 39732 91726 39788
rect 91726 39732 91782 39788
rect 91782 39732 91786 39788
rect 91722 39728 91786 39732
rect 91802 39788 91866 39792
rect 91802 39732 91806 39788
rect 91806 39732 91862 39788
rect 91862 39732 91866 39788
rect 91802 39728 91866 39732
rect 3650 39244 3714 39248
rect 3650 39188 3654 39244
rect 3654 39188 3710 39244
rect 3710 39188 3714 39244
rect 3650 39184 3714 39188
rect 3730 39244 3794 39248
rect 3730 39188 3734 39244
rect 3734 39188 3790 39244
rect 3790 39188 3794 39244
rect 3730 39184 3794 39188
rect 3810 39244 3874 39248
rect 3810 39188 3814 39244
rect 3814 39188 3870 39244
rect 3870 39188 3874 39244
rect 3810 39184 3874 39188
rect 3890 39244 3954 39248
rect 3890 39188 3894 39244
rect 3894 39188 3950 39244
rect 3950 39188 3954 39244
rect 3890 39184 3954 39188
rect 8978 39244 9042 39248
rect 8978 39188 8982 39244
rect 8982 39188 9038 39244
rect 9038 39188 9042 39244
rect 8978 39184 9042 39188
rect 9058 39244 9122 39248
rect 9058 39188 9062 39244
rect 9062 39188 9118 39244
rect 9118 39188 9122 39244
rect 9058 39184 9122 39188
rect 9138 39244 9202 39248
rect 9138 39188 9142 39244
rect 9142 39188 9198 39244
rect 9198 39188 9202 39244
rect 9138 39184 9202 39188
rect 9218 39244 9282 39248
rect 9218 39188 9222 39244
rect 9222 39188 9278 39244
rect 9278 39188 9282 39244
rect 9218 39184 9282 39188
rect 14306 39244 14370 39248
rect 14306 39188 14310 39244
rect 14310 39188 14366 39244
rect 14366 39188 14370 39244
rect 14306 39184 14370 39188
rect 14386 39244 14450 39248
rect 14386 39188 14390 39244
rect 14390 39188 14446 39244
rect 14446 39188 14450 39244
rect 14386 39184 14450 39188
rect 14466 39244 14530 39248
rect 14466 39188 14470 39244
rect 14470 39188 14526 39244
rect 14526 39188 14530 39244
rect 14466 39184 14530 39188
rect 14546 39244 14610 39248
rect 14546 39188 14550 39244
rect 14550 39188 14606 39244
rect 14606 39188 14610 39244
rect 14546 39184 14610 39188
rect 19634 39244 19698 39248
rect 19634 39188 19638 39244
rect 19638 39188 19694 39244
rect 19694 39188 19698 39244
rect 19634 39184 19698 39188
rect 19714 39244 19778 39248
rect 19714 39188 19718 39244
rect 19718 39188 19774 39244
rect 19774 39188 19778 39244
rect 19714 39184 19778 39188
rect 19794 39244 19858 39248
rect 19794 39188 19798 39244
rect 19798 39188 19854 39244
rect 19854 39188 19858 39244
rect 19794 39184 19858 39188
rect 19874 39244 19938 39248
rect 19874 39188 19878 39244
rect 19878 39188 19934 39244
rect 19934 39188 19938 39244
rect 19874 39184 19938 39188
rect 24962 39244 25026 39248
rect 24962 39188 24966 39244
rect 24966 39188 25022 39244
rect 25022 39188 25026 39244
rect 24962 39184 25026 39188
rect 25042 39244 25106 39248
rect 25042 39188 25046 39244
rect 25046 39188 25102 39244
rect 25102 39188 25106 39244
rect 25042 39184 25106 39188
rect 25122 39244 25186 39248
rect 25122 39188 25126 39244
rect 25126 39188 25182 39244
rect 25182 39188 25186 39244
rect 25122 39184 25186 39188
rect 25202 39244 25266 39248
rect 25202 39188 25206 39244
rect 25206 39188 25262 39244
rect 25262 39188 25266 39244
rect 25202 39184 25266 39188
rect 30290 39244 30354 39248
rect 30290 39188 30294 39244
rect 30294 39188 30350 39244
rect 30350 39188 30354 39244
rect 30290 39184 30354 39188
rect 30370 39244 30434 39248
rect 30370 39188 30374 39244
rect 30374 39188 30430 39244
rect 30430 39188 30434 39244
rect 30370 39184 30434 39188
rect 30450 39244 30514 39248
rect 30450 39188 30454 39244
rect 30454 39188 30510 39244
rect 30510 39188 30514 39244
rect 30450 39184 30514 39188
rect 30530 39244 30594 39248
rect 30530 39188 30534 39244
rect 30534 39188 30590 39244
rect 30590 39188 30594 39244
rect 30530 39184 30594 39188
rect 35618 39244 35682 39248
rect 35618 39188 35622 39244
rect 35622 39188 35678 39244
rect 35678 39188 35682 39244
rect 35618 39184 35682 39188
rect 35698 39244 35762 39248
rect 35698 39188 35702 39244
rect 35702 39188 35758 39244
rect 35758 39188 35762 39244
rect 35698 39184 35762 39188
rect 35778 39244 35842 39248
rect 35778 39188 35782 39244
rect 35782 39188 35838 39244
rect 35838 39188 35842 39244
rect 35778 39184 35842 39188
rect 35858 39244 35922 39248
rect 35858 39188 35862 39244
rect 35862 39188 35918 39244
rect 35918 39188 35922 39244
rect 35858 39184 35922 39188
rect 40946 39244 41010 39248
rect 40946 39188 40950 39244
rect 40950 39188 41006 39244
rect 41006 39188 41010 39244
rect 40946 39184 41010 39188
rect 41026 39244 41090 39248
rect 41026 39188 41030 39244
rect 41030 39188 41086 39244
rect 41086 39188 41090 39244
rect 41026 39184 41090 39188
rect 41106 39244 41170 39248
rect 41106 39188 41110 39244
rect 41110 39188 41166 39244
rect 41166 39188 41170 39244
rect 41106 39184 41170 39188
rect 41186 39244 41250 39248
rect 41186 39188 41190 39244
rect 41190 39188 41246 39244
rect 41246 39188 41250 39244
rect 41186 39184 41250 39188
rect 46274 39244 46338 39248
rect 46274 39188 46278 39244
rect 46278 39188 46334 39244
rect 46334 39188 46338 39244
rect 46274 39184 46338 39188
rect 46354 39244 46418 39248
rect 46354 39188 46358 39244
rect 46358 39188 46414 39244
rect 46414 39188 46418 39244
rect 46354 39184 46418 39188
rect 46434 39244 46498 39248
rect 46434 39188 46438 39244
rect 46438 39188 46494 39244
rect 46494 39188 46498 39244
rect 46434 39184 46498 39188
rect 46514 39244 46578 39248
rect 46514 39188 46518 39244
rect 46518 39188 46574 39244
rect 46574 39188 46578 39244
rect 46514 39184 46578 39188
rect 51602 39244 51666 39248
rect 51602 39188 51606 39244
rect 51606 39188 51662 39244
rect 51662 39188 51666 39244
rect 51602 39184 51666 39188
rect 51682 39244 51746 39248
rect 51682 39188 51686 39244
rect 51686 39188 51742 39244
rect 51742 39188 51746 39244
rect 51682 39184 51746 39188
rect 51762 39244 51826 39248
rect 51762 39188 51766 39244
rect 51766 39188 51822 39244
rect 51822 39188 51826 39244
rect 51762 39184 51826 39188
rect 51842 39244 51906 39248
rect 51842 39188 51846 39244
rect 51846 39188 51902 39244
rect 51902 39188 51906 39244
rect 51842 39184 51906 39188
rect 56930 39244 56994 39248
rect 56930 39188 56934 39244
rect 56934 39188 56990 39244
rect 56990 39188 56994 39244
rect 56930 39184 56994 39188
rect 57010 39244 57074 39248
rect 57010 39188 57014 39244
rect 57014 39188 57070 39244
rect 57070 39188 57074 39244
rect 57010 39184 57074 39188
rect 57090 39244 57154 39248
rect 57090 39188 57094 39244
rect 57094 39188 57150 39244
rect 57150 39188 57154 39244
rect 57090 39184 57154 39188
rect 57170 39244 57234 39248
rect 57170 39188 57174 39244
rect 57174 39188 57230 39244
rect 57230 39188 57234 39244
rect 57170 39184 57234 39188
rect 62258 39244 62322 39248
rect 62258 39188 62262 39244
rect 62262 39188 62318 39244
rect 62318 39188 62322 39244
rect 62258 39184 62322 39188
rect 62338 39244 62402 39248
rect 62338 39188 62342 39244
rect 62342 39188 62398 39244
rect 62398 39188 62402 39244
rect 62338 39184 62402 39188
rect 62418 39244 62482 39248
rect 62418 39188 62422 39244
rect 62422 39188 62478 39244
rect 62478 39188 62482 39244
rect 62418 39184 62482 39188
rect 62498 39244 62562 39248
rect 62498 39188 62502 39244
rect 62502 39188 62558 39244
rect 62558 39188 62562 39244
rect 62498 39184 62562 39188
rect 67586 39244 67650 39248
rect 67586 39188 67590 39244
rect 67590 39188 67646 39244
rect 67646 39188 67650 39244
rect 67586 39184 67650 39188
rect 67666 39244 67730 39248
rect 67666 39188 67670 39244
rect 67670 39188 67726 39244
rect 67726 39188 67730 39244
rect 67666 39184 67730 39188
rect 67746 39244 67810 39248
rect 67746 39188 67750 39244
rect 67750 39188 67806 39244
rect 67806 39188 67810 39244
rect 67746 39184 67810 39188
rect 67826 39244 67890 39248
rect 67826 39188 67830 39244
rect 67830 39188 67886 39244
rect 67886 39188 67890 39244
rect 67826 39184 67890 39188
rect 72914 39244 72978 39248
rect 72914 39188 72918 39244
rect 72918 39188 72974 39244
rect 72974 39188 72978 39244
rect 72914 39184 72978 39188
rect 72994 39244 73058 39248
rect 72994 39188 72998 39244
rect 72998 39188 73054 39244
rect 73054 39188 73058 39244
rect 72994 39184 73058 39188
rect 73074 39244 73138 39248
rect 73074 39188 73078 39244
rect 73078 39188 73134 39244
rect 73134 39188 73138 39244
rect 73074 39184 73138 39188
rect 73154 39244 73218 39248
rect 73154 39188 73158 39244
rect 73158 39188 73214 39244
rect 73214 39188 73218 39244
rect 73154 39184 73218 39188
rect 78242 39244 78306 39248
rect 78242 39188 78246 39244
rect 78246 39188 78302 39244
rect 78302 39188 78306 39244
rect 78242 39184 78306 39188
rect 78322 39244 78386 39248
rect 78322 39188 78326 39244
rect 78326 39188 78382 39244
rect 78382 39188 78386 39244
rect 78322 39184 78386 39188
rect 78402 39244 78466 39248
rect 78402 39188 78406 39244
rect 78406 39188 78462 39244
rect 78462 39188 78466 39244
rect 78402 39184 78466 39188
rect 78482 39244 78546 39248
rect 78482 39188 78486 39244
rect 78486 39188 78542 39244
rect 78542 39188 78546 39244
rect 78482 39184 78546 39188
rect 83570 39244 83634 39248
rect 83570 39188 83574 39244
rect 83574 39188 83630 39244
rect 83630 39188 83634 39244
rect 83570 39184 83634 39188
rect 83650 39244 83714 39248
rect 83650 39188 83654 39244
rect 83654 39188 83710 39244
rect 83710 39188 83714 39244
rect 83650 39184 83714 39188
rect 83730 39244 83794 39248
rect 83730 39188 83734 39244
rect 83734 39188 83790 39244
rect 83790 39188 83794 39244
rect 83730 39184 83794 39188
rect 83810 39244 83874 39248
rect 83810 39188 83814 39244
rect 83814 39188 83870 39244
rect 83870 39188 83874 39244
rect 83810 39184 83874 39188
rect 88898 39244 88962 39248
rect 88898 39188 88902 39244
rect 88902 39188 88958 39244
rect 88958 39188 88962 39244
rect 88898 39184 88962 39188
rect 88978 39244 89042 39248
rect 88978 39188 88982 39244
rect 88982 39188 89038 39244
rect 89038 39188 89042 39244
rect 88978 39184 89042 39188
rect 89058 39244 89122 39248
rect 89058 39188 89062 39244
rect 89062 39188 89118 39244
rect 89118 39188 89122 39244
rect 89058 39184 89122 39188
rect 89138 39244 89202 39248
rect 89138 39188 89142 39244
rect 89142 39188 89198 39244
rect 89198 39188 89202 39244
rect 89138 39184 89202 39188
rect 6314 38700 6378 38704
rect 6314 38644 6318 38700
rect 6318 38644 6374 38700
rect 6374 38644 6378 38700
rect 6314 38640 6378 38644
rect 6394 38700 6458 38704
rect 6394 38644 6398 38700
rect 6398 38644 6454 38700
rect 6454 38644 6458 38700
rect 6394 38640 6458 38644
rect 6474 38700 6538 38704
rect 6474 38644 6478 38700
rect 6478 38644 6534 38700
rect 6534 38644 6538 38700
rect 6474 38640 6538 38644
rect 6554 38700 6618 38704
rect 6554 38644 6558 38700
rect 6558 38644 6614 38700
rect 6614 38644 6618 38700
rect 6554 38640 6618 38644
rect 11642 38700 11706 38704
rect 11642 38644 11646 38700
rect 11646 38644 11702 38700
rect 11702 38644 11706 38700
rect 11642 38640 11706 38644
rect 11722 38700 11786 38704
rect 11722 38644 11726 38700
rect 11726 38644 11782 38700
rect 11782 38644 11786 38700
rect 11722 38640 11786 38644
rect 11802 38700 11866 38704
rect 11802 38644 11806 38700
rect 11806 38644 11862 38700
rect 11862 38644 11866 38700
rect 11802 38640 11866 38644
rect 11882 38700 11946 38704
rect 11882 38644 11886 38700
rect 11886 38644 11942 38700
rect 11942 38644 11946 38700
rect 11882 38640 11946 38644
rect 16970 38700 17034 38704
rect 16970 38644 16974 38700
rect 16974 38644 17030 38700
rect 17030 38644 17034 38700
rect 16970 38640 17034 38644
rect 17050 38700 17114 38704
rect 17050 38644 17054 38700
rect 17054 38644 17110 38700
rect 17110 38644 17114 38700
rect 17050 38640 17114 38644
rect 17130 38700 17194 38704
rect 17130 38644 17134 38700
rect 17134 38644 17190 38700
rect 17190 38644 17194 38700
rect 17130 38640 17194 38644
rect 17210 38700 17274 38704
rect 17210 38644 17214 38700
rect 17214 38644 17270 38700
rect 17270 38644 17274 38700
rect 17210 38640 17274 38644
rect 22298 38700 22362 38704
rect 22298 38644 22302 38700
rect 22302 38644 22358 38700
rect 22358 38644 22362 38700
rect 22298 38640 22362 38644
rect 22378 38700 22442 38704
rect 22378 38644 22382 38700
rect 22382 38644 22438 38700
rect 22438 38644 22442 38700
rect 22378 38640 22442 38644
rect 22458 38700 22522 38704
rect 22458 38644 22462 38700
rect 22462 38644 22518 38700
rect 22518 38644 22522 38700
rect 22458 38640 22522 38644
rect 22538 38700 22602 38704
rect 22538 38644 22542 38700
rect 22542 38644 22598 38700
rect 22598 38644 22602 38700
rect 22538 38640 22602 38644
rect 27626 38700 27690 38704
rect 27626 38644 27630 38700
rect 27630 38644 27686 38700
rect 27686 38644 27690 38700
rect 27626 38640 27690 38644
rect 27706 38700 27770 38704
rect 27706 38644 27710 38700
rect 27710 38644 27766 38700
rect 27766 38644 27770 38700
rect 27706 38640 27770 38644
rect 27786 38700 27850 38704
rect 27786 38644 27790 38700
rect 27790 38644 27846 38700
rect 27846 38644 27850 38700
rect 27786 38640 27850 38644
rect 27866 38700 27930 38704
rect 27866 38644 27870 38700
rect 27870 38644 27926 38700
rect 27926 38644 27930 38700
rect 27866 38640 27930 38644
rect 32954 38700 33018 38704
rect 32954 38644 32958 38700
rect 32958 38644 33014 38700
rect 33014 38644 33018 38700
rect 32954 38640 33018 38644
rect 33034 38700 33098 38704
rect 33034 38644 33038 38700
rect 33038 38644 33094 38700
rect 33094 38644 33098 38700
rect 33034 38640 33098 38644
rect 33114 38700 33178 38704
rect 33114 38644 33118 38700
rect 33118 38644 33174 38700
rect 33174 38644 33178 38700
rect 33114 38640 33178 38644
rect 33194 38700 33258 38704
rect 33194 38644 33198 38700
rect 33198 38644 33254 38700
rect 33254 38644 33258 38700
rect 33194 38640 33258 38644
rect 38282 38700 38346 38704
rect 38282 38644 38286 38700
rect 38286 38644 38342 38700
rect 38342 38644 38346 38700
rect 38282 38640 38346 38644
rect 38362 38700 38426 38704
rect 38362 38644 38366 38700
rect 38366 38644 38422 38700
rect 38422 38644 38426 38700
rect 38362 38640 38426 38644
rect 38442 38700 38506 38704
rect 38442 38644 38446 38700
rect 38446 38644 38502 38700
rect 38502 38644 38506 38700
rect 38442 38640 38506 38644
rect 38522 38700 38586 38704
rect 38522 38644 38526 38700
rect 38526 38644 38582 38700
rect 38582 38644 38586 38700
rect 38522 38640 38586 38644
rect 43610 38700 43674 38704
rect 43610 38644 43614 38700
rect 43614 38644 43670 38700
rect 43670 38644 43674 38700
rect 43610 38640 43674 38644
rect 43690 38700 43754 38704
rect 43690 38644 43694 38700
rect 43694 38644 43750 38700
rect 43750 38644 43754 38700
rect 43690 38640 43754 38644
rect 43770 38700 43834 38704
rect 43770 38644 43774 38700
rect 43774 38644 43830 38700
rect 43830 38644 43834 38700
rect 43770 38640 43834 38644
rect 43850 38700 43914 38704
rect 43850 38644 43854 38700
rect 43854 38644 43910 38700
rect 43910 38644 43914 38700
rect 43850 38640 43914 38644
rect 48938 38700 49002 38704
rect 48938 38644 48942 38700
rect 48942 38644 48998 38700
rect 48998 38644 49002 38700
rect 48938 38640 49002 38644
rect 49018 38700 49082 38704
rect 49018 38644 49022 38700
rect 49022 38644 49078 38700
rect 49078 38644 49082 38700
rect 49018 38640 49082 38644
rect 49098 38700 49162 38704
rect 49098 38644 49102 38700
rect 49102 38644 49158 38700
rect 49158 38644 49162 38700
rect 49098 38640 49162 38644
rect 49178 38700 49242 38704
rect 49178 38644 49182 38700
rect 49182 38644 49238 38700
rect 49238 38644 49242 38700
rect 49178 38640 49242 38644
rect 54266 38700 54330 38704
rect 54266 38644 54270 38700
rect 54270 38644 54326 38700
rect 54326 38644 54330 38700
rect 54266 38640 54330 38644
rect 54346 38700 54410 38704
rect 54346 38644 54350 38700
rect 54350 38644 54406 38700
rect 54406 38644 54410 38700
rect 54346 38640 54410 38644
rect 54426 38700 54490 38704
rect 54426 38644 54430 38700
rect 54430 38644 54486 38700
rect 54486 38644 54490 38700
rect 54426 38640 54490 38644
rect 54506 38700 54570 38704
rect 54506 38644 54510 38700
rect 54510 38644 54566 38700
rect 54566 38644 54570 38700
rect 54506 38640 54570 38644
rect 59594 38700 59658 38704
rect 59594 38644 59598 38700
rect 59598 38644 59654 38700
rect 59654 38644 59658 38700
rect 59594 38640 59658 38644
rect 59674 38700 59738 38704
rect 59674 38644 59678 38700
rect 59678 38644 59734 38700
rect 59734 38644 59738 38700
rect 59674 38640 59738 38644
rect 59754 38700 59818 38704
rect 59754 38644 59758 38700
rect 59758 38644 59814 38700
rect 59814 38644 59818 38700
rect 59754 38640 59818 38644
rect 59834 38700 59898 38704
rect 59834 38644 59838 38700
rect 59838 38644 59894 38700
rect 59894 38644 59898 38700
rect 59834 38640 59898 38644
rect 64922 38700 64986 38704
rect 64922 38644 64926 38700
rect 64926 38644 64982 38700
rect 64982 38644 64986 38700
rect 64922 38640 64986 38644
rect 65002 38700 65066 38704
rect 65002 38644 65006 38700
rect 65006 38644 65062 38700
rect 65062 38644 65066 38700
rect 65002 38640 65066 38644
rect 65082 38700 65146 38704
rect 65082 38644 65086 38700
rect 65086 38644 65142 38700
rect 65142 38644 65146 38700
rect 65082 38640 65146 38644
rect 65162 38700 65226 38704
rect 65162 38644 65166 38700
rect 65166 38644 65222 38700
rect 65222 38644 65226 38700
rect 65162 38640 65226 38644
rect 70250 38700 70314 38704
rect 70250 38644 70254 38700
rect 70254 38644 70310 38700
rect 70310 38644 70314 38700
rect 70250 38640 70314 38644
rect 70330 38700 70394 38704
rect 70330 38644 70334 38700
rect 70334 38644 70390 38700
rect 70390 38644 70394 38700
rect 70330 38640 70394 38644
rect 70410 38700 70474 38704
rect 70410 38644 70414 38700
rect 70414 38644 70470 38700
rect 70470 38644 70474 38700
rect 70410 38640 70474 38644
rect 70490 38700 70554 38704
rect 70490 38644 70494 38700
rect 70494 38644 70550 38700
rect 70550 38644 70554 38700
rect 70490 38640 70554 38644
rect 75578 38700 75642 38704
rect 75578 38644 75582 38700
rect 75582 38644 75638 38700
rect 75638 38644 75642 38700
rect 75578 38640 75642 38644
rect 75658 38700 75722 38704
rect 75658 38644 75662 38700
rect 75662 38644 75718 38700
rect 75718 38644 75722 38700
rect 75658 38640 75722 38644
rect 75738 38700 75802 38704
rect 75738 38644 75742 38700
rect 75742 38644 75798 38700
rect 75798 38644 75802 38700
rect 75738 38640 75802 38644
rect 75818 38700 75882 38704
rect 75818 38644 75822 38700
rect 75822 38644 75878 38700
rect 75878 38644 75882 38700
rect 75818 38640 75882 38644
rect 80906 38700 80970 38704
rect 80906 38644 80910 38700
rect 80910 38644 80966 38700
rect 80966 38644 80970 38700
rect 80906 38640 80970 38644
rect 80986 38700 81050 38704
rect 80986 38644 80990 38700
rect 80990 38644 81046 38700
rect 81046 38644 81050 38700
rect 80986 38640 81050 38644
rect 81066 38700 81130 38704
rect 81066 38644 81070 38700
rect 81070 38644 81126 38700
rect 81126 38644 81130 38700
rect 81066 38640 81130 38644
rect 81146 38700 81210 38704
rect 81146 38644 81150 38700
rect 81150 38644 81206 38700
rect 81206 38644 81210 38700
rect 81146 38640 81210 38644
rect 86234 38700 86298 38704
rect 86234 38644 86238 38700
rect 86238 38644 86294 38700
rect 86294 38644 86298 38700
rect 86234 38640 86298 38644
rect 86314 38700 86378 38704
rect 86314 38644 86318 38700
rect 86318 38644 86374 38700
rect 86374 38644 86378 38700
rect 86314 38640 86378 38644
rect 86394 38700 86458 38704
rect 86394 38644 86398 38700
rect 86398 38644 86454 38700
rect 86454 38644 86458 38700
rect 86394 38640 86458 38644
rect 86474 38700 86538 38704
rect 86474 38644 86478 38700
rect 86478 38644 86534 38700
rect 86534 38644 86538 38700
rect 86474 38640 86538 38644
rect 91562 38700 91626 38704
rect 91562 38644 91566 38700
rect 91566 38644 91622 38700
rect 91622 38644 91626 38700
rect 91562 38640 91626 38644
rect 91642 38700 91706 38704
rect 91642 38644 91646 38700
rect 91646 38644 91702 38700
rect 91702 38644 91706 38700
rect 91642 38640 91706 38644
rect 91722 38700 91786 38704
rect 91722 38644 91726 38700
rect 91726 38644 91782 38700
rect 91782 38644 91786 38700
rect 91722 38640 91786 38644
rect 91802 38700 91866 38704
rect 91802 38644 91806 38700
rect 91806 38644 91862 38700
rect 91862 38644 91866 38700
rect 91802 38640 91866 38644
rect 3650 38156 3714 38160
rect 3650 38100 3654 38156
rect 3654 38100 3710 38156
rect 3710 38100 3714 38156
rect 3650 38096 3714 38100
rect 3730 38156 3794 38160
rect 3730 38100 3734 38156
rect 3734 38100 3790 38156
rect 3790 38100 3794 38156
rect 3730 38096 3794 38100
rect 3810 38156 3874 38160
rect 3810 38100 3814 38156
rect 3814 38100 3870 38156
rect 3870 38100 3874 38156
rect 3810 38096 3874 38100
rect 3890 38156 3954 38160
rect 3890 38100 3894 38156
rect 3894 38100 3950 38156
rect 3950 38100 3954 38156
rect 3890 38096 3954 38100
rect 8978 38156 9042 38160
rect 8978 38100 8982 38156
rect 8982 38100 9038 38156
rect 9038 38100 9042 38156
rect 8978 38096 9042 38100
rect 9058 38156 9122 38160
rect 9058 38100 9062 38156
rect 9062 38100 9118 38156
rect 9118 38100 9122 38156
rect 9058 38096 9122 38100
rect 9138 38156 9202 38160
rect 9138 38100 9142 38156
rect 9142 38100 9198 38156
rect 9198 38100 9202 38156
rect 9138 38096 9202 38100
rect 9218 38156 9282 38160
rect 9218 38100 9222 38156
rect 9222 38100 9278 38156
rect 9278 38100 9282 38156
rect 9218 38096 9282 38100
rect 14306 38156 14370 38160
rect 14306 38100 14310 38156
rect 14310 38100 14366 38156
rect 14366 38100 14370 38156
rect 14306 38096 14370 38100
rect 14386 38156 14450 38160
rect 14386 38100 14390 38156
rect 14390 38100 14446 38156
rect 14446 38100 14450 38156
rect 14386 38096 14450 38100
rect 14466 38156 14530 38160
rect 14466 38100 14470 38156
rect 14470 38100 14526 38156
rect 14526 38100 14530 38156
rect 14466 38096 14530 38100
rect 14546 38156 14610 38160
rect 14546 38100 14550 38156
rect 14550 38100 14606 38156
rect 14606 38100 14610 38156
rect 14546 38096 14610 38100
rect 19634 38156 19698 38160
rect 19634 38100 19638 38156
rect 19638 38100 19694 38156
rect 19694 38100 19698 38156
rect 19634 38096 19698 38100
rect 19714 38156 19778 38160
rect 19714 38100 19718 38156
rect 19718 38100 19774 38156
rect 19774 38100 19778 38156
rect 19714 38096 19778 38100
rect 19794 38156 19858 38160
rect 19794 38100 19798 38156
rect 19798 38100 19854 38156
rect 19854 38100 19858 38156
rect 19794 38096 19858 38100
rect 19874 38156 19938 38160
rect 19874 38100 19878 38156
rect 19878 38100 19934 38156
rect 19934 38100 19938 38156
rect 19874 38096 19938 38100
rect 24962 38156 25026 38160
rect 24962 38100 24966 38156
rect 24966 38100 25022 38156
rect 25022 38100 25026 38156
rect 24962 38096 25026 38100
rect 25042 38156 25106 38160
rect 25042 38100 25046 38156
rect 25046 38100 25102 38156
rect 25102 38100 25106 38156
rect 25042 38096 25106 38100
rect 25122 38156 25186 38160
rect 25122 38100 25126 38156
rect 25126 38100 25182 38156
rect 25182 38100 25186 38156
rect 25122 38096 25186 38100
rect 25202 38156 25266 38160
rect 25202 38100 25206 38156
rect 25206 38100 25262 38156
rect 25262 38100 25266 38156
rect 25202 38096 25266 38100
rect 30290 38156 30354 38160
rect 30290 38100 30294 38156
rect 30294 38100 30350 38156
rect 30350 38100 30354 38156
rect 30290 38096 30354 38100
rect 30370 38156 30434 38160
rect 30370 38100 30374 38156
rect 30374 38100 30430 38156
rect 30430 38100 30434 38156
rect 30370 38096 30434 38100
rect 30450 38156 30514 38160
rect 30450 38100 30454 38156
rect 30454 38100 30510 38156
rect 30510 38100 30514 38156
rect 30450 38096 30514 38100
rect 30530 38156 30594 38160
rect 30530 38100 30534 38156
rect 30534 38100 30590 38156
rect 30590 38100 30594 38156
rect 30530 38096 30594 38100
rect 35618 38156 35682 38160
rect 35618 38100 35622 38156
rect 35622 38100 35678 38156
rect 35678 38100 35682 38156
rect 35618 38096 35682 38100
rect 35698 38156 35762 38160
rect 35698 38100 35702 38156
rect 35702 38100 35758 38156
rect 35758 38100 35762 38156
rect 35698 38096 35762 38100
rect 35778 38156 35842 38160
rect 35778 38100 35782 38156
rect 35782 38100 35838 38156
rect 35838 38100 35842 38156
rect 35778 38096 35842 38100
rect 35858 38156 35922 38160
rect 35858 38100 35862 38156
rect 35862 38100 35918 38156
rect 35918 38100 35922 38156
rect 35858 38096 35922 38100
rect 40946 38156 41010 38160
rect 40946 38100 40950 38156
rect 40950 38100 41006 38156
rect 41006 38100 41010 38156
rect 40946 38096 41010 38100
rect 41026 38156 41090 38160
rect 41026 38100 41030 38156
rect 41030 38100 41086 38156
rect 41086 38100 41090 38156
rect 41026 38096 41090 38100
rect 41106 38156 41170 38160
rect 41106 38100 41110 38156
rect 41110 38100 41166 38156
rect 41166 38100 41170 38156
rect 41106 38096 41170 38100
rect 41186 38156 41250 38160
rect 41186 38100 41190 38156
rect 41190 38100 41246 38156
rect 41246 38100 41250 38156
rect 41186 38096 41250 38100
rect 46274 38156 46338 38160
rect 46274 38100 46278 38156
rect 46278 38100 46334 38156
rect 46334 38100 46338 38156
rect 46274 38096 46338 38100
rect 46354 38156 46418 38160
rect 46354 38100 46358 38156
rect 46358 38100 46414 38156
rect 46414 38100 46418 38156
rect 46354 38096 46418 38100
rect 46434 38156 46498 38160
rect 46434 38100 46438 38156
rect 46438 38100 46494 38156
rect 46494 38100 46498 38156
rect 46434 38096 46498 38100
rect 46514 38156 46578 38160
rect 46514 38100 46518 38156
rect 46518 38100 46574 38156
rect 46574 38100 46578 38156
rect 46514 38096 46578 38100
rect 51602 38156 51666 38160
rect 51602 38100 51606 38156
rect 51606 38100 51662 38156
rect 51662 38100 51666 38156
rect 51602 38096 51666 38100
rect 51682 38156 51746 38160
rect 51682 38100 51686 38156
rect 51686 38100 51742 38156
rect 51742 38100 51746 38156
rect 51682 38096 51746 38100
rect 51762 38156 51826 38160
rect 51762 38100 51766 38156
rect 51766 38100 51822 38156
rect 51822 38100 51826 38156
rect 51762 38096 51826 38100
rect 51842 38156 51906 38160
rect 51842 38100 51846 38156
rect 51846 38100 51902 38156
rect 51902 38100 51906 38156
rect 51842 38096 51906 38100
rect 56930 38156 56994 38160
rect 56930 38100 56934 38156
rect 56934 38100 56990 38156
rect 56990 38100 56994 38156
rect 56930 38096 56994 38100
rect 57010 38156 57074 38160
rect 57010 38100 57014 38156
rect 57014 38100 57070 38156
rect 57070 38100 57074 38156
rect 57010 38096 57074 38100
rect 57090 38156 57154 38160
rect 57090 38100 57094 38156
rect 57094 38100 57150 38156
rect 57150 38100 57154 38156
rect 57090 38096 57154 38100
rect 57170 38156 57234 38160
rect 57170 38100 57174 38156
rect 57174 38100 57230 38156
rect 57230 38100 57234 38156
rect 57170 38096 57234 38100
rect 62258 38156 62322 38160
rect 62258 38100 62262 38156
rect 62262 38100 62318 38156
rect 62318 38100 62322 38156
rect 62258 38096 62322 38100
rect 62338 38156 62402 38160
rect 62338 38100 62342 38156
rect 62342 38100 62398 38156
rect 62398 38100 62402 38156
rect 62338 38096 62402 38100
rect 62418 38156 62482 38160
rect 62418 38100 62422 38156
rect 62422 38100 62478 38156
rect 62478 38100 62482 38156
rect 62418 38096 62482 38100
rect 62498 38156 62562 38160
rect 62498 38100 62502 38156
rect 62502 38100 62558 38156
rect 62558 38100 62562 38156
rect 62498 38096 62562 38100
rect 67586 38156 67650 38160
rect 67586 38100 67590 38156
rect 67590 38100 67646 38156
rect 67646 38100 67650 38156
rect 67586 38096 67650 38100
rect 67666 38156 67730 38160
rect 67666 38100 67670 38156
rect 67670 38100 67726 38156
rect 67726 38100 67730 38156
rect 67666 38096 67730 38100
rect 67746 38156 67810 38160
rect 67746 38100 67750 38156
rect 67750 38100 67806 38156
rect 67806 38100 67810 38156
rect 67746 38096 67810 38100
rect 67826 38156 67890 38160
rect 67826 38100 67830 38156
rect 67830 38100 67886 38156
rect 67886 38100 67890 38156
rect 67826 38096 67890 38100
rect 72914 38156 72978 38160
rect 72914 38100 72918 38156
rect 72918 38100 72974 38156
rect 72974 38100 72978 38156
rect 72914 38096 72978 38100
rect 72994 38156 73058 38160
rect 72994 38100 72998 38156
rect 72998 38100 73054 38156
rect 73054 38100 73058 38156
rect 72994 38096 73058 38100
rect 73074 38156 73138 38160
rect 73074 38100 73078 38156
rect 73078 38100 73134 38156
rect 73134 38100 73138 38156
rect 73074 38096 73138 38100
rect 73154 38156 73218 38160
rect 73154 38100 73158 38156
rect 73158 38100 73214 38156
rect 73214 38100 73218 38156
rect 73154 38096 73218 38100
rect 78242 38156 78306 38160
rect 78242 38100 78246 38156
rect 78246 38100 78302 38156
rect 78302 38100 78306 38156
rect 78242 38096 78306 38100
rect 78322 38156 78386 38160
rect 78322 38100 78326 38156
rect 78326 38100 78382 38156
rect 78382 38100 78386 38156
rect 78322 38096 78386 38100
rect 78402 38156 78466 38160
rect 78402 38100 78406 38156
rect 78406 38100 78462 38156
rect 78462 38100 78466 38156
rect 78402 38096 78466 38100
rect 78482 38156 78546 38160
rect 78482 38100 78486 38156
rect 78486 38100 78542 38156
rect 78542 38100 78546 38156
rect 78482 38096 78546 38100
rect 83570 38156 83634 38160
rect 83570 38100 83574 38156
rect 83574 38100 83630 38156
rect 83630 38100 83634 38156
rect 83570 38096 83634 38100
rect 83650 38156 83714 38160
rect 83650 38100 83654 38156
rect 83654 38100 83710 38156
rect 83710 38100 83714 38156
rect 83650 38096 83714 38100
rect 83730 38156 83794 38160
rect 83730 38100 83734 38156
rect 83734 38100 83790 38156
rect 83790 38100 83794 38156
rect 83730 38096 83794 38100
rect 83810 38156 83874 38160
rect 83810 38100 83814 38156
rect 83814 38100 83870 38156
rect 83870 38100 83874 38156
rect 83810 38096 83874 38100
rect 88898 38156 88962 38160
rect 88898 38100 88902 38156
rect 88902 38100 88958 38156
rect 88958 38100 88962 38156
rect 88898 38096 88962 38100
rect 88978 38156 89042 38160
rect 88978 38100 88982 38156
rect 88982 38100 89038 38156
rect 89038 38100 89042 38156
rect 88978 38096 89042 38100
rect 89058 38156 89122 38160
rect 89058 38100 89062 38156
rect 89062 38100 89118 38156
rect 89118 38100 89122 38156
rect 89058 38096 89122 38100
rect 89138 38156 89202 38160
rect 89138 38100 89142 38156
rect 89142 38100 89198 38156
rect 89198 38100 89202 38156
rect 89138 38096 89202 38100
rect 6314 37612 6378 37616
rect 6314 37556 6318 37612
rect 6318 37556 6374 37612
rect 6374 37556 6378 37612
rect 6314 37552 6378 37556
rect 6394 37612 6458 37616
rect 6394 37556 6398 37612
rect 6398 37556 6454 37612
rect 6454 37556 6458 37612
rect 6394 37552 6458 37556
rect 6474 37612 6538 37616
rect 6474 37556 6478 37612
rect 6478 37556 6534 37612
rect 6534 37556 6538 37612
rect 6474 37552 6538 37556
rect 6554 37612 6618 37616
rect 6554 37556 6558 37612
rect 6558 37556 6614 37612
rect 6614 37556 6618 37612
rect 6554 37552 6618 37556
rect 11642 37612 11706 37616
rect 11642 37556 11646 37612
rect 11646 37556 11702 37612
rect 11702 37556 11706 37612
rect 11642 37552 11706 37556
rect 11722 37612 11786 37616
rect 11722 37556 11726 37612
rect 11726 37556 11782 37612
rect 11782 37556 11786 37612
rect 11722 37552 11786 37556
rect 11802 37612 11866 37616
rect 11802 37556 11806 37612
rect 11806 37556 11862 37612
rect 11862 37556 11866 37612
rect 11802 37552 11866 37556
rect 11882 37612 11946 37616
rect 11882 37556 11886 37612
rect 11886 37556 11942 37612
rect 11942 37556 11946 37612
rect 11882 37552 11946 37556
rect 16970 37612 17034 37616
rect 16970 37556 16974 37612
rect 16974 37556 17030 37612
rect 17030 37556 17034 37612
rect 16970 37552 17034 37556
rect 17050 37612 17114 37616
rect 17050 37556 17054 37612
rect 17054 37556 17110 37612
rect 17110 37556 17114 37612
rect 17050 37552 17114 37556
rect 17130 37612 17194 37616
rect 17130 37556 17134 37612
rect 17134 37556 17190 37612
rect 17190 37556 17194 37612
rect 17130 37552 17194 37556
rect 17210 37612 17274 37616
rect 17210 37556 17214 37612
rect 17214 37556 17270 37612
rect 17270 37556 17274 37612
rect 17210 37552 17274 37556
rect 22298 37612 22362 37616
rect 22298 37556 22302 37612
rect 22302 37556 22358 37612
rect 22358 37556 22362 37612
rect 22298 37552 22362 37556
rect 22378 37612 22442 37616
rect 22378 37556 22382 37612
rect 22382 37556 22438 37612
rect 22438 37556 22442 37612
rect 22378 37552 22442 37556
rect 22458 37612 22522 37616
rect 22458 37556 22462 37612
rect 22462 37556 22518 37612
rect 22518 37556 22522 37612
rect 22458 37552 22522 37556
rect 22538 37612 22602 37616
rect 22538 37556 22542 37612
rect 22542 37556 22598 37612
rect 22598 37556 22602 37612
rect 22538 37552 22602 37556
rect 27626 37612 27690 37616
rect 27626 37556 27630 37612
rect 27630 37556 27686 37612
rect 27686 37556 27690 37612
rect 27626 37552 27690 37556
rect 27706 37612 27770 37616
rect 27706 37556 27710 37612
rect 27710 37556 27766 37612
rect 27766 37556 27770 37612
rect 27706 37552 27770 37556
rect 27786 37612 27850 37616
rect 27786 37556 27790 37612
rect 27790 37556 27846 37612
rect 27846 37556 27850 37612
rect 27786 37552 27850 37556
rect 27866 37612 27930 37616
rect 27866 37556 27870 37612
rect 27870 37556 27926 37612
rect 27926 37556 27930 37612
rect 27866 37552 27930 37556
rect 32954 37612 33018 37616
rect 32954 37556 32958 37612
rect 32958 37556 33014 37612
rect 33014 37556 33018 37612
rect 32954 37552 33018 37556
rect 33034 37612 33098 37616
rect 33034 37556 33038 37612
rect 33038 37556 33094 37612
rect 33094 37556 33098 37612
rect 33034 37552 33098 37556
rect 33114 37612 33178 37616
rect 33114 37556 33118 37612
rect 33118 37556 33174 37612
rect 33174 37556 33178 37612
rect 33114 37552 33178 37556
rect 33194 37612 33258 37616
rect 33194 37556 33198 37612
rect 33198 37556 33254 37612
rect 33254 37556 33258 37612
rect 33194 37552 33258 37556
rect 38282 37612 38346 37616
rect 38282 37556 38286 37612
rect 38286 37556 38342 37612
rect 38342 37556 38346 37612
rect 38282 37552 38346 37556
rect 38362 37612 38426 37616
rect 38362 37556 38366 37612
rect 38366 37556 38422 37612
rect 38422 37556 38426 37612
rect 38362 37552 38426 37556
rect 38442 37612 38506 37616
rect 38442 37556 38446 37612
rect 38446 37556 38502 37612
rect 38502 37556 38506 37612
rect 38442 37552 38506 37556
rect 38522 37612 38586 37616
rect 38522 37556 38526 37612
rect 38526 37556 38582 37612
rect 38582 37556 38586 37612
rect 38522 37552 38586 37556
rect 43610 37612 43674 37616
rect 43610 37556 43614 37612
rect 43614 37556 43670 37612
rect 43670 37556 43674 37612
rect 43610 37552 43674 37556
rect 43690 37612 43754 37616
rect 43690 37556 43694 37612
rect 43694 37556 43750 37612
rect 43750 37556 43754 37612
rect 43690 37552 43754 37556
rect 43770 37612 43834 37616
rect 43770 37556 43774 37612
rect 43774 37556 43830 37612
rect 43830 37556 43834 37612
rect 43770 37552 43834 37556
rect 43850 37612 43914 37616
rect 43850 37556 43854 37612
rect 43854 37556 43910 37612
rect 43910 37556 43914 37612
rect 43850 37552 43914 37556
rect 48938 37612 49002 37616
rect 48938 37556 48942 37612
rect 48942 37556 48998 37612
rect 48998 37556 49002 37612
rect 48938 37552 49002 37556
rect 49018 37612 49082 37616
rect 49018 37556 49022 37612
rect 49022 37556 49078 37612
rect 49078 37556 49082 37612
rect 49018 37552 49082 37556
rect 49098 37612 49162 37616
rect 49098 37556 49102 37612
rect 49102 37556 49158 37612
rect 49158 37556 49162 37612
rect 49098 37552 49162 37556
rect 49178 37612 49242 37616
rect 49178 37556 49182 37612
rect 49182 37556 49238 37612
rect 49238 37556 49242 37612
rect 49178 37552 49242 37556
rect 54266 37612 54330 37616
rect 54266 37556 54270 37612
rect 54270 37556 54326 37612
rect 54326 37556 54330 37612
rect 54266 37552 54330 37556
rect 54346 37612 54410 37616
rect 54346 37556 54350 37612
rect 54350 37556 54406 37612
rect 54406 37556 54410 37612
rect 54346 37552 54410 37556
rect 54426 37612 54490 37616
rect 54426 37556 54430 37612
rect 54430 37556 54486 37612
rect 54486 37556 54490 37612
rect 54426 37552 54490 37556
rect 54506 37612 54570 37616
rect 54506 37556 54510 37612
rect 54510 37556 54566 37612
rect 54566 37556 54570 37612
rect 54506 37552 54570 37556
rect 59594 37612 59658 37616
rect 59594 37556 59598 37612
rect 59598 37556 59654 37612
rect 59654 37556 59658 37612
rect 59594 37552 59658 37556
rect 59674 37612 59738 37616
rect 59674 37556 59678 37612
rect 59678 37556 59734 37612
rect 59734 37556 59738 37612
rect 59674 37552 59738 37556
rect 59754 37612 59818 37616
rect 59754 37556 59758 37612
rect 59758 37556 59814 37612
rect 59814 37556 59818 37612
rect 59754 37552 59818 37556
rect 59834 37612 59898 37616
rect 59834 37556 59838 37612
rect 59838 37556 59894 37612
rect 59894 37556 59898 37612
rect 59834 37552 59898 37556
rect 64922 37612 64986 37616
rect 64922 37556 64926 37612
rect 64926 37556 64982 37612
rect 64982 37556 64986 37612
rect 64922 37552 64986 37556
rect 65002 37612 65066 37616
rect 65002 37556 65006 37612
rect 65006 37556 65062 37612
rect 65062 37556 65066 37612
rect 65002 37552 65066 37556
rect 65082 37612 65146 37616
rect 65082 37556 65086 37612
rect 65086 37556 65142 37612
rect 65142 37556 65146 37612
rect 65082 37552 65146 37556
rect 65162 37612 65226 37616
rect 65162 37556 65166 37612
rect 65166 37556 65222 37612
rect 65222 37556 65226 37612
rect 65162 37552 65226 37556
rect 70250 37612 70314 37616
rect 70250 37556 70254 37612
rect 70254 37556 70310 37612
rect 70310 37556 70314 37612
rect 70250 37552 70314 37556
rect 70330 37612 70394 37616
rect 70330 37556 70334 37612
rect 70334 37556 70390 37612
rect 70390 37556 70394 37612
rect 70330 37552 70394 37556
rect 70410 37612 70474 37616
rect 70410 37556 70414 37612
rect 70414 37556 70470 37612
rect 70470 37556 70474 37612
rect 70410 37552 70474 37556
rect 70490 37612 70554 37616
rect 70490 37556 70494 37612
rect 70494 37556 70550 37612
rect 70550 37556 70554 37612
rect 70490 37552 70554 37556
rect 75578 37612 75642 37616
rect 75578 37556 75582 37612
rect 75582 37556 75638 37612
rect 75638 37556 75642 37612
rect 75578 37552 75642 37556
rect 75658 37612 75722 37616
rect 75658 37556 75662 37612
rect 75662 37556 75718 37612
rect 75718 37556 75722 37612
rect 75658 37552 75722 37556
rect 75738 37612 75802 37616
rect 75738 37556 75742 37612
rect 75742 37556 75798 37612
rect 75798 37556 75802 37612
rect 75738 37552 75802 37556
rect 75818 37612 75882 37616
rect 75818 37556 75822 37612
rect 75822 37556 75878 37612
rect 75878 37556 75882 37612
rect 75818 37552 75882 37556
rect 80906 37612 80970 37616
rect 80906 37556 80910 37612
rect 80910 37556 80966 37612
rect 80966 37556 80970 37612
rect 80906 37552 80970 37556
rect 80986 37612 81050 37616
rect 80986 37556 80990 37612
rect 80990 37556 81046 37612
rect 81046 37556 81050 37612
rect 80986 37552 81050 37556
rect 81066 37612 81130 37616
rect 81066 37556 81070 37612
rect 81070 37556 81126 37612
rect 81126 37556 81130 37612
rect 81066 37552 81130 37556
rect 81146 37612 81210 37616
rect 81146 37556 81150 37612
rect 81150 37556 81206 37612
rect 81206 37556 81210 37612
rect 81146 37552 81210 37556
rect 86234 37612 86298 37616
rect 86234 37556 86238 37612
rect 86238 37556 86294 37612
rect 86294 37556 86298 37612
rect 86234 37552 86298 37556
rect 86314 37612 86378 37616
rect 86314 37556 86318 37612
rect 86318 37556 86374 37612
rect 86374 37556 86378 37612
rect 86314 37552 86378 37556
rect 86394 37612 86458 37616
rect 86394 37556 86398 37612
rect 86398 37556 86454 37612
rect 86454 37556 86458 37612
rect 86394 37552 86458 37556
rect 86474 37612 86538 37616
rect 86474 37556 86478 37612
rect 86478 37556 86534 37612
rect 86534 37556 86538 37612
rect 86474 37552 86538 37556
rect 91562 37612 91626 37616
rect 91562 37556 91566 37612
rect 91566 37556 91622 37612
rect 91622 37556 91626 37612
rect 91562 37552 91626 37556
rect 91642 37612 91706 37616
rect 91642 37556 91646 37612
rect 91646 37556 91702 37612
rect 91702 37556 91706 37612
rect 91642 37552 91706 37556
rect 91722 37612 91786 37616
rect 91722 37556 91726 37612
rect 91726 37556 91782 37612
rect 91782 37556 91786 37612
rect 91722 37552 91786 37556
rect 91802 37612 91866 37616
rect 91802 37556 91806 37612
rect 91806 37556 91862 37612
rect 91862 37556 91866 37612
rect 91802 37552 91866 37556
rect 3650 37068 3714 37072
rect 3650 37012 3654 37068
rect 3654 37012 3710 37068
rect 3710 37012 3714 37068
rect 3650 37008 3714 37012
rect 3730 37068 3794 37072
rect 3730 37012 3734 37068
rect 3734 37012 3790 37068
rect 3790 37012 3794 37068
rect 3730 37008 3794 37012
rect 3810 37068 3874 37072
rect 3810 37012 3814 37068
rect 3814 37012 3870 37068
rect 3870 37012 3874 37068
rect 3810 37008 3874 37012
rect 3890 37068 3954 37072
rect 3890 37012 3894 37068
rect 3894 37012 3950 37068
rect 3950 37012 3954 37068
rect 3890 37008 3954 37012
rect 8978 37068 9042 37072
rect 8978 37012 8982 37068
rect 8982 37012 9038 37068
rect 9038 37012 9042 37068
rect 8978 37008 9042 37012
rect 9058 37068 9122 37072
rect 9058 37012 9062 37068
rect 9062 37012 9118 37068
rect 9118 37012 9122 37068
rect 9058 37008 9122 37012
rect 9138 37068 9202 37072
rect 9138 37012 9142 37068
rect 9142 37012 9198 37068
rect 9198 37012 9202 37068
rect 9138 37008 9202 37012
rect 9218 37068 9282 37072
rect 9218 37012 9222 37068
rect 9222 37012 9278 37068
rect 9278 37012 9282 37068
rect 9218 37008 9282 37012
rect 14306 37068 14370 37072
rect 14306 37012 14310 37068
rect 14310 37012 14366 37068
rect 14366 37012 14370 37068
rect 14306 37008 14370 37012
rect 14386 37068 14450 37072
rect 14386 37012 14390 37068
rect 14390 37012 14446 37068
rect 14446 37012 14450 37068
rect 14386 37008 14450 37012
rect 14466 37068 14530 37072
rect 14466 37012 14470 37068
rect 14470 37012 14526 37068
rect 14526 37012 14530 37068
rect 14466 37008 14530 37012
rect 14546 37068 14610 37072
rect 14546 37012 14550 37068
rect 14550 37012 14606 37068
rect 14606 37012 14610 37068
rect 14546 37008 14610 37012
rect 19634 37068 19698 37072
rect 19634 37012 19638 37068
rect 19638 37012 19694 37068
rect 19694 37012 19698 37068
rect 19634 37008 19698 37012
rect 19714 37068 19778 37072
rect 19714 37012 19718 37068
rect 19718 37012 19774 37068
rect 19774 37012 19778 37068
rect 19714 37008 19778 37012
rect 19794 37068 19858 37072
rect 19794 37012 19798 37068
rect 19798 37012 19854 37068
rect 19854 37012 19858 37068
rect 19794 37008 19858 37012
rect 19874 37068 19938 37072
rect 19874 37012 19878 37068
rect 19878 37012 19934 37068
rect 19934 37012 19938 37068
rect 19874 37008 19938 37012
rect 24962 37068 25026 37072
rect 24962 37012 24966 37068
rect 24966 37012 25022 37068
rect 25022 37012 25026 37068
rect 24962 37008 25026 37012
rect 25042 37068 25106 37072
rect 25042 37012 25046 37068
rect 25046 37012 25102 37068
rect 25102 37012 25106 37068
rect 25042 37008 25106 37012
rect 25122 37068 25186 37072
rect 25122 37012 25126 37068
rect 25126 37012 25182 37068
rect 25182 37012 25186 37068
rect 25122 37008 25186 37012
rect 25202 37068 25266 37072
rect 25202 37012 25206 37068
rect 25206 37012 25262 37068
rect 25262 37012 25266 37068
rect 25202 37008 25266 37012
rect 30290 37068 30354 37072
rect 30290 37012 30294 37068
rect 30294 37012 30350 37068
rect 30350 37012 30354 37068
rect 30290 37008 30354 37012
rect 30370 37068 30434 37072
rect 30370 37012 30374 37068
rect 30374 37012 30430 37068
rect 30430 37012 30434 37068
rect 30370 37008 30434 37012
rect 30450 37068 30514 37072
rect 30450 37012 30454 37068
rect 30454 37012 30510 37068
rect 30510 37012 30514 37068
rect 30450 37008 30514 37012
rect 30530 37068 30594 37072
rect 30530 37012 30534 37068
rect 30534 37012 30590 37068
rect 30590 37012 30594 37068
rect 30530 37008 30594 37012
rect 35618 37068 35682 37072
rect 35618 37012 35622 37068
rect 35622 37012 35678 37068
rect 35678 37012 35682 37068
rect 35618 37008 35682 37012
rect 35698 37068 35762 37072
rect 35698 37012 35702 37068
rect 35702 37012 35758 37068
rect 35758 37012 35762 37068
rect 35698 37008 35762 37012
rect 35778 37068 35842 37072
rect 35778 37012 35782 37068
rect 35782 37012 35838 37068
rect 35838 37012 35842 37068
rect 35778 37008 35842 37012
rect 35858 37068 35922 37072
rect 35858 37012 35862 37068
rect 35862 37012 35918 37068
rect 35918 37012 35922 37068
rect 35858 37008 35922 37012
rect 40946 37068 41010 37072
rect 40946 37012 40950 37068
rect 40950 37012 41006 37068
rect 41006 37012 41010 37068
rect 40946 37008 41010 37012
rect 41026 37068 41090 37072
rect 41026 37012 41030 37068
rect 41030 37012 41086 37068
rect 41086 37012 41090 37068
rect 41026 37008 41090 37012
rect 41106 37068 41170 37072
rect 41106 37012 41110 37068
rect 41110 37012 41166 37068
rect 41166 37012 41170 37068
rect 41106 37008 41170 37012
rect 41186 37068 41250 37072
rect 41186 37012 41190 37068
rect 41190 37012 41246 37068
rect 41246 37012 41250 37068
rect 41186 37008 41250 37012
rect 46274 37068 46338 37072
rect 46274 37012 46278 37068
rect 46278 37012 46334 37068
rect 46334 37012 46338 37068
rect 46274 37008 46338 37012
rect 46354 37068 46418 37072
rect 46354 37012 46358 37068
rect 46358 37012 46414 37068
rect 46414 37012 46418 37068
rect 46354 37008 46418 37012
rect 46434 37068 46498 37072
rect 46434 37012 46438 37068
rect 46438 37012 46494 37068
rect 46494 37012 46498 37068
rect 46434 37008 46498 37012
rect 46514 37068 46578 37072
rect 46514 37012 46518 37068
rect 46518 37012 46574 37068
rect 46574 37012 46578 37068
rect 46514 37008 46578 37012
rect 51602 37068 51666 37072
rect 51602 37012 51606 37068
rect 51606 37012 51662 37068
rect 51662 37012 51666 37068
rect 51602 37008 51666 37012
rect 51682 37068 51746 37072
rect 51682 37012 51686 37068
rect 51686 37012 51742 37068
rect 51742 37012 51746 37068
rect 51682 37008 51746 37012
rect 51762 37068 51826 37072
rect 51762 37012 51766 37068
rect 51766 37012 51822 37068
rect 51822 37012 51826 37068
rect 51762 37008 51826 37012
rect 51842 37068 51906 37072
rect 51842 37012 51846 37068
rect 51846 37012 51902 37068
rect 51902 37012 51906 37068
rect 51842 37008 51906 37012
rect 56930 37068 56994 37072
rect 56930 37012 56934 37068
rect 56934 37012 56990 37068
rect 56990 37012 56994 37068
rect 56930 37008 56994 37012
rect 57010 37068 57074 37072
rect 57010 37012 57014 37068
rect 57014 37012 57070 37068
rect 57070 37012 57074 37068
rect 57010 37008 57074 37012
rect 57090 37068 57154 37072
rect 57090 37012 57094 37068
rect 57094 37012 57150 37068
rect 57150 37012 57154 37068
rect 57090 37008 57154 37012
rect 57170 37068 57234 37072
rect 57170 37012 57174 37068
rect 57174 37012 57230 37068
rect 57230 37012 57234 37068
rect 57170 37008 57234 37012
rect 62258 37068 62322 37072
rect 62258 37012 62262 37068
rect 62262 37012 62318 37068
rect 62318 37012 62322 37068
rect 62258 37008 62322 37012
rect 62338 37068 62402 37072
rect 62338 37012 62342 37068
rect 62342 37012 62398 37068
rect 62398 37012 62402 37068
rect 62338 37008 62402 37012
rect 62418 37068 62482 37072
rect 62418 37012 62422 37068
rect 62422 37012 62478 37068
rect 62478 37012 62482 37068
rect 62418 37008 62482 37012
rect 62498 37068 62562 37072
rect 62498 37012 62502 37068
rect 62502 37012 62558 37068
rect 62558 37012 62562 37068
rect 62498 37008 62562 37012
rect 67586 37068 67650 37072
rect 67586 37012 67590 37068
rect 67590 37012 67646 37068
rect 67646 37012 67650 37068
rect 67586 37008 67650 37012
rect 67666 37068 67730 37072
rect 67666 37012 67670 37068
rect 67670 37012 67726 37068
rect 67726 37012 67730 37068
rect 67666 37008 67730 37012
rect 67746 37068 67810 37072
rect 67746 37012 67750 37068
rect 67750 37012 67806 37068
rect 67806 37012 67810 37068
rect 67746 37008 67810 37012
rect 67826 37068 67890 37072
rect 67826 37012 67830 37068
rect 67830 37012 67886 37068
rect 67886 37012 67890 37068
rect 67826 37008 67890 37012
rect 72914 37068 72978 37072
rect 72914 37012 72918 37068
rect 72918 37012 72974 37068
rect 72974 37012 72978 37068
rect 72914 37008 72978 37012
rect 72994 37068 73058 37072
rect 72994 37012 72998 37068
rect 72998 37012 73054 37068
rect 73054 37012 73058 37068
rect 72994 37008 73058 37012
rect 73074 37068 73138 37072
rect 73074 37012 73078 37068
rect 73078 37012 73134 37068
rect 73134 37012 73138 37068
rect 73074 37008 73138 37012
rect 73154 37068 73218 37072
rect 73154 37012 73158 37068
rect 73158 37012 73214 37068
rect 73214 37012 73218 37068
rect 73154 37008 73218 37012
rect 78242 37068 78306 37072
rect 78242 37012 78246 37068
rect 78246 37012 78302 37068
rect 78302 37012 78306 37068
rect 78242 37008 78306 37012
rect 78322 37068 78386 37072
rect 78322 37012 78326 37068
rect 78326 37012 78382 37068
rect 78382 37012 78386 37068
rect 78322 37008 78386 37012
rect 78402 37068 78466 37072
rect 78402 37012 78406 37068
rect 78406 37012 78462 37068
rect 78462 37012 78466 37068
rect 78402 37008 78466 37012
rect 78482 37068 78546 37072
rect 78482 37012 78486 37068
rect 78486 37012 78542 37068
rect 78542 37012 78546 37068
rect 78482 37008 78546 37012
rect 83570 37068 83634 37072
rect 83570 37012 83574 37068
rect 83574 37012 83630 37068
rect 83630 37012 83634 37068
rect 83570 37008 83634 37012
rect 83650 37068 83714 37072
rect 83650 37012 83654 37068
rect 83654 37012 83710 37068
rect 83710 37012 83714 37068
rect 83650 37008 83714 37012
rect 83730 37068 83794 37072
rect 83730 37012 83734 37068
rect 83734 37012 83790 37068
rect 83790 37012 83794 37068
rect 83730 37008 83794 37012
rect 83810 37068 83874 37072
rect 83810 37012 83814 37068
rect 83814 37012 83870 37068
rect 83870 37012 83874 37068
rect 83810 37008 83874 37012
rect 88898 37068 88962 37072
rect 88898 37012 88902 37068
rect 88902 37012 88958 37068
rect 88958 37012 88962 37068
rect 88898 37008 88962 37012
rect 88978 37068 89042 37072
rect 88978 37012 88982 37068
rect 88982 37012 89038 37068
rect 89038 37012 89042 37068
rect 88978 37008 89042 37012
rect 89058 37068 89122 37072
rect 89058 37012 89062 37068
rect 89062 37012 89118 37068
rect 89118 37012 89122 37068
rect 89058 37008 89122 37012
rect 89138 37068 89202 37072
rect 89138 37012 89142 37068
rect 89142 37012 89198 37068
rect 89198 37012 89202 37068
rect 89138 37008 89202 37012
rect 6314 36524 6378 36528
rect 6314 36468 6318 36524
rect 6318 36468 6374 36524
rect 6374 36468 6378 36524
rect 6314 36464 6378 36468
rect 6394 36524 6458 36528
rect 6394 36468 6398 36524
rect 6398 36468 6454 36524
rect 6454 36468 6458 36524
rect 6394 36464 6458 36468
rect 6474 36524 6538 36528
rect 6474 36468 6478 36524
rect 6478 36468 6534 36524
rect 6534 36468 6538 36524
rect 6474 36464 6538 36468
rect 6554 36524 6618 36528
rect 6554 36468 6558 36524
rect 6558 36468 6614 36524
rect 6614 36468 6618 36524
rect 6554 36464 6618 36468
rect 11642 36524 11706 36528
rect 11642 36468 11646 36524
rect 11646 36468 11702 36524
rect 11702 36468 11706 36524
rect 11642 36464 11706 36468
rect 11722 36524 11786 36528
rect 11722 36468 11726 36524
rect 11726 36468 11782 36524
rect 11782 36468 11786 36524
rect 11722 36464 11786 36468
rect 11802 36524 11866 36528
rect 11802 36468 11806 36524
rect 11806 36468 11862 36524
rect 11862 36468 11866 36524
rect 11802 36464 11866 36468
rect 11882 36524 11946 36528
rect 11882 36468 11886 36524
rect 11886 36468 11942 36524
rect 11942 36468 11946 36524
rect 11882 36464 11946 36468
rect 16970 36524 17034 36528
rect 16970 36468 16974 36524
rect 16974 36468 17030 36524
rect 17030 36468 17034 36524
rect 16970 36464 17034 36468
rect 17050 36524 17114 36528
rect 17050 36468 17054 36524
rect 17054 36468 17110 36524
rect 17110 36468 17114 36524
rect 17050 36464 17114 36468
rect 17130 36524 17194 36528
rect 17130 36468 17134 36524
rect 17134 36468 17190 36524
rect 17190 36468 17194 36524
rect 17130 36464 17194 36468
rect 17210 36524 17274 36528
rect 17210 36468 17214 36524
rect 17214 36468 17270 36524
rect 17270 36468 17274 36524
rect 17210 36464 17274 36468
rect 22298 36524 22362 36528
rect 22298 36468 22302 36524
rect 22302 36468 22358 36524
rect 22358 36468 22362 36524
rect 22298 36464 22362 36468
rect 22378 36524 22442 36528
rect 22378 36468 22382 36524
rect 22382 36468 22438 36524
rect 22438 36468 22442 36524
rect 22378 36464 22442 36468
rect 22458 36524 22522 36528
rect 22458 36468 22462 36524
rect 22462 36468 22518 36524
rect 22518 36468 22522 36524
rect 22458 36464 22522 36468
rect 22538 36524 22602 36528
rect 22538 36468 22542 36524
rect 22542 36468 22598 36524
rect 22598 36468 22602 36524
rect 22538 36464 22602 36468
rect 27626 36524 27690 36528
rect 27626 36468 27630 36524
rect 27630 36468 27686 36524
rect 27686 36468 27690 36524
rect 27626 36464 27690 36468
rect 27706 36524 27770 36528
rect 27706 36468 27710 36524
rect 27710 36468 27766 36524
rect 27766 36468 27770 36524
rect 27706 36464 27770 36468
rect 27786 36524 27850 36528
rect 27786 36468 27790 36524
rect 27790 36468 27846 36524
rect 27846 36468 27850 36524
rect 27786 36464 27850 36468
rect 27866 36524 27930 36528
rect 27866 36468 27870 36524
rect 27870 36468 27926 36524
rect 27926 36468 27930 36524
rect 27866 36464 27930 36468
rect 32954 36524 33018 36528
rect 32954 36468 32958 36524
rect 32958 36468 33014 36524
rect 33014 36468 33018 36524
rect 32954 36464 33018 36468
rect 33034 36524 33098 36528
rect 33034 36468 33038 36524
rect 33038 36468 33094 36524
rect 33094 36468 33098 36524
rect 33034 36464 33098 36468
rect 33114 36524 33178 36528
rect 33114 36468 33118 36524
rect 33118 36468 33174 36524
rect 33174 36468 33178 36524
rect 33114 36464 33178 36468
rect 33194 36524 33258 36528
rect 33194 36468 33198 36524
rect 33198 36468 33254 36524
rect 33254 36468 33258 36524
rect 33194 36464 33258 36468
rect 38282 36524 38346 36528
rect 38282 36468 38286 36524
rect 38286 36468 38342 36524
rect 38342 36468 38346 36524
rect 38282 36464 38346 36468
rect 38362 36524 38426 36528
rect 38362 36468 38366 36524
rect 38366 36468 38422 36524
rect 38422 36468 38426 36524
rect 38362 36464 38426 36468
rect 38442 36524 38506 36528
rect 38442 36468 38446 36524
rect 38446 36468 38502 36524
rect 38502 36468 38506 36524
rect 38442 36464 38506 36468
rect 38522 36524 38586 36528
rect 38522 36468 38526 36524
rect 38526 36468 38582 36524
rect 38582 36468 38586 36524
rect 38522 36464 38586 36468
rect 43610 36524 43674 36528
rect 43610 36468 43614 36524
rect 43614 36468 43670 36524
rect 43670 36468 43674 36524
rect 43610 36464 43674 36468
rect 43690 36524 43754 36528
rect 43690 36468 43694 36524
rect 43694 36468 43750 36524
rect 43750 36468 43754 36524
rect 43690 36464 43754 36468
rect 43770 36524 43834 36528
rect 43770 36468 43774 36524
rect 43774 36468 43830 36524
rect 43830 36468 43834 36524
rect 43770 36464 43834 36468
rect 43850 36524 43914 36528
rect 43850 36468 43854 36524
rect 43854 36468 43910 36524
rect 43910 36468 43914 36524
rect 43850 36464 43914 36468
rect 48938 36524 49002 36528
rect 48938 36468 48942 36524
rect 48942 36468 48998 36524
rect 48998 36468 49002 36524
rect 48938 36464 49002 36468
rect 49018 36524 49082 36528
rect 49018 36468 49022 36524
rect 49022 36468 49078 36524
rect 49078 36468 49082 36524
rect 49018 36464 49082 36468
rect 49098 36524 49162 36528
rect 49098 36468 49102 36524
rect 49102 36468 49158 36524
rect 49158 36468 49162 36524
rect 49098 36464 49162 36468
rect 49178 36524 49242 36528
rect 49178 36468 49182 36524
rect 49182 36468 49238 36524
rect 49238 36468 49242 36524
rect 49178 36464 49242 36468
rect 54266 36524 54330 36528
rect 54266 36468 54270 36524
rect 54270 36468 54326 36524
rect 54326 36468 54330 36524
rect 54266 36464 54330 36468
rect 54346 36524 54410 36528
rect 54346 36468 54350 36524
rect 54350 36468 54406 36524
rect 54406 36468 54410 36524
rect 54346 36464 54410 36468
rect 54426 36524 54490 36528
rect 54426 36468 54430 36524
rect 54430 36468 54486 36524
rect 54486 36468 54490 36524
rect 54426 36464 54490 36468
rect 54506 36524 54570 36528
rect 54506 36468 54510 36524
rect 54510 36468 54566 36524
rect 54566 36468 54570 36524
rect 54506 36464 54570 36468
rect 59594 36524 59658 36528
rect 59594 36468 59598 36524
rect 59598 36468 59654 36524
rect 59654 36468 59658 36524
rect 59594 36464 59658 36468
rect 59674 36524 59738 36528
rect 59674 36468 59678 36524
rect 59678 36468 59734 36524
rect 59734 36468 59738 36524
rect 59674 36464 59738 36468
rect 59754 36524 59818 36528
rect 59754 36468 59758 36524
rect 59758 36468 59814 36524
rect 59814 36468 59818 36524
rect 59754 36464 59818 36468
rect 59834 36524 59898 36528
rect 59834 36468 59838 36524
rect 59838 36468 59894 36524
rect 59894 36468 59898 36524
rect 59834 36464 59898 36468
rect 64922 36524 64986 36528
rect 64922 36468 64926 36524
rect 64926 36468 64982 36524
rect 64982 36468 64986 36524
rect 64922 36464 64986 36468
rect 65002 36524 65066 36528
rect 65002 36468 65006 36524
rect 65006 36468 65062 36524
rect 65062 36468 65066 36524
rect 65002 36464 65066 36468
rect 65082 36524 65146 36528
rect 65082 36468 65086 36524
rect 65086 36468 65142 36524
rect 65142 36468 65146 36524
rect 65082 36464 65146 36468
rect 65162 36524 65226 36528
rect 65162 36468 65166 36524
rect 65166 36468 65222 36524
rect 65222 36468 65226 36524
rect 65162 36464 65226 36468
rect 70250 36524 70314 36528
rect 70250 36468 70254 36524
rect 70254 36468 70310 36524
rect 70310 36468 70314 36524
rect 70250 36464 70314 36468
rect 70330 36524 70394 36528
rect 70330 36468 70334 36524
rect 70334 36468 70390 36524
rect 70390 36468 70394 36524
rect 70330 36464 70394 36468
rect 70410 36524 70474 36528
rect 70410 36468 70414 36524
rect 70414 36468 70470 36524
rect 70470 36468 70474 36524
rect 70410 36464 70474 36468
rect 70490 36524 70554 36528
rect 70490 36468 70494 36524
rect 70494 36468 70550 36524
rect 70550 36468 70554 36524
rect 70490 36464 70554 36468
rect 75578 36524 75642 36528
rect 75578 36468 75582 36524
rect 75582 36468 75638 36524
rect 75638 36468 75642 36524
rect 75578 36464 75642 36468
rect 75658 36524 75722 36528
rect 75658 36468 75662 36524
rect 75662 36468 75718 36524
rect 75718 36468 75722 36524
rect 75658 36464 75722 36468
rect 75738 36524 75802 36528
rect 75738 36468 75742 36524
rect 75742 36468 75798 36524
rect 75798 36468 75802 36524
rect 75738 36464 75802 36468
rect 75818 36524 75882 36528
rect 75818 36468 75822 36524
rect 75822 36468 75878 36524
rect 75878 36468 75882 36524
rect 75818 36464 75882 36468
rect 80906 36524 80970 36528
rect 80906 36468 80910 36524
rect 80910 36468 80966 36524
rect 80966 36468 80970 36524
rect 80906 36464 80970 36468
rect 80986 36524 81050 36528
rect 80986 36468 80990 36524
rect 80990 36468 81046 36524
rect 81046 36468 81050 36524
rect 80986 36464 81050 36468
rect 81066 36524 81130 36528
rect 81066 36468 81070 36524
rect 81070 36468 81126 36524
rect 81126 36468 81130 36524
rect 81066 36464 81130 36468
rect 81146 36524 81210 36528
rect 81146 36468 81150 36524
rect 81150 36468 81206 36524
rect 81206 36468 81210 36524
rect 81146 36464 81210 36468
rect 86234 36524 86298 36528
rect 86234 36468 86238 36524
rect 86238 36468 86294 36524
rect 86294 36468 86298 36524
rect 86234 36464 86298 36468
rect 86314 36524 86378 36528
rect 86314 36468 86318 36524
rect 86318 36468 86374 36524
rect 86374 36468 86378 36524
rect 86314 36464 86378 36468
rect 86394 36524 86458 36528
rect 86394 36468 86398 36524
rect 86398 36468 86454 36524
rect 86454 36468 86458 36524
rect 86394 36464 86458 36468
rect 86474 36524 86538 36528
rect 86474 36468 86478 36524
rect 86478 36468 86534 36524
rect 86534 36468 86538 36524
rect 86474 36464 86538 36468
rect 91562 36524 91626 36528
rect 91562 36468 91566 36524
rect 91566 36468 91622 36524
rect 91622 36468 91626 36524
rect 91562 36464 91626 36468
rect 91642 36524 91706 36528
rect 91642 36468 91646 36524
rect 91646 36468 91702 36524
rect 91702 36468 91706 36524
rect 91642 36464 91706 36468
rect 91722 36524 91786 36528
rect 91722 36468 91726 36524
rect 91726 36468 91782 36524
rect 91782 36468 91786 36524
rect 91722 36464 91786 36468
rect 91802 36524 91866 36528
rect 91802 36468 91806 36524
rect 91806 36468 91862 36524
rect 91862 36468 91866 36524
rect 91802 36464 91866 36468
rect 3650 35980 3714 35984
rect 3650 35924 3654 35980
rect 3654 35924 3710 35980
rect 3710 35924 3714 35980
rect 3650 35920 3714 35924
rect 3730 35980 3794 35984
rect 3730 35924 3734 35980
rect 3734 35924 3790 35980
rect 3790 35924 3794 35980
rect 3730 35920 3794 35924
rect 3810 35980 3874 35984
rect 3810 35924 3814 35980
rect 3814 35924 3870 35980
rect 3870 35924 3874 35980
rect 3810 35920 3874 35924
rect 3890 35980 3954 35984
rect 3890 35924 3894 35980
rect 3894 35924 3950 35980
rect 3950 35924 3954 35980
rect 3890 35920 3954 35924
rect 8978 35980 9042 35984
rect 8978 35924 8982 35980
rect 8982 35924 9038 35980
rect 9038 35924 9042 35980
rect 8978 35920 9042 35924
rect 9058 35980 9122 35984
rect 9058 35924 9062 35980
rect 9062 35924 9118 35980
rect 9118 35924 9122 35980
rect 9058 35920 9122 35924
rect 9138 35980 9202 35984
rect 9138 35924 9142 35980
rect 9142 35924 9198 35980
rect 9198 35924 9202 35980
rect 9138 35920 9202 35924
rect 9218 35980 9282 35984
rect 9218 35924 9222 35980
rect 9222 35924 9278 35980
rect 9278 35924 9282 35980
rect 9218 35920 9282 35924
rect 14306 35980 14370 35984
rect 14306 35924 14310 35980
rect 14310 35924 14366 35980
rect 14366 35924 14370 35980
rect 14306 35920 14370 35924
rect 14386 35980 14450 35984
rect 14386 35924 14390 35980
rect 14390 35924 14446 35980
rect 14446 35924 14450 35980
rect 14386 35920 14450 35924
rect 14466 35980 14530 35984
rect 14466 35924 14470 35980
rect 14470 35924 14526 35980
rect 14526 35924 14530 35980
rect 14466 35920 14530 35924
rect 14546 35980 14610 35984
rect 14546 35924 14550 35980
rect 14550 35924 14606 35980
rect 14606 35924 14610 35980
rect 14546 35920 14610 35924
rect 19634 35980 19698 35984
rect 19634 35924 19638 35980
rect 19638 35924 19694 35980
rect 19694 35924 19698 35980
rect 19634 35920 19698 35924
rect 19714 35980 19778 35984
rect 19714 35924 19718 35980
rect 19718 35924 19774 35980
rect 19774 35924 19778 35980
rect 19714 35920 19778 35924
rect 19794 35980 19858 35984
rect 19794 35924 19798 35980
rect 19798 35924 19854 35980
rect 19854 35924 19858 35980
rect 19794 35920 19858 35924
rect 19874 35980 19938 35984
rect 19874 35924 19878 35980
rect 19878 35924 19934 35980
rect 19934 35924 19938 35980
rect 19874 35920 19938 35924
rect 24962 35980 25026 35984
rect 24962 35924 24966 35980
rect 24966 35924 25022 35980
rect 25022 35924 25026 35980
rect 24962 35920 25026 35924
rect 25042 35980 25106 35984
rect 25042 35924 25046 35980
rect 25046 35924 25102 35980
rect 25102 35924 25106 35980
rect 25042 35920 25106 35924
rect 25122 35980 25186 35984
rect 25122 35924 25126 35980
rect 25126 35924 25182 35980
rect 25182 35924 25186 35980
rect 25122 35920 25186 35924
rect 25202 35980 25266 35984
rect 25202 35924 25206 35980
rect 25206 35924 25262 35980
rect 25262 35924 25266 35980
rect 25202 35920 25266 35924
rect 30290 35980 30354 35984
rect 30290 35924 30294 35980
rect 30294 35924 30350 35980
rect 30350 35924 30354 35980
rect 30290 35920 30354 35924
rect 30370 35980 30434 35984
rect 30370 35924 30374 35980
rect 30374 35924 30430 35980
rect 30430 35924 30434 35980
rect 30370 35920 30434 35924
rect 30450 35980 30514 35984
rect 30450 35924 30454 35980
rect 30454 35924 30510 35980
rect 30510 35924 30514 35980
rect 30450 35920 30514 35924
rect 30530 35980 30594 35984
rect 30530 35924 30534 35980
rect 30534 35924 30590 35980
rect 30590 35924 30594 35980
rect 30530 35920 30594 35924
rect 35618 35980 35682 35984
rect 35618 35924 35622 35980
rect 35622 35924 35678 35980
rect 35678 35924 35682 35980
rect 35618 35920 35682 35924
rect 35698 35980 35762 35984
rect 35698 35924 35702 35980
rect 35702 35924 35758 35980
rect 35758 35924 35762 35980
rect 35698 35920 35762 35924
rect 35778 35980 35842 35984
rect 35778 35924 35782 35980
rect 35782 35924 35838 35980
rect 35838 35924 35842 35980
rect 35778 35920 35842 35924
rect 35858 35980 35922 35984
rect 35858 35924 35862 35980
rect 35862 35924 35918 35980
rect 35918 35924 35922 35980
rect 35858 35920 35922 35924
rect 40946 35980 41010 35984
rect 40946 35924 40950 35980
rect 40950 35924 41006 35980
rect 41006 35924 41010 35980
rect 40946 35920 41010 35924
rect 41026 35980 41090 35984
rect 41026 35924 41030 35980
rect 41030 35924 41086 35980
rect 41086 35924 41090 35980
rect 41026 35920 41090 35924
rect 41106 35980 41170 35984
rect 41106 35924 41110 35980
rect 41110 35924 41166 35980
rect 41166 35924 41170 35980
rect 41106 35920 41170 35924
rect 41186 35980 41250 35984
rect 41186 35924 41190 35980
rect 41190 35924 41246 35980
rect 41246 35924 41250 35980
rect 41186 35920 41250 35924
rect 46274 35980 46338 35984
rect 46274 35924 46278 35980
rect 46278 35924 46334 35980
rect 46334 35924 46338 35980
rect 46274 35920 46338 35924
rect 46354 35980 46418 35984
rect 46354 35924 46358 35980
rect 46358 35924 46414 35980
rect 46414 35924 46418 35980
rect 46354 35920 46418 35924
rect 46434 35980 46498 35984
rect 46434 35924 46438 35980
rect 46438 35924 46494 35980
rect 46494 35924 46498 35980
rect 46434 35920 46498 35924
rect 46514 35980 46578 35984
rect 46514 35924 46518 35980
rect 46518 35924 46574 35980
rect 46574 35924 46578 35980
rect 46514 35920 46578 35924
rect 51602 35980 51666 35984
rect 51602 35924 51606 35980
rect 51606 35924 51662 35980
rect 51662 35924 51666 35980
rect 51602 35920 51666 35924
rect 51682 35980 51746 35984
rect 51682 35924 51686 35980
rect 51686 35924 51742 35980
rect 51742 35924 51746 35980
rect 51682 35920 51746 35924
rect 51762 35980 51826 35984
rect 51762 35924 51766 35980
rect 51766 35924 51822 35980
rect 51822 35924 51826 35980
rect 51762 35920 51826 35924
rect 51842 35980 51906 35984
rect 51842 35924 51846 35980
rect 51846 35924 51902 35980
rect 51902 35924 51906 35980
rect 51842 35920 51906 35924
rect 56930 35980 56994 35984
rect 56930 35924 56934 35980
rect 56934 35924 56990 35980
rect 56990 35924 56994 35980
rect 56930 35920 56994 35924
rect 57010 35980 57074 35984
rect 57010 35924 57014 35980
rect 57014 35924 57070 35980
rect 57070 35924 57074 35980
rect 57010 35920 57074 35924
rect 57090 35980 57154 35984
rect 57090 35924 57094 35980
rect 57094 35924 57150 35980
rect 57150 35924 57154 35980
rect 57090 35920 57154 35924
rect 57170 35980 57234 35984
rect 57170 35924 57174 35980
rect 57174 35924 57230 35980
rect 57230 35924 57234 35980
rect 57170 35920 57234 35924
rect 62258 35980 62322 35984
rect 62258 35924 62262 35980
rect 62262 35924 62318 35980
rect 62318 35924 62322 35980
rect 62258 35920 62322 35924
rect 62338 35980 62402 35984
rect 62338 35924 62342 35980
rect 62342 35924 62398 35980
rect 62398 35924 62402 35980
rect 62338 35920 62402 35924
rect 62418 35980 62482 35984
rect 62418 35924 62422 35980
rect 62422 35924 62478 35980
rect 62478 35924 62482 35980
rect 62418 35920 62482 35924
rect 62498 35980 62562 35984
rect 62498 35924 62502 35980
rect 62502 35924 62558 35980
rect 62558 35924 62562 35980
rect 62498 35920 62562 35924
rect 67586 35980 67650 35984
rect 67586 35924 67590 35980
rect 67590 35924 67646 35980
rect 67646 35924 67650 35980
rect 67586 35920 67650 35924
rect 67666 35980 67730 35984
rect 67666 35924 67670 35980
rect 67670 35924 67726 35980
rect 67726 35924 67730 35980
rect 67666 35920 67730 35924
rect 67746 35980 67810 35984
rect 67746 35924 67750 35980
rect 67750 35924 67806 35980
rect 67806 35924 67810 35980
rect 67746 35920 67810 35924
rect 67826 35980 67890 35984
rect 67826 35924 67830 35980
rect 67830 35924 67886 35980
rect 67886 35924 67890 35980
rect 67826 35920 67890 35924
rect 72914 35980 72978 35984
rect 72914 35924 72918 35980
rect 72918 35924 72974 35980
rect 72974 35924 72978 35980
rect 72914 35920 72978 35924
rect 72994 35980 73058 35984
rect 72994 35924 72998 35980
rect 72998 35924 73054 35980
rect 73054 35924 73058 35980
rect 72994 35920 73058 35924
rect 73074 35980 73138 35984
rect 73074 35924 73078 35980
rect 73078 35924 73134 35980
rect 73134 35924 73138 35980
rect 73074 35920 73138 35924
rect 73154 35980 73218 35984
rect 73154 35924 73158 35980
rect 73158 35924 73214 35980
rect 73214 35924 73218 35980
rect 73154 35920 73218 35924
rect 78242 35980 78306 35984
rect 78242 35924 78246 35980
rect 78246 35924 78302 35980
rect 78302 35924 78306 35980
rect 78242 35920 78306 35924
rect 78322 35980 78386 35984
rect 78322 35924 78326 35980
rect 78326 35924 78382 35980
rect 78382 35924 78386 35980
rect 78322 35920 78386 35924
rect 78402 35980 78466 35984
rect 78402 35924 78406 35980
rect 78406 35924 78462 35980
rect 78462 35924 78466 35980
rect 78402 35920 78466 35924
rect 78482 35980 78546 35984
rect 78482 35924 78486 35980
rect 78486 35924 78542 35980
rect 78542 35924 78546 35980
rect 78482 35920 78546 35924
rect 83570 35980 83634 35984
rect 83570 35924 83574 35980
rect 83574 35924 83630 35980
rect 83630 35924 83634 35980
rect 83570 35920 83634 35924
rect 83650 35980 83714 35984
rect 83650 35924 83654 35980
rect 83654 35924 83710 35980
rect 83710 35924 83714 35980
rect 83650 35920 83714 35924
rect 83730 35980 83794 35984
rect 83730 35924 83734 35980
rect 83734 35924 83790 35980
rect 83790 35924 83794 35980
rect 83730 35920 83794 35924
rect 83810 35980 83874 35984
rect 83810 35924 83814 35980
rect 83814 35924 83870 35980
rect 83870 35924 83874 35980
rect 83810 35920 83874 35924
rect 88898 35980 88962 35984
rect 88898 35924 88902 35980
rect 88902 35924 88958 35980
rect 88958 35924 88962 35980
rect 88898 35920 88962 35924
rect 88978 35980 89042 35984
rect 88978 35924 88982 35980
rect 88982 35924 89038 35980
rect 89038 35924 89042 35980
rect 88978 35920 89042 35924
rect 89058 35980 89122 35984
rect 89058 35924 89062 35980
rect 89062 35924 89118 35980
rect 89118 35924 89122 35980
rect 89058 35920 89122 35924
rect 89138 35980 89202 35984
rect 89138 35924 89142 35980
rect 89142 35924 89198 35980
rect 89198 35924 89202 35980
rect 89138 35920 89202 35924
rect 6314 35436 6378 35440
rect 6314 35380 6318 35436
rect 6318 35380 6374 35436
rect 6374 35380 6378 35436
rect 6314 35376 6378 35380
rect 6394 35436 6458 35440
rect 6394 35380 6398 35436
rect 6398 35380 6454 35436
rect 6454 35380 6458 35436
rect 6394 35376 6458 35380
rect 6474 35436 6538 35440
rect 6474 35380 6478 35436
rect 6478 35380 6534 35436
rect 6534 35380 6538 35436
rect 6474 35376 6538 35380
rect 6554 35436 6618 35440
rect 6554 35380 6558 35436
rect 6558 35380 6614 35436
rect 6614 35380 6618 35436
rect 6554 35376 6618 35380
rect 11642 35436 11706 35440
rect 11642 35380 11646 35436
rect 11646 35380 11702 35436
rect 11702 35380 11706 35436
rect 11642 35376 11706 35380
rect 11722 35436 11786 35440
rect 11722 35380 11726 35436
rect 11726 35380 11782 35436
rect 11782 35380 11786 35436
rect 11722 35376 11786 35380
rect 11802 35436 11866 35440
rect 11802 35380 11806 35436
rect 11806 35380 11862 35436
rect 11862 35380 11866 35436
rect 11802 35376 11866 35380
rect 11882 35436 11946 35440
rect 11882 35380 11886 35436
rect 11886 35380 11942 35436
rect 11942 35380 11946 35436
rect 11882 35376 11946 35380
rect 16970 35436 17034 35440
rect 16970 35380 16974 35436
rect 16974 35380 17030 35436
rect 17030 35380 17034 35436
rect 16970 35376 17034 35380
rect 17050 35436 17114 35440
rect 17050 35380 17054 35436
rect 17054 35380 17110 35436
rect 17110 35380 17114 35436
rect 17050 35376 17114 35380
rect 17130 35436 17194 35440
rect 17130 35380 17134 35436
rect 17134 35380 17190 35436
rect 17190 35380 17194 35436
rect 17130 35376 17194 35380
rect 17210 35436 17274 35440
rect 17210 35380 17214 35436
rect 17214 35380 17270 35436
rect 17270 35380 17274 35436
rect 17210 35376 17274 35380
rect 22298 35436 22362 35440
rect 22298 35380 22302 35436
rect 22302 35380 22358 35436
rect 22358 35380 22362 35436
rect 22298 35376 22362 35380
rect 22378 35436 22442 35440
rect 22378 35380 22382 35436
rect 22382 35380 22438 35436
rect 22438 35380 22442 35436
rect 22378 35376 22442 35380
rect 22458 35436 22522 35440
rect 22458 35380 22462 35436
rect 22462 35380 22518 35436
rect 22518 35380 22522 35436
rect 22458 35376 22522 35380
rect 22538 35436 22602 35440
rect 22538 35380 22542 35436
rect 22542 35380 22598 35436
rect 22598 35380 22602 35436
rect 22538 35376 22602 35380
rect 27626 35436 27690 35440
rect 27626 35380 27630 35436
rect 27630 35380 27686 35436
rect 27686 35380 27690 35436
rect 27626 35376 27690 35380
rect 27706 35436 27770 35440
rect 27706 35380 27710 35436
rect 27710 35380 27766 35436
rect 27766 35380 27770 35436
rect 27706 35376 27770 35380
rect 27786 35436 27850 35440
rect 27786 35380 27790 35436
rect 27790 35380 27846 35436
rect 27846 35380 27850 35436
rect 27786 35376 27850 35380
rect 27866 35436 27930 35440
rect 27866 35380 27870 35436
rect 27870 35380 27926 35436
rect 27926 35380 27930 35436
rect 27866 35376 27930 35380
rect 32954 35436 33018 35440
rect 32954 35380 32958 35436
rect 32958 35380 33014 35436
rect 33014 35380 33018 35436
rect 32954 35376 33018 35380
rect 33034 35436 33098 35440
rect 33034 35380 33038 35436
rect 33038 35380 33094 35436
rect 33094 35380 33098 35436
rect 33034 35376 33098 35380
rect 33114 35436 33178 35440
rect 33114 35380 33118 35436
rect 33118 35380 33174 35436
rect 33174 35380 33178 35436
rect 33114 35376 33178 35380
rect 33194 35436 33258 35440
rect 33194 35380 33198 35436
rect 33198 35380 33254 35436
rect 33254 35380 33258 35436
rect 33194 35376 33258 35380
rect 38282 35436 38346 35440
rect 38282 35380 38286 35436
rect 38286 35380 38342 35436
rect 38342 35380 38346 35436
rect 38282 35376 38346 35380
rect 38362 35436 38426 35440
rect 38362 35380 38366 35436
rect 38366 35380 38422 35436
rect 38422 35380 38426 35436
rect 38362 35376 38426 35380
rect 38442 35436 38506 35440
rect 38442 35380 38446 35436
rect 38446 35380 38502 35436
rect 38502 35380 38506 35436
rect 38442 35376 38506 35380
rect 38522 35436 38586 35440
rect 38522 35380 38526 35436
rect 38526 35380 38582 35436
rect 38582 35380 38586 35436
rect 38522 35376 38586 35380
rect 43610 35436 43674 35440
rect 43610 35380 43614 35436
rect 43614 35380 43670 35436
rect 43670 35380 43674 35436
rect 43610 35376 43674 35380
rect 43690 35436 43754 35440
rect 43690 35380 43694 35436
rect 43694 35380 43750 35436
rect 43750 35380 43754 35436
rect 43690 35376 43754 35380
rect 43770 35436 43834 35440
rect 43770 35380 43774 35436
rect 43774 35380 43830 35436
rect 43830 35380 43834 35436
rect 43770 35376 43834 35380
rect 43850 35436 43914 35440
rect 43850 35380 43854 35436
rect 43854 35380 43910 35436
rect 43910 35380 43914 35436
rect 43850 35376 43914 35380
rect 48938 35436 49002 35440
rect 48938 35380 48942 35436
rect 48942 35380 48998 35436
rect 48998 35380 49002 35436
rect 48938 35376 49002 35380
rect 49018 35436 49082 35440
rect 49018 35380 49022 35436
rect 49022 35380 49078 35436
rect 49078 35380 49082 35436
rect 49018 35376 49082 35380
rect 49098 35436 49162 35440
rect 49098 35380 49102 35436
rect 49102 35380 49158 35436
rect 49158 35380 49162 35436
rect 49098 35376 49162 35380
rect 49178 35436 49242 35440
rect 49178 35380 49182 35436
rect 49182 35380 49238 35436
rect 49238 35380 49242 35436
rect 49178 35376 49242 35380
rect 54266 35436 54330 35440
rect 54266 35380 54270 35436
rect 54270 35380 54326 35436
rect 54326 35380 54330 35436
rect 54266 35376 54330 35380
rect 54346 35436 54410 35440
rect 54346 35380 54350 35436
rect 54350 35380 54406 35436
rect 54406 35380 54410 35436
rect 54346 35376 54410 35380
rect 54426 35436 54490 35440
rect 54426 35380 54430 35436
rect 54430 35380 54486 35436
rect 54486 35380 54490 35436
rect 54426 35376 54490 35380
rect 54506 35436 54570 35440
rect 54506 35380 54510 35436
rect 54510 35380 54566 35436
rect 54566 35380 54570 35436
rect 54506 35376 54570 35380
rect 59594 35436 59658 35440
rect 59594 35380 59598 35436
rect 59598 35380 59654 35436
rect 59654 35380 59658 35436
rect 59594 35376 59658 35380
rect 59674 35436 59738 35440
rect 59674 35380 59678 35436
rect 59678 35380 59734 35436
rect 59734 35380 59738 35436
rect 59674 35376 59738 35380
rect 59754 35436 59818 35440
rect 59754 35380 59758 35436
rect 59758 35380 59814 35436
rect 59814 35380 59818 35436
rect 59754 35376 59818 35380
rect 59834 35436 59898 35440
rect 59834 35380 59838 35436
rect 59838 35380 59894 35436
rect 59894 35380 59898 35436
rect 59834 35376 59898 35380
rect 64922 35436 64986 35440
rect 64922 35380 64926 35436
rect 64926 35380 64982 35436
rect 64982 35380 64986 35436
rect 64922 35376 64986 35380
rect 65002 35436 65066 35440
rect 65002 35380 65006 35436
rect 65006 35380 65062 35436
rect 65062 35380 65066 35436
rect 65002 35376 65066 35380
rect 65082 35436 65146 35440
rect 65082 35380 65086 35436
rect 65086 35380 65142 35436
rect 65142 35380 65146 35436
rect 65082 35376 65146 35380
rect 65162 35436 65226 35440
rect 65162 35380 65166 35436
rect 65166 35380 65222 35436
rect 65222 35380 65226 35436
rect 65162 35376 65226 35380
rect 70250 35436 70314 35440
rect 70250 35380 70254 35436
rect 70254 35380 70310 35436
rect 70310 35380 70314 35436
rect 70250 35376 70314 35380
rect 70330 35436 70394 35440
rect 70330 35380 70334 35436
rect 70334 35380 70390 35436
rect 70390 35380 70394 35436
rect 70330 35376 70394 35380
rect 70410 35436 70474 35440
rect 70410 35380 70414 35436
rect 70414 35380 70470 35436
rect 70470 35380 70474 35436
rect 70410 35376 70474 35380
rect 70490 35436 70554 35440
rect 70490 35380 70494 35436
rect 70494 35380 70550 35436
rect 70550 35380 70554 35436
rect 70490 35376 70554 35380
rect 75578 35436 75642 35440
rect 75578 35380 75582 35436
rect 75582 35380 75638 35436
rect 75638 35380 75642 35436
rect 75578 35376 75642 35380
rect 75658 35436 75722 35440
rect 75658 35380 75662 35436
rect 75662 35380 75718 35436
rect 75718 35380 75722 35436
rect 75658 35376 75722 35380
rect 75738 35436 75802 35440
rect 75738 35380 75742 35436
rect 75742 35380 75798 35436
rect 75798 35380 75802 35436
rect 75738 35376 75802 35380
rect 75818 35436 75882 35440
rect 75818 35380 75822 35436
rect 75822 35380 75878 35436
rect 75878 35380 75882 35436
rect 75818 35376 75882 35380
rect 80906 35436 80970 35440
rect 80906 35380 80910 35436
rect 80910 35380 80966 35436
rect 80966 35380 80970 35436
rect 80906 35376 80970 35380
rect 80986 35436 81050 35440
rect 80986 35380 80990 35436
rect 80990 35380 81046 35436
rect 81046 35380 81050 35436
rect 80986 35376 81050 35380
rect 81066 35436 81130 35440
rect 81066 35380 81070 35436
rect 81070 35380 81126 35436
rect 81126 35380 81130 35436
rect 81066 35376 81130 35380
rect 81146 35436 81210 35440
rect 81146 35380 81150 35436
rect 81150 35380 81206 35436
rect 81206 35380 81210 35436
rect 81146 35376 81210 35380
rect 86234 35436 86298 35440
rect 86234 35380 86238 35436
rect 86238 35380 86294 35436
rect 86294 35380 86298 35436
rect 86234 35376 86298 35380
rect 86314 35436 86378 35440
rect 86314 35380 86318 35436
rect 86318 35380 86374 35436
rect 86374 35380 86378 35436
rect 86314 35376 86378 35380
rect 86394 35436 86458 35440
rect 86394 35380 86398 35436
rect 86398 35380 86454 35436
rect 86454 35380 86458 35436
rect 86394 35376 86458 35380
rect 86474 35436 86538 35440
rect 86474 35380 86478 35436
rect 86478 35380 86534 35436
rect 86534 35380 86538 35436
rect 86474 35376 86538 35380
rect 91562 35436 91626 35440
rect 91562 35380 91566 35436
rect 91566 35380 91622 35436
rect 91622 35380 91626 35436
rect 91562 35376 91626 35380
rect 91642 35436 91706 35440
rect 91642 35380 91646 35436
rect 91646 35380 91702 35436
rect 91702 35380 91706 35436
rect 91642 35376 91706 35380
rect 91722 35436 91786 35440
rect 91722 35380 91726 35436
rect 91726 35380 91782 35436
rect 91782 35380 91786 35436
rect 91722 35376 91786 35380
rect 91802 35436 91866 35440
rect 91802 35380 91806 35436
rect 91806 35380 91862 35436
rect 91862 35380 91866 35436
rect 91802 35376 91866 35380
rect 3650 34892 3714 34896
rect 3650 34836 3654 34892
rect 3654 34836 3710 34892
rect 3710 34836 3714 34892
rect 3650 34832 3714 34836
rect 3730 34892 3794 34896
rect 3730 34836 3734 34892
rect 3734 34836 3790 34892
rect 3790 34836 3794 34892
rect 3730 34832 3794 34836
rect 3810 34892 3874 34896
rect 3810 34836 3814 34892
rect 3814 34836 3870 34892
rect 3870 34836 3874 34892
rect 3810 34832 3874 34836
rect 3890 34892 3954 34896
rect 3890 34836 3894 34892
rect 3894 34836 3950 34892
rect 3950 34836 3954 34892
rect 3890 34832 3954 34836
rect 8978 34892 9042 34896
rect 8978 34836 8982 34892
rect 8982 34836 9038 34892
rect 9038 34836 9042 34892
rect 8978 34832 9042 34836
rect 9058 34892 9122 34896
rect 9058 34836 9062 34892
rect 9062 34836 9118 34892
rect 9118 34836 9122 34892
rect 9058 34832 9122 34836
rect 9138 34892 9202 34896
rect 9138 34836 9142 34892
rect 9142 34836 9198 34892
rect 9198 34836 9202 34892
rect 9138 34832 9202 34836
rect 9218 34892 9282 34896
rect 9218 34836 9222 34892
rect 9222 34836 9278 34892
rect 9278 34836 9282 34892
rect 9218 34832 9282 34836
rect 14306 34892 14370 34896
rect 14306 34836 14310 34892
rect 14310 34836 14366 34892
rect 14366 34836 14370 34892
rect 14306 34832 14370 34836
rect 14386 34892 14450 34896
rect 14386 34836 14390 34892
rect 14390 34836 14446 34892
rect 14446 34836 14450 34892
rect 14386 34832 14450 34836
rect 14466 34892 14530 34896
rect 14466 34836 14470 34892
rect 14470 34836 14526 34892
rect 14526 34836 14530 34892
rect 14466 34832 14530 34836
rect 14546 34892 14610 34896
rect 14546 34836 14550 34892
rect 14550 34836 14606 34892
rect 14606 34836 14610 34892
rect 14546 34832 14610 34836
rect 19634 34892 19698 34896
rect 19634 34836 19638 34892
rect 19638 34836 19694 34892
rect 19694 34836 19698 34892
rect 19634 34832 19698 34836
rect 19714 34892 19778 34896
rect 19714 34836 19718 34892
rect 19718 34836 19774 34892
rect 19774 34836 19778 34892
rect 19714 34832 19778 34836
rect 19794 34892 19858 34896
rect 19794 34836 19798 34892
rect 19798 34836 19854 34892
rect 19854 34836 19858 34892
rect 19794 34832 19858 34836
rect 19874 34892 19938 34896
rect 19874 34836 19878 34892
rect 19878 34836 19934 34892
rect 19934 34836 19938 34892
rect 19874 34832 19938 34836
rect 24962 34892 25026 34896
rect 24962 34836 24966 34892
rect 24966 34836 25022 34892
rect 25022 34836 25026 34892
rect 24962 34832 25026 34836
rect 25042 34892 25106 34896
rect 25042 34836 25046 34892
rect 25046 34836 25102 34892
rect 25102 34836 25106 34892
rect 25042 34832 25106 34836
rect 25122 34892 25186 34896
rect 25122 34836 25126 34892
rect 25126 34836 25182 34892
rect 25182 34836 25186 34892
rect 25122 34832 25186 34836
rect 25202 34892 25266 34896
rect 25202 34836 25206 34892
rect 25206 34836 25262 34892
rect 25262 34836 25266 34892
rect 25202 34832 25266 34836
rect 30290 34892 30354 34896
rect 30290 34836 30294 34892
rect 30294 34836 30350 34892
rect 30350 34836 30354 34892
rect 30290 34832 30354 34836
rect 30370 34892 30434 34896
rect 30370 34836 30374 34892
rect 30374 34836 30430 34892
rect 30430 34836 30434 34892
rect 30370 34832 30434 34836
rect 30450 34892 30514 34896
rect 30450 34836 30454 34892
rect 30454 34836 30510 34892
rect 30510 34836 30514 34892
rect 30450 34832 30514 34836
rect 30530 34892 30594 34896
rect 30530 34836 30534 34892
rect 30534 34836 30590 34892
rect 30590 34836 30594 34892
rect 30530 34832 30594 34836
rect 35618 34892 35682 34896
rect 35618 34836 35622 34892
rect 35622 34836 35678 34892
rect 35678 34836 35682 34892
rect 35618 34832 35682 34836
rect 35698 34892 35762 34896
rect 35698 34836 35702 34892
rect 35702 34836 35758 34892
rect 35758 34836 35762 34892
rect 35698 34832 35762 34836
rect 35778 34892 35842 34896
rect 35778 34836 35782 34892
rect 35782 34836 35838 34892
rect 35838 34836 35842 34892
rect 35778 34832 35842 34836
rect 35858 34892 35922 34896
rect 35858 34836 35862 34892
rect 35862 34836 35918 34892
rect 35918 34836 35922 34892
rect 35858 34832 35922 34836
rect 40946 34892 41010 34896
rect 40946 34836 40950 34892
rect 40950 34836 41006 34892
rect 41006 34836 41010 34892
rect 40946 34832 41010 34836
rect 41026 34892 41090 34896
rect 41026 34836 41030 34892
rect 41030 34836 41086 34892
rect 41086 34836 41090 34892
rect 41026 34832 41090 34836
rect 41106 34892 41170 34896
rect 41106 34836 41110 34892
rect 41110 34836 41166 34892
rect 41166 34836 41170 34892
rect 41106 34832 41170 34836
rect 41186 34892 41250 34896
rect 41186 34836 41190 34892
rect 41190 34836 41246 34892
rect 41246 34836 41250 34892
rect 41186 34832 41250 34836
rect 46274 34892 46338 34896
rect 46274 34836 46278 34892
rect 46278 34836 46334 34892
rect 46334 34836 46338 34892
rect 46274 34832 46338 34836
rect 46354 34892 46418 34896
rect 46354 34836 46358 34892
rect 46358 34836 46414 34892
rect 46414 34836 46418 34892
rect 46354 34832 46418 34836
rect 46434 34892 46498 34896
rect 46434 34836 46438 34892
rect 46438 34836 46494 34892
rect 46494 34836 46498 34892
rect 46434 34832 46498 34836
rect 46514 34892 46578 34896
rect 46514 34836 46518 34892
rect 46518 34836 46574 34892
rect 46574 34836 46578 34892
rect 46514 34832 46578 34836
rect 51602 34892 51666 34896
rect 51602 34836 51606 34892
rect 51606 34836 51662 34892
rect 51662 34836 51666 34892
rect 51602 34832 51666 34836
rect 51682 34892 51746 34896
rect 51682 34836 51686 34892
rect 51686 34836 51742 34892
rect 51742 34836 51746 34892
rect 51682 34832 51746 34836
rect 51762 34892 51826 34896
rect 51762 34836 51766 34892
rect 51766 34836 51822 34892
rect 51822 34836 51826 34892
rect 51762 34832 51826 34836
rect 51842 34892 51906 34896
rect 51842 34836 51846 34892
rect 51846 34836 51902 34892
rect 51902 34836 51906 34892
rect 51842 34832 51906 34836
rect 56930 34892 56994 34896
rect 56930 34836 56934 34892
rect 56934 34836 56990 34892
rect 56990 34836 56994 34892
rect 56930 34832 56994 34836
rect 57010 34892 57074 34896
rect 57010 34836 57014 34892
rect 57014 34836 57070 34892
rect 57070 34836 57074 34892
rect 57010 34832 57074 34836
rect 57090 34892 57154 34896
rect 57090 34836 57094 34892
rect 57094 34836 57150 34892
rect 57150 34836 57154 34892
rect 57090 34832 57154 34836
rect 57170 34892 57234 34896
rect 57170 34836 57174 34892
rect 57174 34836 57230 34892
rect 57230 34836 57234 34892
rect 57170 34832 57234 34836
rect 62258 34892 62322 34896
rect 62258 34836 62262 34892
rect 62262 34836 62318 34892
rect 62318 34836 62322 34892
rect 62258 34832 62322 34836
rect 62338 34892 62402 34896
rect 62338 34836 62342 34892
rect 62342 34836 62398 34892
rect 62398 34836 62402 34892
rect 62338 34832 62402 34836
rect 62418 34892 62482 34896
rect 62418 34836 62422 34892
rect 62422 34836 62478 34892
rect 62478 34836 62482 34892
rect 62418 34832 62482 34836
rect 62498 34892 62562 34896
rect 62498 34836 62502 34892
rect 62502 34836 62558 34892
rect 62558 34836 62562 34892
rect 62498 34832 62562 34836
rect 67586 34892 67650 34896
rect 67586 34836 67590 34892
rect 67590 34836 67646 34892
rect 67646 34836 67650 34892
rect 67586 34832 67650 34836
rect 67666 34892 67730 34896
rect 67666 34836 67670 34892
rect 67670 34836 67726 34892
rect 67726 34836 67730 34892
rect 67666 34832 67730 34836
rect 67746 34892 67810 34896
rect 67746 34836 67750 34892
rect 67750 34836 67806 34892
rect 67806 34836 67810 34892
rect 67746 34832 67810 34836
rect 67826 34892 67890 34896
rect 67826 34836 67830 34892
rect 67830 34836 67886 34892
rect 67886 34836 67890 34892
rect 67826 34832 67890 34836
rect 72914 34892 72978 34896
rect 72914 34836 72918 34892
rect 72918 34836 72974 34892
rect 72974 34836 72978 34892
rect 72914 34832 72978 34836
rect 72994 34892 73058 34896
rect 72994 34836 72998 34892
rect 72998 34836 73054 34892
rect 73054 34836 73058 34892
rect 72994 34832 73058 34836
rect 73074 34892 73138 34896
rect 73074 34836 73078 34892
rect 73078 34836 73134 34892
rect 73134 34836 73138 34892
rect 73074 34832 73138 34836
rect 73154 34892 73218 34896
rect 73154 34836 73158 34892
rect 73158 34836 73214 34892
rect 73214 34836 73218 34892
rect 73154 34832 73218 34836
rect 78242 34892 78306 34896
rect 78242 34836 78246 34892
rect 78246 34836 78302 34892
rect 78302 34836 78306 34892
rect 78242 34832 78306 34836
rect 78322 34892 78386 34896
rect 78322 34836 78326 34892
rect 78326 34836 78382 34892
rect 78382 34836 78386 34892
rect 78322 34832 78386 34836
rect 78402 34892 78466 34896
rect 78402 34836 78406 34892
rect 78406 34836 78462 34892
rect 78462 34836 78466 34892
rect 78402 34832 78466 34836
rect 78482 34892 78546 34896
rect 78482 34836 78486 34892
rect 78486 34836 78542 34892
rect 78542 34836 78546 34892
rect 78482 34832 78546 34836
rect 83570 34892 83634 34896
rect 83570 34836 83574 34892
rect 83574 34836 83630 34892
rect 83630 34836 83634 34892
rect 83570 34832 83634 34836
rect 83650 34892 83714 34896
rect 83650 34836 83654 34892
rect 83654 34836 83710 34892
rect 83710 34836 83714 34892
rect 83650 34832 83714 34836
rect 83730 34892 83794 34896
rect 83730 34836 83734 34892
rect 83734 34836 83790 34892
rect 83790 34836 83794 34892
rect 83730 34832 83794 34836
rect 83810 34892 83874 34896
rect 83810 34836 83814 34892
rect 83814 34836 83870 34892
rect 83870 34836 83874 34892
rect 83810 34832 83874 34836
rect 88898 34892 88962 34896
rect 88898 34836 88902 34892
rect 88902 34836 88958 34892
rect 88958 34836 88962 34892
rect 88898 34832 88962 34836
rect 88978 34892 89042 34896
rect 88978 34836 88982 34892
rect 88982 34836 89038 34892
rect 89038 34836 89042 34892
rect 88978 34832 89042 34836
rect 89058 34892 89122 34896
rect 89058 34836 89062 34892
rect 89062 34836 89118 34892
rect 89118 34836 89122 34892
rect 89058 34832 89122 34836
rect 89138 34892 89202 34896
rect 89138 34836 89142 34892
rect 89142 34836 89198 34892
rect 89198 34836 89202 34892
rect 89138 34832 89202 34836
rect 6314 34348 6378 34352
rect 6314 34292 6318 34348
rect 6318 34292 6374 34348
rect 6374 34292 6378 34348
rect 6314 34288 6378 34292
rect 6394 34348 6458 34352
rect 6394 34292 6398 34348
rect 6398 34292 6454 34348
rect 6454 34292 6458 34348
rect 6394 34288 6458 34292
rect 6474 34348 6538 34352
rect 6474 34292 6478 34348
rect 6478 34292 6534 34348
rect 6534 34292 6538 34348
rect 6474 34288 6538 34292
rect 6554 34348 6618 34352
rect 6554 34292 6558 34348
rect 6558 34292 6614 34348
rect 6614 34292 6618 34348
rect 6554 34288 6618 34292
rect 11642 34348 11706 34352
rect 11642 34292 11646 34348
rect 11646 34292 11702 34348
rect 11702 34292 11706 34348
rect 11642 34288 11706 34292
rect 11722 34348 11786 34352
rect 11722 34292 11726 34348
rect 11726 34292 11782 34348
rect 11782 34292 11786 34348
rect 11722 34288 11786 34292
rect 11802 34348 11866 34352
rect 11802 34292 11806 34348
rect 11806 34292 11862 34348
rect 11862 34292 11866 34348
rect 11802 34288 11866 34292
rect 11882 34348 11946 34352
rect 11882 34292 11886 34348
rect 11886 34292 11942 34348
rect 11942 34292 11946 34348
rect 11882 34288 11946 34292
rect 16970 34348 17034 34352
rect 16970 34292 16974 34348
rect 16974 34292 17030 34348
rect 17030 34292 17034 34348
rect 16970 34288 17034 34292
rect 17050 34348 17114 34352
rect 17050 34292 17054 34348
rect 17054 34292 17110 34348
rect 17110 34292 17114 34348
rect 17050 34288 17114 34292
rect 17130 34348 17194 34352
rect 17130 34292 17134 34348
rect 17134 34292 17190 34348
rect 17190 34292 17194 34348
rect 17130 34288 17194 34292
rect 17210 34348 17274 34352
rect 17210 34292 17214 34348
rect 17214 34292 17270 34348
rect 17270 34292 17274 34348
rect 17210 34288 17274 34292
rect 22298 34348 22362 34352
rect 22298 34292 22302 34348
rect 22302 34292 22358 34348
rect 22358 34292 22362 34348
rect 22298 34288 22362 34292
rect 22378 34348 22442 34352
rect 22378 34292 22382 34348
rect 22382 34292 22438 34348
rect 22438 34292 22442 34348
rect 22378 34288 22442 34292
rect 22458 34348 22522 34352
rect 22458 34292 22462 34348
rect 22462 34292 22518 34348
rect 22518 34292 22522 34348
rect 22458 34288 22522 34292
rect 22538 34348 22602 34352
rect 22538 34292 22542 34348
rect 22542 34292 22598 34348
rect 22598 34292 22602 34348
rect 22538 34288 22602 34292
rect 27626 34348 27690 34352
rect 27626 34292 27630 34348
rect 27630 34292 27686 34348
rect 27686 34292 27690 34348
rect 27626 34288 27690 34292
rect 27706 34348 27770 34352
rect 27706 34292 27710 34348
rect 27710 34292 27766 34348
rect 27766 34292 27770 34348
rect 27706 34288 27770 34292
rect 27786 34348 27850 34352
rect 27786 34292 27790 34348
rect 27790 34292 27846 34348
rect 27846 34292 27850 34348
rect 27786 34288 27850 34292
rect 27866 34348 27930 34352
rect 27866 34292 27870 34348
rect 27870 34292 27926 34348
rect 27926 34292 27930 34348
rect 27866 34288 27930 34292
rect 32954 34348 33018 34352
rect 32954 34292 32958 34348
rect 32958 34292 33014 34348
rect 33014 34292 33018 34348
rect 32954 34288 33018 34292
rect 33034 34348 33098 34352
rect 33034 34292 33038 34348
rect 33038 34292 33094 34348
rect 33094 34292 33098 34348
rect 33034 34288 33098 34292
rect 33114 34348 33178 34352
rect 33114 34292 33118 34348
rect 33118 34292 33174 34348
rect 33174 34292 33178 34348
rect 33114 34288 33178 34292
rect 33194 34348 33258 34352
rect 33194 34292 33198 34348
rect 33198 34292 33254 34348
rect 33254 34292 33258 34348
rect 33194 34288 33258 34292
rect 38282 34348 38346 34352
rect 38282 34292 38286 34348
rect 38286 34292 38342 34348
rect 38342 34292 38346 34348
rect 38282 34288 38346 34292
rect 38362 34348 38426 34352
rect 38362 34292 38366 34348
rect 38366 34292 38422 34348
rect 38422 34292 38426 34348
rect 38362 34288 38426 34292
rect 38442 34348 38506 34352
rect 38442 34292 38446 34348
rect 38446 34292 38502 34348
rect 38502 34292 38506 34348
rect 38442 34288 38506 34292
rect 38522 34348 38586 34352
rect 38522 34292 38526 34348
rect 38526 34292 38582 34348
rect 38582 34292 38586 34348
rect 38522 34288 38586 34292
rect 43610 34348 43674 34352
rect 43610 34292 43614 34348
rect 43614 34292 43670 34348
rect 43670 34292 43674 34348
rect 43610 34288 43674 34292
rect 43690 34348 43754 34352
rect 43690 34292 43694 34348
rect 43694 34292 43750 34348
rect 43750 34292 43754 34348
rect 43690 34288 43754 34292
rect 43770 34348 43834 34352
rect 43770 34292 43774 34348
rect 43774 34292 43830 34348
rect 43830 34292 43834 34348
rect 43770 34288 43834 34292
rect 43850 34348 43914 34352
rect 43850 34292 43854 34348
rect 43854 34292 43910 34348
rect 43910 34292 43914 34348
rect 43850 34288 43914 34292
rect 48938 34348 49002 34352
rect 48938 34292 48942 34348
rect 48942 34292 48998 34348
rect 48998 34292 49002 34348
rect 48938 34288 49002 34292
rect 49018 34348 49082 34352
rect 49018 34292 49022 34348
rect 49022 34292 49078 34348
rect 49078 34292 49082 34348
rect 49018 34288 49082 34292
rect 49098 34348 49162 34352
rect 49098 34292 49102 34348
rect 49102 34292 49158 34348
rect 49158 34292 49162 34348
rect 49098 34288 49162 34292
rect 49178 34348 49242 34352
rect 49178 34292 49182 34348
rect 49182 34292 49238 34348
rect 49238 34292 49242 34348
rect 49178 34288 49242 34292
rect 54266 34348 54330 34352
rect 54266 34292 54270 34348
rect 54270 34292 54326 34348
rect 54326 34292 54330 34348
rect 54266 34288 54330 34292
rect 54346 34348 54410 34352
rect 54346 34292 54350 34348
rect 54350 34292 54406 34348
rect 54406 34292 54410 34348
rect 54346 34288 54410 34292
rect 54426 34348 54490 34352
rect 54426 34292 54430 34348
rect 54430 34292 54486 34348
rect 54486 34292 54490 34348
rect 54426 34288 54490 34292
rect 54506 34348 54570 34352
rect 54506 34292 54510 34348
rect 54510 34292 54566 34348
rect 54566 34292 54570 34348
rect 54506 34288 54570 34292
rect 59594 34348 59658 34352
rect 59594 34292 59598 34348
rect 59598 34292 59654 34348
rect 59654 34292 59658 34348
rect 59594 34288 59658 34292
rect 59674 34348 59738 34352
rect 59674 34292 59678 34348
rect 59678 34292 59734 34348
rect 59734 34292 59738 34348
rect 59674 34288 59738 34292
rect 59754 34348 59818 34352
rect 59754 34292 59758 34348
rect 59758 34292 59814 34348
rect 59814 34292 59818 34348
rect 59754 34288 59818 34292
rect 59834 34348 59898 34352
rect 59834 34292 59838 34348
rect 59838 34292 59894 34348
rect 59894 34292 59898 34348
rect 59834 34288 59898 34292
rect 64922 34348 64986 34352
rect 64922 34292 64926 34348
rect 64926 34292 64982 34348
rect 64982 34292 64986 34348
rect 64922 34288 64986 34292
rect 65002 34348 65066 34352
rect 65002 34292 65006 34348
rect 65006 34292 65062 34348
rect 65062 34292 65066 34348
rect 65002 34288 65066 34292
rect 65082 34348 65146 34352
rect 65082 34292 65086 34348
rect 65086 34292 65142 34348
rect 65142 34292 65146 34348
rect 65082 34288 65146 34292
rect 65162 34348 65226 34352
rect 65162 34292 65166 34348
rect 65166 34292 65222 34348
rect 65222 34292 65226 34348
rect 65162 34288 65226 34292
rect 70250 34348 70314 34352
rect 70250 34292 70254 34348
rect 70254 34292 70310 34348
rect 70310 34292 70314 34348
rect 70250 34288 70314 34292
rect 70330 34348 70394 34352
rect 70330 34292 70334 34348
rect 70334 34292 70390 34348
rect 70390 34292 70394 34348
rect 70330 34288 70394 34292
rect 70410 34348 70474 34352
rect 70410 34292 70414 34348
rect 70414 34292 70470 34348
rect 70470 34292 70474 34348
rect 70410 34288 70474 34292
rect 70490 34348 70554 34352
rect 70490 34292 70494 34348
rect 70494 34292 70550 34348
rect 70550 34292 70554 34348
rect 70490 34288 70554 34292
rect 75578 34348 75642 34352
rect 75578 34292 75582 34348
rect 75582 34292 75638 34348
rect 75638 34292 75642 34348
rect 75578 34288 75642 34292
rect 75658 34348 75722 34352
rect 75658 34292 75662 34348
rect 75662 34292 75718 34348
rect 75718 34292 75722 34348
rect 75658 34288 75722 34292
rect 75738 34348 75802 34352
rect 75738 34292 75742 34348
rect 75742 34292 75798 34348
rect 75798 34292 75802 34348
rect 75738 34288 75802 34292
rect 75818 34348 75882 34352
rect 75818 34292 75822 34348
rect 75822 34292 75878 34348
rect 75878 34292 75882 34348
rect 75818 34288 75882 34292
rect 80906 34348 80970 34352
rect 80906 34292 80910 34348
rect 80910 34292 80966 34348
rect 80966 34292 80970 34348
rect 80906 34288 80970 34292
rect 80986 34348 81050 34352
rect 80986 34292 80990 34348
rect 80990 34292 81046 34348
rect 81046 34292 81050 34348
rect 80986 34288 81050 34292
rect 81066 34348 81130 34352
rect 81066 34292 81070 34348
rect 81070 34292 81126 34348
rect 81126 34292 81130 34348
rect 81066 34288 81130 34292
rect 81146 34348 81210 34352
rect 81146 34292 81150 34348
rect 81150 34292 81206 34348
rect 81206 34292 81210 34348
rect 81146 34288 81210 34292
rect 86234 34348 86298 34352
rect 86234 34292 86238 34348
rect 86238 34292 86294 34348
rect 86294 34292 86298 34348
rect 86234 34288 86298 34292
rect 86314 34348 86378 34352
rect 86314 34292 86318 34348
rect 86318 34292 86374 34348
rect 86374 34292 86378 34348
rect 86314 34288 86378 34292
rect 86394 34348 86458 34352
rect 86394 34292 86398 34348
rect 86398 34292 86454 34348
rect 86454 34292 86458 34348
rect 86394 34288 86458 34292
rect 86474 34348 86538 34352
rect 86474 34292 86478 34348
rect 86478 34292 86534 34348
rect 86534 34292 86538 34348
rect 86474 34288 86538 34292
rect 91562 34348 91626 34352
rect 91562 34292 91566 34348
rect 91566 34292 91622 34348
rect 91622 34292 91626 34348
rect 91562 34288 91626 34292
rect 91642 34348 91706 34352
rect 91642 34292 91646 34348
rect 91646 34292 91702 34348
rect 91702 34292 91706 34348
rect 91642 34288 91706 34292
rect 91722 34348 91786 34352
rect 91722 34292 91726 34348
rect 91726 34292 91782 34348
rect 91782 34292 91786 34348
rect 91722 34288 91786 34292
rect 91802 34348 91866 34352
rect 91802 34292 91806 34348
rect 91806 34292 91862 34348
rect 91862 34292 91866 34348
rect 91802 34288 91866 34292
rect 3650 33804 3714 33808
rect 3650 33748 3654 33804
rect 3654 33748 3710 33804
rect 3710 33748 3714 33804
rect 3650 33744 3714 33748
rect 3730 33804 3794 33808
rect 3730 33748 3734 33804
rect 3734 33748 3790 33804
rect 3790 33748 3794 33804
rect 3730 33744 3794 33748
rect 3810 33804 3874 33808
rect 3810 33748 3814 33804
rect 3814 33748 3870 33804
rect 3870 33748 3874 33804
rect 3810 33744 3874 33748
rect 3890 33804 3954 33808
rect 3890 33748 3894 33804
rect 3894 33748 3950 33804
rect 3950 33748 3954 33804
rect 3890 33744 3954 33748
rect 8978 33804 9042 33808
rect 8978 33748 8982 33804
rect 8982 33748 9038 33804
rect 9038 33748 9042 33804
rect 8978 33744 9042 33748
rect 9058 33804 9122 33808
rect 9058 33748 9062 33804
rect 9062 33748 9118 33804
rect 9118 33748 9122 33804
rect 9058 33744 9122 33748
rect 9138 33804 9202 33808
rect 9138 33748 9142 33804
rect 9142 33748 9198 33804
rect 9198 33748 9202 33804
rect 9138 33744 9202 33748
rect 9218 33804 9282 33808
rect 9218 33748 9222 33804
rect 9222 33748 9278 33804
rect 9278 33748 9282 33804
rect 9218 33744 9282 33748
rect 14306 33804 14370 33808
rect 14306 33748 14310 33804
rect 14310 33748 14366 33804
rect 14366 33748 14370 33804
rect 14306 33744 14370 33748
rect 14386 33804 14450 33808
rect 14386 33748 14390 33804
rect 14390 33748 14446 33804
rect 14446 33748 14450 33804
rect 14386 33744 14450 33748
rect 14466 33804 14530 33808
rect 14466 33748 14470 33804
rect 14470 33748 14526 33804
rect 14526 33748 14530 33804
rect 14466 33744 14530 33748
rect 14546 33804 14610 33808
rect 14546 33748 14550 33804
rect 14550 33748 14606 33804
rect 14606 33748 14610 33804
rect 14546 33744 14610 33748
rect 19634 33804 19698 33808
rect 19634 33748 19638 33804
rect 19638 33748 19694 33804
rect 19694 33748 19698 33804
rect 19634 33744 19698 33748
rect 19714 33804 19778 33808
rect 19714 33748 19718 33804
rect 19718 33748 19774 33804
rect 19774 33748 19778 33804
rect 19714 33744 19778 33748
rect 19794 33804 19858 33808
rect 19794 33748 19798 33804
rect 19798 33748 19854 33804
rect 19854 33748 19858 33804
rect 19794 33744 19858 33748
rect 19874 33804 19938 33808
rect 19874 33748 19878 33804
rect 19878 33748 19934 33804
rect 19934 33748 19938 33804
rect 19874 33744 19938 33748
rect 24962 33804 25026 33808
rect 24962 33748 24966 33804
rect 24966 33748 25022 33804
rect 25022 33748 25026 33804
rect 24962 33744 25026 33748
rect 25042 33804 25106 33808
rect 25042 33748 25046 33804
rect 25046 33748 25102 33804
rect 25102 33748 25106 33804
rect 25042 33744 25106 33748
rect 25122 33804 25186 33808
rect 25122 33748 25126 33804
rect 25126 33748 25182 33804
rect 25182 33748 25186 33804
rect 25122 33744 25186 33748
rect 25202 33804 25266 33808
rect 25202 33748 25206 33804
rect 25206 33748 25262 33804
rect 25262 33748 25266 33804
rect 25202 33744 25266 33748
rect 30290 33804 30354 33808
rect 30290 33748 30294 33804
rect 30294 33748 30350 33804
rect 30350 33748 30354 33804
rect 30290 33744 30354 33748
rect 30370 33804 30434 33808
rect 30370 33748 30374 33804
rect 30374 33748 30430 33804
rect 30430 33748 30434 33804
rect 30370 33744 30434 33748
rect 30450 33804 30514 33808
rect 30450 33748 30454 33804
rect 30454 33748 30510 33804
rect 30510 33748 30514 33804
rect 30450 33744 30514 33748
rect 30530 33804 30594 33808
rect 30530 33748 30534 33804
rect 30534 33748 30590 33804
rect 30590 33748 30594 33804
rect 30530 33744 30594 33748
rect 35618 33804 35682 33808
rect 35618 33748 35622 33804
rect 35622 33748 35678 33804
rect 35678 33748 35682 33804
rect 35618 33744 35682 33748
rect 35698 33804 35762 33808
rect 35698 33748 35702 33804
rect 35702 33748 35758 33804
rect 35758 33748 35762 33804
rect 35698 33744 35762 33748
rect 35778 33804 35842 33808
rect 35778 33748 35782 33804
rect 35782 33748 35838 33804
rect 35838 33748 35842 33804
rect 35778 33744 35842 33748
rect 35858 33804 35922 33808
rect 35858 33748 35862 33804
rect 35862 33748 35918 33804
rect 35918 33748 35922 33804
rect 35858 33744 35922 33748
rect 40946 33804 41010 33808
rect 40946 33748 40950 33804
rect 40950 33748 41006 33804
rect 41006 33748 41010 33804
rect 40946 33744 41010 33748
rect 41026 33804 41090 33808
rect 41026 33748 41030 33804
rect 41030 33748 41086 33804
rect 41086 33748 41090 33804
rect 41026 33744 41090 33748
rect 41106 33804 41170 33808
rect 41106 33748 41110 33804
rect 41110 33748 41166 33804
rect 41166 33748 41170 33804
rect 41106 33744 41170 33748
rect 41186 33804 41250 33808
rect 41186 33748 41190 33804
rect 41190 33748 41246 33804
rect 41246 33748 41250 33804
rect 41186 33744 41250 33748
rect 46274 33804 46338 33808
rect 46274 33748 46278 33804
rect 46278 33748 46334 33804
rect 46334 33748 46338 33804
rect 46274 33744 46338 33748
rect 46354 33804 46418 33808
rect 46354 33748 46358 33804
rect 46358 33748 46414 33804
rect 46414 33748 46418 33804
rect 46354 33744 46418 33748
rect 46434 33804 46498 33808
rect 46434 33748 46438 33804
rect 46438 33748 46494 33804
rect 46494 33748 46498 33804
rect 46434 33744 46498 33748
rect 46514 33804 46578 33808
rect 46514 33748 46518 33804
rect 46518 33748 46574 33804
rect 46574 33748 46578 33804
rect 46514 33744 46578 33748
rect 51602 33804 51666 33808
rect 51602 33748 51606 33804
rect 51606 33748 51662 33804
rect 51662 33748 51666 33804
rect 51602 33744 51666 33748
rect 51682 33804 51746 33808
rect 51682 33748 51686 33804
rect 51686 33748 51742 33804
rect 51742 33748 51746 33804
rect 51682 33744 51746 33748
rect 51762 33804 51826 33808
rect 51762 33748 51766 33804
rect 51766 33748 51822 33804
rect 51822 33748 51826 33804
rect 51762 33744 51826 33748
rect 51842 33804 51906 33808
rect 51842 33748 51846 33804
rect 51846 33748 51902 33804
rect 51902 33748 51906 33804
rect 51842 33744 51906 33748
rect 56930 33804 56994 33808
rect 56930 33748 56934 33804
rect 56934 33748 56990 33804
rect 56990 33748 56994 33804
rect 56930 33744 56994 33748
rect 57010 33804 57074 33808
rect 57010 33748 57014 33804
rect 57014 33748 57070 33804
rect 57070 33748 57074 33804
rect 57010 33744 57074 33748
rect 57090 33804 57154 33808
rect 57090 33748 57094 33804
rect 57094 33748 57150 33804
rect 57150 33748 57154 33804
rect 57090 33744 57154 33748
rect 57170 33804 57234 33808
rect 57170 33748 57174 33804
rect 57174 33748 57230 33804
rect 57230 33748 57234 33804
rect 57170 33744 57234 33748
rect 62258 33804 62322 33808
rect 62258 33748 62262 33804
rect 62262 33748 62318 33804
rect 62318 33748 62322 33804
rect 62258 33744 62322 33748
rect 62338 33804 62402 33808
rect 62338 33748 62342 33804
rect 62342 33748 62398 33804
rect 62398 33748 62402 33804
rect 62338 33744 62402 33748
rect 62418 33804 62482 33808
rect 62418 33748 62422 33804
rect 62422 33748 62478 33804
rect 62478 33748 62482 33804
rect 62418 33744 62482 33748
rect 62498 33804 62562 33808
rect 62498 33748 62502 33804
rect 62502 33748 62558 33804
rect 62558 33748 62562 33804
rect 62498 33744 62562 33748
rect 67586 33804 67650 33808
rect 67586 33748 67590 33804
rect 67590 33748 67646 33804
rect 67646 33748 67650 33804
rect 67586 33744 67650 33748
rect 67666 33804 67730 33808
rect 67666 33748 67670 33804
rect 67670 33748 67726 33804
rect 67726 33748 67730 33804
rect 67666 33744 67730 33748
rect 67746 33804 67810 33808
rect 67746 33748 67750 33804
rect 67750 33748 67806 33804
rect 67806 33748 67810 33804
rect 67746 33744 67810 33748
rect 67826 33804 67890 33808
rect 67826 33748 67830 33804
rect 67830 33748 67886 33804
rect 67886 33748 67890 33804
rect 67826 33744 67890 33748
rect 72914 33804 72978 33808
rect 72914 33748 72918 33804
rect 72918 33748 72974 33804
rect 72974 33748 72978 33804
rect 72914 33744 72978 33748
rect 72994 33804 73058 33808
rect 72994 33748 72998 33804
rect 72998 33748 73054 33804
rect 73054 33748 73058 33804
rect 72994 33744 73058 33748
rect 73074 33804 73138 33808
rect 73074 33748 73078 33804
rect 73078 33748 73134 33804
rect 73134 33748 73138 33804
rect 73074 33744 73138 33748
rect 73154 33804 73218 33808
rect 73154 33748 73158 33804
rect 73158 33748 73214 33804
rect 73214 33748 73218 33804
rect 73154 33744 73218 33748
rect 78242 33804 78306 33808
rect 78242 33748 78246 33804
rect 78246 33748 78302 33804
rect 78302 33748 78306 33804
rect 78242 33744 78306 33748
rect 78322 33804 78386 33808
rect 78322 33748 78326 33804
rect 78326 33748 78382 33804
rect 78382 33748 78386 33804
rect 78322 33744 78386 33748
rect 78402 33804 78466 33808
rect 78402 33748 78406 33804
rect 78406 33748 78462 33804
rect 78462 33748 78466 33804
rect 78402 33744 78466 33748
rect 78482 33804 78546 33808
rect 78482 33748 78486 33804
rect 78486 33748 78542 33804
rect 78542 33748 78546 33804
rect 78482 33744 78546 33748
rect 83570 33804 83634 33808
rect 83570 33748 83574 33804
rect 83574 33748 83630 33804
rect 83630 33748 83634 33804
rect 83570 33744 83634 33748
rect 83650 33804 83714 33808
rect 83650 33748 83654 33804
rect 83654 33748 83710 33804
rect 83710 33748 83714 33804
rect 83650 33744 83714 33748
rect 83730 33804 83794 33808
rect 83730 33748 83734 33804
rect 83734 33748 83790 33804
rect 83790 33748 83794 33804
rect 83730 33744 83794 33748
rect 83810 33804 83874 33808
rect 83810 33748 83814 33804
rect 83814 33748 83870 33804
rect 83870 33748 83874 33804
rect 83810 33744 83874 33748
rect 88898 33804 88962 33808
rect 88898 33748 88902 33804
rect 88902 33748 88958 33804
rect 88958 33748 88962 33804
rect 88898 33744 88962 33748
rect 88978 33804 89042 33808
rect 88978 33748 88982 33804
rect 88982 33748 89038 33804
rect 89038 33748 89042 33804
rect 88978 33744 89042 33748
rect 89058 33804 89122 33808
rect 89058 33748 89062 33804
rect 89062 33748 89118 33804
rect 89118 33748 89122 33804
rect 89058 33744 89122 33748
rect 89138 33804 89202 33808
rect 89138 33748 89142 33804
rect 89142 33748 89198 33804
rect 89198 33748 89202 33804
rect 89138 33744 89202 33748
rect 6314 33260 6378 33264
rect 6314 33204 6318 33260
rect 6318 33204 6374 33260
rect 6374 33204 6378 33260
rect 6314 33200 6378 33204
rect 6394 33260 6458 33264
rect 6394 33204 6398 33260
rect 6398 33204 6454 33260
rect 6454 33204 6458 33260
rect 6394 33200 6458 33204
rect 6474 33260 6538 33264
rect 6474 33204 6478 33260
rect 6478 33204 6534 33260
rect 6534 33204 6538 33260
rect 6474 33200 6538 33204
rect 6554 33260 6618 33264
rect 6554 33204 6558 33260
rect 6558 33204 6614 33260
rect 6614 33204 6618 33260
rect 6554 33200 6618 33204
rect 11642 33260 11706 33264
rect 11642 33204 11646 33260
rect 11646 33204 11702 33260
rect 11702 33204 11706 33260
rect 11642 33200 11706 33204
rect 11722 33260 11786 33264
rect 11722 33204 11726 33260
rect 11726 33204 11782 33260
rect 11782 33204 11786 33260
rect 11722 33200 11786 33204
rect 11802 33260 11866 33264
rect 11802 33204 11806 33260
rect 11806 33204 11862 33260
rect 11862 33204 11866 33260
rect 11802 33200 11866 33204
rect 11882 33260 11946 33264
rect 11882 33204 11886 33260
rect 11886 33204 11942 33260
rect 11942 33204 11946 33260
rect 11882 33200 11946 33204
rect 16970 33260 17034 33264
rect 16970 33204 16974 33260
rect 16974 33204 17030 33260
rect 17030 33204 17034 33260
rect 16970 33200 17034 33204
rect 17050 33260 17114 33264
rect 17050 33204 17054 33260
rect 17054 33204 17110 33260
rect 17110 33204 17114 33260
rect 17050 33200 17114 33204
rect 17130 33260 17194 33264
rect 17130 33204 17134 33260
rect 17134 33204 17190 33260
rect 17190 33204 17194 33260
rect 17130 33200 17194 33204
rect 17210 33260 17274 33264
rect 17210 33204 17214 33260
rect 17214 33204 17270 33260
rect 17270 33204 17274 33260
rect 17210 33200 17274 33204
rect 22298 33260 22362 33264
rect 22298 33204 22302 33260
rect 22302 33204 22358 33260
rect 22358 33204 22362 33260
rect 22298 33200 22362 33204
rect 22378 33260 22442 33264
rect 22378 33204 22382 33260
rect 22382 33204 22438 33260
rect 22438 33204 22442 33260
rect 22378 33200 22442 33204
rect 22458 33260 22522 33264
rect 22458 33204 22462 33260
rect 22462 33204 22518 33260
rect 22518 33204 22522 33260
rect 22458 33200 22522 33204
rect 22538 33260 22602 33264
rect 22538 33204 22542 33260
rect 22542 33204 22598 33260
rect 22598 33204 22602 33260
rect 22538 33200 22602 33204
rect 27626 33260 27690 33264
rect 27626 33204 27630 33260
rect 27630 33204 27686 33260
rect 27686 33204 27690 33260
rect 27626 33200 27690 33204
rect 27706 33260 27770 33264
rect 27706 33204 27710 33260
rect 27710 33204 27766 33260
rect 27766 33204 27770 33260
rect 27706 33200 27770 33204
rect 27786 33260 27850 33264
rect 27786 33204 27790 33260
rect 27790 33204 27846 33260
rect 27846 33204 27850 33260
rect 27786 33200 27850 33204
rect 27866 33260 27930 33264
rect 27866 33204 27870 33260
rect 27870 33204 27926 33260
rect 27926 33204 27930 33260
rect 27866 33200 27930 33204
rect 32954 33260 33018 33264
rect 32954 33204 32958 33260
rect 32958 33204 33014 33260
rect 33014 33204 33018 33260
rect 32954 33200 33018 33204
rect 33034 33260 33098 33264
rect 33034 33204 33038 33260
rect 33038 33204 33094 33260
rect 33094 33204 33098 33260
rect 33034 33200 33098 33204
rect 33114 33260 33178 33264
rect 33114 33204 33118 33260
rect 33118 33204 33174 33260
rect 33174 33204 33178 33260
rect 33114 33200 33178 33204
rect 33194 33260 33258 33264
rect 33194 33204 33198 33260
rect 33198 33204 33254 33260
rect 33254 33204 33258 33260
rect 33194 33200 33258 33204
rect 38282 33260 38346 33264
rect 38282 33204 38286 33260
rect 38286 33204 38342 33260
rect 38342 33204 38346 33260
rect 38282 33200 38346 33204
rect 38362 33260 38426 33264
rect 38362 33204 38366 33260
rect 38366 33204 38422 33260
rect 38422 33204 38426 33260
rect 38362 33200 38426 33204
rect 38442 33260 38506 33264
rect 38442 33204 38446 33260
rect 38446 33204 38502 33260
rect 38502 33204 38506 33260
rect 38442 33200 38506 33204
rect 38522 33260 38586 33264
rect 38522 33204 38526 33260
rect 38526 33204 38582 33260
rect 38582 33204 38586 33260
rect 38522 33200 38586 33204
rect 43610 33260 43674 33264
rect 43610 33204 43614 33260
rect 43614 33204 43670 33260
rect 43670 33204 43674 33260
rect 43610 33200 43674 33204
rect 43690 33260 43754 33264
rect 43690 33204 43694 33260
rect 43694 33204 43750 33260
rect 43750 33204 43754 33260
rect 43690 33200 43754 33204
rect 43770 33260 43834 33264
rect 43770 33204 43774 33260
rect 43774 33204 43830 33260
rect 43830 33204 43834 33260
rect 43770 33200 43834 33204
rect 43850 33260 43914 33264
rect 43850 33204 43854 33260
rect 43854 33204 43910 33260
rect 43910 33204 43914 33260
rect 43850 33200 43914 33204
rect 48938 33260 49002 33264
rect 48938 33204 48942 33260
rect 48942 33204 48998 33260
rect 48998 33204 49002 33260
rect 48938 33200 49002 33204
rect 49018 33260 49082 33264
rect 49018 33204 49022 33260
rect 49022 33204 49078 33260
rect 49078 33204 49082 33260
rect 49018 33200 49082 33204
rect 49098 33260 49162 33264
rect 49098 33204 49102 33260
rect 49102 33204 49158 33260
rect 49158 33204 49162 33260
rect 49098 33200 49162 33204
rect 49178 33260 49242 33264
rect 49178 33204 49182 33260
rect 49182 33204 49238 33260
rect 49238 33204 49242 33260
rect 49178 33200 49242 33204
rect 54266 33260 54330 33264
rect 54266 33204 54270 33260
rect 54270 33204 54326 33260
rect 54326 33204 54330 33260
rect 54266 33200 54330 33204
rect 54346 33260 54410 33264
rect 54346 33204 54350 33260
rect 54350 33204 54406 33260
rect 54406 33204 54410 33260
rect 54346 33200 54410 33204
rect 54426 33260 54490 33264
rect 54426 33204 54430 33260
rect 54430 33204 54486 33260
rect 54486 33204 54490 33260
rect 54426 33200 54490 33204
rect 54506 33260 54570 33264
rect 54506 33204 54510 33260
rect 54510 33204 54566 33260
rect 54566 33204 54570 33260
rect 54506 33200 54570 33204
rect 59594 33260 59658 33264
rect 59594 33204 59598 33260
rect 59598 33204 59654 33260
rect 59654 33204 59658 33260
rect 59594 33200 59658 33204
rect 59674 33260 59738 33264
rect 59674 33204 59678 33260
rect 59678 33204 59734 33260
rect 59734 33204 59738 33260
rect 59674 33200 59738 33204
rect 59754 33260 59818 33264
rect 59754 33204 59758 33260
rect 59758 33204 59814 33260
rect 59814 33204 59818 33260
rect 59754 33200 59818 33204
rect 59834 33260 59898 33264
rect 59834 33204 59838 33260
rect 59838 33204 59894 33260
rect 59894 33204 59898 33260
rect 59834 33200 59898 33204
rect 64922 33260 64986 33264
rect 64922 33204 64926 33260
rect 64926 33204 64982 33260
rect 64982 33204 64986 33260
rect 64922 33200 64986 33204
rect 65002 33260 65066 33264
rect 65002 33204 65006 33260
rect 65006 33204 65062 33260
rect 65062 33204 65066 33260
rect 65002 33200 65066 33204
rect 65082 33260 65146 33264
rect 65082 33204 65086 33260
rect 65086 33204 65142 33260
rect 65142 33204 65146 33260
rect 65082 33200 65146 33204
rect 65162 33260 65226 33264
rect 65162 33204 65166 33260
rect 65166 33204 65222 33260
rect 65222 33204 65226 33260
rect 65162 33200 65226 33204
rect 70250 33260 70314 33264
rect 70250 33204 70254 33260
rect 70254 33204 70310 33260
rect 70310 33204 70314 33260
rect 70250 33200 70314 33204
rect 70330 33260 70394 33264
rect 70330 33204 70334 33260
rect 70334 33204 70390 33260
rect 70390 33204 70394 33260
rect 70330 33200 70394 33204
rect 70410 33260 70474 33264
rect 70410 33204 70414 33260
rect 70414 33204 70470 33260
rect 70470 33204 70474 33260
rect 70410 33200 70474 33204
rect 70490 33260 70554 33264
rect 70490 33204 70494 33260
rect 70494 33204 70550 33260
rect 70550 33204 70554 33260
rect 70490 33200 70554 33204
rect 75578 33260 75642 33264
rect 75578 33204 75582 33260
rect 75582 33204 75638 33260
rect 75638 33204 75642 33260
rect 75578 33200 75642 33204
rect 75658 33260 75722 33264
rect 75658 33204 75662 33260
rect 75662 33204 75718 33260
rect 75718 33204 75722 33260
rect 75658 33200 75722 33204
rect 75738 33260 75802 33264
rect 75738 33204 75742 33260
rect 75742 33204 75798 33260
rect 75798 33204 75802 33260
rect 75738 33200 75802 33204
rect 75818 33260 75882 33264
rect 75818 33204 75822 33260
rect 75822 33204 75878 33260
rect 75878 33204 75882 33260
rect 75818 33200 75882 33204
rect 80906 33260 80970 33264
rect 80906 33204 80910 33260
rect 80910 33204 80966 33260
rect 80966 33204 80970 33260
rect 80906 33200 80970 33204
rect 80986 33260 81050 33264
rect 80986 33204 80990 33260
rect 80990 33204 81046 33260
rect 81046 33204 81050 33260
rect 80986 33200 81050 33204
rect 81066 33260 81130 33264
rect 81066 33204 81070 33260
rect 81070 33204 81126 33260
rect 81126 33204 81130 33260
rect 81066 33200 81130 33204
rect 81146 33260 81210 33264
rect 81146 33204 81150 33260
rect 81150 33204 81206 33260
rect 81206 33204 81210 33260
rect 81146 33200 81210 33204
rect 86234 33260 86298 33264
rect 86234 33204 86238 33260
rect 86238 33204 86294 33260
rect 86294 33204 86298 33260
rect 86234 33200 86298 33204
rect 86314 33260 86378 33264
rect 86314 33204 86318 33260
rect 86318 33204 86374 33260
rect 86374 33204 86378 33260
rect 86314 33200 86378 33204
rect 86394 33260 86458 33264
rect 86394 33204 86398 33260
rect 86398 33204 86454 33260
rect 86454 33204 86458 33260
rect 86394 33200 86458 33204
rect 86474 33260 86538 33264
rect 86474 33204 86478 33260
rect 86478 33204 86534 33260
rect 86534 33204 86538 33260
rect 86474 33200 86538 33204
rect 91562 33260 91626 33264
rect 91562 33204 91566 33260
rect 91566 33204 91622 33260
rect 91622 33204 91626 33260
rect 91562 33200 91626 33204
rect 91642 33260 91706 33264
rect 91642 33204 91646 33260
rect 91646 33204 91702 33260
rect 91702 33204 91706 33260
rect 91642 33200 91706 33204
rect 91722 33260 91786 33264
rect 91722 33204 91726 33260
rect 91726 33204 91782 33260
rect 91782 33204 91786 33260
rect 91722 33200 91786 33204
rect 91802 33260 91866 33264
rect 91802 33204 91806 33260
rect 91806 33204 91862 33260
rect 91862 33204 91866 33260
rect 91802 33200 91866 33204
rect 3650 32716 3714 32720
rect 3650 32660 3654 32716
rect 3654 32660 3710 32716
rect 3710 32660 3714 32716
rect 3650 32656 3714 32660
rect 3730 32716 3794 32720
rect 3730 32660 3734 32716
rect 3734 32660 3790 32716
rect 3790 32660 3794 32716
rect 3730 32656 3794 32660
rect 3810 32716 3874 32720
rect 3810 32660 3814 32716
rect 3814 32660 3870 32716
rect 3870 32660 3874 32716
rect 3810 32656 3874 32660
rect 3890 32716 3954 32720
rect 3890 32660 3894 32716
rect 3894 32660 3950 32716
rect 3950 32660 3954 32716
rect 3890 32656 3954 32660
rect 8978 32716 9042 32720
rect 8978 32660 8982 32716
rect 8982 32660 9038 32716
rect 9038 32660 9042 32716
rect 8978 32656 9042 32660
rect 9058 32716 9122 32720
rect 9058 32660 9062 32716
rect 9062 32660 9118 32716
rect 9118 32660 9122 32716
rect 9058 32656 9122 32660
rect 9138 32716 9202 32720
rect 9138 32660 9142 32716
rect 9142 32660 9198 32716
rect 9198 32660 9202 32716
rect 9138 32656 9202 32660
rect 9218 32716 9282 32720
rect 9218 32660 9222 32716
rect 9222 32660 9278 32716
rect 9278 32660 9282 32716
rect 9218 32656 9282 32660
rect 14306 32716 14370 32720
rect 14306 32660 14310 32716
rect 14310 32660 14366 32716
rect 14366 32660 14370 32716
rect 14306 32656 14370 32660
rect 14386 32716 14450 32720
rect 14386 32660 14390 32716
rect 14390 32660 14446 32716
rect 14446 32660 14450 32716
rect 14386 32656 14450 32660
rect 14466 32716 14530 32720
rect 14466 32660 14470 32716
rect 14470 32660 14526 32716
rect 14526 32660 14530 32716
rect 14466 32656 14530 32660
rect 14546 32716 14610 32720
rect 14546 32660 14550 32716
rect 14550 32660 14606 32716
rect 14606 32660 14610 32716
rect 14546 32656 14610 32660
rect 19634 32716 19698 32720
rect 19634 32660 19638 32716
rect 19638 32660 19694 32716
rect 19694 32660 19698 32716
rect 19634 32656 19698 32660
rect 19714 32716 19778 32720
rect 19714 32660 19718 32716
rect 19718 32660 19774 32716
rect 19774 32660 19778 32716
rect 19714 32656 19778 32660
rect 19794 32716 19858 32720
rect 19794 32660 19798 32716
rect 19798 32660 19854 32716
rect 19854 32660 19858 32716
rect 19794 32656 19858 32660
rect 19874 32716 19938 32720
rect 19874 32660 19878 32716
rect 19878 32660 19934 32716
rect 19934 32660 19938 32716
rect 19874 32656 19938 32660
rect 24962 32716 25026 32720
rect 24962 32660 24966 32716
rect 24966 32660 25022 32716
rect 25022 32660 25026 32716
rect 24962 32656 25026 32660
rect 25042 32716 25106 32720
rect 25042 32660 25046 32716
rect 25046 32660 25102 32716
rect 25102 32660 25106 32716
rect 25042 32656 25106 32660
rect 25122 32716 25186 32720
rect 25122 32660 25126 32716
rect 25126 32660 25182 32716
rect 25182 32660 25186 32716
rect 25122 32656 25186 32660
rect 25202 32716 25266 32720
rect 25202 32660 25206 32716
rect 25206 32660 25262 32716
rect 25262 32660 25266 32716
rect 25202 32656 25266 32660
rect 30290 32716 30354 32720
rect 30290 32660 30294 32716
rect 30294 32660 30350 32716
rect 30350 32660 30354 32716
rect 30290 32656 30354 32660
rect 30370 32716 30434 32720
rect 30370 32660 30374 32716
rect 30374 32660 30430 32716
rect 30430 32660 30434 32716
rect 30370 32656 30434 32660
rect 30450 32716 30514 32720
rect 30450 32660 30454 32716
rect 30454 32660 30510 32716
rect 30510 32660 30514 32716
rect 30450 32656 30514 32660
rect 30530 32716 30594 32720
rect 30530 32660 30534 32716
rect 30534 32660 30590 32716
rect 30590 32660 30594 32716
rect 30530 32656 30594 32660
rect 35618 32716 35682 32720
rect 35618 32660 35622 32716
rect 35622 32660 35678 32716
rect 35678 32660 35682 32716
rect 35618 32656 35682 32660
rect 35698 32716 35762 32720
rect 35698 32660 35702 32716
rect 35702 32660 35758 32716
rect 35758 32660 35762 32716
rect 35698 32656 35762 32660
rect 35778 32716 35842 32720
rect 35778 32660 35782 32716
rect 35782 32660 35838 32716
rect 35838 32660 35842 32716
rect 35778 32656 35842 32660
rect 35858 32716 35922 32720
rect 35858 32660 35862 32716
rect 35862 32660 35918 32716
rect 35918 32660 35922 32716
rect 35858 32656 35922 32660
rect 40946 32716 41010 32720
rect 40946 32660 40950 32716
rect 40950 32660 41006 32716
rect 41006 32660 41010 32716
rect 40946 32656 41010 32660
rect 41026 32716 41090 32720
rect 41026 32660 41030 32716
rect 41030 32660 41086 32716
rect 41086 32660 41090 32716
rect 41026 32656 41090 32660
rect 41106 32716 41170 32720
rect 41106 32660 41110 32716
rect 41110 32660 41166 32716
rect 41166 32660 41170 32716
rect 41106 32656 41170 32660
rect 41186 32716 41250 32720
rect 41186 32660 41190 32716
rect 41190 32660 41246 32716
rect 41246 32660 41250 32716
rect 41186 32656 41250 32660
rect 46274 32716 46338 32720
rect 46274 32660 46278 32716
rect 46278 32660 46334 32716
rect 46334 32660 46338 32716
rect 46274 32656 46338 32660
rect 46354 32716 46418 32720
rect 46354 32660 46358 32716
rect 46358 32660 46414 32716
rect 46414 32660 46418 32716
rect 46354 32656 46418 32660
rect 46434 32716 46498 32720
rect 46434 32660 46438 32716
rect 46438 32660 46494 32716
rect 46494 32660 46498 32716
rect 46434 32656 46498 32660
rect 46514 32716 46578 32720
rect 46514 32660 46518 32716
rect 46518 32660 46574 32716
rect 46574 32660 46578 32716
rect 46514 32656 46578 32660
rect 51602 32716 51666 32720
rect 51602 32660 51606 32716
rect 51606 32660 51662 32716
rect 51662 32660 51666 32716
rect 51602 32656 51666 32660
rect 51682 32716 51746 32720
rect 51682 32660 51686 32716
rect 51686 32660 51742 32716
rect 51742 32660 51746 32716
rect 51682 32656 51746 32660
rect 51762 32716 51826 32720
rect 51762 32660 51766 32716
rect 51766 32660 51822 32716
rect 51822 32660 51826 32716
rect 51762 32656 51826 32660
rect 51842 32716 51906 32720
rect 51842 32660 51846 32716
rect 51846 32660 51902 32716
rect 51902 32660 51906 32716
rect 51842 32656 51906 32660
rect 56930 32716 56994 32720
rect 56930 32660 56934 32716
rect 56934 32660 56990 32716
rect 56990 32660 56994 32716
rect 56930 32656 56994 32660
rect 57010 32716 57074 32720
rect 57010 32660 57014 32716
rect 57014 32660 57070 32716
rect 57070 32660 57074 32716
rect 57010 32656 57074 32660
rect 57090 32716 57154 32720
rect 57090 32660 57094 32716
rect 57094 32660 57150 32716
rect 57150 32660 57154 32716
rect 57090 32656 57154 32660
rect 57170 32716 57234 32720
rect 57170 32660 57174 32716
rect 57174 32660 57230 32716
rect 57230 32660 57234 32716
rect 57170 32656 57234 32660
rect 62258 32716 62322 32720
rect 62258 32660 62262 32716
rect 62262 32660 62318 32716
rect 62318 32660 62322 32716
rect 62258 32656 62322 32660
rect 62338 32716 62402 32720
rect 62338 32660 62342 32716
rect 62342 32660 62398 32716
rect 62398 32660 62402 32716
rect 62338 32656 62402 32660
rect 62418 32716 62482 32720
rect 62418 32660 62422 32716
rect 62422 32660 62478 32716
rect 62478 32660 62482 32716
rect 62418 32656 62482 32660
rect 62498 32716 62562 32720
rect 62498 32660 62502 32716
rect 62502 32660 62558 32716
rect 62558 32660 62562 32716
rect 62498 32656 62562 32660
rect 67586 32716 67650 32720
rect 67586 32660 67590 32716
rect 67590 32660 67646 32716
rect 67646 32660 67650 32716
rect 67586 32656 67650 32660
rect 67666 32716 67730 32720
rect 67666 32660 67670 32716
rect 67670 32660 67726 32716
rect 67726 32660 67730 32716
rect 67666 32656 67730 32660
rect 67746 32716 67810 32720
rect 67746 32660 67750 32716
rect 67750 32660 67806 32716
rect 67806 32660 67810 32716
rect 67746 32656 67810 32660
rect 67826 32716 67890 32720
rect 67826 32660 67830 32716
rect 67830 32660 67886 32716
rect 67886 32660 67890 32716
rect 67826 32656 67890 32660
rect 72914 32716 72978 32720
rect 72914 32660 72918 32716
rect 72918 32660 72974 32716
rect 72974 32660 72978 32716
rect 72914 32656 72978 32660
rect 72994 32716 73058 32720
rect 72994 32660 72998 32716
rect 72998 32660 73054 32716
rect 73054 32660 73058 32716
rect 72994 32656 73058 32660
rect 73074 32716 73138 32720
rect 73074 32660 73078 32716
rect 73078 32660 73134 32716
rect 73134 32660 73138 32716
rect 73074 32656 73138 32660
rect 73154 32716 73218 32720
rect 73154 32660 73158 32716
rect 73158 32660 73214 32716
rect 73214 32660 73218 32716
rect 73154 32656 73218 32660
rect 78242 32716 78306 32720
rect 78242 32660 78246 32716
rect 78246 32660 78302 32716
rect 78302 32660 78306 32716
rect 78242 32656 78306 32660
rect 78322 32716 78386 32720
rect 78322 32660 78326 32716
rect 78326 32660 78382 32716
rect 78382 32660 78386 32716
rect 78322 32656 78386 32660
rect 78402 32716 78466 32720
rect 78402 32660 78406 32716
rect 78406 32660 78462 32716
rect 78462 32660 78466 32716
rect 78402 32656 78466 32660
rect 78482 32716 78546 32720
rect 78482 32660 78486 32716
rect 78486 32660 78542 32716
rect 78542 32660 78546 32716
rect 78482 32656 78546 32660
rect 83570 32716 83634 32720
rect 83570 32660 83574 32716
rect 83574 32660 83630 32716
rect 83630 32660 83634 32716
rect 83570 32656 83634 32660
rect 83650 32716 83714 32720
rect 83650 32660 83654 32716
rect 83654 32660 83710 32716
rect 83710 32660 83714 32716
rect 83650 32656 83714 32660
rect 83730 32716 83794 32720
rect 83730 32660 83734 32716
rect 83734 32660 83790 32716
rect 83790 32660 83794 32716
rect 83730 32656 83794 32660
rect 83810 32716 83874 32720
rect 83810 32660 83814 32716
rect 83814 32660 83870 32716
rect 83870 32660 83874 32716
rect 83810 32656 83874 32660
rect 88898 32716 88962 32720
rect 88898 32660 88902 32716
rect 88902 32660 88958 32716
rect 88958 32660 88962 32716
rect 88898 32656 88962 32660
rect 88978 32716 89042 32720
rect 88978 32660 88982 32716
rect 88982 32660 89038 32716
rect 89038 32660 89042 32716
rect 88978 32656 89042 32660
rect 89058 32716 89122 32720
rect 89058 32660 89062 32716
rect 89062 32660 89118 32716
rect 89118 32660 89122 32716
rect 89058 32656 89122 32660
rect 89138 32716 89202 32720
rect 89138 32660 89142 32716
rect 89142 32660 89198 32716
rect 89198 32660 89202 32716
rect 89138 32656 89202 32660
rect 6314 32172 6378 32176
rect 6314 32116 6318 32172
rect 6318 32116 6374 32172
rect 6374 32116 6378 32172
rect 6314 32112 6378 32116
rect 6394 32172 6458 32176
rect 6394 32116 6398 32172
rect 6398 32116 6454 32172
rect 6454 32116 6458 32172
rect 6394 32112 6458 32116
rect 6474 32172 6538 32176
rect 6474 32116 6478 32172
rect 6478 32116 6534 32172
rect 6534 32116 6538 32172
rect 6474 32112 6538 32116
rect 6554 32172 6618 32176
rect 6554 32116 6558 32172
rect 6558 32116 6614 32172
rect 6614 32116 6618 32172
rect 6554 32112 6618 32116
rect 11642 32172 11706 32176
rect 11642 32116 11646 32172
rect 11646 32116 11702 32172
rect 11702 32116 11706 32172
rect 11642 32112 11706 32116
rect 11722 32172 11786 32176
rect 11722 32116 11726 32172
rect 11726 32116 11782 32172
rect 11782 32116 11786 32172
rect 11722 32112 11786 32116
rect 11802 32172 11866 32176
rect 11802 32116 11806 32172
rect 11806 32116 11862 32172
rect 11862 32116 11866 32172
rect 11802 32112 11866 32116
rect 11882 32172 11946 32176
rect 11882 32116 11886 32172
rect 11886 32116 11942 32172
rect 11942 32116 11946 32172
rect 11882 32112 11946 32116
rect 16970 32172 17034 32176
rect 16970 32116 16974 32172
rect 16974 32116 17030 32172
rect 17030 32116 17034 32172
rect 16970 32112 17034 32116
rect 17050 32172 17114 32176
rect 17050 32116 17054 32172
rect 17054 32116 17110 32172
rect 17110 32116 17114 32172
rect 17050 32112 17114 32116
rect 17130 32172 17194 32176
rect 17130 32116 17134 32172
rect 17134 32116 17190 32172
rect 17190 32116 17194 32172
rect 17130 32112 17194 32116
rect 17210 32172 17274 32176
rect 17210 32116 17214 32172
rect 17214 32116 17270 32172
rect 17270 32116 17274 32172
rect 17210 32112 17274 32116
rect 22298 32172 22362 32176
rect 22298 32116 22302 32172
rect 22302 32116 22358 32172
rect 22358 32116 22362 32172
rect 22298 32112 22362 32116
rect 22378 32172 22442 32176
rect 22378 32116 22382 32172
rect 22382 32116 22438 32172
rect 22438 32116 22442 32172
rect 22378 32112 22442 32116
rect 22458 32172 22522 32176
rect 22458 32116 22462 32172
rect 22462 32116 22518 32172
rect 22518 32116 22522 32172
rect 22458 32112 22522 32116
rect 22538 32172 22602 32176
rect 22538 32116 22542 32172
rect 22542 32116 22598 32172
rect 22598 32116 22602 32172
rect 22538 32112 22602 32116
rect 27626 32172 27690 32176
rect 27626 32116 27630 32172
rect 27630 32116 27686 32172
rect 27686 32116 27690 32172
rect 27626 32112 27690 32116
rect 27706 32172 27770 32176
rect 27706 32116 27710 32172
rect 27710 32116 27766 32172
rect 27766 32116 27770 32172
rect 27706 32112 27770 32116
rect 27786 32172 27850 32176
rect 27786 32116 27790 32172
rect 27790 32116 27846 32172
rect 27846 32116 27850 32172
rect 27786 32112 27850 32116
rect 27866 32172 27930 32176
rect 27866 32116 27870 32172
rect 27870 32116 27926 32172
rect 27926 32116 27930 32172
rect 27866 32112 27930 32116
rect 32954 32172 33018 32176
rect 32954 32116 32958 32172
rect 32958 32116 33014 32172
rect 33014 32116 33018 32172
rect 32954 32112 33018 32116
rect 33034 32172 33098 32176
rect 33034 32116 33038 32172
rect 33038 32116 33094 32172
rect 33094 32116 33098 32172
rect 33034 32112 33098 32116
rect 33114 32172 33178 32176
rect 33114 32116 33118 32172
rect 33118 32116 33174 32172
rect 33174 32116 33178 32172
rect 33114 32112 33178 32116
rect 33194 32172 33258 32176
rect 33194 32116 33198 32172
rect 33198 32116 33254 32172
rect 33254 32116 33258 32172
rect 33194 32112 33258 32116
rect 38282 32172 38346 32176
rect 38282 32116 38286 32172
rect 38286 32116 38342 32172
rect 38342 32116 38346 32172
rect 38282 32112 38346 32116
rect 38362 32172 38426 32176
rect 38362 32116 38366 32172
rect 38366 32116 38422 32172
rect 38422 32116 38426 32172
rect 38362 32112 38426 32116
rect 38442 32172 38506 32176
rect 38442 32116 38446 32172
rect 38446 32116 38502 32172
rect 38502 32116 38506 32172
rect 38442 32112 38506 32116
rect 38522 32172 38586 32176
rect 38522 32116 38526 32172
rect 38526 32116 38582 32172
rect 38582 32116 38586 32172
rect 38522 32112 38586 32116
rect 43610 32172 43674 32176
rect 43610 32116 43614 32172
rect 43614 32116 43670 32172
rect 43670 32116 43674 32172
rect 43610 32112 43674 32116
rect 43690 32172 43754 32176
rect 43690 32116 43694 32172
rect 43694 32116 43750 32172
rect 43750 32116 43754 32172
rect 43690 32112 43754 32116
rect 43770 32172 43834 32176
rect 43770 32116 43774 32172
rect 43774 32116 43830 32172
rect 43830 32116 43834 32172
rect 43770 32112 43834 32116
rect 43850 32172 43914 32176
rect 43850 32116 43854 32172
rect 43854 32116 43910 32172
rect 43910 32116 43914 32172
rect 43850 32112 43914 32116
rect 48938 32172 49002 32176
rect 48938 32116 48942 32172
rect 48942 32116 48998 32172
rect 48998 32116 49002 32172
rect 48938 32112 49002 32116
rect 49018 32172 49082 32176
rect 49018 32116 49022 32172
rect 49022 32116 49078 32172
rect 49078 32116 49082 32172
rect 49018 32112 49082 32116
rect 49098 32172 49162 32176
rect 49098 32116 49102 32172
rect 49102 32116 49158 32172
rect 49158 32116 49162 32172
rect 49098 32112 49162 32116
rect 49178 32172 49242 32176
rect 49178 32116 49182 32172
rect 49182 32116 49238 32172
rect 49238 32116 49242 32172
rect 49178 32112 49242 32116
rect 54266 32172 54330 32176
rect 54266 32116 54270 32172
rect 54270 32116 54326 32172
rect 54326 32116 54330 32172
rect 54266 32112 54330 32116
rect 54346 32172 54410 32176
rect 54346 32116 54350 32172
rect 54350 32116 54406 32172
rect 54406 32116 54410 32172
rect 54346 32112 54410 32116
rect 54426 32172 54490 32176
rect 54426 32116 54430 32172
rect 54430 32116 54486 32172
rect 54486 32116 54490 32172
rect 54426 32112 54490 32116
rect 54506 32172 54570 32176
rect 54506 32116 54510 32172
rect 54510 32116 54566 32172
rect 54566 32116 54570 32172
rect 54506 32112 54570 32116
rect 59594 32172 59658 32176
rect 59594 32116 59598 32172
rect 59598 32116 59654 32172
rect 59654 32116 59658 32172
rect 59594 32112 59658 32116
rect 59674 32172 59738 32176
rect 59674 32116 59678 32172
rect 59678 32116 59734 32172
rect 59734 32116 59738 32172
rect 59674 32112 59738 32116
rect 59754 32172 59818 32176
rect 59754 32116 59758 32172
rect 59758 32116 59814 32172
rect 59814 32116 59818 32172
rect 59754 32112 59818 32116
rect 59834 32172 59898 32176
rect 59834 32116 59838 32172
rect 59838 32116 59894 32172
rect 59894 32116 59898 32172
rect 59834 32112 59898 32116
rect 64922 32172 64986 32176
rect 64922 32116 64926 32172
rect 64926 32116 64982 32172
rect 64982 32116 64986 32172
rect 64922 32112 64986 32116
rect 65002 32172 65066 32176
rect 65002 32116 65006 32172
rect 65006 32116 65062 32172
rect 65062 32116 65066 32172
rect 65002 32112 65066 32116
rect 65082 32172 65146 32176
rect 65082 32116 65086 32172
rect 65086 32116 65142 32172
rect 65142 32116 65146 32172
rect 65082 32112 65146 32116
rect 65162 32172 65226 32176
rect 65162 32116 65166 32172
rect 65166 32116 65222 32172
rect 65222 32116 65226 32172
rect 65162 32112 65226 32116
rect 70250 32172 70314 32176
rect 70250 32116 70254 32172
rect 70254 32116 70310 32172
rect 70310 32116 70314 32172
rect 70250 32112 70314 32116
rect 70330 32172 70394 32176
rect 70330 32116 70334 32172
rect 70334 32116 70390 32172
rect 70390 32116 70394 32172
rect 70330 32112 70394 32116
rect 70410 32172 70474 32176
rect 70410 32116 70414 32172
rect 70414 32116 70470 32172
rect 70470 32116 70474 32172
rect 70410 32112 70474 32116
rect 70490 32172 70554 32176
rect 70490 32116 70494 32172
rect 70494 32116 70550 32172
rect 70550 32116 70554 32172
rect 70490 32112 70554 32116
rect 75578 32172 75642 32176
rect 75578 32116 75582 32172
rect 75582 32116 75638 32172
rect 75638 32116 75642 32172
rect 75578 32112 75642 32116
rect 75658 32172 75722 32176
rect 75658 32116 75662 32172
rect 75662 32116 75718 32172
rect 75718 32116 75722 32172
rect 75658 32112 75722 32116
rect 75738 32172 75802 32176
rect 75738 32116 75742 32172
rect 75742 32116 75798 32172
rect 75798 32116 75802 32172
rect 75738 32112 75802 32116
rect 75818 32172 75882 32176
rect 75818 32116 75822 32172
rect 75822 32116 75878 32172
rect 75878 32116 75882 32172
rect 75818 32112 75882 32116
rect 80906 32172 80970 32176
rect 80906 32116 80910 32172
rect 80910 32116 80966 32172
rect 80966 32116 80970 32172
rect 80906 32112 80970 32116
rect 80986 32172 81050 32176
rect 80986 32116 80990 32172
rect 80990 32116 81046 32172
rect 81046 32116 81050 32172
rect 80986 32112 81050 32116
rect 81066 32172 81130 32176
rect 81066 32116 81070 32172
rect 81070 32116 81126 32172
rect 81126 32116 81130 32172
rect 81066 32112 81130 32116
rect 81146 32172 81210 32176
rect 81146 32116 81150 32172
rect 81150 32116 81206 32172
rect 81206 32116 81210 32172
rect 81146 32112 81210 32116
rect 86234 32172 86298 32176
rect 86234 32116 86238 32172
rect 86238 32116 86294 32172
rect 86294 32116 86298 32172
rect 86234 32112 86298 32116
rect 86314 32172 86378 32176
rect 86314 32116 86318 32172
rect 86318 32116 86374 32172
rect 86374 32116 86378 32172
rect 86314 32112 86378 32116
rect 86394 32172 86458 32176
rect 86394 32116 86398 32172
rect 86398 32116 86454 32172
rect 86454 32116 86458 32172
rect 86394 32112 86458 32116
rect 86474 32172 86538 32176
rect 86474 32116 86478 32172
rect 86478 32116 86534 32172
rect 86534 32116 86538 32172
rect 86474 32112 86538 32116
rect 91562 32172 91626 32176
rect 91562 32116 91566 32172
rect 91566 32116 91622 32172
rect 91622 32116 91626 32172
rect 91562 32112 91626 32116
rect 91642 32172 91706 32176
rect 91642 32116 91646 32172
rect 91646 32116 91702 32172
rect 91702 32116 91706 32172
rect 91642 32112 91706 32116
rect 91722 32172 91786 32176
rect 91722 32116 91726 32172
rect 91726 32116 91782 32172
rect 91782 32116 91786 32172
rect 91722 32112 91786 32116
rect 91802 32172 91866 32176
rect 91802 32116 91806 32172
rect 91806 32116 91862 32172
rect 91862 32116 91866 32172
rect 91802 32112 91866 32116
rect 3650 31628 3714 31632
rect 3650 31572 3654 31628
rect 3654 31572 3710 31628
rect 3710 31572 3714 31628
rect 3650 31568 3714 31572
rect 3730 31628 3794 31632
rect 3730 31572 3734 31628
rect 3734 31572 3790 31628
rect 3790 31572 3794 31628
rect 3730 31568 3794 31572
rect 3810 31628 3874 31632
rect 3810 31572 3814 31628
rect 3814 31572 3870 31628
rect 3870 31572 3874 31628
rect 3810 31568 3874 31572
rect 3890 31628 3954 31632
rect 3890 31572 3894 31628
rect 3894 31572 3950 31628
rect 3950 31572 3954 31628
rect 3890 31568 3954 31572
rect 8978 31628 9042 31632
rect 8978 31572 8982 31628
rect 8982 31572 9038 31628
rect 9038 31572 9042 31628
rect 8978 31568 9042 31572
rect 9058 31628 9122 31632
rect 9058 31572 9062 31628
rect 9062 31572 9118 31628
rect 9118 31572 9122 31628
rect 9058 31568 9122 31572
rect 9138 31628 9202 31632
rect 9138 31572 9142 31628
rect 9142 31572 9198 31628
rect 9198 31572 9202 31628
rect 9138 31568 9202 31572
rect 9218 31628 9282 31632
rect 9218 31572 9222 31628
rect 9222 31572 9278 31628
rect 9278 31572 9282 31628
rect 9218 31568 9282 31572
rect 14306 31628 14370 31632
rect 14306 31572 14310 31628
rect 14310 31572 14366 31628
rect 14366 31572 14370 31628
rect 14306 31568 14370 31572
rect 14386 31628 14450 31632
rect 14386 31572 14390 31628
rect 14390 31572 14446 31628
rect 14446 31572 14450 31628
rect 14386 31568 14450 31572
rect 14466 31628 14530 31632
rect 14466 31572 14470 31628
rect 14470 31572 14526 31628
rect 14526 31572 14530 31628
rect 14466 31568 14530 31572
rect 14546 31628 14610 31632
rect 14546 31572 14550 31628
rect 14550 31572 14606 31628
rect 14606 31572 14610 31628
rect 14546 31568 14610 31572
rect 19634 31628 19698 31632
rect 19634 31572 19638 31628
rect 19638 31572 19694 31628
rect 19694 31572 19698 31628
rect 19634 31568 19698 31572
rect 19714 31628 19778 31632
rect 19714 31572 19718 31628
rect 19718 31572 19774 31628
rect 19774 31572 19778 31628
rect 19714 31568 19778 31572
rect 19794 31628 19858 31632
rect 19794 31572 19798 31628
rect 19798 31572 19854 31628
rect 19854 31572 19858 31628
rect 19794 31568 19858 31572
rect 19874 31628 19938 31632
rect 19874 31572 19878 31628
rect 19878 31572 19934 31628
rect 19934 31572 19938 31628
rect 19874 31568 19938 31572
rect 24962 31628 25026 31632
rect 24962 31572 24966 31628
rect 24966 31572 25022 31628
rect 25022 31572 25026 31628
rect 24962 31568 25026 31572
rect 25042 31628 25106 31632
rect 25042 31572 25046 31628
rect 25046 31572 25102 31628
rect 25102 31572 25106 31628
rect 25042 31568 25106 31572
rect 25122 31628 25186 31632
rect 25122 31572 25126 31628
rect 25126 31572 25182 31628
rect 25182 31572 25186 31628
rect 25122 31568 25186 31572
rect 25202 31628 25266 31632
rect 25202 31572 25206 31628
rect 25206 31572 25262 31628
rect 25262 31572 25266 31628
rect 25202 31568 25266 31572
rect 30290 31628 30354 31632
rect 30290 31572 30294 31628
rect 30294 31572 30350 31628
rect 30350 31572 30354 31628
rect 30290 31568 30354 31572
rect 30370 31628 30434 31632
rect 30370 31572 30374 31628
rect 30374 31572 30430 31628
rect 30430 31572 30434 31628
rect 30370 31568 30434 31572
rect 30450 31628 30514 31632
rect 30450 31572 30454 31628
rect 30454 31572 30510 31628
rect 30510 31572 30514 31628
rect 30450 31568 30514 31572
rect 30530 31628 30594 31632
rect 30530 31572 30534 31628
rect 30534 31572 30590 31628
rect 30590 31572 30594 31628
rect 30530 31568 30594 31572
rect 35618 31628 35682 31632
rect 35618 31572 35622 31628
rect 35622 31572 35678 31628
rect 35678 31572 35682 31628
rect 35618 31568 35682 31572
rect 35698 31628 35762 31632
rect 35698 31572 35702 31628
rect 35702 31572 35758 31628
rect 35758 31572 35762 31628
rect 35698 31568 35762 31572
rect 35778 31628 35842 31632
rect 35778 31572 35782 31628
rect 35782 31572 35838 31628
rect 35838 31572 35842 31628
rect 35778 31568 35842 31572
rect 35858 31628 35922 31632
rect 35858 31572 35862 31628
rect 35862 31572 35918 31628
rect 35918 31572 35922 31628
rect 35858 31568 35922 31572
rect 40946 31628 41010 31632
rect 40946 31572 40950 31628
rect 40950 31572 41006 31628
rect 41006 31572 41010 31628
rect 40946 31568 41010 31572
rect 41026 31628 41090 31632
rect 41026 31572 41030 31628
rect 41030 31572 41086 31628
rect 41086 31572 41090 31628
rect 41026 31568 41090 31572
rect 41106 31628 41170 31632
rect 41106 31572 41110 31628
rect 41110 31572 41166 31628
rect 41166 31572 41170 31628
rect 41106 31568 41170 31572
rect 41186 31628 41250 31632
rect 41186 31572 41190 31628
rect 41190 31572 41246 31628
rect 41246 31572 41250 31628
rect 41186 31568 41250 31572
rect 46274 31628 46338 31632
rect 46274 31572 46278 31628
rect 46278 31572 46334 31628
rect 46334 31572 46338 31628
rect 46274 31568 46338 31572
rect 46354 31628 46418 31632
rect 46354 31572 46358 31628
rect 46358 31572 46414 31628
rect 46414 31572 46418 31628
rect 46354 31568 46418 31572
rect 46434 31628 46498 31632
rect 46434 31572 46438 31628
rect 46438 31572 46494 31628
rect 46494 31572 46498 31628
rect 46434 31568 46498 31572
rect 46514 31628 46578 31632
rect 46514 31572 46518 31628
rect 46518 31572 46574 31628
rect 46574 31572 46578 31628
rect 46514 31568 46578 31572
rect 51602 31628 51666 31632
rect 51602 31572 51606 31628
rect 51606 31572 51662 31628
rect 51662 31572 51666 31628
rect 51602 31568 51666 31572
rect 51682 31628 51746 31632
rect 51682 31572 51686 31628
rect 51686 31572 51742 31628
rect 51742 31572 51746 31628
rect 51682 31568 51746 31572
rect 51762 31628 51826 31632
rect 51762 31572 51766 31628
rect 51766 31572 51822 31628
rect 51822 31572 51826 31628
rect 51762 31568 51826 31572
rect 51842 31628 51906 31632
rect 51842 31572 51846 31628
rect 51846 31572 51902 31628
rect 51902 31572 51906 31628
rect 51842 31568 51906 31572
rect 56930 31628 56994 31632
rect 56930 31572 56934 31628
rect 56934 31572 56990 31628
rect 56990 31572 56994 31628
rect 56930 31568 56994 31572
rect 57010 31628 57074 31632
rect 57010 31572 57014 31628
rect 57014 31572 57070 31628
rect 57070 31572 57074 31628
rect 57010 31568 57074 31572
rect 57090 31628 57154 31632
rect 57090 31572 57094 31628
rect 57094 31572 57150 31628
rect 57150 31572 57154 31628
rect 57090 31568 57154 31572
rect 57170 31628 57234 31632
rect 57170 31572 57174 31628
rect 57174 31572 57230 31628
rect 57230 31572 57234 31628
rect 57170 31568 57234 31572
rect 62258 31628 62322 31632
rect 62258 31572 62262 31628
rect 62262 31572 62318 31628
rect 62318 31572 62322 31628
rect 62258 31568 62322 31572
rect 62338 31628 62402 31632
rect 62338 31572 62342 31628
rect 62342 31572 62398 31628
rect 62398 31572 62402 31628
rect 62338 31568 62402 31572
rect 62418 31628 62482 31632
rect 62418 31572 62422 31628
rect 62422 31572 62478 31628
rect 62478 31572 62482 31628
rect 62418 31568 62482 31572
rect 62498 31628 62562 31632
rect 62498 31572 62502 31628
rect 62502 31572 62558 31628
rect 62558 31572 62562 31628
rect 62498 31568 62562 31572
rect 67586 31628 67650 31632
rect 67586 31572 67590 31628
rect 67590 31572 67646 31628
rect 67646 31572 67650 31628
rect 67586 31568 67650 31572
rect 67666 31628 67730 31632
rect 67666 31572 67670 31628
rect 67670 31572 67726 31628
rect 67726 31572 67730 31628
rect 67666 31568 67730 31572
rect 67746 31628 67810 31632
rect 67746 31572 67750 31628
rect 67750 31572 67806 31628
rect 67806 31572 67810 31628
rect 67746 31568 67810 31572
rect 67826 31628 67890 31632
rect 67826 31572 67830 31628
rect 67830 31572 67886 31628
rect 67886 31572 67890 31628
rect 67826 31568 67890 31572
rect 72914 31628 72978 31632
rect 72914 31572 72918 31628
rect 72918 31572 72974 31628
rect 72974 31572 72978 31628
rect 72914 31568 72978 31572
rect 72994 31628 73058 31632
rect 72994 31572 72998 31628
rect 72998 31572 73054 31628
rect 73054 31572 73058 31628
rect 72994 31568 73058 31572
rect 73074 31628 73138 31632
rect 73074 31572 73078 31628
rect 73078 31572 73134 31628
rect 73134 31572 73138 31628
rect 73074 31568 73138 31572
rect 73154 31628 73218 31632
rect 73154 31572 73158 31628
rect 73158 31572 73214 31628
rect 73214 31572 73218 31628
rect 73154 31568 73218 31572
rect 78242 31628 78306 31632
rect 78242 31572 78246 31628
rect 78246 31572 78302 31628
rect 78302 31572 78306 31628
rect 78242 31568 78306 31572
rect 78322 31628 78386 31632
rect 78322 31572 78326 31628
rect 78326 31572 78382 31628
rect 78382 31572 78386 31628
rect 78322 31568 78386 31572
rect 78402 31628 78466 31632
rect 78402 31572 78406 31628
rect 78406 31572 78462 31628
rect 78462 31572 78466 31628
rect 78402 31568 78466 31572
rect 78482 31628 78546 31632
rect 78482 31572 78486 31628
rect 78486 31572 78542 31628
rect 78542 31572 78546 31628
rect 78482 31568 78546 31572
rect 83570 31628 83634 31632
rect 83570 31572 83574 31628
rect 83574 31572 83630 31628
rect 83630 31572 83634 31628
rect 83570 31568 83634 31572
rect 83650 31628 83714 31632
rect 83650 31572 83654 31628
rect 83654 31572 83710 31628
rect 83710 31572 83714 31628
rect 83650 31568 83714 31572
rect 83730 31628 83794 31632
rect 83730 31572 83734 31628
rect 83734 31572 83790 31628
rect 83790 31572 83794 31628
rect 83730 31568 83794 31572
rect 83810 31628 83874 31632
rect 83810 31572 83814 31628
rect 83814 31572 83870 31628
rect 83870 31572 83874 31628
rect 83810 31568 83874 31572
rect 88898 31628 88962 31632
rect 88898 31572 88902 31628
rect 88902 31572 88958 31628
rect 88958 31572 88962 31628
rect 88898 31568 88962 31572
rect 88978 31628 89042 31632
rect 88978 31572 88982 31628
rect 88982 31572 89038 31628
rect 89038 31572 89042 31628
rect 88978 31568 89042 31572
rect 89058 31628 89122 31632
rect 89058 31572 89062 31628
rect 89062 31572 89118 31628
rect 89118 31572 89122 31628
rect 89058 31568 89122 31572
rect 89138 31628 89202 31632
rect 89138 31572 89142 31628
rect 89142 31572 89198 31628
rect 89198 31572 89202 31628
rect 89138 31568 89202 31572
rect 6314 31084 6378 31088
rect 6314 31028 6318 31084
rect 6318 31028 6374 31084
rect 6374 31028 6378 31084
rect 6314 31024 6378 31028
rect 6394 31084 6458 31088
rect 6394 31028 6398 31084
rect 6398 31028 6454 31084
rect 6454 31028 6458 31084
rect 6394 31024 6458 31028
rect 6474 31084 6538 31088
rect 6474 31028 6478 31084
rect 6478 31028 6534 31084
rect 6534 31028 6538 31084
rect 6474 31024 6538 31028
rect 6554 31084 6618 31088
rect 6554 31028 6558 31084
rect 6558 31028 6614 31084
rect 6614 31028 6618 31084
rect 6554 31024 6618 31028
rect 11642 31084 11706 31088
rect 11642 31028 11646 31084
rect 11646 31028 11702 31084
rect 11702 31028 11706 31084
rect 11642 31024 11706 31028
rect 11722 31084 11786 31088
rect 11722 31028 11726 31084
rect 11726 31028 11782 31084
rect 11782 31028 11786 31084
rect 11722 31024 11786 31028
rect 11802 31084 11866 31088
rect 11802 31028 11806 31084
rect 11806 31028 11862 31084
rect 11862 31028 11866 31084
rect 11802 31024 11866 31028
rect 11882 31084 11946 31088
rect 11882 31028 11886 31084
rect 11886 31028 11942 31084
rect 11942 31028 11946 31084
rect 11882 31024 11946 31028
rect 16970 31084 17034 31088
rect 16970 31028 16974 31084
rect 16974 31028 17030 31084
rect 17030 31028 17034 31084
rect 16970 31024 17034 31028
rect 17050 31084 17114 31088
rect 17050 31028 17054 31084
rect 17054 31028 17110 31084
rect 17110 31028 17114 31084
rect 17050 31024 17114 31028
rect 17130 31084 17194 31088
rect 17130 31028 17134 31084
rect 17134 31028 17190 31084
rect 17190 31028 17194 31084
rect 17130 31024 17194 31028
rect 17210 31084 17274 31088
rect 17210 31028 17214 31084
rect 17214 31028 17270 31084
rect 17270 31028 17274 31084
rect 17210 31024 17274 31028
rect 22298 31084 22362 31088
rect 22298 31028 22302 31084
rect 22302 31028 22358 31084
rect 22358 31028 22362 31084
rect 22298 31024 22362 31028
rect 22378 31084 22442 31088
rect 22378 31028 22382 31084
rect 22382 31028 22438 31084
rect 22438 31028 22442 31084
rect 22378 31024 22442 31028
rect 22458 31084 22522 31088
rect 22458 31028 22462 31084
rect 22462 31028 22518 31084
rect 22518 31028 22522 31084
rect 22458 31024 22522 31028
rect 22538 31084 22602 31088
rect 22538 31028 22542 31084
rect 22542 31028 22598 31084
rect 22598 31028 22602 31084
rect 22538 31024 22602 31028
rect 27626 31084 27690 31088
rect 27626 31028 27630 31084
rect 27630 31028 27686 31084
rect 27686 31028 27690 31084
rect 27626 31024 27690 31028
rect 27706 31084 27770 31088
rect 27706 31028 27710 31084
rect 27710 31028 27766 31084
rect 27766 31028 27770 31084
rect 27706 31024 27770 31028
rect 27786 31084 27850 31088
rect 27786 31028 27790 31084
rect 27790 31028 27846 31084
rect 27846 31028 27850 31084
rect 27786 31024 27850 31028
rect 27866 31084 27930 31088
rect 27866 31028 27870 31084
rect 27870 31028 27926 31084
rect 27926 31028 27930 31084
rect 27866 31024 27930 31028
rect 32954 31084 33018 31088
rect 32954 31028 32958 31084
rect 32958 31028 33014 31084
rect 33014 31028 33018 31084
rect 32954 31024 33018 31028
rect 33034 31084 33098 31088
rect 33034 31028 33038 31084
rect 33038 31028 33094 31084
rect 33094 31028 33098 31084
rect 33034 31024 33098 31028
rect 33114 31084 33178 31088
rect 33114 31028 33118 31084
rect 33118 31028 33174 31084
rect 33174 31028 33178 31084
rect 33114 31024 33178 31028
rect 33194 31084 33258 31088
rect 33194 31028 33198 31084
rect 33198 31028 33254 31084
rect 33254 31028 33258 31084
rect 33194 31024 33258 31028
rect 38282 31084 38346 31088
rect 38282 31028 38286 31084
rect 38286 31028 38342 31084
rect 38342 31028 38346 31084
rect 38282 31024 38346 31028
rect 38362 31084 38426 31088
rect 38362 31028 38366 31084
rect 38366 31028 38422 31084
rect 38422 31028 38426 31084
rect 38362 31024 38426 31028
rect 38442 31084 38506 31088
rect 38442 31028 38446 31084
rect 38446 31028 38502 31084
rect 38502 31028 38506 31084
rect 38442 31024 38506 31028
rect 38522 31084 38586 31088
rect 38522 31028 38526 31084
rect 38526 31028 38582 31084
rect 38582 31028 38586 31084
rect 38522 31024 38586 31028
rect 43610 31084 43674 31088
rect 43610 31028 43614 31084
rect 43614 31028 43670 31084
rect 43670 31028 43674 31084
rect 43610 31024 43674 31028
rect 43690 31084 43754 31088
rect 43690 31028 43694 31084
rect 43694 31028 43750 31084
rect 43750 31028 43754 31084
rect 43690 31024 43754 31028
rect 43770 31084 43834 31088
rect 43770 31028 43774 31084
rect 43774 31028 43830 31084
rect 43830 31028 43834 31084
rect 43770 31024 43834 31028
rect 43850 31084 43914 31088
rect 43850 31028 43854 31084
rect 43854 31028 43910 31084
rect 43910 31028 43914 31084
rect 43850 31024 43914 31028
rect 48938 31084 49002 31088
rect 48938 31028 48942 31084
rect 48942 31028 48998 31084
rect 48998 31028 49002 31084
rect 48938 31024 49002 31028
rect 49018 31084 49082 31088
rect 49018 31028 49022 31084
rect 49022 31028 49078 31084
rect 49078 31028 49082 31084
rect 49018 31024 49082 31028
rect 49098 31084 49162 31088
rect 49098 31028 49102 31084
rect 49102 31028 49158 31084
rect 49158 31028 49162 31084
rect 49098 31024 49162 31028
rect 49178 31084 49242 31088
rect 49178 31028 49182 31084
rect 49182 31028 49238 31084
rect 49238 31028 49242 31084
rect 49178 31024 49242 31028
rect 54266 31084 54330 31088
rect 54266 31028 54270 31084
rect 54270 31028 54326 31084
rect 54326 31028 54330 31084
rect 54266 31024 54330 31028
rect 54346 31084 54410 31088
rect 54346 31028 54350 31084
rect 54350 31028 54406 31084
rect 54406 31028 54410 31084
rect 54346 31024 54410 31028
rect 54426 31084 54490 31088
rect 54426 31028 54430 31084
rect 54430 31028 54486 31084
rect 54486 31028 54490 31084
rect 54426 31024 54490 31028
rect 54506 31084 54570 31088
rect 54506 31028 54510 31084
rect 54510 31028 54566 31084
rect 54566 31028 54570 31084
rect 54506 31024 54570 31028
rect 59594 31084 59658 31088
rect 59594 31028 59598 31084
rect 59598 31028 59654 31084
rect 59654 31028 59658 31084
rect 59594 31024 59658 31028
rect 59674 31084 59738 31088
rect 59674 31028 59678 31084
rect 59678 31028 59734 31084
rect 59734 31028 59738 31084
rect 59674 31024 59738 31028
rect 59754 31084 59818 31088
rect 59754 31028 59758 31084
rect 59758 31028 59814 31084
rect 59814 31028 59818 31084
rect 59754 31024 59818 31028
rect 59834 31084 59898 31088
rect 59834 31028 59838 31084
rect 59838 31028 59894 31084
rect 59894 31028 59898 31084
rect 59834 31024 59898 31028
rect 64922 31084 64986 31088
rect 64922 31028 64926 31084
rect 64926 31028 64982 31084
rect 64982 31028 64986 31084
rect 64922 31024 64986 31028
rect 65002 31084 65066 31088
rect 65002 31028 65006 31084
rect 65006 31028 65062 31084
rect 65062 31028 65066 31084
rect 65002 31024 65066 31028
rect 65082 31084 65146 31088
rect 65082 31028 65086 31084
rect 65086 31028 65142 31084
rect 65142 31028 65146 31084
rect 65082 31024 65146 31028
rect 65162 31084 65226 31088
rect 65162 31028 65166 31084
rect 65166 31028 65222 31084
rect 65222 31028 65226 31084
rect 65162 31024 65226 31028
rect 70250 31084 70314 31088
rect 70250 31028 70254 31084
rect 70254 31028 70310 31084
rect 70310 31028 70314 31084
rect 70250 31024 70314 31028
rect 70330 31084 70394 31088
rect 70330 31028 70334 31084
rect 70334 31028 70390 31084
rect 70390 31028 70394 31084
rect 70330 31024 70394 31028
rect 70410 31084 70474 31088
rect 70410 31028 70414 31084
rect 70414 31028 70470 31084
rect 70470 31028 70474 31084
rect 70410 31024 70474 31028
rect 70490 31084 70554 31088
rect 70490 31028 70494 31084
rect 70494 31028 70550 31084
rect 70550 31028 70554 31084
rect 70490 31024 70554 31028
rect 75578 31084 75642 31088
rect 75578 31028 75582 31084
rect 75582 31028 75638 31084
rect 75638 31028 75642 31084
rect 75578 31024 75642 31028
rect 75658 31084 75722 31088
rect 75658 31028 75662 31084
rect 75662 31028 75718 31084
rect 75718 31028 75722 31084
rect 75658 31024 75722 31028
rect 75738 31084 75802 31088
rect 75738 31028 75742 31084
rect 75742 31028 75798 31084
rect 75798 31028 75802 31084
rect 75738 31024 75802 31028
rect 75818 31084 75882 31088
rect 75818 31028 75822 31084
rect 75822 31028 75878 31084
rect 75878 31028 75882 31084
rect 75818 31024 75882 31028
rect 80906 31084 80970 31088
rect 80906 31028 80910 31084
rect 80910 31028 80966 31084
rect 80966 31028 80970 31084
rect 80906 31024 80970 31028
rect 80986 31084 81050 31088
rect 80986 31028 80990 31084
rect 80990 31028 81046 31084
rect 81046 31028 81050 31084
rect 80986 31024 81050 31028
rect 81066 31084 81130 31088
rect 81066 31028 81070 31084
rect 81070 31028 81126 31084
rect 81126 31028 81130 31084
rect 81066 31024 81130 31028
rect 81146 31084 81210 31088
rect 81146 31028 81150 31084
rect 81150 31028 81206 31084
rect 81206 31028 81210 31084
rect 81146 31024 81210 31028
rect 86234 31084 86298 31088
rect 86234 31028 86238 31084
rect 86238 31028 86294 31084
rect 86294 31028 86298 31084
rect 86234 31024 86298 31028
rect 86314 31084 86378 31088
rect 86314 31028 86318 31084
rect 86318 31028 86374 31084
rect 86374 31028 86378 31084
rect 86314 31024 86378 31028
rect 86394 31084 86458 31088
rect 86394 31028 86398 31084
rect 86398 31028 86454 31084
rect 86454 31028 86458 31084
rect 86394 31024 86458 31028
rect 86474 31084 86538 31088
rect 86474 31028 86478 31084
rect 86478 31028 86534 31084
rect 86534 31028 86538 31084
rect 86474 31024 86538 31028
rect 91562 31084 91626 31088
rect 91562 31028 91566 31084
rect 91566 31028 91622 31084
rect 91622 31028 91626 31084
rect 91562 31024 91626 31028
rect 91642 31084 91706 31088
rect 91642 31028 91646 31084
rect 91646 31028 91702 31084
rect 91702 31028 91706 31084
rect 91642 31024 91706 31028
rect 91722 31084 91786 31088
rect 91722 31028 91726 31084
rect 91726 31028 91782 31084
rect 91782 31028 91786 31084
rect 91722 31024 91786 31028
rect 91802 31084 91866 31088
rect 91802 31028 91806 31084
rect 91806 31028 91862 31084
rect 91862 31028 91866 31084
rect 91802 31024 91866 31028
rect 3650 30540 3714 30544
rect 3650 30484 3654 30540
rect 3654 30484 3710 30540
rect 3710 30484 3714 30540
rect 3650 30480 3714 30484
rect 3730 30540 3794 30544
rect 3730 30484 3734 30540
rect 3734 30484 3790 30540
rect 3790 30484 3794 30540
rect 3730 30480 3794 30484
rect 3810 30540 3874 30544
rect 3810 30484 3814 30540
rect 3814 30484 3870 30540
rect 3870 30484 3874 30540
rect 3810 30480 3874 30484
rect 3890 30540 3954 30544
rect 3890 30484 3894 30540
rect 3894 30484 3950 30540
rect 3950 30484 3954 30540
rect 3890 30480 3954 30484
rect 8978 30540 9042 30544
rect 8978 30484 8982 30540
rect 8982 30484 9038 30540
rect 9038 30484 9042 30540
rect 8978 30480 9042 30484
rect 9058 30540 9122 30544
rect 9058 30484 9062 30540
rect 9062 30484 9118 30540
rect 9118 30484 9122 30540
rect 9058 30480 9122 30484
rect 9138 30540 9202 30544
rect 9138 30484 9142 30540
rect 9142 30484 9198 30540
rect 9198 30484 9202 30540
rect 9138 30480 9202 30484
rect 9218 30540 9282 30544
rect 9218 30484 9222 30540
rect 9222 30484 9278 30540
rect 9278 30484 9282 30540
rect 9218 30480 9282 30484
rect 14306 30540 14370 30544
rect 14306 30484 14310 30540
rect 14310 30484 14366 30540
rect 14366 30484 14370 30540
rect 14306 30480 14370 30484
rect 14386 30540 14450 30544
rect 14386 30484 14390 30540
rect 14390 30484 14446 30540
rect 14446 30484 14450 30540
rect 14386 30480 14450 30484
rect 14466 30540 14530 30544
rect 14466 30484 14470 30540
rect 14470 30484 14526 30540
rect 14526 30484 14530 30540
rect 14466 30480 14530 30484
rect 14546 30540 14610 30544
rect 14546 30484 14550 30540
rect 14550 30484 14606 30540
rect 14606 30484 14610 30540
rect 14546 30480 14610 30484
rect 19634 30540 19698 30544
rect 19634 30484 19638 30540
rect 19638 30484 19694 30540
rect 19694 30484 19698 30540
rect 19634 30480 19698 30484
rect 19714 30540 19778 30544
rect 19714 30484 19718 30540
rect 19718 30484 19774 30540
rect 19774 30484 19778 30540
rect 19714 30480 19778 30484
rect 19794 30540 19858 30544
rect 19794 30484 19798 30540
rect 19798 30484 19854 30540
rect 19854 30484 19858 30540
rect 19794 30480 19858 30484
rect 19874 30540 19938 30544
rect 19874 30484 19878 30540
rect 19878 30484 19934 30540
rect 19934 30484 19938 30540
rect 19874 30480 19938 30484
rect 24962 30540 25026 30544
rect 24962 30484 24966 30540
rect 24966 30484 25022 30540
rect 25022 30484 25026 30540
rect 24962 30480 25026 30484
rect 25042 30540 25106 30544
rect 25042 30484 25046 30540
rect 25046 30484 25102 30540
rect 25102 30484 25106 30540
rect 25042 30480 25106 30484
rect 25122 30540 25186 30544
rect 25122 30484 25126 30540
rect 25126 30484 25182 30540
rect 25182 30484 25186 30540
rect 25122 30480 25186 30484
rect 25202 30540 25266 30544
rect 25202 30484 25206 30540
rect 25206 30484 25262 30540
rect 25262 30484 25266 30540
rect 25202 30480 25266 30484
rect 30290 30540 30354 30544
rect 30290 30484 30294 30540
rect 30294 30484 30350 30540
rect 30350 30484 30354 30540
rect 30290 30480 30354 30484
rect 30370 30540 30434 30544
rect 30370 30484 30374 30540
rect 30374 30484 30430 30540
rect 30430 30484 30434 30540
rect 30370 30480 30434 30484
rect 30450 30540 30514 30544
rect 30450 30484 30454 30540
rect 30454 30484 30510 30540
rect 30510 30484 30514 30540
rect 30450 30480 30514 30484
rect 30530 30540 30594 30544
rect 30530 30484 30534 30540
rect 30534 30484 30590 30540
rect 30590 30484 30594 30540
rect 30530 30480 30594 30484
rect 35618 30540 35682 30544
rect 35618 30484 35622 30540
rect 35622 30484 35678 30540
rect 35678 30484 35682 30540
rect 35618 30480 35682 30484
rect 35698 30540 35762 30544
rect 35698 30484 35702 30540
rect 35702 30484 35758 30540
rect 35758 30484 35762 30540
rect 35698 30480 35762 30484
rect 35778 30540 35842 30544
rect 35778 30484 35782 30540
rect 35782 30484 35838 30540
rect 35838 30484 35842 30540
rect 35778 30480 35842 30484
rect 35858 30540 35922 30544
rect 35858 30484 35862 30540
rect 35862 30484 35918 30540
rect 35918 30484 35922 30540
rect 35858 30480 35922 30484
rect 40946 30540 41010 30544
rect 40946 30484 40950 30540
rect 40950 30484 41006 30540
rect 41006 30484 41010 30540
rect 40946 30480 41010 30484
rect 41026 30540 41090 30544
rect 41026 30484 41030 30540
rect 41030 30484 41086 30540
rect 41086 30484 41090 30540
rect 41026 30480 41090 30484
rect 41106 30540 41170 30544
rect 41106 30484 41110 30540
rect 41110 30484 41166 30540
rect 41166 30484 41170 30540
rect 41106 30480 41170 30484
rect 41186 30540 41250 30544
rect 41186 30484 41190 30540
rect 41190 30484 41246 30540
rect 41246 30484 41250 30540
rect 41186 30480 41250 30484
rect 46274 30540 46338 30544
rect 46274 30484 46278 30540
rect 46278 30484 46334 30540
rect 46334 30484 46338 30540
rect 46274 30480 46338 30484
rect 46354 30540 46418 30544
rect 46354 30484 46358 30540
rect 46358 30484 46414 30540
rect 46414 30484 46418 30540
rect 46354 30480 46418 30484
rect 46434 30540 46498 30544
rect 46434 30484 46438 30540
rect 46438 30484 46494 30540
rect 46494 30484 46498 30540
rect 46434 30480 46498 30484
rect 46514 30540 46578 30544
rect 46514 30484 46518 30540
rect 46518 30484 46574 30540
rect 46574 30484 46578 30540
rect 46514 30480 46578 30484
rect 51602 30540 51666 30544
rect 51602 30484 51606 30540
rect 51606 30484 51662 30540
rect 51662 30484 51666 30540
rect 51602 30480 51666 30484
rect 51682 30540 51746 30544
rect 51682 30484 51686 30540
rect 51686 30484 51742 30540
rect 51742 30484 51746 30540
rect 51682 30480 51746 30484
rect 51762 30540 51826 30544
rect 51762 30484 51766 30540
rect 51766 30484 51822 30540
rect 51822 30484 51826 30540
rect 51762 30480 51826 30484
rect 51842 30540 51906 30544
rect 51842 30484 51846 30540
rect 51846 30484 51902 30540
rect 51902 30484 51906 30540
rect 51842 30480 51906 30484
rect 56930 30540 56994 30544
rect 56930 30484 56934 30540
rect 56934 30484 56990 30540
rect 56990 30484 56994 30540
rect 56930 30480 56994 30484
rect 57010 30540 57074 30544
rect 57010 30484 57014 30540
rect 57014 30484 57070 30540
rect 57070 30484 57074 30540
rect 57010 30480 57074 30484
rect 57090 30540 57154 30544
rect 57090 30484 57094 30540
rect 57094 30484 57150 30540
rect 57150 30484 57154 30540
rect 57090 30480 57154 30484
rect 57170 30540 57234 30544
rect 57170 30484 57174 30540
rect 57174 30484 57230 30540
rect 57230 30484 57234 30540
rect 57170 30480 57234 30484
rect 62258 30540 62322 30544
rect 62258 30484 62262 30540
rect 62262 30484 62318 30540
rect 62318 30484 62322 30540
rect 62258 30480 62322 30484
rect 62338 30540 62402 30544
rect 62338 30484 62342 30540
rect 62342 30484 62398 30540
rect 62398 30484 62402 30540
rect 62338 30480 62402 30484
rect 62418 30540 62482 30544
rect 62418 30484 62422 30540
rect 62422 30484 62478 30540
rect 62478 30484 62482 30540
rect 62418 30480 62482 30484
rect 62498 30540 62562 30544
rect 62498 30484 62502 30540
rect 62502 30484 62558 30540
rect 62558 30484 62562 30540
rect 62498 30480 62562 30484
rect 67586 30540 67650 30544
rect 67586 30484 67590 30540
rect 67590 30484 67646 30540
rect 67646 30484 67650 30540
rect 67586 30480 67650 30484
rect 67666 30540 67730 30544
rect 67666 30484 67670 30540
rect 67670 30484 67726 30540
rect 67726 30484 67730 30540
rect 67666 30480 67730 30484
rect 67746 30540 67810 30544
rect 67746 30484 67750 30540
rect 67750 30484 67806 30540
rect 67806 30484 67810 30540
rect 67746 30480 67810 30484
rect 67826 30540 67890 30544
rect 67826 30484 67830 30540
rect 67830 30484 67886 30540
rect 67886 30484 67890 30540
rect 67826 30480 67890 30484
rect 72914 30540 72978 30544
rect 72914 30484 72918 30540
rect 72918 30484 72974 30540
rect 72974 30484 72978 30540
rect 72914 30480 72978 30484
rect 72994 30540 73058 30544
rect 72994 30484 72998 30540
rect 72998 30484 73054 30540
rect 73054 30484 73058 30540
rect 72994 30480 73058 30484
rect 73074 30540 73138 30544
rect 73074 30484 73078 30540
rect 73078 30484 73134 30540
rect 73134 30484 73138 30540
rect 73074 30480 73138 30484
rect 73154 30540 73218 30544
rect 73154 30484 73158 30540
rect 73158 30484 73214 30540
rect 73214 30484 73218 30540
rect 73154 30480 73218 30484
rect 78242 30540 78306 30544
rect 78242 30484 78246 30540
rect 78246 30484 78302 30540
rect 78302 30484 78306 30540
rect 78242 30480 78306 30484
rect 78322 30540 78386 30544
rect 78322 30484 78326 30540
rect 78326 30484 78382 30540
rect 78382 30484 78386 30540
rect 78322 30480 78386 30484
rect 78402 30540 78466 30544
rect 78402 30484 78406 30540
rect 78406 30484 78462 30540
rect 78462 30484 78466 30540
rect 78402 30480 78466 30484
rect 78482 30540 78546 30544
rect 78482 30484 78486 30540
rect 78486 30484 78542 30540
rect 78542 30484 78546 30540
rect 78482 30480 78546 30484
rect 83570 30540 83634 30544
rect 83570 30484 83574 30540
rect 83574 30484 83630 30540
rect 83630 30484 83634 30540
rect 83570 30480 83634 30484
rect 83650 30540 83714 30544
rect 83650 30484 83654 30540
rect 83654 30484 83710 30540
rect 83710 30484 83714 30540
rect 83650 30480 83714 30484
rect 83730 30540 83794 30544
rect 83730 30484 83734 30540
rect 83734 30484 83790 30540
rect 83790 30484 83794 30540
rect 83730 30480 83794 30484
rect 83810 30540 83874 30544
rect 83810 30484 83814 30540
rect 83814 30484 83870 30540
rect 83870 30484 83874 30540
rect 83810 30480 83874 30484
rect 88898 30540 88962 30544
rect 88898 30484 88902 30540
rect 88902 30484 88958 30540
rect 88958 30484 88962 30540
rect 88898 30480 88962 30484
rect 88978 30540 89042 30544
rect 88978 30484 88982 30540
rect 88982 30484 89038 30540
rect 89038 30484 89042 30540
rect 88978 30480 89042 30484
rect 89058 30540 89122 30544
rect 89058 30484 89062 30540
rect 89062 30484 89118 30540
rect 89118 30484 89122 30540
rect 89058 30480 89122 30484
rect 89138 30540 89202 30544
rect 89138 30484 89142 30540
rect 89142 30484 89198 30540
rect 89198 30484 89202 30540
rect 89138 30480 89202 30484
rect 6314 29996 6378 30000
rect 6314 29940 6318 29996
rect 6318 29940 6374 29996
rect 6374 29940 6378 29996
rect 6314 29936 6378 29940
rect 6394 29996 6458 30000
rect 6394 29940 6398 29996
rect 6398 29940 6454 29996
rect 6454 29940 6458 29996
rect 6394 29936 6458 29940
rect 6474 29996 6538 30000
rect 6474 29940 6478 29996
rect 6478 29940 6534 29996
rect 6534 29940 6538 29996
rect 6474 29936 6538 29940
rect 6554 29996 6618 30000
rect 6554 29940 6558 29996
rect 6558 29940 6614 29996
rect 6614 29940 6618 29996
rect 6554 29936 6618 29940
rect 11642 29996 11706 30000
rect 11642 29940 11646 29996
rect 11646 29940 11702 29996
rect 11702 29940 11706 29996
rect 11642 29936 11706 29940
rect 11722 29996 11786 30000
rect 11722 29940 11726 29996
rect 11726 29940 11782 29996
rect 11782 29940 11786 29996
rect 11722 29936 11786 29940
rect 11802 29996 11866 30000
rect 11802 29940 11806 29996
rect 11806 29940 11862 29996
rect 11862 29940 11866 29996
rect 11802 29936 11866 29940
rect 11882 29996 11946 30000
rect 11882 29940 11886 29996
rect 11886 29940 11942 29996
rect 11942 29940 11946 29996
rect 11882 29936 11946 29940
rect 16970 29996 17034 30000
rect 16970 29940 16974 29996
rect 16974 29940 17030 29996
rect 17030 29940 17034 29996
rect 16970 29936 17034 29940
rect 17050 29996 17114 30000
rect 17050 29940 17054 29996
rect 17054 29940 17110 29996
rect 17110 29940 17114 29996
rect 17050 29936 17114 29940
rect 17130 29996 17194 30000
rect 17130 29940 17134 29996
rect 17134 29940 17190 29996
rect 17190 29940 17194 29996
rect 17130 29936 17194 29940
rect 17210 29996 17274 30000
rect 17210 29940 17214 29996
rect 17214 29940 17270 29996
rect 17270 29940 17274 29996
rect 17210 29936 17274 29940
rect 22298 29996 22362 30000
rect 22298 29940 22302 29996
rect 22302 29940 22358 29996
rect 22358 29940 22362 29996
rect 22298 29936 22362 29940
rect 22378 29996 22442 30000
rect 22378 29940 22382 29996
rect 22382 29940 22438 29996
rect 22438 29940 22442 29996
rect 22378 29936 22442 29940
rect 22458 29996 22522 30000
rect 22458 29940 22462 29996
rect 22462 29940 22518 29996
rect 22518 29940 22522 29996
rect 22458 29936 22522 29940
rect 22538 29996 22602 30000
rect 22538 29940 22542 29996
rect 22542 29940 22598 29996
rect 22598 29940 22602 29996
rect 22538 29936 22602 29940
rect 27626 29996 27690 30000
rect 27626 29940 27630 29996
rect 27630 29940 27686 29996
rect 27686 29940 27690 29996
rect 27626 29936 27690 29940
rect 27706 29996 27770 30000
rect 27706 29940 27710 29996
rect 27710 29940 27766 29996
rect 27766 29940 27770 29996
rect 27706 29936 27770 29940
rect 27786 29996 27850 30000
rect 27786 29940 27790 29996
rect 27790 29940 27846 29996
rect 27846 29940 27850 29996
rect 27786 29936 27850 29940
rect 27866 29996 27930 30000
rect 27866 29940 27870 29996
rect 27870 29940 27926 29996
rect 27926 29940 27930 29996
rect 27866 29936 27930 29940
rect 32954 29996 33018 30000
rect 32954 29940 32958 29996
rect 32958 29940 33014 29996
rect 33014 29940 33018 29996
rect 32954 29936 33018 29940
rect 33034 29996 33098 30000
rect 33034 29940 33038 29996
rect 33038 29940 33094 29996
rect 33094 29940 33098 29996
rect 33034 29936 33098 29940
rect 33114 29996 33178 30000
rect 33114 29940 33118 29996
rect 33118 29940 33174 29996
rect 33174 29940 33178 29996
rect 33114 29936 33178 29940
rect 33194 29996 33258 30000
rect 33194 29940 33198 29996
rect 33198 29940 33254 29996
rect 33254 29940 33258 29996
rect 33194 29936 33258 29940
rect 38282 29996 38346 30000
rect 38282 29940 38286 29996
rect 38286 29940 38342 29996
rect 38342 29940 38346 29996
rect 38282 29936 38346 29940
rect 38362 29996 38426 30000
rect 38362 29940 38366 29996
rect 38366 29940 38422 29996
rect 38422 29940 38426 29996
rect 38362 29936 38426 29940
rect 38442 29996 38506 30000
rect 38442 29940 38446 29996
rect 38446 29940 38502 29996
rect 38502 29940 38506 29996
rect 38442 29936 38506 29940
rect 38522 29996 38586 30000
rect 38522 29940 38526 29996
rect 38526 29940 38582 29996
rect 38582 29940 38586 29996
rect 38522 29936 38586 29940
rect 43610 29996 43674 30000
rect 43610 29940 43614 29996
rect 43614 29940 43670 29996
rect 43670 29940 43674 29996
rect 43610 29936 43674 29940
rect 43690 29996 43754 30000
rect 43690 29940 43694 29996
rect 43694 29940 43750 29996
rect 43750 29940 43754 29996
rect 43690 29936 43754 29940
rect 43770 29996 43834 30000
rect 43770 29940 43774 29996
rect 43774 29940 43830 29996
rect 43830 29940 43834 29996
rect 43770 29936 43834 29940
rect 43850 29996 43914 30000
rect 43850 29940 43854 29996
rect 43854 29940 43910 29996
rect 43910 29940 43914 29996
rect 43850 29936 43914 29940
rect 48938 29996 49002 30000
rect 48938 29940 48942 29996
rect 48942 29940 48998 29996
rect 48998 29940 49002 29996
rect 48938 29936 49002 29940
rect 49018 29996 49082 30000
rect 49018 29940 49022 29996
rect 49022 29940 49078 29996
rect 49078 29940 49082 29996
rect 49018 29936 49082 29940
rect 49098 29996 49162 30000
rect 49098 29940 49102 29996
rect 49102 29940 49158 29996
rect 49158 29940 49162 29996
rect 49098 29936 49162 29940
rect 49178 29996 49242 30000
rect 49178 29940 49182 29996
rect 49182 29940 49238 29996
rect 49238 29940 49242 29996
rect 49178 29936 49242 29940
rect 54266 29996 54330 30000
rect 54266 29940 54270 29996
rect 54270 29940 54326 29996
rect 54326 29940 54330 29996
rect 54266 29936 54330 29940
rect 54346 29996 54410 30000
rect 54346 29940 54350 29996
rect 54350 29940 54406 29996
rect 54406 29940 54410 29996
rect 54346 29936 54410 29940
rect 54426 29996 54490 30000
rect 54426 29940 54430 29996
rect 54430 29940 54486 29996
rect 54486 29940 54490 29996
rect 54426 29936 54490 29940
rect 54506 29996 54570 30000
rect 54506 29940 54510 29996
rect 54510 29940 54566 29996
rect 54566 29940 54570 29996
rect 54506 29936 54570 29940
rect 59594 29996 59658 30000
rect 59594 29940 59598 29996
rect 59598 29940 59654 29996
rect 59654 29940 59658 29996
rect 59594 29936 59658 29940
rect 59674 29996 59738 30000
rect 59674 29940 59678 29996
rect 59678 29940 59734 29996
rect 59734 29940 59738 29996
rect 59674 29936 59738 29940
rect 59754 29996 59818 30000
rect 59754 29940 59758 29996
rect 59758 29940 59814 29996
rect 59814 29940 59818 29996
rect 59754 29936 59818 29940
rect 59834 29996 59898 30000
rect 59834 29940 59838 29996
rect 59838 29940 59894 29996
rect 59894 29940 59898 29996
rect 59834 29936 59898 29940
rect 64922 29996 64986 30000
rect 64922 29940 64926 29996
rect 64926 29940 64982 29996
rect 64982 29940 64986 29996
rect 64922 29936 64986 29940
rect 65002 29996 65066 30000
rect 65002 29940 65006 29996
rect 65006 29940 65062 29996
rect 65062 29940 65066 29996
rect 65002 29936 65066 29940
rect 65082 29996 65146 30000
rect 65082 29940 65086 29996
rect 65086 29940 65142 29996
rect 65142 29940 65146 29996
rect 65082 29936 65146 29940
rect 65162 29996 65226 30000
rect 65162 29940 65166 29996
rect 65166 29940 65222 29996
rect 65222 29940 65226 29996
rect 65162 29936 65226 29940
rect 70250 29996 70314 30000
rect 70250 29940 70254 29996
rect 70254 29940 70310 29996
rect 70310 29940 70314 29996
rect 70250 29936 70314 29940
rect 70330 29996 70394 30000
rect 70330 29940 70334 29996
rect 70334 29940 70390 29996
rect 70390 29940 70394 29996
rect 70330 29936 70394 29940
rect 70410 29996 70474 30000
rect 70410 29940 70414 29996
rect 70414 29940 70470 29996
rect 70470 29940 70474 29996
rect 70410 29936 70474 29940
rect 70490 29996 70554 30000
rect 70490 29940 70494 29996
rect 70494 29940 70550 29996
rect 70550 29940 70554 29996
rect 70490 29936 70554 29940
rect 75578 29996 75642 30000
rect 75578 29940 75582 29996
rect 75582 29940 75638 29996
rect 75638 29940 75642 29996
rect 75578 29936 75642 29940
rect 75658 29996 75722 30000
rect 75658 29940 75662 29996
rect 75662 29940 75718 29996
rect 75718 29940 75722 29996
rect 75658 29936 75722 29940
rect 75738 29996 75802 30000
rect 75738 29940 75742 29996
rect 75742 29940 75798 29996
rect 75798 29940 75802 29996
rect 75738 29936 75802 29940
rect 75818 29996 75882 30000
rect 75818 29940 75822 29996
rect 75822 29940 75878 29996
rect 75878 29940 75882 29996
rect 75818 29936 75882 29940
rect 80906 29996 80970 30000
rect 80906 29940 80910 29996
rect 80910 29940 80966 29996
rect 80966 29940 80970 29996
rect 80906 29936 80970 29940
rect 80986 29996 81050 30000
rect 80986 29940 80990 29996
rect 80990 29940 81046 29996
rect 81046 29940 81050 29996
rect 80986 29936 81050 29940
rect 81066 29996 81130 30000
rect 81066 29940 81070 29996
rect 81070 29940 81126 29996
rect 81126 29940 81130 29996
rect 81066 29936 81130 29940
rect 81146 29996 81210 30000
rect 81146 29940 81150 29996
rect 81150 29940 81206 29996
rect 81206 29940 81210 29996
rect 81146 29936 81210 29940
rect 86234 29996 86298 30000
rect 86234 29940 86238 29996
rect 86238 29940 86294 29996
rect 86294 29940 86298 29996
rect 86234 29936 86298 29940
rect 86314 29996 86378 30000
rect 86314 29940 86318 29996
rect 86318 29940 86374 29996
rect 86374 29940 86378 29996
rect 86314 29936 86378 29940
rect 86394 29996 86458 30000
rect 86394 29940 86398 29996
rect 86398 29940 86454 29996
rect 86454 29940 86458 29996
rect 86394 29936 86458 29940
rect 86474 29996 86538 30000
rect 86474 29940 86478 29996
rect 86478 29940 86534 29996
rect 86534 29940 86538 29996
rect 86474 29936 86538 29940
rect 91562 29996 91626 30000
rect 91562 29940 91566 29996
rect 91566 29940 91622 29996
rect 91622 29940 91626 29996
rect 91562 29936 91626 29940
rect 91642 29996 91706 30000
rect 91642 29940 91646 29996
rect 91646 29940 91702 29996
rect 91702 29940 91706 29996
rect 91642 29936 91706 29940
rect 91722 29996 91786 30000
rect 91722 29940 91726 29996
rect 91726 29940 91782 29996
rect 91782 29940 91786 29996
rect 91722 29936 91786 29940
rect 91802 29996 91866 30000
rect 91802 29940 91806 29996
rect 91806 29940 91862 29996
rect 91862 29940 91866 29996
rect 91802 29936 91866 29940
rect 3650 29452 3714 29456
rect 3650 29396 3654 29452
rect 3654 29396 3710 29452
rect 3710 29396 3714 29452
rect 3650 29392 3714 29396
rect 3730 29452 3794 29456
rect 3730 29396 3734 29452
rect 3734 29396 3790 29452
rect 3790 29396 3794 29452
rect 3730 29392 3794 29396
rect 3810 29452 3874 29456
rect 3810 29396 3814 29452
rect 3814 29396 3870 29452
rect 3870 29396 3874 29452
rect 3810 29392 3874 29396
rect 3890 29452 3954 29456
rect 3890 29396 3894 29452
rect 3894 29396 3950 29452
rect 3950 29396 3954 29452
rect 3890 29392 3954 29396
rect 8978 29452 9042 29456
rect 8978 29396 8982 29452
rect 8982 29396 9038 29452
rect 9038 29396 9042 29452
rect 8978 29392 9042 29396
rect 9058 29452 9122 29456
rect 9058 29396 9062 29452
rect 9062 29396 9118 29452
rect 9118 29396 9122 29452
rect 9058 29392 9122 29396
rect 9138 29452 9202 29456
rect 9138 29396 9142 29452
rect 9142 29396 9198 29452
rect 9198 29396 9202 29452
rect 9138 29392 9202 29396
rect 9218 29452 9282 29456
rect 9218 29396 9222 29452
rect 9222 29396 9278 29452
rect 9278 29396 9282 29452
rect 9218 29392 9282 29396
rect 14306 29452 14370 29456
rect 14306 29396 14310 29452
rect 14310 29396 14366 29452
rect 14366 29396 14370 29452
rect 14306 29392 14370 29396
rect 14386 29452 14450 29456
rect 14386 29396 14390 29452
rect 14390 29396 14446 29452
rect 14446 29396 14450 29452
rect 14386 29392 14450 29396
rect 14466 29452 14530 29456
rect 14466 29396 14470 29452
rect 14470 29396 14526 29452
rect 14526 29396 14530 29452
rect 14466 29392 14530 29396
rect 14546 29452 14610 29456
rect 14546 29396 14550 29452
rect 14550 29396 14606 29452
rect 14606 29396 14610 29452
rect 14546 29392 14610 29396
rect 19634 29452 19698 29456
rect 19634 29396 19638 29452
rect 19638 29396 19694 29452
rect 19694 29396 19698 29452
rect 19634 29392 19698 29396
rect 19714 29452 19778 29456
rect 19714 29396 19718 29452
rect 19718 29396 19774 29452
rect 19774 29396 19778 29452
rect 19714 29392 19778 29396
rect 19794 29452 19858 29456
rect 19794 29396 19798 29452
rect 19798 29396 19854 29452
rect 19854 29396 19858 29452
rect 19794 29392 19858 29396
rect 19874 29452 19938 29456
rect 19874 29396 19878 29452
rect 19878 29396 19934 29452
rect 19934 29396 19938 29452
rect 19874 29392 19938 29396
rect 24962 29452 25026 29456
rect 24962 29396 24966 29452
rect 24966 29396 25022 29452
rect 25022 29396 25026 29452
rect 24962 29392 25026 29396
rect 25042 29452 25106 29456
rect 25042 29396 25046 29452
rect 25046 29396 25102 29452
rect 25102 29396 25106 29452
rect 25042 29392 25106 29396
rect 25122 29452 25186 29456
rect 25122 29396 25126 29452
rect 25126 29396 25182 29452
rect 25182 29396 25186 29452
rect 25122 29392 25186 29396
rect 25202 29452 25266 29456
rect 25202 29396 25206 29452
rect 25206 29396 25262 29452
rect 25262 29396 25266 29452
rect 25202 29392 25266 29396
rect 30290 29452 30354 29456
rect 30290 29396 30294 29452
rect 30294 29396 30350 29452
rect 30350 29396 30354 29452
rect 30290 29392 30354 29396
rect 30370 29452 30434 29456
rect 30370 29396 30374 29452
rect 30374 29396 30430 29452
rect 30430 29396 30434 29452
rect 30370 29392 30434 29396
rect 30450 29452 30514 29456
rect 30450 29396 30454 29452
rect 30454 29396 30510 29452
rect 30510 29396 30514 29452
rect 30450 29392 30514 29396
rect 30530 29452 30594 29456
rect 30530 29396 30534 29452
rect 30534 29396 30590 29452
rect 30590 29396 30594 29452
rect 30530 29392 30594 29396
rect 35618 29452 35682 29456
rect 35618 29396 35622 29452
rect 35622 29396 35678 29452
rect 35678 29396 35682 29452
rect 35618 29392 35682 29396
rect 35698 29452 35762 29456
rect 35698 29396 35702 29452
rect 35702 29396 35758 29452
rect 35758 29396 35762 29452
rect 35698 29392 35762 29396
rect 35778 29452 35842 29456
rect 35778 29396 35782 29452
rect 35782 29396 35838 29452
rect 35838 29396 35842 29452
rect 35778 29392 35842 29396
rect 35858 29452 35922 29456
rect 35858 29396 35862 29452
rect 35862 29396 35918 29452
rect 35918 29396 35922 29452
rect 35858 29392 35922 29396
rect 40946 29452 41010 29456
rect 40946 29396 40950 29452
rect 40950 29396 41006 29452
rect 41006 29396 41010 29452
rect 40946 29392 41010 29396
rect 41026 29452 41090 29456
rect 41026 29396 41030 29452
rect 41030 29396 41086 29452
rect 41086 29396 41090 29452
rect 41026 29392 41090 29396
rect 41106 29452 41170 29456
rect 41106 29396 41110 29452
rect 41110 29396 41166 29452
rect 41166 29396 41170 29452
rect 41106 29392 41170 29396
rect 41186 29452 41250 29456
rect 41186 29396 41190 29452
rect 41190 29396 41246 29452
rect 41246 29396 41250 29452
rect 41186 29392 41250 29396
rect 46274 29452 46338 29456
rect 46274 29396 46278 29452
rect 46278 29396 46334 29452
rect 46334 29396 46338 29452
rect 46274 29392 46338 29396
rect 46354 29452 46418 29456
rect 46354 29396 46358 29452
rect 46358 29396 46414 29452
rect 46414 29396 46418 29452
rect 46354 29392 46418 29396
rect 46434 29452 46498 29456
rect 46434 29396 46438 29452
rect 46438 29396 46494 29452
rect 46494 29396 46498 29452
rect 46434 29392 46498 29396
rect 46514 29452 46578 29456
rect 46514 29396 46518 29452
rect 46518 29396 46574 29452
rect 46574 29396 46578 29452
rect 46514 29392 46578 29396
rect 51602 29452 51666 29456
rect 51602 29396 51606 29452
rect 51606 29396 51662 29452
rect 51662 29396 51666 29452
rect 51602 29392 51666 29396
rect 51682 29452 51746 29456
rect 51682 29396 51686 29452
rect 51686 29396 51742 29452
rect 51742 29396 51746 29452
rect 51682 29392 51746 29396
rect 51762 29452 51826 29456
rect 51762 29396 51766 29452
rect 51766 29396 51822 29452
rect 51822 29396 51826 29452
rect 51762 29392 51826 29396
rect 51842 29452 51906 29456
rect 51842 29396 51846 29452
rect 51846 29396 51902 29452
rect 51902 29396 51906 29452
rect 51842 29392 51906 29396
rect 56930 29452 56994 29456
rect 56930 29396 56934 29452
rect 56934 29396 56990 29452
rect 56990 29396 56994 29452
rect 56930 29392 56994 29396
rect 57010 29452 57074 29456
rect 57010 29396 57014 29452
rect 57014 29396 57070 29452
rect 57070 29396 57074 29452
rect 57010 29392 57074 29396
rect 57090 29452 57154 29456
rect 57090 29396 57094 29452
rect 57094 29396 57150 29452
rect 57150 29396 57154 29452
rect 57090 29392 57154 29396
rect 57170 29452 57234 29456
rect 57170 29396 57174 29452
rect 57174 29396 57230 29452
rect 57230 29396 57234 29452
rect 57170 29392 57234 29396
rect 62258 29452 62322 29456
rect 62258 29396 62262 29452
rect 62262 29396 62318 29452
rect 62318 29396 62322 29452
rect 62258 29392 62322 29396
rect 62338 29452 62402 29456
rect 62338 29396 62342 29452
rect 62342 29396 62398 29452
rect 62398 29396 62402 29452
rect 62338 29392 62402 29396
rect 62418 29452 62482 29456
rect 62418 29396 62422 29452
rect 62422 29396 62478 29452
rect 62478 29396 62482 29452
rect 62418 29392 62482 29396
rect 62498 29452 62562 29456
rect 62498 29396 62502 29452
rect 62502 29396 62558 29452
rect 62558 29396 62562 29452
rect 62498 29392 62562 29396
rect 67586 29452 67650 29456
rect 67586 29396 67590 29452
rect 67590 29396 67646 29452
rect 67646 29396 67650 29452
rect 67586 29392 67650 29396
rect 67666 29452 67730 29456
rect 67666 29396 67670 29452
rect 67670 29396 67726 29452
rect 67726 29396 67730 29452
rect 67666 29392 67730 29396
rect 67746 29452 67810 29456
rect 67746 29396 67750 29452
rect 67750 29396 67806 29452
rect 67806 29396 67810 29452
rect 67746 29392 67810 29396
rect 67826 29452 67890 29456
rect 67826 29396 67830 29452
rect 67830 29396 67886 29452
rect 67886 29396 67890 29452
rect 67826 29392 67890 29396
rect 72914 29452 72978 29456
rect 72914 29396 72918 29452
rect 72918 29396 72974 29452
rect 72974 29396 72978 29452
rect 72914 29392 72978 29396
rect 72994 29452 73058 29456
rect 72994 29396 72998 29452
rect 72998 29396 73054 29452
rect 73054 29396 73058 29452
rect 72994 29392 73058 29396
rect 73074 29452 73138 29456
rect 73074 29396 73078 29452
rect 73078 29396 73134 29452
rect 73134 29396 73138 29452
rect 73074 29392 73138 29396
rect 73154 29452 73218 29456
rect 73154 29396 73158 29452
rect 73158 29396 73214 29452
rect 73214 29396 73218 29452
rect 73154 29392 73218 29396
rect 78242 29452 78306 29456
rect 78242 29396 78246 29452
rect 78246 29396 78302 29452
rect 78302 29396 78306 29452
rect 78242 29392 78306 29396
rect 78322 29452 78386 29456
rect 78322 29396 78326 29452
rect 78326 29396 78382 29452
rect 78382 29396 78386 29452
rect 78322 29392 78386 29396
rect 78402 29452 78466 29456
rect 78402 29396 78406 29452
rect 78406 29396 78462 29452
rect 78462 29396 78466 29452
rect 78402 29392 78466 29396
rect 78482 29452 78546 29456
rect 78482 29396 78486 29452
rect 78486 29396 78542 29452
rect 78542 29396 78546 29452
rect 78482 29392 78546 29396
rect 83570 29452 83634 29456
rect 83570 29396 83574 29452
rect 83574 29396 83630 29452
rect 83630 29396 83634 29452
rect 83570 29392 83634 29396
rect 83650 29452 83714 29456
rect 83650 29396 83654 29452
rect 83654 29396 83710 29452
rect 83710 29396 83714 29452
rect 83650 29392 83714 29396
rect 83730 29452 83794 29456
rect 83730 29396 83734 29452
rect 83734 29396 83790 29452
rect 83790 29396 83794 29452
rect 83730 29392 83794 29396
rect 83810 29452 83874 29456
rect 83810 29396 83814 29452
rect 83814 29396 83870 29452
rect 83870 29396 83874 29452
rect 83810 29392 83874 29396
rect 88898 29452 88962 29456
rect 88898 29396 88902 29452
rect 88902 29396 88958 29452
rect 88958 29396 88962 29452
rect 88898 29392 88962 29396
rect 88978 29452 89042 29456
rect 88978 29396 88982 29452
rect 88982 29396 89038 29452
rect 89038 29396 89042 29452
rect 88978 29392 89042 29396
rect 89058 29452 89122 29456
rect 89058 29396 89062 29452
rect 89062 29396 89118 29452
rect 89118 29396 89122 29452
rect 89058 29392 89122 29396
rect 89138 29452 89202 29456
rect 89138 29396 89142 29452
rect 89142 29396 89198 29452
rect 89198 29396 89202 29452
rect 89138 29392 89202 29396
rect 6314 28908 6378 28912
rect 6314 28852 6318 28908
rect 6318 28852 6374 28908
rect 6374 28852 6378 28908
rect 6314 28848 6378 28852
rect 6394 28908 6458 28912
rect 6394 28852 6398 28908
rect 6398 28852 6454 28908
rect 6454 28852 6458 28908
rect 6394 28848 6458 28852
rect 6474 28908 6538 28912
rect 6474 28852 6478 28908
rect 6478 28852 6534 28908
rect 6534 28852 6538 28908
rect 6474 28848 6538 28852
rect 6554 28908 6618 28912
rect 6554 28852 6558 28908
rect 6558 28852 6614 28908
rect 6614 28852 6618 28908
rect 6554 28848 6618 28852
rect 11642 28908 11706 28912
rect 11642 28852 11646 28908
rect 11646 28852 11702 28908
rect 11702 28852 11706 28908
rect 11642 28848 11706 28852
rect 11722 28908 11786 28912
rect 11722 28852 11726 28908
rect 11726 28852 11782 28908
rect 11782 28852 11786 28908
rect 11722 28848 11786 28852
rect 11802 28908 11866 28912
rect 11802 28852 11806 28908
rect 11806 28852 11862 28908
rect 11862 28852 11866 28908
rect 11802 28848 11866 28852
rect 11882 28908 11946 28912
rect 11882 28852 11886 28908
rect 11886 28852 11942 28908
rect 11942 28852 11946 28908
rect 11882 28848 11946 28852
rect 16970 28908 17034 28912
rect 16970 28852 16974 28908
rect 16974 28852 17030 28908
rect 17030 28852 17034 28908
rect 16970 28848 17034 28852
rect 17050 28908 17114 28912
rect 17050 28852 17054 28908
rect 17054 28852 17110 28908
rect 17110 28852 17114 28908
rect 17050 28848 17114 28852
rect 17130 28908 17194 28912
rect 17130 28852 17134 28908
rect 17134 28852 17190 28908
rect 17190 28852 17194 28908
rect 17130 28848 17194 28852
rect 17210 28908 17274 28912
rect 17210 28852 17214 28908
rect 17214 28852 17270 28908
rect 17270 28852 17274 28908
rect 17210 28848 17274 28852
rect 22298 28908 22362 28912
rect 22298 28852 22302 28908
rect 22302 28852 22358 28908
rect 22358 28852 22362 28908
rect 22298 28848 22362 28852
rect 22378 28908 22442 28912
rect 22378 28852 22382 28908
rect 22382 28852 22438 28908
rect 22438 28852 22442 28908
rect 22378 28848 22442 28852
rect 22458 28908 22522 28912
rect 22458 28852 22462 28908
rect 22462 28852 22518 28908
rect 22518 28852 22522 28908
rect 22458 28848 22522 28852
rect 22538 28908 22602 28912
rect 22538 28852 22542 28908
rect 22542 28852 22598 28908
rect 22598 28852 22602 28908
rect 22538 28848 22602 28852
rect 27626 28908 27690 28912
rect 27626 28852 27630 28908
rect 27630 28852 27686 28908
rect 27686 28852 27690 28908
rect 27626 28848 27690 28852
rect 27706 28908 27770 28912
rect 27706 28852 27710 28908
rect 27710 28852 27766 28908
rect 27766 28852 27770 28908
rect 27706 28848 27770 28852
rect 27786 28908 27850 28912
rect 27786 28852 27790 28908
rect 27790 28852 27846 28908
rect 27846 28852 27850 28908
rect 27786 28848 27850 28852
rect 27866 28908 27930 28912
rect 27866 28852 27870 28908
rect 27870 28852 27926 28908
rect 27926 28852 27930 28908
rect 27866 28848 27930 28852
rect 32954 28908 33018 28912
rect 32954 28852 32958 28908
rect 32958 28852 33014 28908
rect 33014 28852 33018 28908
rect 32954 28848 33018 28852
rect 33034 28908 33098 28912
rect 33034 28852 33038 28908
rect 33038 28852 33094 28908
rect 33094 28852 33098 28908
rect 33034 28848 33098 28852
rect 33114 28908 33178 28912
rect 33114 28852 33118 28908
rect 33118 28852 33174 28908
rect 33174 28852 33178 28908
rect 33114 28848 33178 28852
rect 33194 28908 33258 28912
rect 33194 28852 33198 28908
rect 33198 28852 33254 28908
rect 33254 28852 33258 28908
rect 33194 28848 33258 28852
rect 38282 28908 38346 28912
rect 38282 28852 38286 28908
rect 38286 28852 38342 28908
rect 38342 28852 38346 28908
rect 38282 28848 38346 28852
rect 38362 28908 38426 28912
rect 38362 28852 38366 28908
rect 38366 28852 38422 28908
rect 38422 28852 38426 28908
rect 38362 28848 38426 28852
rect 38442 28908 38506 28912
rect 38442 28852 38446 28908
rect 38446 28852 38502 28908
rect 38502 28852 38506 28908
rect 38442 28848 38506 28852
rect 38522 28908 38586 28912
rect 38522 28852 38526 28908
rect 38526 28852 38582 28908
rect 38582 28852 38586 28908
rect 38522 28848 38586 28852
rect 43610 28908 43674 28912
rect 43610 28852 43614 28908
rect 43614 28852 43670 28908
rect 43670 28852 43674 28908
rect 43610 28848 43674 28852
rect 43690 28908 43754 28912
rect 43690 28852 43694 28908
rect 43694 28852 43750 28908
rect 43750 28852 43754 28908
rect 43690 28848 43754 28852
rect 43770 28908 43834 28912
rect 43770 28852 43774 28908
rect 43774 28852 43830 28908
rect 43830 28852 43834 28908
rect 43770 28848 43834 28852
rect 43850 28908 43914 28912
rect 43850 28852 43854 28908
rect 43854 28852 43910 28908
rect 43910 28852 43914 28908
rect 43850 28848 43914 28852
rect 48938 28908 49002 28912
rect 48938 28852 48942 28908
rect 48942 28852 48998 28908
rect 48998 28852 49002 28908
rect 48938 28848 49002 28852
rect 49018 28908 49082 28912
rect 49018 28852 49022 28908
rect 49022 28852 49078 28908
rect 49078 28852 49082 28908
rect 49018 28848 49082 28852
rect 49098 28908 49162 28912
rect 49098 28852 49102 28908
rect 49102 28852 49158 28908
rect 49158 28852 49162 28908
rect 49098 28848 49162 28852
rect 49178 28908 49242 28912
rect 49178 28852 49182 28908
rect 49182 28852 49238 28908
rect 49238 28852 49242 28908
rect 49178 28848 49242 28852
rect 54266 28908 54330 28912
rect 54266 28852 54270 28908
rect 54270 28852 54326 28908
rect 54326 28852 54330 28908
rect 54266 28848 54330 28852
rect 54346 28908 54410 28912
rect 54346 28852 54350 28908
rect 54350 28852 54406 28908
rect 54406 28852 54410 28908
rect 54346 28848 54410 28852
rect 54426 28908 54490 28912
rect 54426 28852 54430 28908
rect 54430 28852 54486 28908
rect 54486 28852 54490 28908
rect 54426 28848 54490 28852
rect 54506 28908 54570 28912
rect 54506 28852 54510 28908
rect 54510 28852 54566 28908
rect 54566 28852 54570 28908
rect 54506 28848 54570 28852
rect 59594 28908 59658 28912
rect 59594 28852 59598 28908
rect 59598 28852 59654 28908
rect 59654 28852 59658 28908
rect 59594 28848 59658 28852
rect 59674 28908 59738 28912
rect 59674 28852 59678 28908
rect 59678 28852 59734 28908
rect 59734 28852 59738 28908
rect 59674 28848 59738 28852
rect 59754 28908 59818 28912
rect 59754 28852 59758 28908
rect 59758 28852 59814 28908
rect 59814 28852 59818 28908
rect 59754 28848 59818 28852
rect 59834 28908 59898 28912
rect 59834 28852 59838 28908
rect 59838 28852 59894 28908
rect 59894 28852 59898 28908
rect 59834 28848 59898 28852
rect 64922 28908 64986 28912
rect 64922 28852 64926 28908
rect 64926 28852 64982 28908
rect 64982 28852 64986 28908
rect 64922 28848 64986 28852
rect 65002 28908 65066 28912
rect 65002 28852 65006 28908
rect 65006 28852 65062 28908
rect 65062 28852 65066 28908
rect 65002 28848 65066 28852
rect 65082 28908 65146 28912
rect 65082 28852 65086 28908
rect 65086 28852 65142 28908
rect 65142 28852 65146 28908
rect 65082 28848 65146 28852
rect 65162 28908 65226 28912
rect 65162 28852 65166 28908
rect 65166 28852 65222 28908
rect 65222 28852 65226 28908
rect 65162 28848 65226 28852
rect 70250 28908 70314 28912
rect 70250 28852 70254 28908
rect 70254 28852 70310 28908
rect 70310 28852 70314 28908
rect 70250 28848 70314 28852
rect 70330 28908 70394 28912
rect 70330 28852 70334 28908
rect 70334 28852 70390 28908
rect 70390 28852 70394 28908
rect 70330 28848 70394 28852
rect 70410 28908 70474 28912
rect 70410 28852 70414 28908
rect 70414 28852 70470 28908
rect 70470 28852 70474 28908
rect 70410 28848 70474 28852
rect 70490 28908 70554 28912
rect 70490 28852 70494 28908
rect 70494 28852 70550 28908
rect 70550 28852 70554 28908
rect 70490 28848 70554 28852
rect 75578 28908 75642 28912
rect 75578 28852 75582 28908
rect 75582 28852 75638 28908
rect 75638 28852 75642 28908
rect 75578 28848 75642 28852
rect 75658 28908 75722 28912
rect 75658 28852 75662 28908
rect 75662 28852 75718 28908
rect 75718 28852 75722 28908
rect 75658 28848 75722 28852
rect 75738 28908 75802 28912
rect 75738 28852 75742 28908
rect 75742 28852 75798 28908
rect 75798 28852 75802 28908
rect 75738 28848 75802 28852
rect 75818 28908 75882 28912
rect 75818 28852 75822 28908
rect 75822 28852 75878 28908
rect 75878 28852 75882 28908
rect 75818 28848 75882 28852
rect 80906 28908 80970 28912
rect 80906 28852 80910 28908
rect 80910 28852 80966 28908
rect 80966 28852 80970 28908
rect 80906 28848 80970 28852
rect 80986 28908 81050 28912
rect 80986 28852 80990 28908
rect 80990 28852 81046 28908
rect 81046 28852 81050 28908
rect 80986 28848 81050 28852
rect 81066 28908 81130 28912
rect 81066 28852 81070 28908
rect 81070 28852 81126 28908
rect 81126 28852 81130 28908
rect 81066 28848 81130 28852
rect 81146 28908 81210 28912
rect 81146 28852 81150 28908
rect 81150 28852 81206 28908
rect 81206 28852 81210 28908
rect 81146 28848 81210 28852
rect 86234 28908 86298 28912
rect 86234 28852 86238 28908
rect 86238 28852 86294 28908
rect 86294 28852 86298 28908
rect 86234 28848 86298 28852
rect 86314 28908 86378 28912
rect 86314 28852 86318 28908
rect 86318 28852 86374 28908
rect 86374 28852 86378 28908
rect 86314 28848 86378 28852
rect 86394 28908 86458 28912
rect 86394 28852 86398 28908
rect 86398 28852 86454 28908
rect 86454 28852 86458 28908
rect 86394 28848 86458 28852
rect 86474 28908 86538 28912
rect 86474 28852 86478 28908
rect 86478 28852 86534 28908
rect 86534 28852 86538 28908
rect 86474 28848 86538 28852
rect 91562 28908 91626 28912
rect 91562 28852 91566 28908
rect 91566 28852 91622 28908
rect 91622 28852 91626 28908
rect 91562 28848 91626 28852
rect 91642 28908 91706 28912
rect 91642 28852 91646 28908
rect 91646 28852 91702 28908
rect 91702 28852 91706 28908
rect 91642 28848 91706 28852
rect 91722 28908 91786 28912
rect 91722 28852 91726 28908
rect 91726 28852 91782 28908
rect 91782 28852 91786 28908
rect 91722 28848 91786 28852
rect 91802 28908 91866 28912
rect 91802 28852 91806 28908
rect 91806 28852 91862 28908
rect 91862 28852 91866 28908
rect 91802 28848 91866 28852
rect 3650 28364 3714 28368
rect 3650 28308 3654 28364
rect 3654 28308 3710 28364
rect 3710 28308 3714 28364
rect 3650 28304 3714 28308
rect 3730 28364 3794 28368
rect 3730 28308 3734 28364
rect 3734 28308 3790 28364
rect 3790 28308 3794 28364
rect 3730 28304 3794 28308
rect 3810 28364 3874 28368
rect 3810 28308 3814 28364
rect 3814 28308 3870 28364
rect 3870 28308 3874 28364
rect 3810 28304 3874 28308
rect 3890 28364 3954 28368
rect 3890 28308 3894 28364
rect 3894 28308 3950 28364
rect 3950 28308 3954 28364
rect 3890 28304 3954 28308
rect 8978 28364 9042 28368
rect 8978 28308 8982 28364
rect 8982 28308 9038 28364
rect 9038 28308 9042 28364
rect 8978 28304 9042 28308
rect 9058 28364 9122 28368
rect 9058 28308 9062 28364
rect 9062 28308 9118 28364
rect 9118 28308 9122 28364
rect 9058 28304 9122 28308
rect 9138 28364 9202 28368
rect 9138 28308 9142 28364
rect 9142 28308 9198 28364
rect 9198 28308 9202 28364
rect 9138 28304 9202 28308
rect 9218 28364 9282 28368
rect 9218 28308 9222 28364
rect 9222 28308 9278 28364
rect 9278 28308 9282 28364
rect 9218 28304 9282 28308
rect 14306 28364 14370 28368
rect 14306 28308 14310 28364
rect 14310 28308 14366 28364
rect 14366 28308 14370 28364
rect 14306 28304 14370 28308
rect 14386 28364 14450 28368
rect 14386 28308 14390 28364
rect 14390 28308 14446 28364
rect 14446 28308 14450 28364
rect 14386 28304 14450 28308
rect 14466 28364 14530 28368
rect 14466 28308 14470 28364
rect 14470 28308 14526 28364
rect 14526 28308 14530 28364
rect 14466 28304 14530 28308
rect 14546 28364 14610 28368
rect 14546 28308 14550 28364
rect 14550 28308 14606 28364
rect 14606 28308 14610 28364
rect 14546 28304 14610 28308
rect 19634 28364 19698 28368
rect 19634 28308 19638 28364
rect 19638 28308 19694 28364
rect 19694 28308 19698 28364
rect 19634 28304 19698 28308
rect 19714 28364 19778 28368
rect 19714 28308 19718 28364
rect 19718 28308 19774 28364
rect 19774 28308 19778 28364
rect 19714 28304 19778 28308
rect 19794 28364 19858 28368
rect 19794 28308 19798 28364
rect 19798 28308 19854 28364
rect 19854 28308 19858 28364
rect 19794 28304 19858 28308
rect 19874 28364 19938 28368
rect 19874 28308 19878 28364
rect 19878 28308 19934 28364
rect 19934 28308 19938 28364
rect 19874 28304 19938 28308
rect 24962 28364 25026 28368
rect 24962 28308 24966 28364
rect 24966 28308 25022 28364
rect 25022 28308 25026 28364
rect 24962 28304 25026 28308
rect 25042 28364 25106 28368
rect 25042 28308 25046 28364
rect 25046 28308 25102 28364
rect 25102 28308 25106 28364
rect 25042 28304 25106 28308
rect 25122 28364 25186 28368
rect 25122 28308 25126 28364
rect 25126 28308 25182 28364
rect 25182 28308 25186 28364
rect 25122 28304 25186 28308
rect 25202 28364 25266 28368
rect 25202 28308 25206 28364
rect 25206 28308 25262 28364
rect 25262 28308 25266 28364
rect 25202 28304 25266 28308
rect 30290 28364 30354 28368
rect 30290 28308 30294 28364
rect 30294 28308 30350 28364
rect 30350 28308 30354 28364
rect 30290 28304 30354 28308
rect 30370 28364 30434 28368
rect 30370 28308 30374 28364
rect 30374 28308 30430 28364
rect 30430 28308 30434 28364
rect 30370 28304 30434 28308
rect 30450 28364 30514 28368
rect 30450 28308 30454 28364
rect 30454 28308 30510 28364
rect 30510 28308 30514 28364
rect 30450 28304 30514 28308
rect 30530 28364 30594 28368
rect 30530 28308 30534 28364
rect 30534 28308 30590 28364
rect 30590 28308 30594 28364
rect 30530 28304 30594 28308
rect 35618 28364 35682 28368
rect 35618 28308 35622 28364
rect 35622 28308 35678 28364
rect 35678 28308 35682 28364
rect 35618 28304 35682 28308
rect 35698 28364 35762 28368
rect 35698 28308 35702 28364
rect 35702 28308 35758 28364
rect 35758 28308 35762 28364
rect 35698 28304 35762 28308
rect 35778 28364 35842 28368
rect 35778 28308 35782 28364
rect 35782 28308 35838 28364
rect 35838 28308 35842 28364
rect 35778 28304 35842 28308
rect 35858 28364 35922 28368
rect 35858 28308 35862 28364
rect 35862 28308 35918 28364
rect 35918 28308 35922 28364
rect 35858 28304 35922 28308
rect 40946 28364 41010 28368
rect 40946 28308 40950 28364
rect 40950 28308 41006 28364
rect 41006 28308 41010 28364
rect 40946 28304 41010 28308
rect 41026 28364 41090 28368
rect 41026 28308 41030 28364
rect 41030 28308 41086 28364
rect 41086 28308 41090 28364
rect 41026 28304 41090 28308
rect 41106 28364 41170 28368
rect 41106 28308 41110 28364
rect 41110 28308 41166 28364
rect 41166 28308 41170 28364
rect 41106 28304 41170 28308
rect 41186 28364 41250 28368
rect 41186 28308 41190 28364
rect 41190 28308 41246 28364
rect 41246 28308 41250 28364
rect 41186 28304 41250 28308
rect 46274 28364 46338 28368
rect 46274 28308 46278 28364
rect 46278 28308 46334 28364
rect 46334 28308 46338 28364
rect 46274 28304 46338 28308
rect 46354 28364 46418 28368
rect 46354 28308 46358 28364
rect 46358 28308 46414 28364
rect 46414 28308 46418 28364
rect 46354 28304 46418 28308
rect 46434 28364 46498 28368
rect 46434 28308 46438 28364
rect 46438 28308 46494 28364
rect 46494 28308 46498 28364
rect 46434 28304 46498 28308
rect 46514 28364 46578 28368
rect 46514 28308 46518 28364
rect 46518 28308 46574 28364
rect 46574 28308 46578 28364
rect 46514 28304 46578 28308
rect 51602 28364 51666 28368
rect 51602 28308 51606 28364
rect 51606 28308 51662 28364
rect 51662 28308 51666 28364
rect 51602 28304 51666 28308
rect 51682 28364 51746 28368
rect 51682 28308 51686 28364
rect 51686 28308 51742 28364
rect 51742 28308 51746 28364
rect 51682 28304 51746 28308
rect 51762 28364 51826 28368
rect 51762 28308 51766 28364
rect 51766 28308 51822 28364
rect 51822 28308 51826 28364
rect 51762 28304 51826 28308
rect 51842 28364 51906 28368
rect 51842 28308 51846 28364
rect 51846 28308 51902 28364
rect 51902 28308 51906 28364
rect 51842 28304 51906 28308
rect 56930 28364 56994 28368
rect 56930 28308 56934 28364
rect 56934 28308 56990 28364
rect 56990 28308 56994 28364
rect 56930 28304 56994 28308
rect 57010 28364 57074 28368
rect 57010 28308 57014 28364
rect 57014 28308 57070 28364
rect 57070 28308 57074 28364
rect 57010 28304 57074 28308
rect 57090 28364 57154 28368
rect 57090 28308 57094 28364
rect 57094 28308 57150 28364
rect 57150 28308 57154 28364
rect 57090 28304 57154 28308
rect 57170 28364 57234 28368
rect 57170 28308 57174 28364
rect 57174 28308 57230 28364
rect 57230 28308 57234 28364
rect 57170 28304 57234 28308
rect 62258 28364 62322 28368
rect 62258 28308 62262 28364
rect 62262 28308 62318 28364
rect 62318 28308 62322 28364
rect 62258 28304 62322 28308
rect 62338 28364 62402 28368
rect 62338 28308 62342 28364
rect 62342 28308 62398 28364
rect 62398 28308 62402 28364
rect 62338 28304 62402 28308
rect 62418 28364 62482 28368
rect 62418 28308 62422 28364
rect 62422 28308 62478 28364
rect 62478 28308 62482 28364
rect 62418 28304 62482 28308
rect 62498 28364 62562 28368
rect 62498 28308 62502 28364
rect 62502 28308 62558 28364
rect 62558 28308 62562 28364
rect 62498 28304 62562 28308
rect 67586 28364 67650 28368
rect 67586 28308 67590 28364
rect 67590 28308 67646 28364
rect 67646 28308 67650 28364
rect 67586 28304 67650 28308
rect 67666 28364 67730 28368
rect 67666 28308 67670 28364
rect 67670 28308 67726 28364
rect 67726 28308 67730 28364
rect 67666 28304 67730 28308
rect 67746 28364 67810 28368
rect 67746 28308 67750 28364
rect 67750 28308 67806 28364
rect 67806 28308 67810 28364
rect 67746 28304 67810 28308
rect 67826 28364 67890 28368
rect 67826 28308 67830 28364
rect 67830 28308 67886 28364
rect 67886 28308 67890 28364
rect 67826 28304 67890 28308
rect 72914 28364 72978 28368
rect 72914 28308 72918 28364
rect 72918 28308 72974 28364
rect 72974 28308 72978 28364
rect 72914 28304 72978 28308
rect 72994 28364 73058 28368
rect 72994 28308 72998 28364
rect 72998 28308 73054 28364
rect 73054 28308 73058 28364
rect 72994 28304 73058 28308
rect 73074 28364 73138 28368
rect 73074 28308 73078 28364
rect 73078 28308 73134 28364
rect 73134 28308 73138 28364
rect 73074 28304 73138 28308
rect 73154 28364 73218 28368
rect 73154 28308 73158 28364
rect 73158 28308 73214 28364
rect 73214 28308 73218 28364
rect 73154 28304 73218 28308
rect 78242 28364 78306 28368
rect 78242 28308 78246 28364
rect 78246 28308 78302 28364
rect 78302 28308 78306 28364
rect 78242 28304 78306 28308
rect 78322 28364 78386 28368
rect 78322 28308 78326 28364
rect 78326 28308 78382 28364
rect 78382 28308 78386 28364
rect 78322 28304 78386 28308
rect 78402 28364 78466 28368
rect 78402 28308 78406 28364
rect 78406 28308 78462 28364
rect 78462 28308 78466 28364
rect 78402 28304 78466 28308
rect 78482 28364 78546 28368
rect 78482 28308 78486 28364
rect 78486 28308 78542 28364
rect 78542 28308 78546 28364
rect 78482 28304 78546 28308
rect 83570 28364 83634 28368
rect 83570 28308 83574 28364
rect 83574 28308 83630 28364
rect 83630 28308 83634 28364
rect 83570 28304 83634 28308
rect 83650 28364 83714 28368
rect 83650 28308 83654 28364
rect 83654 28308 83710 28364
rect 83710 28308 83714 28364
rect 83650 28304 83714 28308
rect 83730 28364 83794 28368
rect 83730 28308 83734 28364
rect 83734 28308 83790 28364
rect 83790 28308 83794 28364
rect 83730 28304 83794 28308
rect 83810 28364 83874 28368
rect 83810 28308 83814 28364
rect 83814 28308 83870 28364
rect 83870 28308 83874 28364
rect 83810 28304 83874 28308
rect 88898 28364 88962 28368
rect 88898 28308 88902 28364
rect 88902 28308 88958 28364
rect 88958 28308 88962 28364
rect 88898 28304 88962 28308
rect 88978 28364 89042 28368
rect 88978 28308 88982 28364
rect 88982 28308 89038 28364
rect 89038 28308 89042 28364
rect 88978 28304 89042 28308
rect 89058 28364 89122 28368
rect 89058 28308 89062 28364
rect 89062 28308 89118 28364
rect 89118 28308 89122 28364
rect 89058 28304 89122 28308
rect 89138 28364 89202 28368
rect 89138 28308 89142 28364
rect 89142 28308 89198 28364
rect 89198 28308 89202 28364
rect 89138 28304 89202 28308
rect 6314 27820 6378 27824
rect 6314 27764 6318 27820
rect 6318 27764 6374 27820
rect 6374 27764 6378 27820
rect 6314 27760 6378 27764
rect 6394 27820 6458 27824
rect 6394 27764 6398 27820
rect 6398 27764 6454 27820
rect 6454 27764 6458 27820
rect 6394 27760 6458 27764
rect 6474 27820 6538 27824
rect 6474 27764 6478 27820
rect 6478 27764 6534 27820
rect 6534 27764 6538 27820
rect 6474 27760 6538 27764
rect 6554 27820 6618 27824
rect 6554 27764 6558 27820
rect 6558 27764 6614 27820
rect 6614 27764 6618 27820
rect 6554 27760 6618 27764
rect 11642 27820 11706 27824
rect 11642 27764 11646 27820
rect 11646 27764 11702 27820
rect 11702 27764 11706 27820
rect 11642 27760 11706 27764
rect 11722 27820 11786 27824
rect 11722 27764 11726 27820
rect 11726 27764 11782 27820
rect 11782 27764 11786 27820
rect 11722 27760 11786 27764
rect 11802 27820 11866 27824
rect 11802 27764 11806 27820
rect 11806 27764 11862 27820
rect 11862 27764 11866 27820
rect 11802 27760 11866 27764
rect 11882 27820 11946 27824
rect 11882 27764 11886 27820
rect 11886 27764 11942 27820
rect 11942 27764 11946 27820
rect 11882 27760 11946 27764
rect 16970 27820 17034 27824
rect 16970 27764 16974 27820
rect 16974 27764 17030 27820
rect 17030 27764 17034 27820
rect 16970 27760 17034 27764
rect 17050 27820 17114 27824
rect 17050 27764 17054 27820
rect 17054 27764 17110 27820
rect 17110 27764 17114 27820
rect 17050 27760 17114 27764
rect 17130 27820 17194 27824
rect 17130 27764 17134 27820
rect 17134 27764 17190 27820
rect 17190 27764 17194 27820
rect 17130 27760 17194 27764
rect 17210 27820 17274 27824
rect 17210 27764 17214 27820
rect 17214 27764 17270 27820
rect 17270 27764 17274 27820
rect 17210 27760 17274 27764
rect 22298 27820 22362 27824
rect 22298 27764 22302 27820
rect 22302 27764 22358 27820
rect 22358 27764 22362 27820
rect 22298 27760 22362 27764
rect 22378 27820 22442 27824
rect 22378 27764 22382 27820
rect 22382 27764 22438 27820
rect 22438 27764 22442 27820
rect 22378 27760 22442 27764
rect 22458 27820 22522 27824
rect 22458 27764 22462 27820
rect 22462 27764 22518 27820
rect 22518 27764 22522 27820
rect 22458 27760 22522 27764
rect 22538 27820 22602 27824
rect 22538 27764 22542 27820
rect 22542 27764 22598 27820
rect 22598 27764 22602 27820
rect 22538 27760 22602 27764
rect 27626 27820 27690 27824
rect 27626 27764 27630 27820
rect 27630 27764 27686 27820
rect 27686 27764 27690 27820
rect 27626 27760 27690 27764
rect 27706 27820 27770 27824
rect 27706 27764 27710 27820
rect 27710 27764 27766 27820
rect 27766 27764 27770 27820
rect 27706 27760 27770 27764
rect 27786 27820 27850 27824
rect 27786 27764 27790 27820
rect 27790 27764 27846 27820
rect 27846 27764 27850 27820
rect 27786 27760 27850 27764
rect 27866 27820 27930 27824
rect 27866 27764 27870 27820
rect 27870 27764 27926 27820
rect 27926 27764 27930 27820
rect 27866 27760 27930 27764
rect 32954 27820 33018 27824
rect 32954 27764 32958 27820
rect 32958 27764 33014 27820
rect 33014 27764 33018 27820
rect 32954 27760 33018 27764
rect 33034 27820 33098 27824
rect 33034 27764 33038 27820
rect 33038 27764 33094 27820
rect 33094 27764 33098 27820
rect 33034 27760 33098 27764
rect 33114 27820 33178 27824
rect 33114 27764 33118 27820
rect 33118 27764 33174 27820
rect 33174 27764 33178 27820
rect 33114 27760 33178 27764
rect 33194 27820 33258 27824
rect 33194 27764 33198 27820
rect 33198 27764 33254 27820
rect 33254 27764 33258 27820
rect 33194 27760 33258 27764
rect 38282 27820 38346 27824
rect 38282 27764 38286 27820
rect 38286 27764 38342 27820
rect 38342 27764 38346 27820
rect 38282 27760 38346 27764
rect 38362 27820 38426 27824
rect 38362 27764 38366 27820
rect 38366 27764 38422 27820
rect 38422 27764 38426 27820
rect 38362 27760 38426 27764
rect 38442 27820 38506 27824
rect 38442 27764 38446 27820
rect 38446 27764 38502 27820
rect 38502 27764 38506 27820
rect 38442 27760 38506 27764
rect 38522 27820 38586 27824
rect 38522 27764 38526 27820
rect 38526 27764 38582 27820
rect 38582 27764 38586 27820
rect 38522 27760 38586 27764
rect 43610 27820 43674 27824
rect 43610 27764 43614 27820
rect 43614 27764 43670 27820
rect 43670 27764 43674 27820
rect 43610 27760 43674 27764
rect 43690 27820 43754 27824
rect 43690 27764 43694 27820
rect 43694 27764 43750 27820
rect 43750 27764 43754 27820
rect 43690 27760 43754 27764
rect 43770 27820 43834 27824
rect 43770 27764 43774 27820
rect 43774 27764 43830 27820
rect 43830 27764 43834 27820
rect 43770 27760 43834 27764
rect 43850 27820 43914 27824
rect 43850 27764 43854 27820
rect 43854 27764 43910 27820
rect 43910 27764 43914 27820
rect 43850 27760 43914 27764
rect 48938 27820 49002 27824
rect 48938 27764 48942 27820
rect 48942 27764 48998 27820
rect 48998 27764 49002 27820
rect 48938 27760 49002 27764
rect 49018 27820 49082 27824
rect 49018 27764 49022 27820
rect 49022 27764 49078 27820
rect 49078 27764 49082 27820
rect 49018 27760 49082 27764
rect 49098 27820 49162 27824
rect 49098 27764 49102 27820
rect 49102 27764 49158 27820
rect 49158 27764 49162 27820
rect 49098 27760 49162 27764
rect 49178 27820 49242 27824
rect 49178 27764 49182 27820
rect 49182 27764 49238 27820
rect 49238 27764 49242 27820
rect 49178 27760 49242 27764
rect 54266 27820 54330 27824
rect 54266 27764 54270 27820
rect 54270 27764 54326 27820
rect 54326 27764 54330 27820
rect 54266 27760 54330 27764
rect 54346 27820 54410 27824
rect 54346 27764 54350 27820
rect 54350 27764 54406 27820
rect 54406 27764 54410 27820
rect 54346 27760 54410 27764
rect 54426 27820 54490 27824
rect 54426 27764 54430 27820
rect 54430 27764 54486 27820
rect 54486 27764 54490 27820
rect 54426 27760 54490 27764
rect 54506 27820 54570 27824
rect 54506 27764 54510 27820
rect 54510 27764 54566 27820
rect 54566 27764 54570 27820
rect 54506 27760 54570 27764
rect 59594 27820 59658 27824
rect 59594 27764 59598 27820
rect 59598 27764 59654 27820
rect 59654 27764 59658 27820
rect 59594 27760 59658 27764
rect 59674 27820 59738 27824
rect 59674 27764 59678 27820
rect 59678 27764 59734 27820
rect 59734 27764 59738 27820
rect 59674 27760 59738 27764
rect 59754 27820 59818 27824
rect 59754 27764 59758 27820
rect 59758 27764 59814 27820
rect 59814 27764 59818 27820
rect 59754 27760 59818 27764
rect 59834 27820 59898 27824
rect 59834 27764 59838 27820
rect 59838 27764 59894 27820
rect 59894 27764 59898 27820
rect 59834 27760 59898 27764
rect 64922 27820 64986 27824
rect 64922 27764 64926 27820
rect 64926 27764 64982 27820
rect 64982 27764 64986 27820
rect 64922 27760 64986 27764
rect 65002 27820 65066 27824
rect 65002 27764 65006 27820
rect 65006 27764 65062 27820
rect 65062 27764 65066 27820
rect 65002 27760 65066 27764
rect 65082 27820 65146 27824
rect 65082 27764 65086 27820
rect 65086 27764 65142 27820
rect 65142 27764 65146 27820
rect 65082 27760 65146 27764
rect 65162 27820 65226 27824
rect 65162 27764 65166 27820
rect 65166 27764 65222 27820
rect 65222 27764 65226 27820
rect 65162 27760 65226 27764
rect 70250 27820 70314 27824
rect 70250 27764 70254 27820
rect 70254 27764 70310 27820
rect 70310 27764 70314 27820
rect 70250 27760 70314 27764
rect 70330 27820 70394 27824
rect 70330 27764 70334 27820
rect 70334 27764 70390 27820
rect 70390 27764 70394 27820
rect 70330 27760 70394 27764
rect 70410 27820 70474 27824
rect 70410 27764 70414 27820
rect 70414 27764 70470 27820
rect 70470 27764 70474 27820
rect 70410 27760 70474 27764
rect 70490 27820 70554 27824
rect 70490 27764 70494 27820
rect 70494 27764 70550 27820
rect 70550 27764 70554 27820
rect 70490 27760 70554 27764
rect 75578 27820 75642 27824
rect 75578 27764 75582 27820
rect 75582 27764 75638 27820
rect 75638 27764 75642 27820
rect 75578 27760 75642 27764
rect 75658 27820 75722 27824
rect 75658 27764 75662 27820
rect 75662 27764 75718 27820
rect 75718 27764 75722 27820
rect 75658 27760 75722 27764
rect 75738 27820 75802 27824
rect 75738 27764 75742 27820
rect 75742 27764 75798 27820
rect 75798 27764 75802 27820
rect 75738 27760 75802 27764
rect 75818 27820 75882 27824
rect 75818 27764 75822 27820
rect 75822 27764 75878 27820
rect 75878 27764 75882 27820
rect 75818 27760 75882 27764
rect 80906 27820 80970 27824
rect 80906 27764 80910 27820
rect 80910 27764 80966 27820
rect 80966 27764 80970 27820
rect 80906 27760 80970 27764
rect 80986 27820 81050 27824
rect 80986 27764 80990 27820
rect 80990 27764 81046 27820
rect 81046 27764 81050 27820
rect 80986 27760 81050 27764
rect 81066 27820 81130 27824
rect 81066 27764 81070 27820
rect 81070 27764 81126 27820
rect 81126 27764 81130 27820
rect 81066 27760 81130 27764
rect 81146 27820 81210 27824
rect 81146 27764 81150 27820
rect 81150 27764 81206 27820
rect 81206 27764 81210 27820
rect 81146 27760 81210 27764
rect 86234 27820 86298 27824
rect 86234 27764 86238 27820
rect 86238 27764 86294 27820
rect 86294 27764 86298 27820
rect 86234 27760 86298 27764
rect 86314 27820 86378 27824
rect 86314 27764 86318 27820
rect 86318 27764 86374 27820
rect 86374 27764 86378 27820
rect 86314 27760 86378 27764
rect 86394 27820 86458 27824
rect 86394 27764 86398 27820
rect 86398 27764 86454 27820
rect 86454 27764 86458 27820
rect 86394 27760 86458 27764
rect 86474 27820 86538 27824
rect 86474 27764 86478 27820
rect 86478 27764 86534 27820
rect 86534 27764 86538 27820
rect 86474 27760 86538 27764
rect 91562 27820 91626 27824
rect 91562 27764 91566 27820
rect 91566 27764 91622 27820
rect 91622 27764 91626 27820
rect 91562 27760 91626 27764
rect 91642 27820 91706 27824
rect 91642 27764 91646 27820
rect 91646 27764 91702 27820
rect 91702 27764 91706 27820
rect 91642 27760 91706 27764
rect 91722 27820 91786 27824
rect 91722 27764 91726 27820
rect 91726 27764 91782 27820
rect 91782 27764 91786 27820
rect 91722 27760 91786 27764
rect 91802 27820 91866 27824
rect 91802 27764 91806 27820
rect 91806 27764 91862 27820
rect 91862 27764 91866 27820
rect 91802 27760 91866 27764
rect 3650 27276 3714 27280
rect 3650 27220 3654 27276
rect 3654 27220 3710 27276
rect 3710 27220 3714 27276
rect 3650 27216 3714 27220
rect 3730 27276 3794 27280
rect 3730 27220 3734 27276
rect 3734 27220 3790 27276
rect 3790 27220 3794 27276
rect 3730 27216 3794 27220
rect 3810 27276 3874 27280
rect 3810 27220 3814 27276
rect 3814 27220 3870 27276
rect 3870 27220 3874 27276
rect 3810 27216 3874 27220
rect 3890 27276 3954 27280
rect 3890 27220 3894 27276
rect 3894 27220 3950 27276
rect 3950 27220 3954 27276
rect 3890 27216 3954 27220
rect 8978 27276 9042 27280
rect 8978 27220 8982 27276
rect 8982 27220 9038 27276
rect 9038 27220 9042 27276
rect 8978 27216 9042 27220
rect 9058 27276 9122 27280
rect 9058 27220 9062 27276
rect 9062 27220 9118 27276
rect 9118 27220 9122 27276
rect 9058 27216 9122 27220
rect 9138 27276 9202 27280
rect 9138 27220 9142 27276
rect 9142 27220 9198 27276
rect 9198 27220 9202 27276
rect 9138 27216 9202 27220
rect 9218 27276 9282 27280
rect 9218 27220 9222 27276
rect 9222 27220 9278 27276
rect 9278 27220 9282 27276
rect 9218 27216 9282 27220
rect 14306 27276 14370 27280
rect 14306 27220 14310 27276
rect 14310 27220 14366 27276
rect 14366 27220 14370 27276
rect 14306 27216 14370 27220
rect 14386 27276 14450 27280
rect 14386 27220 14390 27276
rect 14390 27220 14446 27276
rect 14446 27220 14450 27276
rect 14386 27216 14450 27220
rect 14466 27276 14530 27280
rect 14466 27220 14470 27276
rect 14470 27220 14526 27276
rect 14526 27220 14530 27276
rect 14466 27216 14530 27220
rect 14546 27276 14610 27280
rect 14546 27220 14550 27276
rect 14550 27220 14606 27276
rect 14606 27220 14610 27276
rect 14546 27216 14610 27220
rect 19634 27276 19698 27280
rect 19634 27220 19638 27276
rect 19638 27220 19694 27276
rect 19694 27220 19698 27276
rect 19634 27216 19698 27220
rect 19714 27276 19778 27280
rect 19714 27220 19718 27276
rect 19718 27220 19774 27276
rect 19774 27220 19778 27276
rect 19714 27216 19778 27220
rect 19794 27276 19858 27280
rect 19794 27220 19798 27276
rect 19798 27220 19854 27276
rect 19854 27220 19858 27276
rect 19794 27216 19858 27220
rect 19874 27276 19938 27280
rect 19874 27220 19878 27276
rect 19878 27220 19934 27276
rect 19934 27220 19938 27276
rect 19874 27216 19938 27220
rect 24962 27276 25026 27280
rect 24962 27220 24966 27276
rect 24966 27220 25022 27276
rect 25022 27220 25026 27276
rect 24962 27216 25026 27220
rect 25042 27276 25106 27280
rect 25042 27220 25046 27276
rect 25046 27220 25102 27276
rect 25102 27220 25106 27276
rect 25042 27216 25106 27220
rect 25122 27276 25186 27280
rect 25122 27220 25126 27276
rect 25126 27220 25182 27276
rect 25182 27220 25186 27276
rect 25122 27216 25186 27220
rect 25202 27276 25266 27280
rect 25202 27220 25206 27276
rect 25206 27220 25262 27276
rect 25262 27220 25266 27276
rect 25202 27216 25266 27220
rect 30290 27276 30354 27280
rect 30290 27220 30294 27276
rect 30294 27220 30350 27276
rect 30350 27220 30354 27276
rect 30290 27216 30354 27220
rect 30370 27276 30434 27280
rect 30370 27220 30374 27276
rect 30374 27220 30430 27276
rect 30430 27220 30434 27276
rect 30370 27216 30434 27220
rect 30450 27276 30514 27280
rect 30450 27220 30454 27276
rect 30454 27220 30510 27276
rect 30510 27220 30514 27276
rect 30450 27216 30514 27220
rect 30530 27276 30594 27280
rect 30530 27220 30534 27276
rect 30534 27220 30590 27276
rect 30590 27220 30594 27276
rect 30530 27216 30594 27220
rect 35618 27276 35682 27280
rect 35618 27220 35622 27276
rect 35622 27220 35678 27276
rect 35678 27220 35682 27276
rect 35618 27216 35682 27220
rect 35698 27276 35762 27280
rect 35698 27220 35702 27276
rect 35702 27220 35758 27276
rect 35758 27220 35762 27276
rect 35698 27216 35762 27220
rect 35778 27276 35842 27280
rect 35778 27220 35782 27276
rect 35782 27220 35838 27276
rect 35838 27220 35842 27276
rect 35778 27216 35842 27220
rect 35858 27276 35922 27280
rect 35858 27220 35862 27276
rect 35862 27220 35918 27276
rect 35918 27220 35922 27276
rect 35858 27216 35922 27220
rect 40946 27276 41010 27280
rect 40946 27220 40950 27276
rect 40950 27220 41006 27276
rect 41006 27220 41010 27276
rect 40946 27216 41010 27220
rect 41026 27276 41090 27280
rect 41026 27220 41030 27276
rect 41030 27220 41086 27276
rect 41086 27220 41090 27276
rect 41026 27216 41090 27220
rect 41106 27276 41170 27280
rect 41106 27220 41110 27276
rect 41110 27220 41166 27276
rect 41166 27220 41170 27276
rect 41106 27216 41170 27220
rect 41186 27276 41250 27280
rect 41186 27220 41190 27276
rect 41190 27220 41246 27276
rect 41246 27220 41250 27276
rect 41186 27216 41250 27220
rect 46274 27276 46338 27280
rect 46274 27220 46278 27276
rect 46278 27220 46334 27276
rect 46334 27220 46338 27276
rect 46274 27216 46338 27220
rect 46354 27276 46418 27280
rect 46354 27220 46358 27276
rect 46358 27220 46414 27276
rect 46414 27220 46418 27276
rect 46354 27216 46418 27220
rect 46434 27276 46498 27280
rect 46434 27220 46438 27276
rect 46438 27220 46494 27276
rect 46494 27220 46498 27276
rect 46434 27216 46498 27220
rect 46514 27276 46578 27280
rect 46514 27220 46518 27276
rect 46518 27220 46574 27276
rect 46574 27220 46578 27276
rect 46514 27216 46578 27220
rect 51602 27276 51666 27280
rect 51602 27220 51606 27276
rect 51606 27220 51662 27276
rect 51662 27220 51666 27276
rect 51602 27216 51666 27220
rect 51682 27276 51746 27280
rect 51682 27220 51686 27276
rect 51686 27220 51742 27276
rect 51742 27220 51746 27276
rect 51682 27216 51746 27220
rect 51762 27276 51826 27280
rect 51762 27220 51766 27276
rect 51766 27220 51822 27276
rect 51822 27220 51826 27276
rect 51762 27216 51826 27220
rect 51842 27276 51906 27280
rect 51842 27220 51846 27276
rect 51846 27220 51902 27276
rect 51902 27220 51906 27276
rect 51842 27216 51906 27220
rect 56930 27276 56994 27280
rect 56930 27220 56934 27276
rect 56934 27220 56990 27276
rect 56990 27220 56994 27276
rect 56930 27216 56994 27220
rect 57010 27276 57074 27280
rect 57010 27220 57014 27276
rect 57014 27220 57070 27276
rect 57070 27220 57074 27276
rect 57010 27216 57074 27220
rect 57090 27276 57154 27280
rect 57090 27220 57094 27276
rect 57094 27220 57150 27276
rect 57150 27220 57154 27276
rect 57090 27216 57154 27220
rect 57170 27276 57234 27280
rect 57170 27220 57174 27276
rect 57174 27220 57230 27276
rect 57230 27220 57234 27276
rect 57170 27216 57234 27220
rect 62258 27276 62322 27280
rect 62258 27220 62262 27276
rect 62262 27220 62318 27276
rect 62318 27220 62322 27276
rect 62258 27216 62322 27220
rect 62338 27276 62402 27280
rect 62338 27220 62342 27276
rect 62342 27220 62398 27276
rect 62398 27220 62402 27276
rect 62338 27216 62402 27220
rect 62418 27276 62482 27280
rect 62418 27220 62422 27276
rect 62422 27220 62478 27276
rect 62478 27220 62482 27276
rect 62418 27216 62482 27220
rect 62498 27276 62562 27280
rect 62498 27220 62502 27276
rect 62502 27220 62558 27276
rect 62558 27220 62562 27276
rect 62498 27216 62562 27220
rect 67586 27276 67650 27280
rect 67586 27220 67590 27276
rect 67590 27220 67646 27276
rect 67646 27220 67650 27276
rect 67586 27216 67650 27220
rect 67666 27276 67730 27280
rect 67666 27220 67670 27276
rect 67670 27220 67726 27276
rect 67726 27220 67730 27276
rect 67666 27216 67730 27220
rect 67746 27276 67810 27280
rect 67746 27220 67750 27276
rect 67750 27220 67806 27276
rect 67806 27220 67810 27276
rect 67746 27216 67810 27220
rect 67826 27276 67890 27280
rect 67826 27220 67830 27276
rect 67830 27220 67886 27276
rect 67886 27220 67890 27276
rect 67826 27216 67890 27220
rect 72914 27276 72978 27280
rect 72914 27220 72918 27276
rect 72918 27220 72974 27276
rect 72974 27220 72978 27276
rect 72914 27216 72978 27220
rect 72994 27276 73058 27280
rect 72994 27220 72998 27276
rect 72998 27220 73054 27276
rect 73054 27220 73058 27276
rect 72994 27216 73058 27220
rect 73074 27276 73138 27280
rect 73074 27220 73078 27276
rect 73078 27220 73134 27276
rect 73134 27220 73138 27276
rect 73074 27216 73138 27220
rect 73154 27276 73218 27280
rect 73154 27220 73158 27276
rect 73158 27220 73214 27276
rect 73214 27220 73218 27276
rect 73154 27216 73218 27220
rect 78242 27276 78306 27280
rect 78242 27220 78246 27276
rect 78246 27220 78302 27276
rect 78302 27220 78306 27276
rect 78242 27216 78306 27220
rect 78322 27276 78386 27280
rect 78322 27220 78326 27276
rect 78326 27220 78382 27276
rect 78382 27220 78386 27276
rect 78322 27216 78386 27220
rect 78402 27276 78466 27280
rect 78402 27220 78406 27276
rect 78406 27220 78462 27276
rect 78462 27220 78466 27276
rect 78402 27216 78466 27220
rect 78482 27276 78546 27280
rect 78482 27220 78486 27276
rect 78486 27220 78542 27276
rect 78542 27220 78546 27276
rect 78482 27216 78546 27220
rect 83570 27276 83634 27280
rect 83570 27220 83574 27276
rect 83574 27220 83630 27276
rect 83630 27220 83634 27276
rect 83570 27216 83634 27220
rect 83650 27276 83714 27280
rect 83650 27220 83654 27276
rect 83654 27220 83710 27276
rect 83710 27220 83714 27276
rect 83650 27216 83714 27220
rect 83730 27276 83794 27280
rect 83730 27220 83734 27276
rect 83734 27220 83790 27276
rect 83790 27220 83794 27276
rect 83730 27216 83794 27220
rect 83810 27276 83874 27280
rect 83810 27220 83814 27276
rect 83814 27220 83870 27276
rect 83870 27220 83874 27276
rect 83810 27216 83874 27220
rect 88898 27276 88962 27280
rect 88898 27220 88902 27276
rect 88902 27220 88958 27276
rect 88958 27220 88962 27276
rect 88898 27216 88962 27220
rect 88978 27276 89042 27280
rect 88978 27220 88982 27276
rect 88982 27220 89038 27276
rect 89038 27220 89042 27276
rect 88978 27216 89042 27220
rect 89058 27276 89122 27280
rect 89058 27220 89062 27276
rect 89062 27220 89118 27276
rect 89118 27220 89122 27276
rect 89058 27216 89122 27220
rect 89138 27276 89202 27280
rect 89138 27220 89142 27276
rect 89142 27220 89198 27276
rect 89198 27220 89202 27276
rect 89138 27216 89202 27220
rect 6314 26732 6378 26736
rect 6314 26676 6318 26732
rect 6318 26676 6374 26732
rect 6374 26676 6378 26732
rect 6314 26672 6378 26676
rect 6394 26732 6458 26736
rect 6394 26676 6398 26732
rect 6398 26676 6454 26732
rect 6454 26676 6458 26732
rect 6394 26672 6458 26676
rect 6474 26732 6538 26736
rect 6474 26676 6478 26732
rect 6478 26676 6534 26732
rect 6534 26676 6538 26732
rect 6474 26672 6538 26676
rect 6554 26732 6618 26736
rect 6554 26676 6558 26732
rect 6558 26676 6614 26732
rect 6614 26676 6618 26732
rect 6554 26672 6618 26676
rect 11642 26732 11706 26736
rect 11642 26676 11646 26732
rect 11646 26676 11702 26732
rect 11702 26676 11706 26732
rect 11642 26672 11706 26676
rect 11722 26732 11786 26736
rect 11722 26676 11726 26732
rect 11726 26676 11782 26732
rect 11782 26676 11786 26732
rect 11722 26672 11786 26676
rect 11802 26732 11866 26736
rect 11802 26676 11806 26732
rect 11806 26676 11862 26732
rect 11862 26676 11866 26732
rect 11802 26672 11866 26676
rect 11882 26732 11946 26736
rect 11882 26676 11886 26732
rect 11886 26676 11942 26732
rect 11942 26676 11946 26732
rect 11882 26672 11946 26676
rect 16970 26732 17034 26736
rect 16970 26676 16974 26732
rect 16974 26676 17030 26732
rect 17030 26676 17034 26732
rect 16970 26672 17034 26676
rect 17050 26732 17114 26736
rect 17050 26676 17054 26732
rect 17054 26676 17110 26732
rect 17110 26676 17114 26732
rect 17050 26672 17114 26676
rect 17130 26732 17194 26736
rect 17130 26676 17134 26732
rect 17134 26676 17190 26732
rect 17190 26676 17194 26732
rect 17130 26672 17194 26676
rect 17210 26732 17274 26736
rect 17210 26676 17214 26732
rect 17214 26676 17270 26732
rect 17270 26676 17274 26732
rect 17210 26672 17274 26676
rect 22298 26732 22362 26736
rect 22298 26676 22302 26732
rect 22302 26676 22358 26732
rect 22358 26676 22362 26732
rect 22298 26672 22362 26676
rect 22378 26732 22442 26736
rect 22378 26676 22382 26732
rect 22382 26676 22438 26732
rect 22438 26676 22442 26732
rect 22378 26672 22442 26676
rect 22458 26732 22522 26736
rect 22458 26676 22462 26732
rect 22462 26676 22518 26732
rect 22518 26676 22522 26732
rect 22458 26672 22522 26676
rect 22538 26732 22602 26736
rect 22538 26676 22542 26732
rect 22542 26676 22598 26732
rect 22598 26676 22602 26732
rect 22538 26672 22602 26676
rect 27626 26732 27690 26736
rect 27626 26676 27630 26732
rect 27630 26676 27686 26732
rect 27686 26676 27690 26732
rect 27626 26672 27690 26676
rect 27706 26732 27770 26736
rect 27706 26676 27710 26732
rect 27710 26676 27766 26732
rect 27766 26676 27770 26732
rect 27706 26672 27770 26676
rect 27786 26732 27850 26736
rect 27786 26676 27790 26732
rect 27790 26676 27846 26732
rect 27846 26676 27850 26732
rect 27786 26672 27850 26676
rect 27866 26732 27930 26736
rect 27866 26676 27870 26732
rect 27870 26676 27926 26732
rect 27926 26676 27930 26732
rect 27866 26672 27930 26676
rect 32954 26732 33018 26736
rect 32954 26676 32958 26732
rect 32958 26676 33014 26732
rect 33014 26676 33018 26732
rect 32954 26672 33018 26676
rect 33034 26732 33098 26736
rect 33034 26676 33038 26732
rect 33038 26676 33094 26732
rect 33094 26676 33098 26732
rect 33034 26672 33098 26676
rect 33114 26732 33178 26736
rect 33114 26676 33118 26732
rect 33118 26676 33174 26732
rect 33174 26676 33178 26732
rect 33114 26672 33178 26676
rect 33194 26732 33258 26736
rect 33194 26676 33198 26732
rect 33198 26676 33254 26732
rect 33254 26676 33258 26732
rect 33194 26672 33258 26676
rect 38282 26732 38346 26736
rect 38282 26676 38286 26732
rect 38286 26676 38342 26732
rect 38342 26676 38346 26732
rect 38282 26672 38346 26676
rect 38362 26732 38426 26736
rect 38362 26676 38366 26732
rect 38366 26676 38422 26732
rect 38422 26676 38426 26732
rect 38362 26672 38426 26676
rect 38442 26732 38506 26736
rect 38442 26676 38446 26732
rect 38446 26676 38502 26732
rect 38502 26676 38506 26732
rect 38442 26672 38506 26676
rect 38522 26732 38586 26736
rect 38522 26676 38526 26732
rect 38526 26676 38582 26732
rect 38582 26676 38586 26732
rect 38522 26672 38586 26676
rect 43610 26732 43674 26736
rect 43610 26676 43614 26732
rect 43614 26676 43670 26732
rect 43670 26676 43674 26732
rect 43610 26672 43674 26676
rect 43690 26732 43754 26736
rect 43690 26676 43694 26732
rect 43694 26676 43750 26732
rect 43750 26676 43754 26732
rect 43690 26672 43754 26676
rect 43770 26732 43834 26736
rect 43770 26676 43774 26732
rect 43774 26676 43830 26732
rect 43830 26676 43834 26732
rect 43770 26672 43834 26676
rect 43850 26732 43914 26736
rect 43850 26676 43854 26732
rect 43854 26676 43910 26732
rect 43910 26676 43914 26732
rect 43850 26672 43914 26676
rect 48938 26732 49002 26736
rect 48938 26676 48942 26732
rect 48942 26676 48998 26732
rect 48998 26676 49002 26732
rect 48938 26672 49002 26676
rect 49018 26732 49082 26736
rect 49018 26676 49022 26732
rect 49022 26676 49078 26732
rect 49078 26676 49082 26732
rect 49018 26672 49082 26676
rect 49098 26732 49162 26736
rect 49098 26676 49102 26732
rect 49102 26676 49158 26732
rect 49158 26676 49162 26732
rect 49098 26672 49162 26676
rect 49178 26732 49242 26736
rect 49178 26676 49182 26732
rect 49182 26676 49238 26732
rect 49238 26676 49242 26732
rect 49178 26672 49242 26676
rect 54266 26732 54330 26736
rect 54266 26676 54270 26732
rect 54270 26676 54326 26732
rect 54326 26676 54330 26732
rect 54266 26672 54330 26676
rect 54346 26732 54410 26736
rect 54346 26676 54350 26732
rect 54350 26676 54406 26732
rect 54406 26676 54410 26732
rect 54346 26672 54410 26676
rect 54426 26732 54490 26736
rect 54426 26676 54430 26732
rect 54430 26676 54486 26732
rect 54486 26676 54490 26732
rect 54426 26672 54490 26676
rect 54506 26732 54570 26736
rect 54506 26676 54510 26732
rect 54510 26676 54566 26732
rect 54566 26676 54570 26732
rect 54506 26672 54570 26676
rect 59594 26732 59658 26736
rect 59594 26676 59598 26732
rect 59598 26676 59654 26732
rect 59654 26676 59658 26732
rect 59594 26672 59658 26676
rect 59674 26732 59738 26736
rect 59674 26676 59678 26732
rect 59678 26676 59734 26732
rect 59734 26676 59738 26732
rect 59674 26672 59738 26676
rect 59754 26732 59818 26736
rect 59754 26676 59758 26732
rect 59758 26676 59814 26732
rect 59814 26676 59818 26732
rect 59754 26672 59818 26676
rect 59834 26732 59898 26736
rect 59834 26676 59838 26732
rect 59838 26676 59894 26732
rect 59894 26676 59898 26732
rect 59834 26672 59898 26676
rect 64922 26732 64986 26736
rect 64922 26676 64926 26732
rect 64926 26676 64982 26732
rect 64982 26676 64986 26732
rect 64922 26672 64986 26676
rect 65002 26732 65066 26736
rect 65002 26676 65006 26732
rect 65006 26676 65062 26732
rect 65062 26676 65066 26732
rect 65002 26672 65066 26676
rect 65082 26732 65146 26736
rect 65082 26676 65086 26732
rect 65086 26676 65142 26732
rect 65142 26676 65146 26732
rect 65082 26672 65146 26676
rect 65162 26732 65226 26736
rect 65162 26676 65166 26732
rect 65166 26676 65222 26732
rect 65222 26676 65226 26732
rect 65162 26672 65226 26676
rect 70250 26732 70314 26736
rect 70250 26676 70254 26732
rect 70254 26676 70310 26732
rect 70310 26676 70314 26732
rect 70250 26672 70314 26676
rect 70330 26732 70394 26736
rect 70330 26676 70334 26732
rect 70334 26676 70390 26732
rect 70390 26676 70394 26732
rect 70330 26672 70394 26676
rect 70410 26732 70474 26736
rect 70410 26676 70414 26732
rect 70414 26676 70470 26732
rect 70470 26676 70474 26732
rect 70410 26672 70474 26676
rect 70490 26732 70554 26736
rect 70490 26676 70494 26732
rect 70494 26676 70550 26732
rect 70550 26676 70554 26732
rect 70490 26672 70554 26676
rect 75578 26732 75642 26736
rect 75578 26676 75582 26732
rect 75582 26676 75638 26732
rect 75638 26676 75642 26732
rect 75578 26672 75642 26676
rect 75658 26732 75722 26736
rect 75658 26676 75662 26732
rect 75662 26676 75718 26732
rect 75718 26676 75722 26732
rect 75658 26672 75722 26676
rect 75738 26732 75802 26736
rect 75738 26676 75742 26732
rect 75742 26676 75798 26732
rect 75798 26676 75802 26732
rect 75738 26672 75802 26676
rect 75818 26732 75882 26736
rect 75818 26676 75822 26732
rect 75822 26676 75878 26732
rect 75878 26676 75882 26732
rect 75818 26672 75882 26676
rect 80906 26732 80970 26736
rect 80906 26676 80910 26732
rect 80910 26676 80966 26732
rect 80966 26676 80970 26732
rect 80906 26672 80970 26676
rect 80986 26732 81050 26736
rect 80986 26676 80990 26732
rect 80990 26676 81046 26732
rect 81046 26676 81050 26732
rect 80986 26672 81050 26676
rect 81066 26732 81130 26736
rect 81066 26676 81070 26732
rect 81070 26676 81126 26732
rect 81126 26676 81130 26732
rect 81066 26672 81130 26676
rect 81146 26732 81210 26736
rect 81146 26676 81150 26732
rect 81150 26676 81206 26732
rect 81206 26676 81210 26732
rect 81146 26672 81210 26676
rect 86234 26732 86298 26736
rect 86234 26676 86238 26732
rect 86238 26676 86294 26732
rect 86294 26676 86298 26732
rect 86234 26672 86298 26676
rect 86314 26732 86378 26736
rect 86314 26676 86318 26732
rect 86318 26676 86374 26732
rect 86374 26676 86378 26732
rect 86314 26672 86378 26676
rect 86394 26732 86458 26736
rect 86394 26676 86398 26732
rect 86398 26676 86454 26732
rect 86454 26676 86458 26732
rect 86394 26672 86458 26676
rect 86474 26732 86538 26736
rect 86474 26676 86478 26732
rect 86478 26676 86534 26732
rect 86534 26676 86538 26732
rect 86474 26672 86538 26676
rect 91562 26732 91626 26736
rect 91562 26676 91566 26732
rect 91566 26676 91622 26732
rect 91622 26676 91626 26732
rect 91562 26672 91626 26676
rect 91642 26732 91706 26736
rect 91642 26676 91646 26732
rect 91646 26676 91702 26732
rect 91702 26676 91706 26732
rect 91642 26672 91706 26676
rect 91722 26732 91786 26736
rect 91722 26676 91726 26732
rect 91726 26676 91782 26732
rect 91782 26676 91786 26732
rect 91722 26672 91786 26676
rect 91802 26732 91866 26736
rect 91802 26676 91806 26732
rect 91806 26676 91862 26732
rect 91862 26676 91866 26732
rect 91802 26672 91866 26676
rect 3650 26188 3714 26192
rect 3650 26132 3654 26188
rect 3654 26132 3710 26188
rect 3710 26132 3714 26188
rect 3650 26128 3714 26132
rect 3730 26188 3794 26192
rect 3730 26132 3734 26188
rect 3734 26132 3790 26188
rect 3790 26132 3794 26188
rect 3730 26128 3794 26132
rect 3810 26188 3874 26192
rect 3810 26132 3814 26188
rect 3814 26132 3870 26188
rect 3870 26132 3874 26188
rect 3810 26128 3874 26132
rect 3890 26188 3954 26192
rect 3890 26132 3894 26188
rect 3894 26132 3950 26188
rect 3950 26132 3954 26188
rect 3890 26128 3954 26132
rect 35618 26188 35682 26192
rect 35618 26132 35622 26188
rect 35622 26132 35678 26188
rect 35678 26132 35682 26188
rect 35618 26128 35682 26132
rect 35698 26188 35762 26192
rect 35698 26132 35702 26188
rect 35702 26132 35758 26188
rect 35758 26132 35762 26188
rect 35698 26128 35762 26132
rect 35778 26188 35842 26192
rect 35778 26132 35782 26188
rect 35782 26132 35838 26188
rect 35838 26132 35842 26188
rect 35778 26128 35842 26132
rect 35858 26188 35922 26192
rect 35858 26132 35862 26188
rect 35862 26132 35918 26188
rect 35918 26132 35922 26188
rect 35858 26128 35922 26132
rect 40946 26188 41010 26192
rect 40946 26132 40950 26188
rect 40950 26132 41006 26188
rect 41006 26132 41010 26188
rect 40946 26128 41010 26132
rect 41026 26188 41090 26192
rect 41026 26132 41030 26188
rect 41030 26132 41086 26188
rect 41086 26132 41090 26188
rect 41026 26128 41090 26132
rect 41106 26188 41170 26192
rect 41106 26132 41110 26188
rect 41110 26132 41166 26188
rect 41166 26132 41170 26188
rect 41106 26128 41170 26132
rect 41186 26188 41250 26192
rect 41186 26132 41190 26188
rect 41190 26132 41246 26188
rect 41246 26132 41250 26188
rect 41186 26128 41250 26132
rect 6314 25644 6378 25648
rect 6314 25588 6318 25644
rect 6318 25588 6374 25644
rect 6374 25588 6378 25644
rect 6314 25584 6378 25588
rect 6394 25644 6458 25648
rect 6394 25588 6398 25644
rect 6398 25588 6454 25644
rect 6454 25588 6458 25644
rect 6394 25584 6458 25588
rect 6474 25644 6538 25648
rect 6474 25588 6478 25644
rect 6478 25588 6534 25644
rect 6534 25588 6538 25644
rect 6474 25584 6538 25588
rect 6554 25644 6618 25648
rect 6554 25588 6558 25644
rect 6558 25588 6614 25644
rect 6614 25588 6618 25644
rect 6554 25584 6618 25588
rect 38282 25644 38346 25648
rect 38282 25588 38286 25644
rect 38286 25588 38342 25644
rect 38342 25588 38346 25644
rect 38282 25584 38346 25588
rect 38362 25644 38426 25648
rect 38362 25588 38366 25644
rect 38366 25588 38422 25644
rect 38422 25588 38426 25644
rect 38362 25584 38426 25588
rect 38442 25644 38506 25648
rect 38442 25588 38446 25644
rect 38446 25588 38502 25644
rect 38502 25588 38506 25644
rect 38442 25584 38506 25588
rect 38522 25644 38586 25648
rect 38522 25588 38526 25644
rect 38526 25588 38582 25644
rect 38582 25588 38586 25644
rect 38522 25584 38586 25588
rect 3650 25100 3714 25104
rect 3650 25044 3654 25100
rect 3654 25044 3710 25100
rect 3710 25044 3714 25100
rect 3650 25040 3714 25044
rect 3730 25100 3794 25104
rect 3730 25044 3734 25100
rect 3734 25044 3790 25100
rect 3790 25044 3794 25100
rect 3730 25040 3794 25044
rect 3810 25100 3874 25104
rect 3810 25044 3814 25100
rect 3814 25044 3870 25100
rect 3870 25044 3874 25100
rect 3810 25040 3874 25044
rect 3890 25100 3954 25104
rect 3890 25044 3894 25100
rect 3894 25044 3950 25100
rect 3950 25044 3954 25100
rect 3890 25040 3954 25044
rect 35618 25100 35682 25104
rect 35618 25044 35622 25100
rect 35622 25044 35678 25100
rect 35678 25044 35682 25100
rect 35618 25040 35682 25044
rect 35698 25100 35762 25104
rect 35698 25044 35702 25100
rect 35702 25044 35758 25100
rect 35758 25044 35762 25100
rect 35698 25040 35762 25044
rect 35778 25100 35842 25104
rect 35778 25044 35782 25100
rect 35782 25044 35838 25100
rect 35838 25044 35842 25100
rect 35778 25040 35842 25044
rect 35858 25100 35922 25104
rect 35858 25044 35862 25100
rect 35862 25044 35918 25100
rect 35918 25044 35922 25100
rect 35858 25040 35922 25044
rect 40946 25100 41010 25104
rect 40946 25044 40950 25100
rect 40950 25044 41006 25100
rect 41006 25044 41010 25100
rect 40946 25040 41010 25044
rect 41026 25100 41090 25104
rect 41026 25044 41030 25100
rect 41030 25044 41086 25100
rect 41086 25044 41090 25100
rect 41026 25040 41090 25044
rect 41106 25100 41170 25104
rect 41106 25044 41110 25100
rect 41110 25044 41166 25100
rect 41166 25044 41170 25100
rect 41106 25040 41170 25044
rect 41186 25100 41250 25104
rect 41186 25044 41190 25100
rect 41190 25044 41246 25100
rect 41246 25044 41250 25100
rect 41186 25040 41250 25044
rect 6314 24556 6378 24560
rect 6314 24500 6318 24556
rect 6318 24500 6374 24556
rect 6374 24500 6378 24556
rect 6314 24496 6378 24500
rect 6394 24556 6458 24560
rect 6394 24500 6398 24556
rect 6398 24500 6454 24556
rect 6454 24500 6458 24556
rect 6394 24496 6458 24500
rect 6474 24556 6538 24560
rect 6474 24500 6478 24556
rect 6478 24500 6534 24556
rect 6534 24500 6538 24556
rect 6474 24496 6538 24500
rect 6554 24556 6618 24560
rect 6554 24500 6558 24556
rect 6558 24500 6614 24556
rect 6614 24500 6618 24556
rect 6554 24496 6618 24500
rect 38282 24556 38346 24560
rect 38282 24500 38286 24556
rect 38286 24500 38342 24556
rect 38342 24500 38346 24556
rect 38282 24496 38346 24500
rect 38362 24556 38426 24560
rect 38362 24500 38366 24556
rect 38366 24500 38422 24556
rect 38422 24500 38426 24556
rect 38362 24496 38426 24500
rect 38442 24556 38506 24560
rect 38442 24500 38446 24556
rect 38446 24500 38502 24556
rect 38502 24500 38506 24556
rect 38442 24496 38506 24500
rect 38522 24556 38586 24560
rect 38522 24500 38526 24556
rect 38526 24500 38582 24556
rect 38582 24500 38586 24556
rect 38522 24496 38586 24500
rect 3650 24012 3714 24016
rect 3650 23956 3654 24012
rect 3654 23956 3710 24012
rect 3710 23956 3714 24012
rect 3650 23952 3714 23956
rect 3730 24012 3794 24016
rect 3730 23956 3734 24012
rect 3734 23956 3790 24012
rect 3790 23956 3794 24012
rect 3730 23952 3794 23956
rect 3810 24012 3874 24016
rect 3810 23956 3814 24012
rect 3814 23956 3870 24012
rect 3870 23956 3874 24012
rect 3810 23952 3874 23956
rect 3890 24012 3954 24016
rect 3890 23956 3894 24012
rect 3894 23956 3950 24012
rect 3950 23956 3954 24012
rect 3890 23952 3954 23956
rect 35618 24012 35682 24016
rect 35618 23956 35622 24012
rect 35622 23956 35678 24012
rect 35678 23956 35682 24012
rect 35618 23952 35682 23956
rect 35698 24012 35762 24016
rect 35698 23956 35702 24012
rect 35702 23956 35758 24012
rect 35758 23956 35762 24012
rect 35698 23952 35762 23956
rect 35778 24012 35842 24016
rect 35778 23956 35782 24012
rect 35782 23956 35838 24012
rect 35838 23956 35842 24012
rect 35778 23952 35842 23956
rect 35858 24012 35922 24016
rect 35858 23956 35862 24012
rect 35862 23956 35918 24012
rect 35918 23956 35922 24012
rect 35858 23952 35922 23956
rect 40946 24012 41010 24016
rect 40946 23956 40950 24012
rect 40950 23956 41006 24012
rect 41006 23956 41010 24012
rect 40946 23952 41010 23956
rect 41026 24012 41090 24016
rect 41026 23956 41030 24012
rect 41030 23956 41086 24012
rect 41086 23956 41090 24012
rect 41026 23952 41090 23956
rect 41106 24012 41170 24016
rect 41106 23956 41110 24012
rect 41110 23956 41166 24012
rect 41166 23956 41170 24012
rect 41106 23952 41170 23956
rect 41186 24012 41250 24016
rect 41186 23956 41190 24012
rect 41190 23956 41246 24012
rect 41246 23956 41250 24012
rect 41186 23952 41250 23956
rect 6314 23468 6378 23472
rect 6314 23412 6318 23468
rect 6318 23412 6374 23468
rect 6374 23412 6378 23468
rect 6314 23408 6378 23412
rect 6394 23468 6458 23472
rect 6394 23412 6398 23468
rect 6398 23412 6454 23468
rect 6454 23412 6458 23468
rect 6394 23408 6458 23412
rect 6474 23468 6538 23472
rect 6474 23412 6478 23468
rect 6478 23412 6534 23468
rect 6534 23412 6538 23468
rect 6474 23408 6538 23412
rect 6554 23468 6618 23472
rect 6554 23412 6558 23468
rect 6558 23412 6614 23468
rect 6614 23412 6618 23468
rect 6554 23408 6618 23412
rect 38282 23468 38346 23472
rect 38282 23412 38286 23468
rect 38286 23412 38342 23468
rect 38342 23412 38346 23468
rect 38282 23408 38346 23412
rect 38362 23468 38426 23472
rect 38362 23412 38366 23468
rect 38366 23412 38422 23468
rect 38422 23412 38426 23468
rect 38362 23408 38426 23412
rect 38442 23468 38506 23472
rect 38442 23412 38446 23468
rect 38446 23412 38502 23468
rect 38502 23412 38506 23468
rect 38442 23408 38506 23412
rect 38522 23468 38586 23472
rect 38522 23412 38526 23468
rect 38526 23412 38582 23468
rect 38582 23412 38586 23468
rect 38522 23408 38586 23412
rect 3650 22924 3714 22928
rect 3650 22868 3654 22924
rect 3654 22868 3710 22924
rect 3710 22868 3714 22924
rect 3650 22864 3714 22868
rect 3730 22924 3794 22928
rect 3730 22868 3734 22924
rect 3734 22868 3790 22924
rect 3790 22868 3794 22924
rect 3730 22864 3794 22868
rect 3810 22924 3874 22928
rect 3810 22868 3814 22924
rect 3814 22868 3870 22924
rect 3870 22868 3874 22924
rect 3810 22864 3874 22868
rect 3890 22924 3954 22928
rect 3890 22868 3894 22924
rect 3894 22868 3950 22924
rect 3950 22868 3954 22924
rect 3890 22864 3954 22868
rect 35618 22924 35682 22928
rect 35618 22868 35622 22924
rect 35622 22868 35678 22924
rect 35678 22868 35682 22924
rect 35618 22864 35682 22868
rect 35698 22924 35762 22928
rect 35698 22868 35702 22924
rect 35702 22868 35758 22924
rect 35758 22868 35762 22924
rect 35698 22864 35762 22868
rect 35778 22924 35842 22928
rect 35778 22868 35782 22924
rect 35782 22868 35838 22924
rect 35838 22868 35842 22924
rect 35778 22864 35842 22868
rect 35858 22924 35922 22928
rect 35858 22868 35862 22924
rect 35862 22868 35918 22924
rect 35918 22868 35922 22924
rect 35858 22864 35922 22868
rect 40946 22924 41010 22928
rect 40946 22868 40950 22924
rect 40950 22868 41006 22924
rect 41006 22868 41010 22924
rect 40946 22864 41010 22868
rect 41026 22924 41090 22928
rect 41026 22868 41030 22924
rect 41030 22868 41086 22924
rect 41086 22868 41090 22924
rect 41026 22864 41090 22868
rect 41106 22924 41170 22928
rect 41106 22868 41110 22924
rect 41110 22868 41166 22924
rect 41166 22868 41170 22924
rect 41106 22864 41170 22868
rect 41186 22924 41250 22928
rect 41186 22868 41190 22924
rect 41190 22868 41246 22924
rect 41246 22868 41250 22924
rect 41186 22864 41250 22868
rect 3358 22660 3422 22724
rect 31510 22388 31574 22452
rect 6314 22380 6378 22384
rect 6314 22324 6318 22380
rect 6318 22324 6374 22380
rect 6374 22324 6378 22380
rect 6314 22320 6378 22324
rect 6394 22380 6458 22384
rect 6394 22324 6398 22380
rect 6398 22324 6454 22380
rect 6454 22324 6458 22380
rect 6394 22320 6458 22324
rect 6474 22380 6538 22384
rect 6474 22324 6478 22380
rect 6478 22324 6534 22380
rect 6534 22324 6538 22380
rect 6474 22320 6538 22324
rect 6554 22380 6618 22384
rect 6554 22324 6558 22380
rect 6558 22324 6614 22380
rect 6614 22324 6618 22380
rect 6554 22320 6618 22324
rect 38282 22380 38346 22384
rect 38282 22324 38286 22380
rect 38286 22324 38342 22380
rect 38342 22324 38346 22380
rect 38282 22320 38346 22324
rect 38362 22380 38426 22384
rect 38362 22324 38366 22380
rect 38366 22324 38422 22380
rect 38422 22324 38426 22380
rect 38362 22320 38426 22324
rect 38442 22380 38506 22384
rect 38442 22324 38446 22380
rect 38446 22324 38502 22380
rect 38502 22324 38506 22380
rect 38442 22320 38506 22324
rect 38522 22380 38586 22384
rect 38522 22324 38526 22380
rect 38526 22324 38582 22380
rect 38582 22324 38586 22380
rect 38522 22320 38586 22324
rect 3650 21836 3714 21840
rect 3650 21780 3654 21836
rect 3654 21780 3710 21836
rect 3710 21780 3714 21836
rect 3650 21776 3714 21780
rect 3730 21836 3794 21840
rect 3730 21780 3734 21836
rect 3734 21780 3790 21836
rect 3790 21780 3794 21836
rect 3730 21776 3794 21780
rect 3810 21836 3874 21840
rect 3810 21780 3814 21836
rect 3814 21780 3870 21836
rect 3870 21780 3874 21836
rect 3810 21776 3874 21780
rect 3890 21836 3954 21840
rect 3890 21780 3894 21836
rect 3894 21780 3950 21836
rect 3950 21780 3954 21836
rect 3890 21776 3954 21780
rect 35618 21836 35682 21840
rect 35618 21780 35622 21836
rect 35622 21780 35678 21836
rect 35678 21780 35682 21836
rect 35618 21776 35682 21780
rect 35698 21836 35762 21840
rect 35698 21780 35702 21836
rect 35702 21780 35758 21836
rect 35758 21780 35762 21836
rect 35698 21776 35762 21780
rect 35778 21836 35842 21840
rect 35778 21780 35782 21836
rect 35782 21780 35838 21836
rect 35838 21780 35842 21836
rect 35778 21776 35842 21780
rect 35858 21836 35922 21840
rect 35858 21780 35862 21836
rect 35862 21780 35918 21836
rect 35918 21780 35922 21836
rect 35858 21776 35922 21780
rect 40946 21836 41010 21840
rect 40946 21780 40950 21836
rect 40950 21780 41006 21836
rect 41006 21780 41010 21836
rect 40946 21776 41010 21780
rect 41026 21836 41090 21840
rect 41026 21780 41030 21836
rect 41030 21780 41086 21836
rect 41086 21780 41090 21836
rect 41026 21776 41090 21780
rect 41106 21836 41170 21840
rect 41106 21780 41110 21836
rect 41110 21780 41166 21836
rect 41166 21780 41170 21836
rect 41106 21776 41170 21780
rect 41186 21836 41250 21840
rect 41186 21780 41190 21836
rect 41190 21780 41246 21836
rect 41246 21780 41250 21836
rect 41186 21776 41250 21780
rect 37950 21436 38014 21500
rect 6314 21292 6378 21296
rect 6314 21236 6318 21292
rect 6318 21236 6374 21292
rect 6374 21236 6378 21292
rect 6314 21232 6378 21236
rect 6394 21292 6458 21296
rect 6394 21236 6398 21292
rect 6398 21236 6454 21292
rect 6454 21236 6458 21292
rect 6394 21232 6458 21236
rect 6474 21292 6538 21296
rect 6474 21236 6478 21292
rect 6478 21236 6534 21292
rect 6534 21236 6538 21292
rect 6474 21232 6538 21236
rect 6554 21292 6618 21296
rect 6554 21236 6558 21292
rect 6558 21236 6614 21292
rect 6614 21236 6618 21292
rect 6554 21232 6618 21236
rect 38282 21292 38346 21296
rect 38282 21236 38286 21292
rect 38286 21236 38342 21292
rect 38342 21236 38346 21292
rect 38282 21232 38346 21236
rect 38362 21292 38426 21296
rect 38362 21236 38366 21292
rect 38366 21236 38422 21292
rect 38422 21236 38426 21292
rect 38362 21232 38426 21236
rect 38442 21292 38506 21296
rect 38442 21236 38446 21292
rect 38446 21236 38502 21292
rect 38502 21236 38506 21292
rect 38442 21232 38506 21236
rect 38522 21292 38586 21296
rect 38522 21236 38526 21292
rect 38526 21236 38582 21292
rect 38582 21236 38586 21292
rect 38522 21232 38586 21236
rect 3650 20748 3714 20752
rect 3650 20692 3654 20748
rect 3654 20692 3710 20748
rect 3710 20692 3714 20748
rect 3650 20688 3714 20692
rect 3730 20748 3794 20752
rect 3730 20692 3734 20748
rect 3734 20692 3790 20748
rect 3790 20692 3794 20748
rect 3730 20688 3794 20692
rect 3810 20748 3874 20752
rect 3810 20692 3814 20748
rect 3814 20692 3870 20748
rect 3870 20692 3874 20748
rect 3810 20688 3874 20692
rect 3890 20748 3954 20752
rect 3890 20692 3894 20748
rect 3894 20692 3950 20748
rect 3950 20692 3954 20748
rect 3890 20688 3954 20692
rect 35618 20748 35682 20752
rect 35618 20692 35622 20748
rect 35622 20692 35678 20748
rect 35678 20692 35682 20748
rect 35618 20688 35682 20692
rect 35698 20748 35762 20752
rect 35698 20692 35702 20748
rect 35702 20692 35758 20748
rect 35758 20692 35762 20748
rect 35698 20688 35762 20692
rect 35778 20748 35842 20752
rect 35778 20692 35782 20748
rect 35782 20692 35838 20748
rect 35838 20692 35842 20748
rect 35778 20688 35842 20692
rect 35858 20748 35922 20752
rect 35858 20692 35862 20748
rect 35862 20692 35918 20748
rect 35918 20692 35922 20748
rect 35858 20688 35922 20692
rect 40946 20748 41010 20752
rect 40946 20692 40950 20748
rect 40950 20692 41006 20748
rect 41006 20692 41010 20748
rect 40946 20688 41010 20692
rect 41026 20748 41090 20752
rect 41026 20692 41030 20748
rect 41030 20692 41086 20748
rect 41086 20692 41090 20748
rect 41026 20688 41090 20692
rect 41106 20748 41170 20752
rect 41106 20692 41110 20748
rect 41110 20692 41166 20748
rect 41166 20692 41170 20748
rect 41106 20688 41170 20692
rect 41186 20748 41250 20752
rect 41186 20692 41190 20748
rect 41190 20692 41246 20748
rect 41246 20692 41250 20748
rect 41186 20688 41250 20692
rect 66838 20620 66902 20684
rect 31510 20212 31574 20276
rect 6314 20204 6378 20208
rect 6314 20148 6318 20204
rect 6318 20148 6374 20204
rect 6374 20148 6378 20204
rect 6314 20144 6378 20148
rect 6394 20204 6458 20208
rect 6394 20148 6398 20204
rect 6398 20148 6454 20204
rect 6454 20148 6458 20204
rect 6394 20144 6458 20148
rect 6474 20204 6538 20208
rect 6474 20148 6478 20204
rect 6478 20148 6534 20204
rect 6534 20148 6538 20204
rect 6474 20144 6538 20148
rect 6554 20204 6618 20208
rect 6554 20148 6558 20204
rect 6558 20148 6614 20204
rect 6614 20148 6618 20204
rect 6554 20144 6618 20148
rect 38282 20204 38346 20208
rect 38282 20148 38286 20204
rect 38286 20148 38342 20204
rect 38342 20148 38346 20204
rect 38282 20144 38346 20148
rect 38362 20204 38426 20208
rect 38362 20148 38366 20204
rect 38366 20148 38422 20204
rect 38422 20148 38426 20204
rect 38362 20144 38426 20148
rect 38442 20204 38506 20208
rect 38442 20148 38446 20204
rect 38446 20148 38502 20204
rect 38502 20148 38506 20204
rect 38442 20144 38506 20148
rect 38522 20204 38586 20208
rect 38522 20148 38526 20204
rect 38526 20148 38582 20204
rect 38582 20148 38586 20204
rect 38522 20144 38586 20148
rect 6854 20000 6918 20004
rect 6854 19944 6868 20000
rect 6868 19944 6918 20000
rect 6854 19940 6918 19944
rect 41630 19940 41694 20004
rect 67022 19940 67086 20004
rect 3650 19660 3714 19664
rect 3650 19604 3654 19660
rect 3654 19604 3710 19660
rect 3710 19604 3714 19660
rect 3650 19600 3714 19604
rect 3730 19660 3794 19664
rect 3730 19604 3734 19660
rect 3734 19604 3790 19660
rect 3790 19604 3794 19660
rect 3730 19600 3794 19604
rect 3810 19660 3874 19664
rect 3810 19604 3814 19660
rect 3814 19604 3870 19660
rect 3870 19604 3874 19660
rect 3810 19600 3874 19604
rect 3890 19660 3954 19664
rect 3890 19604 3894 19660
rect 3894 19604 3950 19660
rect 3950 19604 3954 19660
rect 3890 19600 3954 19604
rect 35618 19660 35682 19664
rect 35618 19604 35622 19660
rect 35622 19604 35678 19660
rect 35678 19604 35682 19660
rect 35618 19600 35682 19604
rect 35698 19660 35762 19664
rect 35698 19604 35702 19660
rect 35702 19604 35758 19660
rect 35758 19604 35762 19660
rect 35698 19600 35762 19604
rect 35778 19660 35842 19664
rect 35778 19604 35782 19660
rect 35782 19604 35838 19660
rect 35838 19604 35842 19660
rect 35778 19600 35842 19604
rect 35858 19660 35922 19664
rect 35858 19604 35862 19660
rect 35862 19604 35918 19660
rect 35918 19604 35922 19660
rect 35858 19600 35922 19604
rect 40946 19660 41010 19664
rect 40946 19604 40950 19660
rect 40950 19604 41006 19660
rect 41006 19604 41010 19660
rect 40946 19600 41010 19604
rect 41026 19660 41090 19664
rect 41026 19604 41030 19660
rect 41030 19604 41086 19660
rect 41086 19604 41090 19660
rect 41026 19600 41090 19604
rect 41106 19660 41170 19664
rect 41106 19604 41110 19660
rect 41110 19604 41166 19660
rect 41166 19604 41170 19660
rect 41106 19600 41170 19604
rect 41186 19660 41250 19664
rect 41186 19604 41190 19660
rect 41190 19604 41246 19660
rect 41246 19604 41250 19660
rect 41186 19600 41250 19604
rect 4278 19260 4342 19324
rect 31510 19124 31574 19188
rect 6314 19116 6378 19120
rect 6314 19060 6318 19116
rect 6318 19060 6374 19116
rect 6374 19060 6378 19116
rect 6314 19056 6378 19060
rect 6394 19116 6458 19120
rect 6394 19060 6398 19116
rect 6398 19060 6454 19116
rect 6454 19060 6458 19116
rect 6394 19056 6458 19060
rect 6474 19116 6538 19120
rect 6474 19060 6478 19116
rect 6478 19060 6534 19116
rect 6534 19060 6538 19116
rect 6474 19056 6538 19060
rect 6554 19116 6618 19120
rect 6554 19060 6558 19116
rect 6558 19060 6614 19116
rect 6614 19060 6618 19116
rect 6554 19056 6618 19060
rect 38282 19116 38346 19120
rect 38282 19060 38286 19116
rect 38286 19060 38342 19116
rect 38342 19060 38346 19116
rect 38282 19056 38346 19060
rect 38362 19116 38426 19120
rect 38362 19060 38366 19116
rect 38366 19060 38422 19116
rect 38422 19060 38426 19116
rect 38362 19056 38426 19060
rect 38442 19116 38506 19120
rect 38442 19060 38446 19116
rect 38446 19060 38502 19116
rect 38502 19060 38506 19116
rect 38442 19056 38506 19060
rect 38522 19116 38586 19120
rect 38522 19060 38526 19116
rect 38526 19060 38582 19116
rect 38582 19060 38586 19116
rect 38522 19056 38586 19060
rect 3650 18572 3714 18576
rect 3650 18516 3654 18572
rect 3654 18516 3710 18572
rect 3710 18516 3714 18572
rect 3650 18512 3714 18516
rect 3730 18572 3794 18576
rect 3730 18516 3734 18572
rect 3734 18516 3790 18572
rect 3790 18516 3794 18572
rect 3730 18512 3794 18516
rect 3810 18572 3874 18576
rect 3810 18516 3814 18572
rect 3814 18516 3870 18572
rect 3870 18516 3874 18572
rect 3810 18512 3874 18516
rect 3890 18572 3954 18576
rect 3890 18516 3894 18572
rect 3894 18516 3950 18572
rect 3950 18516 3954 18572
rect 3890 18512 3954 18516
rect 35618 18572 35682 18576
rect 35618 18516 35622 18572
rect 35622 18516 35678 18572
rect 35678 18516 35682 18572
rect 35618 18512 35682 18516
rect 35698 18572 35762 18576
rect 35698 18516 35702 18572
rect 35702 18516 35758 18572
rect 35758 18516 35762 18572
rect 35698 18512 35762 18516
rect 35778 18572 35842 18576
rect 35778 18516 35782 18572
rect 35782 18516 35838 18572
rect 35838 18516 35842 18572
rect 35778 18512 35842 18516
rect 35858 18572 35922 18576
rect 35858 18516 35862 18572
rect 35862 18516 35918 18572
rect 35918 18516 35922 18572
rect 35858 18512 35922 18516
rect 40946 18572 41010 18576
rect 40946 18516 40950 18572
rect 40950 18516 41006 18572
rect 41006 18516 41010 18572
rect 40946 18512 41010 18516
rect 41026 18572 41090 18576
rect 41026 18516 41030 18572
rect 41030 18516 41086 18572
rect 41086 18516 41090 18572
rect 41026 18512 41090 18516
rect 41106 18572 41170 18576
rect 41106 18516 41110 18572
rect 41110 18516 41166 18572
rect 41166 18516 41170 18572
rect 41106 18512 41170 18516
rect 41186 18572 41250 18576
rect 41186 18516 41190 18572
rect 41190 18516 41246 18572
rect 41246 18516 41250 18572
rect 41186 18512 41250 18516
rect 31510 18036 31574 18100
rect 6314 18028 6378 18032
rect 6314 17972 6318 18028
rect 6318 17972 6374 18028
rect 6374 17972 6378 18028
rect 6314 17968 6378 17972
rect 6394 18028 6458 18032
rect 6394 17972 6398 18028
rect 6398 17972 6454 18028
rect 6454 17972 6458 18028
rect 6394 17968 6458 17972
rect 6474 18028 6538 18032
rect 6474 17972 6478 18028
rect 6478 17972 6534 18028
rect 6534 17972 6538 18028
rect 6474 17968 6538 17972
rect 6554 18028 6618 18032
rect 6554 17972 6558 18028
rect 6558 17972 6614 18028
rect 6614 17972 6618 18028
rect 6554 17968 6618 17972
rect 38282 18028 38346 18032
rect 38282 17972 38286 18028
rect 38286 17972 38342 18028
rect 38342 17972 38346 18028
rect 38282 17968 38346 17972
rect 38362 18028 38426 18032
rect 38362 17972 38366 18028
rect 38366 17972 38422 18028
rect 38422 17972 38426 18028
rect 38362 17968 38426 17972
rect 38442 18028 38506 18032
rect 38442 17972 38446 18028
rect 38446 17972 38502 18028
rect 38502 17972 38506 18028
rect 38442 17968 38506 17972
rect 38522 18028 38586 18032
rect 38522 17972 38526 18028
rect 38526 17972 38582 18028
rect 38582 17972 38586 18028
rect 38522 17968 38586 17972
rect 41998 17960 42062 17964
rect 41998 17904 42048 17960
rect 42048 17904 42062 17960
rect 41998 17900 42062 17904
rect 67758 17900 67822 17964
rect 7406 17492 7470 17556
rect 3650 17484 3714 17488
rect 3650 17428 3654 17484
rect 3654 17428 3710 17484
rect 3710 17428 3714 17484
rect 3650 17424 3714 17428
rect 3730 17484 3794 17488
rect 3730 17428 3734 17484
rect 3734 17428 3790 17484
rect 3790 17428 3794 17484
rect 3730 17424 3794 17428
rect 3810 17484 3874 17488
rect 3810 17428 3814 17484
rect 3814 17428 3870 17484
rect 3870 17428 3874 17484
rect 3810 17424 3874 17428
rect 3890 17484 3954 17488
rect 3890 17428 3894 17484
rect 3894 17428 3950 17484
rect 3950 17428 3954 17484
rect 3890 17424 3954 17428
rect 35618 17484 35682 17488
rect 35618 17428 35622 17484
rect 35622 17428 35678 17484
rect 35678 17428 35682 17484
rect 35618 17424 35682 17428
rect 35698 17484 35762 17488
rect 35698 17428 35702 17484
rect 35702 17428 35758 17484
rect 35758 17428 35762 17484
rect 35698 17424 35762 17428
rect 35778 17484 35842 17488
rect 35778 17428 35782 17484
rect 35782 17428 35838 17484
rect 35838 17428 35842 17484
rect 35778 17424 35842 17428
rect 35858 17484 35922 17488
rect 35858 17428 35862 17484
rect 35862 17428 35918 17484
rect 35918 17428 35922 17484
rect 35858 17424 35922 17428
rect 40946 17484 41010 17488
rect 40946 17428 40950 17484
rect 40950 17428 41006 17484
rect 41006 17428 41010 17484
rect 40946 17424 41010 17428
rect 41026 17484 41090 17488
rect 41026 17428 41030 17484
rect 41030 17428 41086 17484
rect 41086 17428 41090 17484
rect 41026 17424 41090 17428
rect 41106 17484 41170 17488
rect 41106 17428 41110 17484
rect 41110 17428 41166 17484
rect 41166 17428 41170 17484
rect 41106 17424 41170 17428
rect 41186 17484 41250 17488
rect 41186 17428 41190 17484
rect 41190 17428 41246 17484
rect 41246 17428 41250 17484
rect 41186 17424 41250 17428
rect 5198 17220 5262 17284
rect 31510 16948 31574 17012
rect 6314 16940 6378 16944
rect 6314 16884 6318 16940
rect 6318 16884 6374 16940
rect 6374 16884 6378 16940
rect 6314 16880 6378 16884
rect 6394 16940 6458 16944
rect 6394 16884 6398 16940
rect 6398 16884 6454 16940
rect 6454 16884 6458 16940
rect 6394 16880 6458 16884
rect 6474 16940 6538 16944
rect 6474 16884 6478 16940
rect 6478 16884 6534 16940
rect 6534 16884 6538 16940
rect 6474 16880 6538 16884
rect 6554 16940 6618 16944
rect 6554 16884 6558 16940
rect 6558 16884 6614 16940
rect 6614 16884 6618 16940
rect 6554 16880 6618 16884
rect 38282 16940 38346 16944
rect 38282 16884 38286 16940
rect 38286 16884 38342 16940
rect 38342 16884 38346 16940
rect 38282 16880 38346 16884
rect 38362 16940 38426 16944
rect 38362 16884 38366 16940
rect 38366 16884 38422 16940
rect 38422 16884 38426 16940
rect 38362 16880 38426 16884
rect 38442 16940 38506 16944
rect 38442 16884 38446 16940
rect 38446 16884 38502 16940
rect 38502 16884 38506 16940
rect 38442 16880 38506 16884
rect 38522 16940 38586 16944
rect 38522 16884 38526 16940
rect 38526 16884 38582 16940
rect 38582 16884 38586 16940
rect 38522 16880 38586 16884
rect 5750 16600 5814 16604
rect 5750 16544 5764 16600
rect 5764 16544 5814 16600
rect 5750 16540 5814 16544
rect 36294 16600 36358 16604
rect 36294 16544 36344 16600
rect 36344 16544 36358 16600
rect 36294 16540 36358 16544
rect 41814 16540 41878 16604
rect 68310 16600 68374 16604
rect 68310 16544 68360 16600
rect 68360 16544 68374 16600
rect 68310 16540 68374 16544
rect 3650 16396 3714 16400
rect 3650 16340 3654 16396
rect 3654 16340 3710 16396
rect 3710 16340 3714 16396
rect 3650 16336 3714 16340
rect 3730 16396 3794 16400
rect 3730 16340 3734 16396
rect 3734 16340 3790 16396
rect 3790 16340 3794 16396
rect 3730 16336 3794 16340
rect 3810 16396 3874 16400
rect 3810 16340 3814 16396
rect 3814 16340 3870 16396
rect 3870 16340 3874 16396
rect 3810 16336 3874 16340
rect 3890 16396 3954 16400
rect 3890 16340 3894 16396
rect 3894 16340 3950 16396
rect 3950 16340 3954 16396
rect 3890 16336 3954 16340
rect 35618 16396 35682 16400
rect 35618 16340 35622 16396
rect 35622 16340 35678 16396
rect 35678 16340 35682 16396
rect 35618 16336 35682 16340
rect 35698 16396 35762 16400
rect 35698 16340 35702 16396
rect 35702 16340 35758 16396
rect 35758 16340 35762 16396
rect 35698 16336 35762 16340
rect 35778 16396 35842 16400
rect 35778 16340 35782 16396
rect 35782 16340 35838 16396
rect 35838 16340 35842 16396
rect 35778 16336 35842 16340
rect 35858 16396 35922 16400
rect 35858 16340 35862 16396
rect 35862 16340 35918 16396
rect 35918 16340 35922 16396
rect 35858 16336 35922 16340
rect 40946 16396 41010 16400
rect 40946 16340 40950 16396
rect 40950 16340 41006 16396
rect 41006 16340 41010 16396
rect 40946 16336 41010 16340
rect 41026 16396 41090 16400
rect 41026 16340 41030 16396
rect 41030 16340 41086 16396
rect 41086 16340 41090 16396
rect 41026 16336 41090 16340
rect 41106 16396 41170 16400
rect 41106 16340 41110 16396
rect 41110 16340 41166 16396
rect 41166 16340 41170 16396
rect 41106 16336 41170 16340
rect 41186 16396 41250 16400
rect 41186 16340 41190 16396
rect 41190 16340 41246 16396
rect 41246 16340 41250 16396
rect 41186 16336 41250 16340
rect 6314 15852 6378 15856
rect 6314 15796 6318 15852
rect 6318 15796 6374 15852
rect 6374 15796 6378 15852
rect 6314 15792 6378 15796
rect 6394 15852 6458 15856
rect 6394 15796 6398 15852
rect 6398 15796 6454 15852
rect 6454 15796 6458 15852
rect 6394 15792 6458 15796
rect 6474 15852 6538 15856
rect 6474 15796 6478 15852
rect 6478 15796 6534 15852
rect 6534 15796 6538 15852
rect 6474 15792 6538 15796
rect 6554 15852 6618 15856
rect 6554 15796 6558 15852
rect 6558 15796 6614 15852
rect 6614 15796 6618 15852
rect 6554 15792 6618 15796
rect 38282 15852 38346 15856
rect 38282 15796 38286 15852
rect 38286 15796 38342 15852
rect 38342 15796 38346 15852
rect 38282 15792 38346 15796
rect 38362 15852 38426 15856
rect 38362 15796 38366 15852
rect 38366 15796 38422 15852
rect 38422 15796 38426 15852
rect 38362 15792 38426 15796
rect 38442 15852 38506 15856
rect 38442 15796 38446 15852
rect 38446 15796 38502 15852
rect 38502 15796 38506 15852
rect 38442 15792 38506 15796
rect 38522 15852 38586 15856
rect 38522 15796 38526 15852
rect 38526 15796 38582 15852
rect 38582 15796 38586 15852
rect 38522 15792 38586 15796
rect 3650 15308 3714 15312
rect 3650 15252 3654 15308
rect 3654 15252 3710 15308
rect 3710 15252 3714 15308
rect 3650 15248 3714 15252
rect 3730 15308 3794 15312
rect 3730 15252 3734 15308
rect 3734 15252 3790 15308
rect 3790 15252 3794 15308
rect 3730 15248 3794 15252
rect 3810 15308 3874 15312
rect 3810 15252 3814 15308
rect 3814 15252 3870 15308
rect 3870 15252 3874 15308
rect 3810 15248 3874 15252
rect 3890 15308 3954 15312
rect 3890 15252 3894 15308
rect 3894 15252 3950 15308
rect 3950 15252 3954 15308
rect 3890 15248 3954 15252
rect 35618 15308 35682 15312
rect 35618 15252 35622 15308
rect 35622 15252 35678 15308
rect 35678 15252 35682 15308
rect 35618 15248 35682 15252
rect 35698 15308 35762 15312
rect 35698 15252 35702 15308
rect 35702 15252 35758 15308
rect 35758 15252 35762 15308
rect 35698 15248 35762 15252
rect 35778 15308 35842 15312
rect 35778 15252 35782 15308
rect 35782 15252 35838 15308
rect 35838 15252 35842 15308
rect 35778 15248 35842 15252
rect 35858 15308 35922 15312
rect 35858 15252 35862 15308
rect 35862 15252 35918 15308
rect 35918 15252 35922 15308
rect 35858 15248 35922 15252
rect 40946 15308 41010 15312
rect 40946 15252 40950 15308
rect 40950 15252 41006 15308
rect 41006 15252 41010 15308
rect 40946 15248 41010 15252
rect 41026 15308 41090 15312
rect 41026 15252 41030 15308
rect 41030 15252 41086 15308
rect 41086 15252 41090 15308
rect 41026 15248 41090 15252
rect 41106 15308 41170 15312
rect 41106 15252 41110 15308
rect 41110 15252 41166 15308
rect 41166 15252 41170 15308
rect 41106 15248 41170 15252
rect 41186 15308 41250 15312
rect 41186 15252 41190 15308
rect 41190 15252 41246 15308
rect 41246 15252 41250 15308
rect 41186 15248 41250 15252
rect 7222 15180 7286 15244
rect 31510 14772 31574 14836
rect 6314 14764 6378 14768
rect 6314 14708 6318 14764
rect 6318 14708 6374 14764
rect 6374 14708 6378 14764
rect 6314 14704 6378 14708
rect 6394 14764 6458 14768
rect 6394 14708 6398 14764
rect 6398 14708 6454 14764
rect 6454 14708 6458 14764
rect 6394 14704 6458 14708
rect 6474 14764 6538 14768
rect 6474 14708 6478 14764
rect 6478 14708 6534 14764
rect 6534 14708 6538 14764
rect 6474 14704 6538 14708
rect 6554 14764 6618 14768
rect 6554 14708 6558 14764
rect 6558 14708 6614 14764
rect 6614 14708 6618 14764
rect 6554 14704 6618 14708
rect 38282 14764 38346 14768
rect 38282 14708 38286 14764
rect 38286 14708 38342 14764
rect 38342 14708 38346 14764
rect 38282 14704 38346 14708
rect 38362 14764 38426 14768
rect 38362 14708 38366 14764
rect 38366 14708 38422 14764
rect 38422 14708 38426 14764
rect 38362 14704 38426 14708
rect 38442 14764 38506 14768
rect 38442 14708 38446 14764
rect 38446 14708 38502 14764
rect 38502 14708 38506 14764
rect 38442 14704 38506 14708
rect 38522 14764 38586 14768
rect 38522 14708 38526 14764
rect 38526 14708 38582 14764
rect 38582 14708 38586 14764
rect 38522 14704 38586 14708
rect 7406 14560 7470 14564
rect 7406 14504 7420 14560
rect 7420 14504 7470 14560
rect 7406 14500 7470 14504
rect 3650 14220 3714 14224
rect 3650 14164 3654 14220
rect 3654 14164 3710 14220
rect 3710 14164 3714 14220
rect 3650 14160 3714 14164
rect 3730 14220 3794 14224
rect 3730 14164 3734 14220
rect 3734 14164 3790 14220
rect 3790 14164 3794 14220
rect 3730 14160 3794 14164
rect 3810 14220 3874 14224
rect 3810 14164 3814 14220
rect 3814 14164 3870 14220
rect 3870 14164 3874 14220
rect 3810 14160 3874 14164
rect 3890 14220 3954 14224
rect 3890 14164 3894 14220
rect 3894 14164 3950 14220
rect 3950 14164 3954 14220
rect 3890 14160 3954 14164
rect 35618 14220 35682 14224
rect 35618 14164 35622 14220
rect 35622 14164 35678 14220
rect 35678 14164 35682 14220
rect 35618 14160 35682 14164
rect 35698 14220 35762 14224
rect 35698 14164 35702 14220
rect 35702 14164 35758 14220
rect 35758 14164 35762 14220
rect 35698 14160 35762 14164
rect 35778 14220 35842 14224
rect 35778 14164 35782 14220
rect 35782 14164 35838 14220
rect 35838 14164 35842 14220
rect 35778 14160 35842 14164
rect 35858 14220 35922 14224
rect 35858 14164 35862 14220
rect 35862 14164 35918 14220
rect 35918 14164 35922 14220
rect 35858 14160 35922 14164
rect 40946 14220 41010 14224
rect 40946 14164 40950 14220
rect 40950 14164 41006 14220
rect 41006 14164 41010 14220
rect 40946 14160 41010 14164
rect 41026 14220 41090 14224
rect 41026 14164 41030 14220
rect 41030 14164 41086 14220
rect 41086 14164 41090 14220
rect 41026 14160 41090 14164
rect 41106 14220 41170 14224
rect 41106 14164 41110 14220
rect 41110 14164 41166 14220
rect 41166 14164 41170 14220
rect 41106 14160 41170 14164
rect 41186 14220 41250 14224
rect 41186 14164 41190 14220
rect 41190 14164 41246 14220
rect 41246 14164 41250 14220
rect 41186 14160 41250 14164
rect 6314 13676 6378 13680
rect 6314 13620 6318 13676
rect 6318 13620 6374 13676
rect 6374 13620 6378 13676
rect 6314 13616 6378 13620
rect 6394 13676 6458 13680
rect 6394 13620 6398 13676
rect 6398 13620 6454 13676
rect 6454 13620 6458 13676
rect 6394 13616 6458 13620
rect 6474 13676 6538 13680
rect 6474 13620 6478 13676
rect 6478 13620 6534 13676
rect 6534 13620 6538 13676
rect 6474 13616 6538 13620
rect 6554 13676 6618 13680
rect 6554 13620 6558 13676
rect 6558 13620 6614 13676
rect 6614 13620 6618 13676
rect 6554 13616 6618 13620
rect 38282 13676 38346 13680
rect 38282 13620 38286 13676
rect 38286 13620 38342 13676
rect 38342 13620 38346 13676
rect 38282 13616 38346 13620
rect 38362 13676 38426 13680
rect 38362 13620 38366 13676
rect 38366 13620 38422 13676
rect 38422 13620 38426 13676
rect 38362 13616 38426 13620
rect 38442 13676 38506 13680
rect 38442 13620 38446 13676
rect 38446 13620 38502 13676
rect 38502 13620 38506 13676
rect 38442 13616 38506 13620
rect 38522 13676 38586 13680
rect 38522 13620 38526 13676
rect 38526 13620 38582 13676
rect 38582 13620 38586 13676
rect 38522 13616 38586 13620
rect 3650 13132 3714 13136
rect 3650 13076 3654 13132
rect 3654 13076 3710 13132
rect 3710 13076 3714 13132
rect 3650 13072 3714 13076
rect 3730 13132 3794 13136
rect 3730 13076 3734 13132
rect 3734 13076 3790 13132
rect 3790 13076 3794 13132
rect 3730 13072 3794 13076
rect 3810 13132 3874 13136
rect 3810 13076 3814 13132
rect 3814 13076 3870 13132
rect 3870 13076 3874 13132
rect 3810 13072 3874 13076
rect 3890 13132 3954 13136
rect 3890 13076 3894 13132
rect 3894 13076 3950 13132
rect 3950 13076 3954 13132
rect 3890 13072 3954 13076
rect 35618 13132 35682 13136
rect 35618 13076 35622 13132
rect 35622 13076 35678 13132
rect 35678 13076 35682 13132
rect 35618 13072 35682 13076
rect 35698 13132 35762 13136
rect 35698 13076 35702 13132
rect 35702 13076 35758 13132
rect 35758 13076 35762 13132
rect 35698 13072 35762 13076
rect 35778 13132 35842 13136
rect 35778 13076 35782 13132
rect 35782 13076 35838 13132
rect 35838 13076 35842 13132
rect 35778 13072 35842 13076
rect 35858 13132 35922 13136
rect 35858 13076 35862 13132
rect 35862 13076 35918 13132
rect 35918 13076 35922 13132
rect 35858 13072 35922 13076
rect 40946 13132 41010 13136
rect 40946 13076 40950 13132
rect 40950 13076 41006 13132
rect 41006 13076 41010 13132
rect 40946 13072 41010 13076
rect 41026 13132 41090 13136
rect 41026 13076 41030 13132
rect 41030 13076 41086 13132
rect 41086 13076 41090 13132
rect 41026 13072 41090 13076
rect 41106 13132 41170 13136
rect 41106 13076 41110 13132
rect 41110 13076 41166 13132
rect 41166 13076 41170 13132
rect 41106 13072 41170 13076
rect 41186 13132 41250 13136
rect 41186 13076 41190 13132
rect 41190 13076 41246 13132
rect 41246 13076 41250 13132
rect 41186 13072 41250 13076
rect 6314 12588 6378 12592
rect 6314 12532 6318 12588
rect 6318 12532 6374 12588
rect 6374 12532 6378 12588
rect 6314 12528 6378 12532
rect 6394 12588 6458 12592
rect 6394 12532 6398 12588
rect 6398 12532 6454 12588
rect 6454 12532 6458 12588
rect 6394 12528 6458 12532
rect 6474 12588 6538 12592
rect 6474 12532 6478 12588
rect 6478 12532 6534 12588
rect 6534 12532 6538 12588
rect 6474 12528 6538 12532
rect 6554 12588 6618 12592
rect 6554 12532 6558 12588
rect 6558 12532 6614 12588
rect 6614 12532 6618 12588
rect 6554 12528 6618 12532
rect 38282 12588 38346 12592
rect 38282 12532 38286 12588
rect 38286 12532 38342 12588
rect 38342 12532 38346 12588
rect 38282 12528 38346 12532
rect 38362 12588 38426 12592
rect 38362 12532 38366 12588
rect 38366 12532 38422 12588
rect 38422 12532 38426 12588
rect 38362 12528 38426 12532
rect 38442 12588 38506 12592
rect 38442 12532 38446 12588
rect 38446 12532 38502 12588
rect 38502 12532 38506 12588
rect 38442 12528 38506 12532
rect 38522 12588 38586 12592
rect 38522 12532 38526 12588
rect 38526 12532 38582 12588
rect 38582 12532 38586 12588
rect 38522 12528 38586 12532
rect 3650 12044 3714 12048
rect 3650 11988 3654 12044
rect 3654 11988 3710 12044
rect 3710 11988 3714 12044
rect 3650 11984 3714 11988
rect 3730 12044 3794 12048
rect 3730 11988 3734 12044
rect 3734 11988 3790 12044
rect 3790 11988 3794 12044
rect 3730 11984 3794 11988
rect 3810 12044 3874 12048
rect 3810 11988 3814 12044
rect 3814 11988 3870 12044
rect 3870 11988 3874 12044
rect 3810 11984 3874 11988
rect 3890 12044 3954 12048
rect 3890 11988 3894 12044
rect 3894 11988 3950 12044
rect 3950 11988 3954 12044
rect 3890 11984 3954 11988
rect 35618 12044 35682 12048
rect 35618 11988 35622 12044
rect 35622 11988 35678 12044
rect 35678 11988 35682 12044
rect 35618 11984 35682 11988
rect 35698 12044 35762 12048
rect 35698 11988 35702 12044
rect 35702 11988 35758 12044
rect 35758 11988 35762 12044
rect 35698 11984 35762 11988
rect 35778 12044 35842 12048
rect 35778 11988 35782 12044
rect 35782 11988 35838 12044
rect 35838 11988 35842 12044
rect 35778 11984 35842 11988
rect 35858 12044 35922 12048
rect 35858 11988 35862 12044
rect 35862 11988 35918 12044
rect 35918 11988 35922 12044
rect 35858 11984 35922 11988
rect 40946 12044 41010 12048
rect 40946 11988 40950 12044
rect 40950 11988 41006 12044
rect 41006 11988 41010 12044
rect 40946 11984 41010 11988
rect 41026 12044 41090 12048
rect 41026 11988 41030 12044
rect 41030 11988 41086 12044
rect 41086 11988 41090 12044
rect 41026 11984 41090 11988
rect 41106 12044 41170 12048
rect 41106 11988 41110 12044
rect 41110 11988 41166 12044
rect 41166 11988 41170 12044
rect 41106 11984 41170 11988
rect 41186 12044 41250 12048
rect 41186 11988 41190 12044
rect 41190 11988 41246 12044
rect 41246 11988 41250 12044
rect 41186 11984 41250 11988
rect 6314 11500 6378 11504
rect 6314 11444 6318 11500
rect 6318 11444 6374 11500
rect 6374 11444 6378 11500
rect 6314 11440 6378 11444
rect 6394 11500 6458 11504
rect 6394 11444 6398 11500
rect 6398 11444 6454 11500
rect 6454 11444 6458 11500
rect 6394 11440 6458 11444
rect 6474 11500 6538 11504
rect 6474 11444 6478 11500
rect 6478 11444 6534 11500
rect 6534 11444 6538 11500
rect 6474 11440 6538 11444
rect 6554 11500 6618 11504
rect 6554 11444 6558 11500
rect 6558 11444 6614 11500
rect 6614 11444 6618 11500
rect 6554 11440 6618 11444
rect 38282 11500 38346 11504
rect 38282 11444 38286 11500
rect 38286 11444 38342 11500
rect 38342 11444 38346 11500
rect 38282 11440 38346 11444
rect 38362 11500 38426 11504
rect 38362 11444 38366 11500
rect 38366 11444 38422 11500
rect 38422 11444 38426 11500
rect 38362 11440 38426 11444
rect 38442 11500 38506 11504
rect 38442 11444 38446 11500
rect 38446 11444 38502 11500
rect 38502 11444 38506 11500
rect 38442 11440 38506 11444
rect 38522 11500 38586 11504
rect 38522 11444 38526 11500
rect 38526 11444 38582 11500
rect 38582 11444 38586 11500
rect 38522 11440 38586 11444
rect 3650 10956 3714 10960
rect 3650 10900 3654 10956
rect 3654 10900 3710 10956
rect 3710 10900 3714 10956
rect 3650 10896 3714 10900
rect 3730 10956 3794 10960
rect 3730 10900 3734 10956
rect 3734 10900 3790 10956
rect 3790 10900 3794 10956
rect 3730 10896 3794 10900
rect 3810 10956 3874 10960
rect 3810 10900 3814 10956
rect 3814 10900 3870 10956
rect 3870 10900 3874 10956
rect 3810 10896 3874 10900
rect 3890 10956 3954 10960
rect 3890 10900 3894 10956
rect 3894 10900 3950 10956
rect 3950 10900 3954 10956
rect 3890 10896 3954 10900
rect 35618 10956 35682 10960
rect 35618 10900 35622 10956
rect 35622 10900 35678 10956
rect 35678 10900 35682 10956
rect 35618 10896 35682 10900
rect 35698 10956 35762 10960
rect 35698 10900 35702 10956
rect 35702 10900 35758 10956
rect 35758 10900 35762 10956
rect 35698 10896 35762 10900
rect 35778 10956 35842 10960
rect 35778 10900 35782 10956
rect 35782 10900 35838 10956
rect 35838 10900 35842 10956
rect 35778 10896 35842 10900
rect 35858 10956 35922 10960
rect 35858 10900 35862 10956
rect 35862 10900 35918 10956
rect 35918 10900 35922 10956
rect 35858 10896 35922 10900
rect 40946 10956 41010 10960
rect 40946 10900 40950 10956
rect 40950 10900 41006 10956
rect 41006 10900 41010 10956
rect 40946 10896 41010 10900
rect 41026 10956 41090 10960
rect 41026 10900 41030 10956
rect 41030 10900 41086 10956
rect 41086 10900 41090 10956
rect 41026 10896 41090 10900
rect 41106 10956 41170 10960
rect 41106 10900 41110 10956
rect 41110 10900 41166 10956
rect 41166 10900 41170 10956
rect 41106 10896 41170 10900
rect 41186 10956 41250 10960
rect 41186 10900 41190 10956
rect 41190 10900 41246 10956
rect 41246 10900 41250 10956
rect 41186 10896 41250 10900
rect 31510 10420 31574 10484
rect 6314 10412 6378 10416
rect 6314 10356 6318 10412
rect 6318 10356 6374 10412
rect 6374 10356 6378 10412
rect 6314 10352 6378 10356
rect 6394 10412 6458 10416
rect 6394 10356 6398 10412
rect 6398 10356 6454 10412
rect 6454 10356 6458 10412
rect 6394 10352 6458 10356
rect 6474 10412 6538 10416
rect 6474 10356 6478 10412
rect 6478 10356 6534 10412
rect 6534 10356 6538 10412
rect 6474 10352 6538 10356
rect 6554 10412 6618 10416
rect 6554 10356 6558 10412
rect 6558 10356 6614 10412
rect 6614 10356 6618 10412
rect 6554 10352 6618 10356
rect 38282 10412 38346 10416
rect 38282 10356 38286 10412
rect 38286 10356 38342 10412
rect 38342 10356 38346 10412
rect 38282 10352 38346 10356
rect 38362 10412 38426 10416
rect 38362 10356 38366 10412
rect 38366 10356 38422 10412
rect 38422 10356 38426 10412
rect 38362 10352 38426 10356
rect 38442 10412 38506 10416
rect 38442 10356 38446 10412
rect 38446 10356 38502 10412
rect 38502 10356 38506 10412
rect 38442 10352 38506 10356
rect 38522 10412 38586 10416
rect 38522 10356 38526 10412
rect 38526 10356 38582 10412
rect 38582 10356 38586 10412
rect 38522 10352 38586 10356
rect 3650 9868 3714 9872
rect 3650 9812 3654 9868
rect 3654 9812 3710 9868
rect 3710 9812 3714 9868
rect 3650 9808 3714 9812
rect 3730 9868 3794 9872
rect 3730 9812 3734 9868
rect 3734 9812 3790 9868
rect 3790 9812 3794 9868
rect 3730 9808 3794 9812
rect 3810 9868 3874 9872
rect 3810 9812 3814 9868
rect 3814 9812 3870 9868
rect 3870 9812 3874 9868
rect 3810 9808 3874 9812
rect 3890 9868 3954 9872
rect 3890 9812 3894 9868
rect 3894 9812 3950 9868
rect 3950 9812 3954 9868
rect 3890 9808 3954 9812
rect 35618 9868 35682 9872
rect 35618 9812 35622 9868
rect 35622 9812 35678 9868
rect 35678 9812 35682 9868
rect 35618 9808 35682 9812
rect 35698 9868 35762 9872
rect 35698 9812 35702 9868
rect 35702 9812 35758 9868
rect 35758 9812 35762 9868
rect 35698 9808 35762 9812
rect 35778 9868 35842 9872
rect 35778 9812 35782 9868
rect 35782 9812 35838 9868
rect 35838 9812 35842 9868
rect 35778 9808 35842 9812
rect 35858 9868 35922 9872
rect 35858 9812 35862 9868
rect 35862 9812 35918 9868
rect 35918 9812 35922 9868
rect 35858 9808 35922 9812
rect 40946 9868 41010 9872
rect 40946 9812 40950 9868
rect 40950 9812 41006 9868
rect 41006 9812 41010 9868
rect 40946 9808 41010 9812
rect 41026 9868 41090 9872
rect 41026 9812 41030 9868
rect 41030 9812 41086 9868
rect 41086 9812 41090 9868
rect 41026 9808 41090 9812
rect 41106 9868 41170 9872
rect 41106 9812 41110 9868
rect 41110 9812 41166 9868
rect 41166 9812 41170 9868
rect 41106 9808 41170 9812
rect 41186 9868 41250 9872
rect 41186 9812 41190 9868
rect 41190 9812 41246 9868
rect 41246 9812 41250 9868
rect 41186 9808 41250 9812
rect 6314 9324 6378 9328
rect 6314 9268 6318 9324
rect 6318 9268 6374 9324
rect 6374 9268 6378 9324
rect 6314 9264 6378 9268
rect 6394 9324 6458 9328
rect 6394 9268 6398 9324
rect 6398 9268 6454 9324
rect 6454 9268 6458 9324
rect 6394 9264 6458 9268
rect 6474 9324 6538 9328
rect 6474 9268 6478 9324
rect 6478 9268 6534 9324
rect 6534 9268 6538 9324
rect 6474 9264 6538 9268
rect 6554 9324 6618 9328
rect 6554 9268 6558 9324
rect 6558 9268 6614 9324
rect 6614 9268 6618 9324
rect 6554 9264 6618 9268
rect 38282 9324 38346 9328
rect 38282 9268 38286 9324
rect 38286 9268 38342 9324
rect 38342 9268 38346 9324
rect 38282 9264 38346 9268
rect 38362 9324 38426 9328
rect 38362 9268 38366 9324
rect 38366 9268 38422 9324
rect 38422 9268 38426 9324
rect 38362 9264 38426 9268
rect 38442 9324 38506 9328
rect 38442 9268 38446 9324
rect 38446 9268 38502 9324
rect 38502 9268 38506 9324
rect 38442 9264 38506 9268
rect 38522 9324 38586 9328
rect 38522 9268 38526 9324
rect 38526 9268 38582 9324
rect 38582 9268 38586 9324
rect 38522 9264 38586 9268
rect 3650 8780 3714 8784
rect 3650 8724 3654 8780
rect 3654 8724 3710 8780
rect 3710 8724 3714 8780
rect 3650 8720 3714 8724
rect 3730 8780 3794 8784
rect 3730 8724 3734 8780
rect 3734 8724 3790 8780
rect 3790 8724 3794 8780
rect 3730 8720 3794 8724
rect 3810 8780 3874 8784
rect 3810 8724 3814 8780
rect 3814 8724 3870 8780
rect 3870 8724 3874 8780
rect 3810 8720 3874 8724
rect 3890 8780 3954 8784
rect 3890 8724 3894 8780
rect 3894 8724 3950 8780
rect 3950 8724 3954 8780
rect 3890 8720 3954 8724
rect 35618 8780 35682 8784
rect 35618 8724 35622 8780
rect 35622 8724 35678 8780
rect 35678 8724 35682 8780
rect 35618 8720 35682 8724
rect 35698 8780 35762 8784
rect 35698 8724 35702 8780
rect 35702 8724 35758 8780
rect 35758 8724 35762 8780
rect 35698 8720 35762 8724
rect 35778 8780 35842 8784
rect 35778 8724 35782 8780
rect 35782 8724 35838 8780
rect 35838 8724 35842 8780
rect 35778 8720 35842 8724
rect 35858 8780 35922 8784
rect 35858 8724 35862 8780
rect 35862 8724 35918 8780
rect 35918 8724 35922 8780
rect 35858 8720 35922 8724
rect 40946 8780 41010 8784
rect 40946 8724 40950 8780
rect 40950 8724 41006 8780
rect 41006 8724 41010 8780
rect 40946 8720 41010 8724
rect 41026 8780 41090 8784
rect 41026 8724 41030 8780
rect 41030 8724 41086 8780
rect 41086 8724 41090 8780
rect 41026 8720 41090 8724
rect 41106 8780 41170 8784
rect 41106 8724 41110 8780
rect 41110 8724 41166 8780
rect 41166 8724 41170 8780
rect 41106 8720 41170 8724
rect 41186 8780 41250 8784
rect 41186 8724 41190 8780
rect 41190 8724 41246 8780
rect 41246 8724 41250 8780
rect 41186 8720 41250 8724
rect 6314 8236 6378 8240
rect 6314 8180 6318 8236
rect 6318 8180 6374 8236
rect 6374 8180 6378 8236
rect 6314 8176 6378 8180
rect 6394 8236 6458 8240
rect 6394 8180 6398 8236
rect 6398 8180 6454 8236
rect 6454 8180 6458 8236
rect 6394 8176 6458 8180
rect 6474 8236 6538 8240
rect 6474 8180 6478 8236
rect 6478 8180 6534 8236
rect 6534 8180 6538 8236
rect 6474 8176 6538 8180
rect 6554 8236 6618 8240
rect 6554 8180 6558 8236
rect 6558 8180 6614 8236
rect 6614 8180 6618 8236
rect 6554 8176 6618 8180
rect 38282 8236 38346 8240
rect 38282 8180 38286 8236
rect 38286 8180 38342 8236
rect 38342 8180 38346 8236
rect 38282 8176 38346 8180
rect 38362 8236 38426 8240
rect 38362 8180 38366 8236
rect 38366 8180 38422 8236
rect 38422 8180 38426 8236
rect 38362 8176 38426 8180
rect 38442 8236 38506 8240
rect 38442 8180 38446 8236
rect 38446 8180 38502 8236
rect 38502 8180 38506 8236
rect 38442 8176 38506 8180
rect 38522 8236 38586 8240
rect 38522 8180 38526 8236
rect 38526 8180 38582 8236
rect 38582 8180 38586 8236
rect 38522 8176 38586 8180
rect 3650 7692 3714 7696
rect 3650 7636 3654 7692
rect 3654 7636 3710 7692
rect 3710 7636 3714 7692
rect 3650 7632 3714 7636
rect 3730 7692 3794 7696
rect 3730 7636 3734 7692
rect 3734 7636 3790 7692
rect 3790 7636 3794 7692
rect 3730 7632 3794 7636
rect 3810 7692 3874 7696
rect 3810 7636 3814 7692
rect 3814 7636 3870 7692
rect 3870 7636 3874 7692
rect 3810 7632 3874 7636
rect 3890 7692 3954 7696
rect 3890 7636 3894 7692
rect 3894 7636 3950 7692
rect 3950 7636 3954 7692
rect 3890 7632 3954 7636
rect 35618 7692 35682 7696
rect 35618 7636 35622 7692
rect 35622 7636 35678 7692
rect 35678 7636 35682 7692
rect 35618 7632 35682 7636
rect 35698 7692 35762 7696
rect 35698 7636 35702 7692
rect 35702 7636 35758 7692
rect 35758 7636 35762 7692
rect 35698 7632 35762 7636
rect 35778 7692 35842 7696
rect 35778 7636 35782 7692
rect 35782 7636 35838 7692
rect 35838 7636 35842 7692
rect 35778 7632 35842 7636
rect 35858 7692 35922 7696
rect 35858 7636 35862 7692
rect 35862 7636 35918 7692
rect 35918 7636 35922 7692
rect 35858 7632 35922 7636
rect 40946 7692 41010 7696
rect 40946 7636 40950 7692
rect 40950 7636 41006 7692
rect 41006 7636 41010 7692
rect 40946 7632 41010 7636
rect 41026 7692 41090 7696
rect 41026 7636 41030 7692
rect 41030 7636 41086 7692
rect 41086 7636 41090 7692
rect 41026 7632 41090 7636
rect 41106 7692 41170 7696
rect 41106 7636 41110 7692
rect 41110 7636 41166 7692
rect 41166 7636 41170 7692
rect 41106 7632 41170 7636
rect 41186 7692 41250 7696
rect 41186 7636 41190 7692
rect 41190 7636 41246 7692
rect 41246 7636 41250 7692
rect 41186 7632 41250 7636
rect 6314 7148 6378 7152
rect 6314 7092 6318 7148
rect 6318 7092 6374 7148
rect 6374 7092 6378 7148
rect 6314 7088 6378 7092
rect 6394 7148 6458 7152
rect 6394 7092 6398 7148
rect 6398 7092 6454 7148
rect 6454 7092 6458 7148
rect 6394 7088 6458 7092
rect 6474 7148 6538 7152
rect 6474 7092 6478 7148
rect 6478 7092 6534 7148
rect 6534 7092 6538 7148
rect 6474 7088 6538 7092
rect 6554 7148 6618 7152
rect 6554 7092 6558 7148
rect 6558 7092 6614 7148
rect 6614 7092 6618 7148
rect 6554 7088 6618 7092
rect 38282 7148 38346 7152
rect 38282 7092 38286 7148
rect 38286 7092 38342 7148
rect 38342 7092 38346 7148
rect 38282 7088 38346 7092
rect 38362 7148 38426 7152
rect 38362 7092 38366 7148
rect 38366 7092 38422 7148
rect 38422 7092 38426 7148
rect 38362 7088 38426 7092
rect 38442 7148 38506 7152
rect 38442 7092 38446 7148
rect 38446 7092 38502 7148
rect 38502 7092 38506 7148
rect 38442 7088 38506 7092
rect 38522 7148 38586 7152
rect 38522 7092 38526 7148
rect 38526 7092 38582 7148
rect 38582 7092 38586 7148
rect 38522 7088 38586 7092
rect 3650 6604 3714 6608
rect 3650 6548 3654 6604
rect 3654 6548 3710 6604
rect 3710 6548 3714 6604
rect 3650 6544 3714 6548
rect 3730 6604 3794 6608
rect 3730 6548 3734 6604
rect 3734 6548 3790 6604
rect 3790 6548 3794 6604
rect 3730 6544 3794 6548
rect 3810 6604 3874 6608
rect 3810 6548 3814 6604
rect 3814 6548 3870 6604
rect 3870 6548 3874 6604
rect 3810 6544 3874 6548
rect 3890 6604 3954 6608
rect 3890 6548 3894 6604
rect 3894 6548 3950 6604
rect 3950 6548 3954 6604
rect 3890 6544 3954 6548
rect 35618 6604 35682 6608
rect 35618 6548 35622 6604
rect 35622 6548 35678 6604
rect 35678 6548 35682 6604
rect 35618 6544 35682 6548
rect 35698 6604 35762 6608
rect 35698 6548 35702 6604
rect 35702 6548 35758 6604
rect 35758 6548 35762 6604
rect 35698 6544 35762 6548
rect 35778 6604 35842 6608
rect 35778 6548 35782 6604
rect 35782 6548 35838 6604
rect 35838 6548 35842 6604
rect 35778 6544 35842 6548
rect 35858 6604 35922 6608
rect 35858 6548 35862 6604
rect 35862 6548 35918 6604
rect 35918 6548 35922 6604
rect 35858 6544 35922 6548
rect 40946 6604 41010 6608
rect 40946 6548 40950 6604
rect 40950 6548 41006 6604
rect 41006 6548 41010 6604
rect 40946 6544 41010 6548
rect 41026 6604 41090 6608
rect 41026 6548 41030 6604
rect 41030 6548 41086 6604
rect 41086 6548 41090 6604
rect 41026 6544 41090 6548
rect 41106 6604 41170 6608
rect 41106 6548 41110 6604
rect 41110 6548 41166 6604
rect 41166 6548 41170 6604
rect 41106 6544 41170 6548
rect 41186 6604 41250 6608
rect 41186 6548 41190 6604
rect 41190 6548 41246 6604
rect 41246 6548 41250 6604
rect 41186 6544 41250 6548
rect 6314 6060 6378 6064
rect 6314 6004 6318 6060
rect 6318 6004 6374 6060
rect 6374 6004 6378 6060
rect 6314 6000 6378 6004
rect 6394 6060 6458 6064
rect 6394 6004 6398 6060
rect 6398 6004 6454 6060
rect 6454 6004 6458 6060
rect 6394 6000 6458 6004
rect 6474 6060 6538 6064
rect 6474 6004 6478 6060
rect 6478 6004 6534 6060
rect 6534 6004 6538 6060
rect 6474 6000 6538 6004
rect 6554 6060 6618 6064
rect 6554 6004 6558 6060
rect 6558 6004 6614 6060
rect 6614 6004 6618 6060
rect 6554 6000 6618 6004
rect 38282 6060 38346 6064
rect 38282 6004 38286 6060
rect 38286 6004 38342 6060
rect 38342 6004 38346 6060
rect 38282 6000 38346 6004
rect 38362 6060 38426 6064
rect 38362 6004 38366 6060
rect 38366 6004 38422 6060
rect 38422 6004 38426 6060
rect 38362 6000 38426 6004
rect 38442 6060 38506 6064
rect 38442 6004 38446 6060
rect 38446 6004 38502 6060
rect 38502 6004 38506 6060
rect 38442 6000 38506 6004
rect 38522 6060 38586 6064
rect 38522 6004 38526 6060
rect 38526 6004 38582 6060
rect 38582 6004 38586 6060
rect 38522 6000 38586 6004
rect 3650 5516 3714 5520
rect 3650 5460 3654 5516
rect 3654 5460 3710 5516
rect 3710 5460 3714 5516
rect 3650 5456 3714 5460
rect 3730 5516 3794 5520
rect 3730 5460 3734 5516
rect 3734 5460 3790 5516
rect 3790 5460 3794 5516
rect 3730 5456 3794 5460
rect 3810 5516 3874 5520
rect 3810 5460 3814 5516
rect 3814 5460 3870 5516
rect 3870 5460 3874 5516
rect 3810 5456 3874 5460
rect 3890 5516 3954 5520
rect 3890 5460 3894 5516
rect 3894 5460 3950 5516
rect 3950 5460 3954 5516
rect 3890 5456 3954 5460
rect 35618 5516 35682 5520
rect 35618 5460 35622 5516
rect 35622 5460 35678 5516
rect 35678 5460 35682 5516
rect 35618 5456 35682 5460
rect 35698 5516 35762 5520
rect 35698 5460 35702 5516
rect 35702 5460 35758 5516
rect 35758 5460 35762 5516
rect 35698 5456 35762 5460
rect 35778 5516 35842 5520
rect 35778 5460 35782 5516
rect 35782 5460 35838 5516
rect 35838 5460 35842 5516
rect 35778 5456 35842 5460
rect 35858 5516 35922 5520
rect 35858 5460 35862 5516
rect 35862 5460 35918 5516
rect 35918 5460 35922 5516
rect 35858 5456 35922 5460
rect 40946 5516 41010 5520
rect 40946 5460 40950 5516
rect 40950 5460 41006 5516
rect 41006 5460 41010 5516
rect 40946 5456 41010 5460
rect 41026 5516 41090 5520
rect 41026 5460 41030 5516
rect 41030 5460 41086 5516
rect 41086 5460 41090 5516
rect 41026 5456 41090 5460
rect 41106 5516 41170 5520
rect 41106 5460 41110 5516
rect 41110 5460 41166 5516
rect 41166 5460 41170 5516
rect 41106 5456 41170 5460
rect 41186 5516 41250 5520
rect 41186 5460 41190 5516
rect 41190 5460 41246 5516
rect 41246 5460 41250 5516
rect 41186 5456 41250 5460
rect 6314 4972 6378 4976
rect 6314 4916 6318 4972
rect 6318 4916 6374 4972
rect 6374 4916 6378 4972
rect 6314 4912 6378 4916
rect 6394 4972 6458 4976
rect 6394 4916 6398 4972
rect 6398 4916 6454 4972
rect 6454 4916 6458 4972
rect 6394 4912 6458 4916
rect 6474 4972 6538 4976
rect 6474 4916 6478 4972
rect 6478 4916 6534 4972
rect 6534 4916 6538 4972
rect 6474 4912 6538 4916
rect 6554 4972 6618 4976
rect 6554 4916 6558 4972
rect 6558 4916 6614 4972
rect 6614 4916 6618 4972
rect 6554 4912 6618 4916
rect 38282 4972 38346 4976
rect 38282 4916 38286 4972
rect 38286 4916 38342 4972
rect 38342 4916 38346 4972
rect 38282 4912 38346 4916
rect 38362 4972 38426 4976
rect 38362 4916 38366 4972
rect 38366 4916 38422 4972
rect 38422 4916 38426 4972
rect 38362 4912 38426 4916
rect 38442 4972 38506 4976
rect 38442 4916 38446 4972
rect 38446 4916 38502 4972
rect 38502 4916 38506 4972
rect 38442 4912 38506 4916
rect 38522 4972 38586 4976
rect 38522 4916 38526 4972
rect 38526 4916 38582 4972
rect 38582 4916 38586 4972
rect 38522 4912 38586 4916
rect 3650 4428 3714 4432
rect 3650 4372 3654 4428
rect 3654 4372 3710 4428
rect 3710 4372 3714 4428
rect 3650 4368 3714 4372
rect 3730 4428 3794 4432
rect 3730 4372 3734 4428
rect 3734 4372 3790 4428
rect 3790 4372 3794 4428
rect 3730 4368 3794 4372
rect 3810 4428 3874 4432
rect 3810 4372 3814 4428
rect 3814 4372 3870 4428
rect 3870 4372 3874 4428
rect 3810 4368 3874 4372
rect 3890 4428 3954 4432
rect 3890 4372 3894 4428
rect 3894 4372 3950 4428
rect 3950 4372 3954 4428
rect 3890 4368 3954 4372
rect 35618 4428 35682 4432
rect 35618 4372 35622 4428
rect 35622 4372 35678 4428
rect 35678 4372 35682 4428
rect 35618 4368 35682 4372
rect 35698 4428 35762 4432
rect 35698 4372 35702 4428
rect 35702 4372 35758 4428
rect 35758 4372 35762 4428
rect 35698 4368 35762 4372
rect 35778 4428 35842 4432
rect 35778 4372 35782 4428
rect 35782 4372 35838 4428
rect 35838 4372 35842 4428
rect 35778 4368 35842 4372
rect 35858 4428 35922 4432
rect 35858 4372 35862 4428
rect 35862 4372 35918 4428
rect 35918 4372 35922 4428
rect 35858 4368 35922 4372
rect 40946 4428 41010 4432
rect 40946 4372 40950 4428
rect 40950 4372 41006 4428
rect 41006 4372 41010 4428
rect 40946 4368 41010 4372
rect 41026 4428 41090 4432
rect 41026 4372 41030 4428
rect 41030 4372 41086 4428
rect 41086 4372 41090 4428
rect 41026 4368 41090 4372
rect 41106 4428 41170 4432
rect 41106 4372 41110 4428
rect 41110 4372 41166 4428
rect 41166 4372 41170 4428
rect 41106 4368 41170 4372
rect 41186 4428 41250 4432
rect 41186 4372 41190 4428
rect 41190 4372 41246 4428
rect 41246 4372 41250 4428
rect 41186 4368 41250 4372
rect 6314 3884 6378 3888
rect 6314 3828 6318 3884
rect 6318 3828 6374 3884
rect 6374 3828 6378 3884
rect 6314 3824 6378 3828
rect 6394 3884 6458 3888
rect 6394 3828 6398 3884
rect 6398 3828 6454 3884
rect 6454 3828 6458 3884
rect 6394 3824 6458 3828
rect 6474 3884 6538 3888
rect 6474 3828 6478 3884
rect 6478 3828 6534 3884
rect 6534 3828 6538 3884
rect 6474 3824 6538 3828
rect 6554 3884 6618 3888
rect 6554 3828 6558 3884
rect 6558 3828 6614 3884
rect 6614 3828 6618 3884
rect 6554 3824 6618 3828
rect 38282 3884 38346 3888
rect 38282 3828 38286 3884
rect 38286 3828 38342 3884
rect 38342 3828 38346 3884
rect 38282 3824 38346 3828
rect 38362 3884 38426 3888
rect 38362 3828 38366 3884
rect 38366 3828 38422 3884
rect 38422 3828 38426 3884
rect 38362 3824 38426 3828
rect 38442 3884 38506 3888
rect 38442 3828 38446 3884
rect 38446 3828 38502 3884
rect 38502 3828 38506 3884
rect 38442 3824 38506 3828
rect 38522 3884 38586 3888
rect 38522 3828 38526 3884
rect 38526 3828 38582 3884
rect 38582 3828 38586 3884
rect 38522 3824 38586 3828
rect 3650 3340 3714 3344
rect 3650 3284 3654 3340
rect 3654 3284 3710 3340
rect 3710 3284 3714 3340
rect 3650 3280 3714 3284
rect 3730 3340 3794 3344
rect 3730 3284 3734 3340
rect 3734 3284 3790 3340
rect 3790 3284 3794 3340
rect 3730 3280 3794 3284
rect 3810 3340 3874 3344
rect 3810 3284 3814 3340
rect 3814 3284 3870 3340
rect 3870 3284 3874 3340
rect 3810 3280 3874 3284
rect 3890 3340 3954 3344
rect 3890 3284 3894 3340
rect 3894 3284 3950 3340
rect 3950 3284 3954 3340
rect 3890 3280 3954 3284
rect 35618 3340 35682 3344
rect 35618 3284 35622 3340
rect 35622 3284 35678 3340
rect 35678 3284 35682 3340
rect 35618 3280 35682 3284
rect 35698 3340 35762 3344
rect 35698 3284 35702 3340
rect 35702 3284 35758 3340
rect 35758 3284 35762 3340
rect 35698 3280 35762 3284
rect 35778 3340 35842 3344
rect 35778 3284 35782 3340
rect 35782 3284 35838 3340
rect 35838 3284 35842 3340
rect 35778 3280 35842 3284
rect 35858 3340 35922 3344
rect 35858 3284 35862 3340
rect 35862 3284 35918 3340
rect 35918 3284 35922 3340
rect 35858 3280 35922 3284
rect 40946 3340 41010 3344
rect 40946 3284 40950 3340
rect 40950 3284 41006 3340
rect 41006 3284 41010 3340
rect 40946 3280 41010 3284
rect 41026 3340 41090 3344
rect 41026 3284 41030 3340
rect 41030 3284 41086 3340
rect 41086 3284 41090 3340
rect 41026 3280 41090 3284
rect 41106 3340 41170 3344
rect 41106 3284 41110 3340
rect 41110 3284 41166 3340
rect 41166 3284 41170 3340
rect 41106 3280 41170 3284
rect 41186 3340 41250 3344
rect 41186 3284 41190 3340
rect 41190 3284 41246 3340
rect 41246 3284 41250 3340
rect 41186 3280 41250 3284
rect 6314 2796 6378 2800
rect 6314 2740 6318 2796
rect 6318 2740 6374 2796
rect 6374 2740 6378 2796
rect 6314 2736 6378 2740
rect 6394 2796 6458 2800
rect 6394 2740 6398 2796
rect 6398 2740 6454 2796
rect 6454 2740 6458 2796
rect 6394 2736 6458 2740
rect 6474 2796 6538 2800
rect 6474 2740 6478 2796
rect 6478 2740 6534 2796
rect 6534 2740 6538 2796
rect 6474 2736 6538 2740
rect 6554 2796 6618 2800
rect 6554 2740 6558 2796
rect 6558 2740 6614 2796
rect 6614 2740 6618 2796
rect 6554 2736 6618 2740
rect 38282 2796 38346 2800
rect 38282 2740 38286 2796
rect 38286 2740 38342 2796
rect 38342 2740 38346 2796
rect 38282 2736 38346 2740
rect 38362 2796 38426 2800
rect 38362 2740 38366 2796
rect 38366 2740 38422 2796
rect 38422 2740 38426 2796
rect 38362 2736 38426 2740
rect 38442 2796 38506 2800
rect 38442 2740 38446 2796
rect 38446 2740 38502 2796
rect 38502 2740 38506 2796
rect 38442 2736 38506 2740
rect 38522 2796 38586 2800
rect 38522 2740 38526 2796
rect 38526 2740 38582 2796
rect 38582 2740 38586 2796
rect 38522 2736 38586 2740
rect 3650 2252 3714 2256
rect 3650 2196 3654 2252
rect 3654 2196 3710 2252
rect 3710 2196 3714 2252
rect 3650 2192 3714 2196
rect 3730 2252 3794 2256
rect 3730 2196 3734 2252
rect 3734 2196 3790 2252
rect 3790 2196 3794 2252
rect 3730 2192 3794 2196
rect 3810 2252 3874 2256
rect 3810 2196 3814 2252
rect 3814 2196 3870 2252
rect 3870 2196 3874 2252
rect 3810 2192 3874 2196
rect 3890 2252 3954 2256
rect 3890 2196 3894 2252
rect 3894 2196 3950 2252
rect 3950 2196 3954 2252
rect 3890 2192 3954 2196
rect 35618 2252 35682 2256
rect 35618 2196 35622 2252
rect 35622 2196 35678 2252
rect 35678 2196 35682 2252
rect 35618 2192 35682 2196
rect 35698 2252 35762 2256
rect 35698 2196 35702 2252
rect 35702 2196 35758 2252
rect 35758 2196 35762 2252
rect 35698 2192 35762 2196
rect 35778 2252 35842 2256
rect 35778 2196 35782 2252
rect 35782 2196 35838 2252
rect 35838 2196 35842 2252
rect 35778 2192 35842 2196
rect 35858 2252 35922 2256
rect 35858 2196 35862 2252
rect 35862 2196 35918 2252
rect 35918 2196 35922 2252
rect 35858 2192 35922 2196
rect 40946 2252 41010 2256
rect 40946 2196 40950 2252
rect 40950 2196 41006 2252
rect 41006 2196 41010 2252
rect 40946 2192 41010 2196
rect 41026 2252 41090 2256
rect 41026 2196 41030 2252
rect 41030 2196 41086 2252
rect 41086 2196 41090 2252
rect 41026 2192 41090 2196
rect 41106 2252 41170 2256
rect 41106 2196 41110 2252
rect 41110 2196 41166 2252
rect 41166 2196 41170 2252
rect 41106 2192 41170 2196
rect 41186 2252 41250 2256
rect 41186 2196 41190 2252
rect 41190 2196 41246 2252
rect 41246 2196 41250 2252
rect 41186 2192 41250 2196
rect 6314 1708 6378 1712
rect 6314 1652 6318 1708
rect 6318 1652 6374 1708
rect 6374 1652 6378 1708
rect 6314 1648 6378 1652
rect 6394 1708 6458 1712
rect 6394 1652 6398 1708
rect 6398 1652 6454 1708
rect 6454 1652 6458 1708
rect 6394 1648 6458 1652
rect 6474 1708 6538 1712
rect 6474 1652 6478 1708
rect 6478 1652 6534 1708
rect 6534 1652 6538 1708
rect 6474 1648 6538 1652
rect 6554 1708 6618 1712
rect 6554 1652 6558 1708
rect 6558 1652 6614 1708
rect 6614 1652 6618 1708
rect 6554 1648 6618 1652
rect 38282 1708 38346 1712
rect 38282 1652 38286 1708
rect 38286 1652 38342 1708
rect 38342 1652 38346 1708
rect 38282 1648 38346 1652
rect 38362 1708 38426 1712
rect 38362 1652 38366 1708
rect 38366 1652 38422 1708
rect 38422 1652 38426 1708
rect 38362 1648 38426 1652
rect 38442 1708 38506 1712
rect 38442 1652 38446 1708
rect 38446 1652 38502 1708
rect 38502 1652 38506 1708
rect 38442 1648 38506 1652
rect 38522 1708 38586 1712
rect 38522 1652 38526 1708
rect 38526 1652 38582 1708
rect 38582 1652 38586 1708
rect 38522 1648 38586 1652
rect 3650 1164 3714 1168
rect 3650 1108 3654 1164
rect 3654 1108 3710 1164
rect 3710 1108 3714 1164
rect 3650 1104 3714 1108
rect 3730 1164 3794 1168
rect 3730 1108 3734 1164
rect 3734 1108 3790 1164
rect 3790 1108 3794 1164
rect 3730 1104 3794 1108
rect 3810 1164 3874 1168
rect 3810 1108 3814 1164
rect 3814 1108 3870 1164
rect 3870 1108 3874 1164
rect 3810 1104 3874 1108
rect 3890 1164 3954 1168
rect 3890 1108 3894 1164
rect 3894 1108 3950 1164
rect 3950 1108 3954 1164
rect 3890 1104 3954 1108
rect 35618 1164 35682 1168
rect 35618 1108 35622 1164
rect 35622 1108 35678 1164
rect 35678 1108 35682 1164
rect 35618 1104 35682 1108
rect 35698 1164 35762 1168
rect 35698 1108 35702 1164
rect 35702 1108 35758 1164
rect 35758 1108 35762 1164
rect 35698 1104 35762 1108
rect 35778 1164 35842 1168
rect 35778 1108 35782 1164
rect 35782 1108 35838 1164
rect 35838 1108 35842 1164
rect 35778 1104 35842 1108
rect 35858 1164 35922 1168
rect 35858 1108 35862 1164
rect 35862 1108 35918 1164
rect 35918 1108 35922 1164
rect 35858 1104 35922 1108
rect 40946 1164 41010 1168
rect 40946 1108 40950 1164
rect 40950 1108 41006 1164
rect 41006 1108 41010 1164
rect 40946 1104 41010 1108
rect 41026 1164 41090 1168
rect 41026 1108 41030 1164
rect 41030 1108 41086 1164
rect 41086 1108 41090 1164
rect 41026 1104 41090 1108
rect 41106 1164 41170 1168
rect 41106 1108 41110 1164
rect 41110 1108 41166 1164
rect 41166 1108 41170 1164
rect 41106 1104 41170 1108
rect 41186 1164 41250 1168
rect 41186 1108 41190 1164
rect 41190 1108 41246 1164
rect 41246 1108 41250 1164
rect 41186 1104 41250 1108
rect 6314 620 6378 624
rect 6314 564 6318 620
rect 6318 564 6374 620
rect 6374 564 6378 620
rect 6314 560 6378 564
rect 6394 620 6458 624
rect 6394 564 6398 620
rect 6398 564 6454 620
rect 6454 564 6458 620
rect 6394 560 6458 564
rect 6474 620 6538 624
rect 6474 564 6478 620
rect 6478 564 6534 620
rect 6534 564 6538 620
rect 6474 560 6538 564
rect 6554 620 6618 624
rect 6554 564 6558 620
rect 6558 564 6614 620
rect 6614 564 6618 620
rect 6554 560 6618 564
rect 38282 620 38346 624
rect 38282 564 38286 620
rect 38286 564 38342 620
rect 38342 564 38346 620
rect 38282 560 38346 564
rect 38362 620 38426 624
rect 38362 564 38366 620
rect 38366 564 38422 620
rect 38422 564 38426 620
rect 38362 560 38426 564
rect 38442 620 38506 624
rect 38442 564 38446 620
rect 38446 564 38502 620
rect 38502 564 38506 620
rect 38442 560 38506 564
rect 38522 620 38586 624
rect 38522 564 38526 620
rect 38526 564 38582 620
rect 38582 564 38586 620
rect 38522 560 38586 564
rect 3650 76 3714 80
rect 3650 20 3654 76
rect 3654 20 3710 76
rect 3710 20 3714 76
rect 3650 16 3714 20
rect 3730 76 3794 80
rect 3730 20 3734 76
rect 3734 20 3790 76
rect 3790 20 3794 76
rect 3730 16 3794 20
rect 3810 76 3874 80
rect 3810 20 3814 76
rect 3814 20 3870 76
rect 3870 20 3874 76
rect 3810 16 3874 20
rect 3890 76 3954 80
rect 3890 20 3894 76
rect 3894 20 3950 76
rect 3950 20 3954 76
rect 3890 16 3954 20
rect 35618 76 35682 80
rect 35618 20 35622 76
rect 35622 20 35678 76
rect 35678 20 35682 76
rect 35618 16 35682 20
rect 35698 76 35762 80
rect 35698 20 35702 76
rect 35702 20 35758 76
rect 35758 20 35762 76
rect 35698 16 35762 20
rect 35778 76 35842 80
rect 35778 20 35782 76
rect 35782 20 35838 76
rect 35838 20 35842 76
rect 35778 16 35842 20
rect 35858 76 35922 80
rect 35858 20 35862 76
rect 35862 20 35918 76
rect 35918 20 35922 76
rect 35858 16 35922 20
rect 40946 76 41010 80
rect 40946 20 40950 76
rect 40950 20 41006 76
rect 41006 20 41010 76
rect 40946 16 41010 20
rect 41026 76 41090 80
rect 41026 20 41030 76
rect 41030 20 41086 76
rect 41086 20 41090 76
rect 41026 16 41090 20
rect 41106 76 41170 80
rect 41106 20 41110 76
rect 41110 20 41166 76
rect 41166 20 41170 76
rect 41106 16 41170 20
rect 41186 76 41250 80
rect 41186 20 41190 76
rect 41190 20 41246 76
rect 41246 20 41250 76
rect 41186 16 41250 20
<< metal4 >>
rect 3642 41424 3962 41984
rect 3642 41360 3650 41424
rect 3714 41360 3730 41424
rect 3794 41360 3810 41424
rect 3874 41360 3890 41424
rect 3954 41360 3962 41424
rect 3642 40336 3962 41360
rect 3642 40272 3650 40336
rect 3714 40326 3730 40336
rect 3794 40326 3810 40336
rect 3874 40326 3890 40336
rect 3954 40272 3962 40336
rect 3642 40090 3684 40272
rect 3920 40090 3962 40272
rect 3642 40006 3962 40090
rect 3642 39770 3684 40006
rect 3920 39770 3962 40006
rect 3642 39248 3962 39770
rect 3642 39184 3650 39248
rect 3714 39184 3730 39248
rect 3794 39184 3810 39248
rect 3874 39184 3890 39248
rect 3954 39184 3962 39248
rect 3642 38160 3962 39184
rect 3642 38096 3650 38160
rect 3714 38096 3730 38160
rect 3794 38096 3810 38160
rect 3874 38096 3890 38160
rect 3954 38096 3962 38160
rect 3642 37072 3962 38096
rect 3642 37008 3650 37072
rect 3714 37008 3730 37072
rect 3794 37008 3810 37072
rect 3874 37008 3890 37072
rect 3954 37008 3962 37072
rect 3642 35984 3962 37008
rect 3642 35920 3650 35984
rect 3714 35920 3730 35984
rect 3794 35920 3810 35984
rect 3874 35920 3890 35984
rect 3954 35920 3962 35984
rect 3642 34896 3962 35920
rect 3642 34832 3650 34896
rect 3714 34832 3730 34896
rect 3794 34832 3810 34896
rect 3874 34832 3890 34896
rect 3954 34832 3962 34896
rect 3642 33808 3962 34832
rect 3642 33744 3650 33808
rect 3714 33744 3730 33808
rect 3794 33744 3810 33808
rect 3874 33744 3890 33808
rect 3954 33744 3962 33808
rect 3642 32720 3962 33744
rect 3642 32656 3650 32720
rect 3714 32656 3730 32720
rect 3794 32656 3810 32720
rect 3874 32656 3890 32720
rect 3954 32656 3962 32720
rect 3642 31632 3962 32656
rect 3642 31568 3650 31632
rect 3714 31568 3730 31632
rect 3794 31568 3810 31632
rect 3874 31568 3890 31632
rect 3954 31568 3962 31632
rect 3642 30544 3962 31568
rect 3642 30480 3650 30544
rect 3714 30480 3730 30544
rect 3794 30480 3810 30544
rect 3874 30480 3890 30544
rect 3954 30480 3962 30544
rect 3642 29456 3962 30480
rect 3642 29392 3650 29456
rect 3714 29392 3730 29456
rect 3794 29392 3810 29456
rect 3874 29392 3890 29456
rect 3954 29392 3962 29456
rect 3642 28368 3962 29392
rect 3642 28304 3650 28368
rect 3714 28304 3730 28368
rect 3794 28304 3810 28368
rect 3874 28304 3890 28368
rect 3954 28304 3962 28368
rect 3642 27280 3962 28304
rect 3642 27216 3650 27280
rect 3714 27216 3730 27280
rect 3794 27216 3810 27280
rect 3874 27216 3890 27280
rect 3954 27216 3962 27280
rect 3642 26192 3962 27216
rect 3642 26128 3650 26192
rect 3714 26128 3730 26192
rect 3794 26128 3810 26192
rect 3874 26128 3890 26192
rect 3954 26128 3962 26192
rect 3642 25104 3962 26128
rect 3642 25040 3650 25104
rect 3714 25040 3730 25104
rect 3794 25040 3810 25104
rect 3874 25040 3890 25104
rect 3954 25040 3962 25104
rect 3642 24016 3962 25040
rect 3642 23952 3650 24016
rect 3714 23952 3730 24016
rect 3794 23952 3810 24016
rect 3874 23952 3890 24016
rect 3954 23952 3962 24016
rect 3642 22928 3962 23952
rect 3642 22864 3650 22928
rect 3714 22864 3730 22928
rect 3794 22864 3810 22928
rect 3874 22864 3890 22928
rect 3954 22864 3962 22928
rect 3357 22724 3423 22725
rect 3357 22660 3358 22724
rect 3422 22660 3423 22724
rect 3357 22659 3423 22660
rect 3360 20770 3420 22659
rect 3642 21840 3962 22864
rect 3642 21776 3650 21840
rect 3714 21776 3730 21840
rect 3794 21776 3810 21840
rect 3874 21776 3890 21840
rect 3954 21776 3962 21840
rect 3642 20752 3962 21776
rect 3642 20688 3650 20752
rect 3714 20688 3730 20752
rect 3794 20688 3810 20752
rect 3874 20688 3890 20752
rect 3954 20688 3962 20752
rect 3642 19664 3962 20688
rect 3642 19600 3650 19664
rect 3714 19600 3730 19664
rect 3794 19600 3810 19664
rect 3874 19600 3890 19664
rect 3954 19600 3962 19664
rect 3642 18576 3962 19600
rect 6306 41968 6626 41984
rect 6306 41904 6314 41968
rect 6378 41904 6394 41968
rect 6458 41904 6474 41968
rect 6538 41904 6554 41968
rect 6618 41904 6626 41968
rect 6306 40880 6626 41904
rect 6306 40816 6314 40880
rect 6378 40816 6394 40880
rect 6458 40816 6474 40880
rect 6538 40816 6554 40880
rect 6618 40816 6626 40880
rect 6306 39792 6626 40816
rect 6306 39728 6314 39792
rect 6378 39728 6394 39792
rect 6458 39728 6474 39792
rect 6538 39728 6554 39792
rect 6618 39728 6626 39792
rect 6306 38704 6626 39728
rect 6306 38640 6314 38704
rect 6378 38640 6394 38704
rect 6458 38640 6474 38704
rect 6538 38640 6554 38704
rect 6618 38640 6626 38704
rect 6306 37616 6626 38640
rect 6306 37552 6314 37616
rect 6378 37552 6394 37616
rect 6458 37552 6474 37616
rect 6538 37552 6554 37616
rect 6618 37552 6626 37616
rect 6306 36528 6626 37552
rect 6306 36464 6314 36528
rect 6378 36464 6394 36528
rect 6458 36464 6474 36528
rect 6538 36464 6554 36528
rect 6618 36464 6626 36528
rect 6306 35440 6626 36464
rect 6306 35376 6314 35440
rect 6378 35376 6394 35440
rect 6458 35376 6474 35440
rect 6538 35376 6554 35440
rect 6618 35376 6626 35440
rect 6306 34352 6626 35376
rect 6306 34288 6314 34352
rect 6378 34288 6394 34352
rect 6458 34288 6474 34352
rect 6538 34288 6554 34352
rect 6618 34288 6626 34352
rect 6306 33264 6626 34288
rect 6306 33200 6314 33264
rect 6378 33200 6394 33264
rect 6458 33200 6474 33264
rect 6538 33200 6554 33264
rect 6618 33200 6626 33264
rect 6306 32176 6626 33200
rect 6306 32112 6314 32176
rect 6378 32112 6394 32176
rect 6458 32112 6474 32176
rect 6538 32112 6554 32176
rect 6618 32112 6626 32176
rect 6306 31088 6626 32112
rect 6306 31024 6314 31088
rect 6378 31024 6394 31088
rect 6458 31024 6474 31088
rect 6538 31024 6554 31088
rect 6618 31024 6626 31088
rect 6306 30000 6626 31024
rect 6306 29936 6314 30000
rect 6378 29936 6394 30000
rect 6458 29936 6474 30000
rect 6538 29936 6554 30000
rect 6618 29936 6626 30000
rect 6306 28912 6626 29936
rect 6306 28848 6314 28912
rect 6378 28848 6394 28912
rect 6458 28848 6474 28912
rect 6538 28848 6554 28912
rect 6618 28848 6626 28912
rect 6306 27824 6626 28848
rect 6306 27760 6314 27824
rect 6378 27760 6394 27824
rect 6458 27760 6474 27824
rect 6538 27760 6554 27824
rect 6618 27760 6626 27824
rect 6306 26736 6626 27760
rect 6306 26672 6314 26736
rect 6378 26672 6394 26736
rect 6458 26672 6474 26736
rect 6538 26672 6554 26736
rect 6618 26672 6626 26736
rect 6306 25648 6626 26672
rect 8970 41424 9290 41984
rect 8970 41360 8978 41424
rect 9042 41360 9058 41424
rect 9122 41360 9138 41424
rect 9202 41360 9218 41424
rect 9282 41360 9290 41424
rect 8970 40336 9290 41360
rect 8970 40272 8978 40336
rect 9042 40326 9058 40336
rect 9122 40326 9138 40336
rect 9202 40326 9218 40336
rect 9282 40272 9290 40336
rect 8970 40090 9012 40272
rect 9248 40090 9290 40272
rect 8970 40006 9290 40090
rect 8970 39770 9012 40006
rect 9248 39770 9290 40006
rect 8970 39248 9290 39770
rect 8970 39184 8978 39248
rect 9042 39184 9058 39248
rect 9122 39184 9138 39248
rect 9202 39184 9218 39248
rect 9282 39184 9290 39248
rect 8970 38160 9290 39184
rect 8970 38096 8978 38160
rect 9042 38096 9058 38160
rect 9122 38096 9138 38160
rect 9202 38096 9218 38160
rect 9282 38096 9290 38160
rect 8970 37072 9290 38096
rect 8970 37008 8978 37072
rect 9042 37008 9058 37072
rect 9122 37008 9138 37072
rect 9202 37008 9218 37072
rect 9282 37008 9290 37072
rect 8970 35984 9290 37008
rect 8970 35920 8978 35984
rect 9042 35920 9058 35984
rect 9122 35920 9138 35984
rect 9202 35920 9218 35984
rect 9282 35920 9290 35984
rect 8970 34896 9290 35920
rect 8970 34832 8978 34896
rect 9042 34832 9058 34896
rect 9122 34832 9138 34896
rect 9202 34832 9218 34896
rect 9282 34832 9290 34896
rect 8970 33808 9290 34832
rect 8970 33744 8978 33808
rect 9042 33744 9058 33808
rect 9122 33744 9138 33808
rect 9202 33744 9218 33808
rect 9282 33744 9290 33808
rect 8970 32720 9290 33744
rect 8970 32656 8978 32720
rect 9042 32656 9058 32720
rect 9122 32656 9138 32720
rect 9202 32656 9218 32720
rect 9282 32656 9290 32720
rect 8970 31632 9290 32656
rect 8970 31568 8978 31632
rect 9042 31568 9058 31632
rect 9122 31568 9138 31632
rect 9202 31568 9218 31632
rect 9282 31568 9290 31632
rect 8970 30544 9290 31568
rect 8970 30480 8978 30544
rect 9042 30480 9058 30544
rect 9122 30480 9138 30544
rect 9202 30480 9218 30544
rect 9282 30480 9290 30544
rect 8970 29456 9290 30480
rect 8970 29392 8978 29456
rect 9042 29392 9058 29456
rect 9122 29392 9138 29456
rect 9202 29392 9218 29456
rect 9282 29392 9290 29456
rect 8970 28368 9290 29392
rect 8970 28304 8978 28368
rect 9042 28304 9058 28368
rect 9122 28304 9138 28368
rect 9202 28304 9218 28368
rect 9282 28304 9290 28368
rect 8970 27280 9290 28304
rect 8970 27216 8978 27280
rect 9042 27216 9058 27280
rect 9122 27216 9138 27280
rect 9202 27216 9218 27280
rect 9282 27216 9290 27280
rect 8970 26609 9290 27216
rect 11634 41968 11954 41984
rect 11634 41904 11642 41968
rect 11706 41904 11722 41968
rect 11786 41904 11802 41968
rect 11866 41904 11882 41968
rect 11946 41904 11954 41968
rect 11634 40880 11954 41904
rect 11634 40816 11642 40880
rect 11706 40816 11722 40880
rect 11786 40816 11802 40880
rect 11866 40816 11882 40880
rect 11946 40816 11954 40880
rect 11634 39792 11954 40816
rect 11634 39728 11642 39792
rect 11706 39728 11722 39792
rect 11786 39728 11802 39792
rect 11866 39728 11882 39792
rect 11946 39728 11954 39792
rect 11634 38704 11954 39728
rect 11634 38640 11642 38704
rect 11706 38640 11722 38704
rect 11786 38640 11802 38704
rect 11866 38640 11882 38704
rect 11946 38640 11954 38704
rect 11634 37616 11954 38640
rect 11634 37552 11642 37616
rect 11706 37552 11722 37616
rect 11786 37552 11802 37616
rect 11866 37552 11882 37616
rect 11946 37552 11954 37616
rect 11634 36528 11954 37552
rect 11634 36464 11642 36528
rect 11706 36464 11722 36528
rect 11786 36464 11802 36528
rect 11866 36464 11882 36528
rect 11946 36464 11954 36528
rect 11634 35440 11954 36464
rect 11634 35376 11642 35440
rect 11706 35376 11722 35440
rect 11786 35376 11802 35440
rect 11866 35376 11882 35440
rect 11946 35376 11954 35440
rect 11634 34352 11954 35376
rect 11634 34288 11642 34352
rect 11706 34288 11722 34352
rect 11786 34288 11802 34352
rect 11866 34288 11882 34352
rect 11946 34288 11954 34352
rect 11634 33264 11954 34288
rect 11634 33200 11642 33264
rect 11706 33200 11722 33264
rect 11786 33200 11802 33264
rect 11866 33200 11882 33264
rect 11946 33200 11954 33264
rect 11634 32176 11954 33200
rect 11634 32112 11642 32176
rect 11706 32112 11722 32176
rect 11786 32112 11802 32176
rect 11866 32112 11882 32176
rect 11946 32112 11954 32176
rect 11634 31088 11954 32112
rect 11634 31024 11642 31088
rect 11706 31024 11722 31088
rect 11786 31024 11802 31088
rect 11866 31024 11882 31088
rect 11946 31024 11954 31088
rect 11634 30000 11954 31024
rect 11634 29936 11642 30000
rect 11706 29936 11722 30000
rect 11786 29936 11802 30000
rect 11866 29936 11882 30000
rect 11946 29936 11954 30000
rect 11634 28912 11954 29936
rect 11634 28848 11642 28912
rect 11706 28848 11722 28912
rect 11786 28848 11802 28912
rect 11866 28848 11882 28912
rect 11946 28848 11954 28912
rect 11634 27824 11954 28848
rect 11634 27760 11642 27824
rect 11706 27760 11722 27824
rect 11786 27760 11802 27824
rect 11866 27760 11882 27824
rect 11946 27760 11954 27824
rect 11634 26736 11954 27760
rect 11634 26672 11642 26736
rect 11706 26672 11722 26736
rect 11786 26672 11802 26736
rect 11866 26672 11882 26736
rect 11946 26672 11954 26736
rect 11634 26609 11954 26672
rect 14298 41424 14618 41984
rect 14298 41360 14306 41424
rect 14370 41360 14386 41424
rect 14450 41360 14466 41424
rect 14530 41360 14546 41424
rect 14610 41360 14618 41424
rect 14298 40336 14618 41360
rect 14298 40272 14306 40336
rect 14370 40326 14386 40336
rect 14450 40326 14466 40336
rect 14530 40326 14546 40336
rect 14610 40272 14618 40336
rect 14298 40090 14340 40272
rect 14576 40090 14618 40272
rect 14298 40006 14618 40090
rect 14298 39770 14340 40006
rect 14576 39770 14618 40006
rect 14298 39248 14618 39770
rect 14298 39184 14306 39248
rect 14370 39184 14386 39248
rect 14450 39184 14466 39248
rect 14530 39184 14546 39248
rect 14610 39184 14618 39248
rect 14298 38160 14618 39184
rect 14298 38096 14306 38160
rect 14370 38096 14386 38160
rect 14450 38096 14466 38160
rect 14530 38096 14546 38160
rect 14610 38096 14618 38160
rect 14298 37072 14618 38096
rect 14298 37008 14306 37072
rect 14370 37008 14386 37072
rect 14450 37008 14466 37072
rect 14530 37008 14546 37072
rect 14610 37008 14618 37072
rect 14298 35984 14618 37008
rect 14298 35920 14306 35984
rect 14370 35920 14386 35984
rect 14450 35920 14466 35984
rect 14530 35920 14546 35984
rect 14610 35920 14618 35984
rect 14298 34896 14618 35920
rect 14298 34832 14306 34896
rect 14370 34832 14386 34896
rect 14450 34832 14466 34896
rect 14530 34832 14546 34896
rect 14610 34832 14618 34896
rect 14298 33808 14618 34832
rect 14298 33744 14306 33808
rect 14370 33744 14386 33808
rect 14450 33744 14466 33808
rect 14530 33744 14546 33808
rect 14610 33744 14618 33808
rect 14298 32720 14618 33744
rect 14298 32656 14306 32720
rect 14370 32656 14386 32720
rect 14450 32656 14466 32720
rect 14530 32656 14546 32720
rect 14610 32656 14618 32720
rect 14298 31632 14618 32656
rect 14298 31568 14306 31632
rect 14370 31568 14386 31632
rect 14450 31568 14466 31632
rect 14530 31568 14546 31632
rect 14610 31568 14618 31632
rect 14298 30544 14618 31568
rect 14298 30480 14306 30544
rect 14370 30480 14386 30544
rect 14450 30480 14466 30544
rect 14530 30480 14546 30544
rect 14610 30480 14618 30544
rect 14298 29456 14618 30480
rect 14298 29392 14306 29456
rect 14370 29392 14386 29456
rect 14450 29392 14466 29456
rect 14530 29392 14546 29456
rect 14610 29392 14618 29456
rect 14298 28368 14618 29392
rect 14298 28304 14306 28368
rect 14370 28304 14386 28368
rect 14450 28304 14466 28368
rect 14530 28304 14546 28368
rect 14610 28304 14618 28368
rect 14298 27280 14618 28304
rect 14298 27216 14306 27280
rect 14370 27216 14386 27280
rect 14450 27216 14466 27280
rect 14530 27216 14546 27280
rect 14610 27216 14618 27280
rect 14298 26609 14618 27216
rect 16962 41968 17282 41984
rect 16962 41904 16970 41968
rect 17034 41904 17050 41968
rect 17114 41904 17130 41968
rect 17194 41904 17210 41968
rect 17274 41904 17282 41968
rect 16962 40880 17282 41904
rect 16962 40816 16970 40880
rect 17034 40816 17050 40880
rect 17114 40816 17130 40880
rect 17194 40816 17210 40880
rect 17274 40816 17282 40880
rect 16962 39792 17282 40816
rect 16962 39728 16970 39792
rect 17034 39728 17050 39792
rect 17114 39728 17130 39792
rect 17194 39728 17210 39792
rect 17274 39728 17282 39792
rect 16962 38704 17282 39728
rect 16962 38640 16970 38704
rect 17034 38640 17050 38704
rect 17114 38640 17130 38704
rect 17194 38640 17210 38704
rect 17274 38640 17282 38704
rect 16962 37616 17282 38640
rect 16962 37552 16970 37616
rect 17034 37552 17050 37616
rect 17114 37552 17130 37616
rect 17194 37552 17210 37616
rect 17274 37552 17282 37616
rect 16962 36528 17282 37552
rect 16962 36464 16970 36528
rect 17034 36464 17050 36528
rect 17114 36464 17130 36528
rect 17194 36464 17210 36528
rect 17274 36464 17282 36528
rect 16962 35440 17282 36464
rect 16962 35376 16970 35440
rect 17034 35376 17050 35440
rect 17114 35376 17130 35440
rect 17194 35376 17210 35440
rect 17274 35376 17282 35440
rect 16962 34352 17282 35376
rect 16962 34288 16970 34352
rect 17034 34288 17050 34352
rect 17114 34288 17130 34352
rect 17194 34288 17210 34352
rect 17274 34288 17282 34352
rect 16962 33264 17282 34288
rect 16962 33200 16970 33264
rect 17034 33200 17050 33264
rect 17114 33200 17130 33264
rect 17194 33200 17210 33264
rect 17274 33200 17282 33264
rect 16962 32176 17282 33200
rect 16962 32112 16970 32176
rect 17034 32112 17050 32176
rect 17114 32112 17130 32176
rect 17194 32112 17210 32176
rect 17274 32112 17282 32176
rect 16962 31088 17282 32112
rect 16962 31024 16970 31088
rect 17034 31024 17050 31088
rect 17114 31024 17130 31088
rect 17194 31024 17210 31088
rect 17274 31024 17282 31088
rect 16962 30000 17282 31024
rect 16962 29936 16970 30000
rect 17034 29936 17050 30000
rect 17114 29936 17130 30000
rect 17194 29936 17210 30000
rect 17274 29936 17282 30000
rect 16962 28912 17282 29936
rect 16962 28848 16970 28912
rect 17034 28848 17050 28912
rect 17114 28848 17130 28912
rect 17194 28848 17210 28912
rect 17274 28848 17282 28912
rect 16962 27824 17282 28848
rect 16962 27760 16970 27824
rect 17034 27760 17050 27824
rect 17114 27760 17130 27824
rect 17194 27760 17210 27824
rect 17274 27760 17282 27824
rect 16962 26736 17282 27760
rect 16962 26672 16970 26736
rect 17034 26672 17050 26736
rect 17114 26672 17130 26736
rect 17194 26672 17210 26736
rect 17274 26672 17282 26736
rect 16962 26609 17282 26672
rect 19626 41424 19946 41984
rect 19626 41360 19634 41424
rect 19698 41360 19714 41424
rect 19778 41360 19794 41424
rect 19858 41360 19874 41424
rect 19938 41360 19946 41424
rect 19626 40336 19946 41360
rect 19626 40272 19634 40336
rect 19698 40326 19714 40336
rect 19778 40326 19794 40336
rect 19858 40326 19874 40336
rect 19938 40272 19946 40336
rect 19626 40090 19668 40272
rect 19904 40090 19946 40272
rect 19626 40006 19946 40090
rect 19626 39770 19668 40006
rect 19904 39770 19946 40006
rect 19626 39248 19946 39770
rect 19626 39184 19634 39248
rect 19698 39184 19714 39248
rect 19778 39184 19794 39248
rect 19858 39184 19874 39248
rect 19938 39184 19946 39248
rect 19626 38160 19946 39184
rect 19626 38096 19634 38160
rect 19698 38096 19714 38160
rect 19778 38096 19794 38160
rect 19858 38096 19874 38160
rect 19938 38096 19946 38160
rect 19626 37072 19946 38096
rect 19626 37008 19634 37072
rect 19698 37008 19714 37072
rect 19778 37008 19794 37072
rect 19858 37008 19874 37072
rect 19938 37008 19946 37072
rect 19626 35984 19946 37008
rect 19626 35920 19634 35984
rect 19698 35920 19714 35984
rect 19778 35920 19794 35984
rect 19858 35920 19874 35984
rect 19938 35920 19946 35984
rect 19626 34896 19946 35920
rect 19626 34832 19634 34896
rect 19698 34832 19714 34896
rect 19778 34832 19794 34896
rect 19858 34832 19874 34896
rect 19938 34832 19946 34896
rect 19626 33808 19946 34832
rect 19626 33744 19634 33808
rect 19698 33744 19714 33808
rect 19778 33744 19794 33808
rect 19858 33744 19874 33808
rect 19938 33744 19946 33808
rect 19626 32720 19946 33744
rect 19626 32656 19634 32720
rect 19698 32656 19714 32720
rect 19778 32656 19794 32720
rect 19858 32656 19874 32720
rect 19938 32656 19946 32720
rect 19626 31632 19946 32656
rect 19626 31568 19634 31632
rect 19698 31568 19714 31632
rect 19778 31568 19794 31632
rect 19858 31568 19874 31632
rect 19938 31568 19946 31632
rect 19626 30544 19946 31568
rect 19626 30480 19634 30544
rect 19698 30480 19714 30544
rect 19778 30480 19794 30544
rect 19858 30480 19874 30544
rect 19938 30480 19946 30544
rect 19626 29456 19946 30480
rect 19626 29392 19634 29456
rect 19698 29392 19714 29456
rect 19778 29392 19794 29456
rect 19858 29392 19874 29456
rect 19938 29392 19946 29456
rect 19626 28368 19946 29392
rect 19626 28304 19634 28368
rect 19698 28304 19714 28368
rect 19778 28304 19794 28368
rect 19858 28304 19874 28368
rect 19938 28304 19946 28368
rect 19626 27280 19946 28304
rect 19626 27216 19634 27280
rect 19698 27216 19714 27280
rect 19778 27216 19794 27280
rect 19858 27216 19874 27280
rect 19938 27216 19946 27280
rect 19626 26609 19946 27216
rect 22290 41968 22610 41984
rect 22290 41904 22298 41968
rect 22362 41904 22378 41968
rect 22442 41904 22458 41968
rect 22522 41904 22538 41968
rect 22602 41904 22610 41968
rect 22290 40880 22610 41904
rect 22290 40816 22298 40880
rect 22362 40816 22378 40880
rect 22442 40816 22458 40880
rect 22522 40816 22538 40880
rect 22602 40816 22610 40880
rect 22290 39792 22610 40816
rect 22290 39728 22298 39792
rect 22362 39728 22378 39792
rect 22442 39728 22458 39792
rect 22522 39728 22538 39792
rect 22602 39728 22610 39792
rect 22290 38704 22610 39728
rect 22290 38640 22298 38704
rect 22362 38640 22378 38704
rect 22442 38640 22458 38704
rect 22522 38640 22538 38704
rect 22602 38640 22610 38704
rect 22290 37616 22610 38640
rect 22290 37552 22298 37616
rect 22362 37552 22378 37616
rect 22442 37552 22458 37616
rect 22522 37552 22538 37616
rect 22602 37552 22610 37616
rect 22290 36528 22610 37552
rect 22290 36464 22298 36528
rect 22362 36464 22378 36528
rect 22442 36464 22458 36528
rect 22522 36464 22538 36528
rect 22602 36464 22610 36528
rect 22290 35440 22610 36464
rect 22290 35376 22298 35440
rect 22362 35376 22378 35440
rect 22442 35376 22458 35440
rect 22522 35376 22538 35440
rect 22602 35376 22610 35440
rect 22290 34352 22610 35376
rect 22290 34288 22298 34352
rect 22362 34288 22378 34352
rect 22442 34288 22458 34352
rect 22522 34288 22538 34352
rect 22602 34288 22610 34352
rect 22290 33264 22610 34288
rect 22290 33200 22298 33264
rect 22362 33200 22378 33264
rect 22442 33200 22458 33264
rect 22522 33200 22538 33264
rect 22602 33200 22610 33264
rect 22290 32176 22610 33200
rect 22290 32112 22298 32176
rect 22362 32112 22378 32176
rect 22442 32112 22458 32176
rect 22522 32112 22538 32176
rect 22602 32112 22610 32176
rect 22290 31088 22610 32112
rect 22290 31024 22298 31088
rect 22362 31024 22378 31088
rect 22442 31024 22458 31088
rect 22522 31024 22538 31088
rect 22602 31024 22610 31088
rect 22290 30000 22610 31024
rect 22290 29936 22298 30000
rect 22362 29936 22378 30000
rect 22442 29936 22458 30000
rect 22522 29936 22538 30000
rect 22602 29936 22610 30000
rect 22290 28912 22610 29936
rect 22290 28848 22298 28912
rect 22362 28848 22378 28912
rect 22442 28848 22458 28912
rect 22522 28848 22538 28912
rect 22602 28848 22610 28912
rect 22290 27824 22610 28848
rect 22290 27760 22298 27824
rect 22362 27760 22378 27824
rect 22442 27760 22458 27824
rect 22522 27760 22538 27824
rect 22602 27760 22610 27824
rect 22290 26736 22610 27760
rect 22290 26672 22298 26736
rect 22362 26672 22378 26736
rect 22442 26672 22458 26736
rect 22522 26672 22538 26736
rect 22602 26672 22610 26736
rect 22290 26609 22610 26672
rect 24954 41424 25274 41984
rect 24954 41360 24962 41424
rect 25026 41360 25042 41424
rect 25106 41360 25122 41424
rect 25186 41360 25202 41424
rect 25266 41360 25274 41424
rect 24954 40336 25274 41360
rect 24954 40272 24962 40336
rect 25026 40326 25042 40336
rect 25106 40326 25122 40336
rect 25186 40326 25202 40336
rect 25266 40272 25274 40336
rect 24954 40090 24996 40272
rect 25232 40090 25274 40272
rect 24954 40006 25274 40090
rect 24954 39770 24996 40006
rect 25232 39770 25274 40006
rect 24954 39248 25274 39770
rect 24954 39184 24962 39248
rect 25026 39184 25042 39248
rect 25106 39184 25122 39248
rect 25186 39184 25202 39248
rect 25266 39184 25274 39248
rect 24954 38160 25274 39184
rect 24954 38096 24962 38160
rect 25026 38096 25042 38160
rect 25106 38096 25122 38160
rect 25186 38096 25202 38160
rect 25266 38096 25274 38160
rect 24954 37072 25274 38096
rect 24954 37008 24962 37072
rect 25026 37008 25042 37072
rect 25106 37008 25122 37072
rect 25186 37008 25202 37072
rect 25266 37008 25274 37072
rect 24954 35984 25274 37008
rect 24954 35920 24962 35984
rect 25026 35920 25042 35984
rect 25106 35920 25122 35984
rect 25186 35920 25202 35984
rect 25266 35920 25274 35984
rect 24954 34896 25274 35920
rect 24954 34832 24962 34896
rect 25026 34832 25042 34896
rect 25106 34832 25122 34896
rect 25186 34832 25202 34896
rect 25266 34832 25274 34896
rect 24954 33808 25274 34832
rect 24954 33744 24962 33808
rect 25026 33744 25042 33808
rect 25106 33744 25122 33808
rect 25186 33744 25202 33808
rect 25266 33744 25274 33808
rect 24954 32720 25274 33744
rect 24954 32656 24962 32720
rect 25026 32656 25042 32720
rect 25106 32656 25122 32720
rect 25186 32656 25202 32720
rect 25266 32656 25274 32720
rect 24954 31632 25274 32656
rect 24954 31568 24962 31632
rect 25026 31568 25042 31632
rect 25106 31568 25122 31632
rect 25186 31568 25202 31632
rect 25266 31568 25274 31632
rect 24954 30544 25274 31568
rect 24954 30480 24962 30544
rect 25026 30480 25042 30544
rect 25106 30480 25122 30544
rect 25186 30480 25202 30544
rect 25266 30480 25274 30544
rect 24954 29456 25274 30480
rect 24954 29392 24962 29456
rect 25026 29392 25042 29456
rect 25106 29392 25122 29456
rect 25186 29392 25202 29456
rect 25266 29392 25274 29456
rect 24954 28368 25274 29392
rect 24954 28304 24962 28368
rect 25026 28304 25042 28368
rect 25106 28304 25122 28368
rect 25186 28304 25202 28368
rect 25266 28304 25274 28368
rect 24954 27280 25274 28304
rect 24954 27216 24962 27280
rect 25026 27216 25042 27280
rect 25106 27216 25122 27280
rect 25186 27216 25202 27280
rect 25266 27216 25274 27280
rect 24954 26609 25274 27216
rect 27618 41968 27938 41984
rect 27618 41904 27626 41968
rect 27690 41904 27706 41968
rect 27770 41904 27786 41968
rect 27850 41904 27866 41968
rect 27930 41904 27938 41968
rect 27618 40880 27938 41904
rect 27618 40816 27626 40880
rect 27690 40816 27706 40880
rect 27770 40816 27786 40880
rect 27850 40816 27866 40880
rect 27930 40816 27938 40880
rect 27618 39792 27938 40816
rect 27618 39728 27626 39792
rect 27690 39728 27706 39792
rect 27770 39728 27786 39792
rect 27850 39728 27866 39792
rect 27930 39728 27938 39792
rect 27618 38704 27938 39728
rect 27618 38640 27626 38704
rect 27690 38640 27706 38704
rect 27770 38640 27786 38704
rect 27850 38640 27866 38704
rect 27930 38640 27938 38704
rect 27618 37616 27938 38640
rect 27618 37552 27626 37616
rect 27690 37552 27706 37616
rect 27770 37552 27786 37616
rect 27850 37552 27866 37616
rect 27930 37552 27938 37616
rect 27618 36528 27938 37552
rect 27618 36464 27626 36528
rect 27690 36464 27706 36528
rect 27770 36464 27786 36528
rect 27850 36464 27866 36528
rect 27930 36464 27938 36528
rect 27618 35440 27938 36464
rect 27618 35376 27626 35440
rect 27690 35376 27706 35440
rect 27770 35376 27786 35440
rect 27850 35376 27866 35440
rect 27930 35376 27938 35440
rect 27618 34352 27938 35376
rect 27618 34288 27626 34352
rect 27690 34288 27706 34352
rect 27770 34288 27786 34352
rect 27850 34288 27866 34352
rect 27930 34288 27938 34352
rect 27618 33264 27938 34288
rect 27618 33200 27626 33264
rect 27690 33200 27706 33264
rect 27770 33200 27786 33264
rect 27850 33200 27866 33264
rect 27930 33200 27938 33264
rect 27618 32176 27938 33200
rect 27618 32112 27626 32176
rect 27690 32112 27706 32176
rect 27770 32112 27786 32176
rect 27850 32112 27866 32176
rect 27930 32112 27938 32176
rect 27618 31088 27938 32112
rect 27618 31024 27626 31088
rect 27690 31024 27706 31088
rect 27770 31024 27786 31088
rect 27850 31024 27866 31088
rect 27930 31024 27938 31088
rect 27618 30000 27938 31024
rect 27618 29936 27626 30000
rect 27690 29936 27706 30000
rect 27770 29936 27786 30000
rect 27850 29936 27866 30000
rect 27930 29936 27938 30000
rect 27618 28912 27938 29936
rect 27618 28848 27626 28912
rect 27690 28848 27706 28912
rect 27770 28848 27786 28912
rect 27850 28848 27866 28912
rect 27930 28848 27938 28912
rect 27618 27824 27938 28848
rect 27618 27760 27626 27824
rect 27690 27760 27706 27824
rect 27770 27760 27786 27824
rect 27850 27760 27866 27824
rect 27930 27760 27938 27824
rect 27618 26736 27938 27760
rect 27618 26672 27626 26736
rect 27690 26672 27706 26736
rect 27770 26672 27786 26736
rect 27850 26672 27866 26736
rect 27930 26672 27938 26736
rect 27618 26609 27938 26672
rect 30282 41424 30602 41984
rect 30282 41360 30290 41424
rect 30354 41360 30370 41424
rect 30434 41360 30450 41424
rect 30514 41360 30530 41424
rect 30594 41360 30602 41424
rect 30282 40336 30602 41360
rect 30282 40272 30290 40336
rect 30354 40326 30370 40336
rect 30434 40326 30450 40336
rect 30514 40326 30530 40336
rect 30594 40272 30602 40336
rect 30282 40090 30324 40272
rect 30560 40090 30602 40272
rect 30282 40006 30602 40090
rect 30282 39770 30324 40006
rect 30560 39770 30602 40006
rect 30282 39248 30602 39770
rect 30282 39184 30290 39248
rect 30354 39184 30370 39248
rect 30434 39184 30450 39248
rect 30514 39184 30530 39248
rect 30594 39184 30602 39248
rect 30282 38160 30602 39184
rect 30282 38096 30290 38160
rect 30354 38096 30370 38160
rect 30434 38096 30450 38160
rect 30514 38096 30530 38160
rect 30594 38096 30602 38160
rect 30282 37072 30602 38096
rect 30282 37008 30290 37072
rect 30354 37008 30370 37072
rect 30434 37008 30450 37072
rect 30514 37008 30530 37072
rect 30594 37008 30602 37072
rect 30282 35984 30602 37008
rect 30282 35920 30290 35984
rect 30354 35920 30370 35984
rect 30434 35920 30450 35984
rect 30514 35920 30530 35984
rect 30594 35920 30602 35984
rect 30282 34896 30602 35920
rect 30282 34832 30290 34896
rect 30354 34832 30370 34896
rect 30434 34832 30450 34896
rect 30514 34832 30530 34896
rect 30594 34832 30602 34896
rect 30282 33808 30602 34832
rect 30282 33744 30290 33808
rect 30354 33744 30370 33808
rect 30434 33744 30450 33808
rect 30514 33744 30530 33808
rect 30594 33744 30602 33808
rect 30282 32720 30602 33744
rect 30282 32656 30290 32720
rect 30354 32656 30370 32720
rect 30434 32656 30450 32720
rect 30514 32656 30530 32720
rect 30594 32656 30602 32720
rect 30282 31632 30602 32656
rect 30282 31568 30290 31632
rect 30354 31568 30370 31632
rect 30434 31568 30450 31632
rect 30514 31568 30530 31632
rect 30594 31568 30602 31632
rect 30282 30544 30602 31568
rect 30282 30480 30290 30544
rect 30354 30480 30370 30544
rect 30434 30480 30450 30544
rect 30514 30480 30530 30544
rect 30594 30480 30602 30544
rect 30282 29456 30602 30480
rect 30282 29392 30290 29456
rect 30354 29392 30370 29456
rect 30434 29392 30450 29456
rect 30514 29392 30530 29456
rect 30594 29392 30602 29456
rect 30282 28368 30602 29392
rect 30282 28304 30290 28368
rect 30354 28304 30370 28368
rect 30434 28304 30450 28368
rect 30514 28304 30530 28368
rect 30594 28304 30602 28368
rect 30282 27280 30602 28304
rect 30282 27216 30290 27280
rect 30354 27216 30370 27280
rect 30434 27216 30450 27280
rect 30514 27216 30530 27280
rect 30594 27216 30602 27280
rect 30282 26609 30602 27216
rect 32946 41968 33266 41984
rect 32946 41904 32954 41968
rect 33018 41904 33034 41968
rect 33098 41904 33114 41968
rect 33178 41904 33194 41968
rect 33258 41904 33266 41968
rect 32946 40880 33266 41904
rect 32946 40816 32954 40880
rect 33018 40816 33034 40880
rect 33098 40816 33114 40880
rect 33178 40816 33194 40880
rect 33258 40816 33266 40880
rect 32946 39792 33266 40816
rect 32946 39728 32954 39792
rect 33018 39728 33034 39792
rect 33098 39728 33114 39792
rect 33178 39728 33194 39792
rect 33258 39728 33266 39792
rect 32946 38704 33266 39728
rect 32946 38640 32954 38704
rect 33018 38640 33034 38704
rect 33098 38640 33114 38704
rect 33178 38640 33194 38704
rect 33258 38640 33266 38704
rect 32946 37616 33266 38640
rect 32946 37552 32954 37616
rect 33018 37552 33034 37616
rect 33098 37552 33114 37616
rect 33178 37552 33194 37616
rect 33258 37552 33266 37616
rect 32946 36528 33266 37552
rect 32946 36464 32954 36528
rect 33018 36464 33034 36528
rect 33098 36464 33114 36528
rect 33178 36464 33194 36528
rect 33258 36464 33266 36528
rect 32946 35440 33266 36464
rect 32946 35376 32954 35440
rect 33018 35376 33034 35440
rect 33098 35376 33114 35440
rect 33178 35376 33194 35440
rect 33258 35376 33266 35440
rect 32946 34352 33266 35376
rect 32946 34288 32954 34352
rect 33018 34288 33034 34352
rect 33098 34288 33114 34352
rect 33178 34288 33194 34352
rect 33258 34288 33266 34352
rect 32946 33264 33266 34288
rect 32946 33200 32954 33264
rect 33018 33200 33034 33264
rect 33098 33200 33114 33264
rect 33178 33200 33194 33264
rect 33258 33200 33266 33264
rect 32946 32176 33266 33200
rect 32946 32112 32954 32176
rect 33018 32112 33034 32176
rect 33098 32112 33114 32176
rect 33178 32112 33194 32176
rect 33258 32112 33266 32176
rect 32946 31088 33266 32112
rect 32946 31024 32954 31088
rect 33018 31024 33034 31088
rect 33098 31024 33114 31088
rect 33178 31024 33194 31088
rect 33258 31024 33266 31088
rect 32946 30000 33266 31024
rect 32946 29936 32954 30000
rect 33018 29936 33034 30000
rect 33098 29936 33114 30000
rect 33178 29936 33194 30000
rect 33258 29936 33266 30000
rect 32946 28912 33266 29936
rect 32946 28848 32954 28912
rect 33018 28848 33034 28912
rect 33098 28848 33114 28912
rect 33178 28848 33194 28912
rect 33258 28848 33266 28912
rect 32946 27824 33266 28848
rect 32946 27760 32954 27824
rect 33018 27760 33034 27824
rect 33098 27760 33114 27824
rect 33178 27760 33194 27824
rect 33258 27760 33266 27824
rect 32946 26736 33266 27760
rect 32946 26672 32954 26736
rect 33018 26672 33034 26736
rect 33098 26672 33114 26736
rect 33178 26672 33194 26736
rect 33258 26672 33266 26736
rect 32946 26609 33266 26672
rect 35610 41424 35930 41984
rect 35610 41360 35618 41424
rect 35682 41360 35698 41424
rect 35762 41360 35778 41424
rect 35842 41360 35858 41424
rect 35922 41360 35930 41424
rect 35610 40336 35930 41360
rect 35610 40272 35618 40336
rect 35682 40326 35698 40336
rect 35762 40326 35778 40336
rect 35842 40326 35858 40336
rect 35922 40272 35930 40336
rect 35610 40090 35652 40272
rect 35888 40090 35930 40272
rect 35610 40006 35930 40090
rect 35610 39770 35652 40006
rect 35888 39770 35930 40006
rect 35610 39248 35930 39770
rect 35610 39184 35618 39248
rect 35682 39184 35698 39248
rect 35762 39184 35778 39248
rect 35842 39184 35858 39248
rect 35922 39184 35930 39248
rect 35610 38160 35930 39184
rect 35610 38096 35618 38160
rect 35682 38096 35698 38160
rect 35762 38096 35778 38160
rect 35842 38096 35858 38160
rect 35922 38096 35930 38160
rect 35610 37072 35930 38096
rect 35610 37008 35618 37072
rect 35682 37008 35698 37072
rect 35762 37008 35778 37072
rect 35842 37008 35858 37072
rect 35922 37008 35930 37072
rect 35610 35984 35930 37008
rect 35610 35920 35618 35984
rect 35682 35920 35698 35984
rect 35762 35920 35778 35984
rect 35842 35920 35858 35984
rect 35922 35920 35930 35984
rect 35610 34896 35930 35920
rect 35610 34832 35618 34896
rect 35682 34832 35698 34896
rect 35762 34832 35778 34896
rect 35842 34832 35858 34896
rect 35922 34832 35930 34896
rect 35610 33808 35930 34832
rect 35610 33744 35618 33808
rect 35682 33744 35698 33808
rect 35762 33744 35778 33808
rect 35842 33744 35858 33808
rect 35922 33744 35930 33808
rect 35610 32720 35930 33744
rect 35610 32656 35618 32720
rect 35682 32656 35698 32720
rect 35762 32656 35778 32720
rect 35842 32656 35858 32720
rect 35922 32656 35930 32720
rect 35610 31632 35930 32656
rect 35610 31568 35618 31632
rect 35682 31568 35698 31632
rect 35762 31568 35778 31632
rect 35842 31568 35858 31632
rect 35922 31568 35930 31632
rect 35610 30544 35930 31568
rect 35610 30480 35618 30544
rect 35682 30480 35698 30544
rect 35762 30480 35778 30544
rect 35842 30480 35858 30544
rect 35922 30480 35930 30544
rect 35610 29456 35930 30480
rect 35610 29392 35618 29456
rect 35682 29392 35698 29456
rect 35762 29392 35778 29456
rect 35842 29392 35858 29456
rect 35922 29392 35930 29456
rect 35610 28368 35930 29392
rect 35610 28304 35618 28368
rect 35682 28304 35698 28368
rect 35762 28304 35778 28368
rect 35842 28304 35858 28368
rect 35922 28304 35930 28368
rect 35610 27280 35930 28304
rect 35610 27216 35618 27280
rect 35682 27216 35698 27280
rect 35762 27216 35778 27280
rect 35842 27216 35858 27280
rect 35922 27216 35930 27280
rect 6306 25584 6314 25648
rect 6378 25584 6394 25648
rect 6458 25584 6474 25648
rect 6538 25584 6554 25648
rect 6618 25584 6626 25648
rect 6306 24560 6626 25584
rect 6306 24496 6314 24560
rect 6378 24496 6394 24560
rect 6458 24496 6474 24560
rect 6538 24496 6554 24560
rect 6618 24496 6626 24560
rect 6306 23472 6626 24496
rect 6306 23408 6314 23472
rect 6378 23408 6394 23472
rect 6458 23408 6474 23472
rect 6538 23408 6554 23472
rect 6618 23408 6626 23472
rect 6306 22384 6626 23408
rect 35610 26192 35930 27216
rect 35610 26128 35618 26192
rect 35682 26128 35698 26192
rect 35762 26128 35778 26192
rect 35842 26128 35858 26192
rect 35922 26128 35930 26192
rect 35610 25104 35930 26128
rect 35610 25040 35618 25104
rect 35682 25040 35698 25104
rect 35762 25040 35778 25104
rect 35842 25040 35858 25104
rect 35922 25040 35930 25104
rect 35610 24016 35930 25040
rect 35610 23952 35618 24016
rect 35682 23952 35698 24016
rect 35762 23952 35778 24016
rect 35842 23952 35858 24016
rect 35922 23952 35930 24016
rect 35610 22928 35930 23952
rect 35610 22864 35618 22928
rect 35682 22864 35698 22928
rect 35762 22864 35778 22928
rect 35842 22864 35858 22928
rect 35922 22864 35930 22928
rect 31509 22452 31575 22453
rect 31509 22388 31510 22452
rect 31574 22388 31575 22452
rect 31509 22387 31575 22388
rect 6306 22320 6314 22384
rect 6378 22326 6394 22384
rect 6458 22326 6474 22384
rect 6538 22326 6554 22384
rect 6618 22320 6626 22384
rect 6306 22090 6348 22320
rect 6584 22090 6626 22320
rect 6306 22006 6626 22090
rect 6306 21770 6348 22006
rect 6584 21770 6626 22006
rect 6306 21296 6626 21770
rect 6306 21232 6314 21296
rect 6378 21232 6394 21296
rect 6458 21232 6474 21296
rect 6538 21232 6554 21296
rect 6618 21232 6626 21296
rect 6306 20208 6626 21232
rect 31512 20770 31572 22387
rect 35610 21840 35930 22864
rect 35610 21776 35618 21840
rect 35682 21776 35698 21840
rect 35762 21776 35778 21840
rect 35842 21776 35858 21840
rect 35922 21776 35930 21840
rect 35610 20752 35930 21776
rect 38274 41968 38594 41984
rect 38274 41904 38282 41968
rect 38346 41904 38362 41968
rect 38426 41904 38442 41968
rect 38506 41904 38522 41968
rect 38586 41904 38594 41968
rect 38274 40880 38594 41904
rect 38274 40816 38282 40880
rect 38346 40816 38362 40880
rect 38426 40816 38442 40880
rect 38506 40816 38522 40880
rect 38586 40816 38594 40880
rect 38274 39792 38594 40816
rect 38274 39728 38282 39792
rect 38346 39728 38362 39792
rect 38426 39728 38442 39792
rect 38506 39728 38522 39792
rect 38586 39728 38594 39792
rect 38274 38704 38594 39728
rect 38274 38640 38282 38704
rect 38346 38640 38362 38704
rect 38426 38640 38442 38704
rect 38506 38640 38522 38704
rect 38586 38640 38594 38704
rect 38274 37616 38594 38640
rect 38274 37552 38282 37616
rect 38346 37552 38362 37616
rect 38426 37552 38442 37616
rect 38506 37552 38522 37616
rect 38586 37552 38594 37616
rect 38274 36528 38594 37552
rect 38274 36464 38282 36528
rect 38346 36464 38362 36528
rect 38426 36464 38442 36528
rect 38506 36464 38522 36528
rect 38586 36464 38594 36528
rect 38274 35440 38594 36464
rect 38274 35376 38282 35440
rect 38346 35376 38362 35440
rect 38426 35376 38442 35440
rect 38506 35376 38522 35440
rect 38586 35376 38594 35440
rect 38274 34352 38594 35376
rect 38274 34288 38282 34352
rect 38346 34288 38362 34352
rect 38426 34288 38442 34352
rect 38506 34288 38522 34352
rect 38586 34288 38594 34352
rect 38274 33264 38594 34288
rect 38274 33200 38282 33264
rect 38346 33200 38362 33264
rect 38426 33200 38442 33264
rect 38506 33200 38522 33264
rect 38586 33200 38594 33264
rect 38274 32176 38594 33200
rect 38274 32112 38282 32176
rect 38346 32112 38362 32176
rect 38426 32112 38442 32176
rect 38506 32112 38522 32176
rect 38586 32112 38594 32176
rect 38274 31088 38594 32112
rect 38274 31024 38282 31088
rect 38346 31024 38362 31088
rect 38426 31024 38442 31088
rect 38506 31024 38522 31088
rect 38586 31024 38594 31088
rect 38274 30000 38594 31024
rect 38274 29936 38282 30000
rect 38346 29936 38362 30000
rect 38426 29936 38442 30000
rect 38506 29936 38522 30000
rect 38586 29936 38594 30000
rect 38274 28912 38594 29936
rect 38274 28848 38282 28912
rect 38346 28848 38362 28912
rect 38426 28848 38442 28912
rect 38506 28848 38522 28912
rect 38586 28848 38594 28912
rect 38274 27824 38594 28848
rect 38274 27760 38282 27824
rect 38346 27760 38362 27824
rect 38426 27760 38442 27824
rect 38506 27760 38522 27824
rect 38586 27760 38594 27824
rect 38274 26736 38594 27760
rect 38274 26672 38282 26736
rect 38346 26672 38362 26736
rect 38426 26672 38442 26736
rect 38506 26672 38522 26736
rect 38586 26672 38594 26736
rect 38274 25648 38594 26672
rect 38274 25584 38282 25648
rect 38346 25584 38362 25648
rect 38426 25584 38442 25648
rect 38506 25584 38522 25648
rect 38586 25584 38594 25648
rect 38274 24560 38594 25584
rect 38274 24496 38282 24560
rect 38346 24496 38362 24560
rect 38426 24496 38442 24560
rect 38506 24496 38522 24560
rect 38586 24496 38594 24560
rect 38274 23472 38594 24496
rect 38274 23408 38282 23472
rect 38346 23408 38362 23472
rect 38426 23408 38442 23472
rect 38506 23408 38522 23472
rect 38586 23408 38594 23472
rect 38274 22384 38594 23408
rect 38274 22320 38282 22384
rect 38346 22326 38362 22384
rect 38426 22326 38442 22384
rect 38506 22326 38522 22384
rect 38586 22320 38594 22384
rect 38274 22090 38316 22320
rect 38552 22090 38594 22320
rect 38274 22006 38594 22090
rect 38274 21770 38316 22006
rect 38552 21770 38594 22006
rect 37949 21500 38015 21501
rect 37949 21436 37950 21500
rect 38014 21436 38015 21500
rect 37949 21435 38015 21436
rect 37952 20770 38012 21435
rect 38274 21296 38594 21770
rect 38274 21232 38282 21296
rect 38346 21232 38362 21296
rect 38426 21232 38442 21296
rect 38506 21232 38522 21296
rect 38586 21232 38594 21296
rect 35610 20688 35618 20752
rect 35682 20688 35698 20752
rect 35762 20688 35778 20752
rect 35842 20688 35858 20752
rect 35922 20688 35930 20752
rect 31509 20276 31575 20277
rect 31509 20212 31510 20276
rect 31574 20212 31575 20276
rect 31509 20211 31575 20212
rect 6306 20144 6314 20208
rect 6378 20144 6394 20208
rect 6458 20144 6474 20208
rect 6538 20144 6554 20208
rect 6618 20144 6626 20208
rect 3642 18512 3650 18576
rect 3714 18512 3730 18576
rect 3794 18512 3810 18576
rect 3874 18512 3890 18576
rect 3954 18512 3962 18576
rect 3642 17488 3962 18512
rect 3642 17424 3650 17488
rect 3714 17424 3730 17488
rect 3794 17424 3810 17488
rect 3874 17424 3890 17488
rect 3954 17424 3962 17488
rect 3642 16400 3962 17424
rect 6306 19120 6626 20144
rect 31512 20090 31572 20211
rect 6306 19056 6314 19120
rect 6378 19056 6394 19120
rect 6458 19056 6474 19120
rect 6538 19056 6554 19120
rect 6618 19056 6626 19120
rect 6306 18032 6626 19056
rect 6306 17968 6314 18032
rect 6378 17968 6394 18032
rect 6458 17968 6474 18032
rect 6538 17968 6554 18032
rect 6618 17968 6626 18032
rect 6306 16944 6626 17968
rect 7405 17556 7471 17557
rect 7405 17492 7406 17556
rect 7470 17492 7471 17556
rect 7405 17491 7471 17492
rect 6306 16880 6314 16944
rect 6378 16880 6394 16944
rect 6458 16880 6474 16944
rect 6538 16880 6554 16944
rect 6618 16880 6626 16944
rect 3642 16336 3650 16400
rect 3714 16336 3730 16400
rect 3794 16336 3810 16400
rect 3874 16336 3890 16400
rect 3954 16336 3962 16400
rect 3642 15312 3962 16336
rect 3642 15248 3650 15312
rect 3714 15248 3730 15312
rect 3794 15248 3810 15312
rect 3874 15248 3890 15312
rect 3954 15248 3962 15312
rect 3642 14224 3962 15248
rect 3642 14160 3650 14224
rect 3714 14160 3730 14224
rect 3794 14160 3810 14224
rect 3874 14160 3890 14224
rect 3954 14160 3962 14224
rect 3642 13136 3962 14160
rect 3642 13072 3650 13136
rect 3714 13072 3730 13136
rect 3794 13072 3810 13136
rect 3874 13072 3890 13136
rect 3954 13072 3962 13136
rect 3642 12048 3962 13072
rect 3642 11984 3650 12048
rect 3714 11984 3730 12048
rect 3794 11984 3810 12048
rect 3874 11984 3890 12048
rect 3954 11984 3962 12048
rect 3642 10960 3962 11984
rect 3642 10896 3650 10960
rect 3714 10896 3730 10960
rect 3794 10896 3810 10960
rect 3874 10896 3890 10960
rect 3954 10896 3962 10960
rect 3642 9872 3962 10896
rect 3642 9808 3650 9872
rect 3714 9808 3730 9872
rect 3794 9808 3810 9872
rect 3874 9808 3890 9872
rect 3954 9808 3962 9872
rect 3642 8784 3962 9808
rect 3642 8720 3650 8784
rect 3714 8720 3730 8784
rect 3794 8720 3810 8784
rect 3874 8720 3890 8784
rect 3954 8720 3962 8784
rect 3642 7696 3962 8720
rect 3642 7632 3650 7696
rect 3714 7632 3730 7696
rect 3794 7632 3810 7696
rect 3874 7632 3890 7696
rect 3954 7632 3962 7696
rect 3642 6608 3962 7632
rect 3642 6544 3650 6608
rect 3714 6544 3730 6608
rect 3794 6544 3810 6608
rect 3874 6544 3890 6608
rect 3954 6544 3962 6608
rect 3642 5520 3962 6544
rect 3642 5456 3650 5520
rect 3714 5456 3730 5520
rect 3794 5456 3810 5520
rect 3874 5456 3890 5520
rect 3954 5456 3962 5520
rect 3642 4432 3962 5456
rect 3642 4368 3650 4432
rect 3714 4368 3730 4432
rect 3794 4368 3810 4432
rect 3874 4368 3890 4432
rect 3954 4368 3962 4432
rect 3642 4326 3962 4368
rect 3642 4090 3684 4326
rect 3920 4090 3962 4326
rect 3642 4006 3962 4090
rect 3642 3770 3684 4006
rect 3920 3770 3962 4006
rect 3642 3344 3962 3770
rect 3642 3280 3650 3344
rect 3714 3280 3730 3344
rect 3794 3280 3810 3344
rect 3874 3280 3890 3344
rect 3954 3280 3962 3344
rect 3642 2256 3962 3280
rect 3642 2192 3650 2256
rect 3714 2192 3730 2256
rect 3794 2192 3810 2256
rect 3874 2192 3890 2256
rect 3954 2192 3962 2256
rect 3642 1168 3962 2192
rect 3642 1104 3650 1168
rect 3714 1104 3730 1168
rect 3794 1104 3810 1168
rect 3874 1104 3890 1168
rect 3954 1104 3962 1168
rect 3642 80 3962 1104
rect 3642 16 3650 80
rect 3714 16 3730 80
rect 3794 16 3810 80
rect 3874 16 3890 80
rect 3954 16 3962 80
rect 3642 0 3962 16
rect 6306 15856 6626 16880
rect 7408 16010 7468 17491
rect 13664 17370 13724 19854
rect 28016 17370 28076 19854
rect 35610 19664 35930 20688
rect 35610 19600 35618 19664
rect 35682 19600 35698 19664
rect 35762 19600 35778 19664
rect 35842 19600 35858 19664
rect 35922 19600 35930 19664
rect 31509 19124 31510 19174
rect 31574 19124 31575 19174
rect 31509 19123 31575 19124
rect 35610 18576 35930 19600
rect 35610 18512 35618 18576
rect 35682 18512 35698 18576
rect 35762 18512 35778 18576
rect 35842 18512 35858 18576
rect 35922 18512 35930 18576
rect 31509 18100 31575 18101
rect 31509 18050 31510 18100
rect 31574 18050 31575 18100
rect 35610 17488 35930 18512
rect 35610 17424 35618 17488
rect 35682 17424 35698 17488
rect 35762 17424 35778 17488
rect 35842 17424 35858 17488
rect 35922 17424 35930 17488
rect 31509 17012 31575 17013
rect 31509 16948 31510 17012
rect 31574 16948 31575 17012
rect 31509 16947 31575 16948
rect 31512 16010 31572 16947
rect 35610 16400 35930 17424
rect 38274 20208 38594 21232
rect 38274 20144 38282 20208
rect 38346 20144 38362 20208
rect 38426 20144 38442 20208
rect 38506 20144 38522 20208
rect 38586 20144 38594 20208
rect 38274 19120 38594 20144
rect 38274 19056 38282 19120
rect 38346 19056 38362 19120
rect 38426 19056 38442 19120
rect 38506 19056 38522 19120
rect 38586 19056 38594 19120
rect 38274 18032 38594 19056
rect 38274 17968 38282 18032
rect 38346 17968 38362 18032
rect 38426 17968 38442 18032
rect 38506 17968 38522 18032
rect 38586 17968 38594 18032
rect 38274 16944 38594 17968
rect 38274 16880 38282 16944
rect 38346 16880 38362 16944
rect 38426 16880 38442 16944
rect 38506 16880 38522 16944
rect 38586 16880 38594 16944
rect 35610 16336 35618 16400
rect 35682 16336 35698 16400
rect 35762 16336 35778 16400
rect 35842 16336 35858 16400
rect 35922 16336 35930 16400
rect 6306 15792 6314 15856
rect 6378 15792 6394 15856
rect 6458 15792 6474 15856
rect 6538 15792 6554 15856
rect 6618 15792 6626 15856
rect 6306 14768 6626 15792
rect 35610 15312 35930 16336
rect 35610 15248 35618 15312
rect 35682 15248 35698 15312
rect 35762 15248 35778 15312
rect 35842 15248 35858 15312
rect 35922 15248 35930 15312
rect 31512 14837 31572 15094
rect 31509 14836 31575 14837
rect 31509 14772 31510 14836
rect 31574 14772 31575 14836
rect 31509 14771 31575 14772
rect 6306 14704 6314 14768
rect 6378 14704 6394 14768
rect 6458 14704 6474 14768
rect 6538 14704 6554 14768
rect 6618 14704 6626 14768
rect 6306 13680 6626 14704
rect 7405 14564 7471 14565
rect 7405 14500 7406 14564
rect 7470 14500 7471 14564
rect 7405 14499 7471 14500
rect 6306 13616 6314 13680
rect 6378 13616 6394 13680
rect 6458 13616 6474 13680
rect 6538 13616 6554 13680
rect 6618 13616 6626 13680
rect 6306 12592 6626 13616
rect 6306 12528 6314 12592
rect 6378 12528 6394 12592
rect 6458 12528 6474 12592
rect 6538 12528 6554 12592
rect 6618 12528 6626 12592
rect 6306 11504 6626 12528
rect 6306 11440 6314 11504
rect 6378 11440 6394 11504
rect 6458 11440 6474 11504
rect 6538 11440 6554 11504
rect 6618 11440 6626 11504
rect 6306 10416 6626 11440
rect 7408 11250 7468 14499
rect 35610 14224 35930 15248
rect 35610 14160 35618 14224
rect 35682 14160 35698 14224
rect 35762 14160 35778 14224
rect 35842 14160 35858 14224
rect 35922 14160 35930 14224
rect 35610 13136 35930 14160
rect 35610 13072 35618 13136
rect 35682 13072 35698 13136
rect 35762 13072 35778 13136
rect 35842 13072 35858 13136
rect 35922 13072 35930 13136
rect 35610 12048 35930 13072
rect 35610 11984 35618 12048
rect 35682 11984 35698 12048
rect 35762 11984 35778 12048
rect 35842 11984 35858 12048
rect 35922 11984 35930 12048
rect 31512 10485 31572 11014
rect 35610 10960 35930 11984
rect 35610 10896 35618 10960
rect 35682 10896 35698 10960
rect 35762 10896 35778 10960
rect 35842 10896 35858 10960
rect 35922 10896 35930 10960
rect 31509 10484 31575 10485
rect 31509 10420 31510 10484
rect 31574 10420 31575 10484
rect 31509 10419 31575 10420
rect 6306 10352 6314 10416
rect 6378 10352 6394 10416
rect 6458 10352 6474 10416
rect 6538 10352 6554 10416
rect 6618 10352 6626 10416
rect 6306 9328 6626 10352
rect 6306 9264 6314 9328
rect 6378 9264 6394 9328
rect 6458 9264 6474 9328
rect 6538 9264 6554 9328
rect 6618 9264 6626 9328
rect 6306 8240 6626 9264
rect 6306 8176 6314 8240
rect 6378 8176 6394 8240
rect 6458 8176 6474 8240
rect 6538 8176 6554 8240
rect 6618 8176 6626 8240
rect 6306 7152 6626 8176
rect 6306 7088 6314 7152
rect 6378 7088 6394 7152
rect 6458 7088 6474 7152
rect 6538 7088 6554 7152
rect 6618 7088 6626 7152
rect 6306 6064 6626 7088
rect 6306 6000 6314 6064
rect 6378 6000 6394 6064
rect 6458 6000 6474 6064
rect 6538 6000 6554 6064
rect 6618 6000 6626 6064
rect 6306 4976 6626 6000
rect 6306 4912 6314 4976
rect 6378 4912 6394 4976
rect 6458 4912 6474 4976
rect 6538 4912 6554 4976
rect 6618 4912 6626 4976
rect 6306 3888 6626 4912
rect 6306 3824 6314 3888
rect 6378 3824 6394 3888
rect 6458 3824 6474 3888
rect 6538 3824 6554 3888
rect 6618 3824 6626 3888
rect 6306 2800 6626 3824
rect 6306 2736 6314 2800
rect 6378 2736 6394 2800
rect 6458 2736 6474 2800
rect 6538 2736 6554 2800
rect 6618 2736 6626 2800
rect 6306 1712 6626 2736
rect 6306 1648 6314 1712
rect 6378 1648 6394 1712
rect 6458 1648 6474 1712
rect 6538 1648 6554 1712
rect 6618 1648 6626 1712
rect 6306 624 6626 1648
rect 6306 560 6314 624
rect 6378 560 6394 624
rect 6458 560 6474 624
rect 6538 560 6554 624
rect 6618 560 6626 624
rect 6306 0 6626 560
rect 35610 9872 35930 10896
rect 35610 9808 35618 9872
rect 35682 9808 35698 9872
rect 35762 9808 35778 9872
rect 35842 9808 35858 9872
rect 35922 9808 35930 9872
rect 35610 8784 35930 9808
rect 35610 8720 35618 8784
rect 35682 8720 35698 8784
rect 35762 8720 35778 8784
rect 35842 8720 35858 8784
rect 35922 8720 35930 8784
rect 35610 7696 35930 8720
rect 35610 7632 35618 7696
rect 35682 7632 35698 7696
rect 35762 7632 35778 7696
rect 35842 7632 35858 7696
rect 35922 7632 35930 7696
rect 35610 6608 35930 7632
rect 35610 6544 35618 6608
rect 35682 6544 35698 6608
rect 35762 6544 35778 6608
rect 35842 6544 35858 6608
rect 35922 6544 35930 6608
rect 35610 5520 35930 6544
rect 35610 5456 35618 5520
rect 35682 5456 35698 5520
rect 35762 5456 35778 5520
rect 35842 5456 35858 5520
rect 35922 5456 35930 5520
rect 35610 4432 35930 5456
rect 35610 4368 35618 4432
rect 35682 4368 35698 4432
rect 35762 4368 35778 4432
rect 35842 4368 35858 4432
rect 35922 4368 35930 4432
rect 35610 4326 35930 4368
rect 35610 4090 35652 4326
rect 35888 4090 35930 4326
rect 35610 4006 35930 4090
rect 35610 3770 35652 4006
rect 35888 3770 35930 4006
rect 35610 3344 35930 3770
rect 35610 3280 35618 3344
rect 35682 3280 35698 3344
rect 35762 3280 35778 3344
rect 35842 3280 35858 3344
rect 35922 3280 35930 3344
rect 35610 2256 35930 3280
rect 35610 2192 35618 2256
rect 35682 2192 35698 2256
rect 35762 2192 35778 2256
rect 35842 2192 35858 2256
rect 35922 2192 35930 2256
rect 35610 1168 35930 2192
rect 35610 1104 35618 1168
rect 35682 1104 35698 1168
rect 35762 1104 35778 1168
rect 35842 1104 35858 1168
rect 35922 1104 35930 1168
rect 35610 80 35930 1104
rect 35610 16 35618 80
rect 35682 16 35698 80
rect 35762 16 35778 80
rect 35842 16 35858 80
rect 35922 16 35930 80
rect 35610 0 35930 16
rect 38274 15856 38594 16880
rect 38274 15792 38282 15856
rect 38346 15792 38362 15856
rect 38426 15792 38442 15856
rect 38506 15792 38522 15856
rect 38586 15792 38594 15856
rect 38274 14768 38594 15792
rect 38274 14704 38282 14768
rect 38346 14704 38362 14768
rect 38426 14704 38442 14768
rect 38506 14704 38522 14768
rect 38586 14704 38594 14768
rect 38274 13680 38594 14704
rect 38274 13616 38282 13680
rect 38346 13616 38362 13680
rect 38426 13616 38442 13680
rect 38506 13616 38522 13680
rect 38586 13616 38594 13680
rect 38274 12592 38594 13616
rect 38274 12528 38282 12592
rect 38346 12528 38362 12592
rect 38426 12528 38442 12592
rect 38506 12528 38522 12592
rect 38586 12528 38594 12592
rect 38274 11504 38594 12528
rect 38274 11440 38282 11504
rect 38346 11440 38362 11504
rect 38426 11440 38442 11504
rect 38506 11440 38522 11504
rect 38586 11440 38594 11504
rect 38274 10416 38594 11440
rect 38274 10352 38282 10416
rect 38346 10352 38362 10416
rect 38426 10352 38442 10416
rect 38506 10352 38522 10416
rect 38586 10352 38594 10416
rect 38274 9328 38594 10352
rect 38274 9264 38282 9328
rect 38346 9264 38362 9328
rect 38426 9264 38442 9328
rect 38506 9264 38522 9328
rect 38586 9264 38594 9328
rect 38274 8240 38594 9264
rect 38274 8176 38282 8240
rect 38346 8176 38362 8240
rect 38426 8176 38442 8240
rect 38506 8176 38522 8240
rect 38586 8176 38594 8240
rect 38274 7152 38594 8176
rect 38274 7088 38282 7152
rect 38346 7088 38362 7152
rect 38426 7088 38442 7152
rect 38506 7088 38522 7152
rect 38586 7088 38594 7152
rect 38274 6064 38594 7088
rect 38274 6000 38282 6064
rect 38346 6000 38362 6064
rect 38426 6000 38442 6064
rect 38506 6000 38522 6064
rect 38586 6000 38594 6064
rect 38274 4976 38594 6000
rect 38274 4912 38282 4976
rect 38346 4912 38362 4976
rect 38426 4912 38442 4976
rect 38506 4912 38522 4976
rect 38586 4912 38594 4976
rect 38274 3888 38594 4912
rect 38274 3824 38282 3888
rect 38346 3824 38362 3888
rect 38426 3824 38442 3888
rect 38506 3824 38522 3888
rect 38586 3824 38594 3888
rect 38274 2800 38594 3824
rect 38274 2736 38282 2800
rect 38346 2736 38362 2800
rect 38426 2736 38442 2800
rect 38506 2736 38522 2800
rect 38586 2736 38594 2800
rect 38274 1712 38594 2736
rect 38274 1648 38282 1712
rect 38346 1648 38362 1712
rect 38426 1648 38442 1712
rect 38506 1648 38522 1712
rect 38586 1648 38594 1712
rect 38274 624 38594 1648
rect 38274 560 38282 624
rect 38346 560 38362 624
rect 38426 560 38442 624
rect 38506 560 38522 624
rect 38586 560 38594 624
rect 38274 0 38594 560
rect 40938 41424 41258 41984
rect 40938 41360 40946 41424
rect 41010 41360 41026 41424
rect 41090 41360 41106 41424
rect 41170 41360 41186 41424
rect 41250 41360 41258 41424
rect 40938 40336 41258 41360
rect 40938 40272 40946 40336
rect 41010 40326 41026 40336
rect 41090 40326 41106 40336
rect 41170 40326 41186 40336
rect 41250 40272 41258 40336
rect 40938 40090 40980 40272
rect 41216 40090 41258 40272
rect 40938 40006 41258 40090
rect 40938 39770 40980 40006
rect 41216 39770 41258 40006
rect 40938 39248 41258 39770
rect 40938 39184 40946 39248
rect 41010 39184 41026 39248
rect 41090 39184 41106 39248
rect 41170 39184 41186 39248
rect 41250 39184 41258 39248
rect 40938 38160 41258 39184
rect 40938 38096 40946 38160
rect 41010 38096 41026 38160
rect 41090 38096 41106 38160
rect 41170 38096 41186 38160
rect 41250 38096 41258 38160
rect 40938 37072 41258 38096
rect 40938 37008 40946 37072
rect 41010 37008 41026 37072
rect 41090 37008 41106 37072
rect 41170 37008 41186 37072
rect 41250 37008 41258 37072
rect 40938 35984 41258 37008
rect 40938 35920 40946 35984
rect 41010 35920 41026 35984
rect 41090 35920 41106 35984
rect 41170 35920 41186 35984
rect 41250 35920 41258 35984
rect 40938 34896 41258 35920
rect 40938 34832 40946 34896
rect 41010 34832 41026 34896
rect 41090 34832 41106 34896
rect 41170 34832 41186 34896
rect 41250 34832 41258 34896
rect 40938 33808 41258 34832
rect 40938 33744 40946 33808
rect 41010 33744 41026 33808
rect 41090 33744 41106 33808
rect 41170 33744 41186 33808
rect 41250 33744 41258 33808
rect 40938 32720 41258 33744
rect 40938 32656 40946 32720
rect 41010 32656 41026 32720
rect 41090 32656 41106 32720
rect 41170 32656 41186 32720
rect 41250 32656 41258 32720
rect 40938 31632 41258 32656
rect 40938 31568 40946 31632
rect 41010 31568 41026 31632
rect 41090 31568 41106 31632
rect 41170 31568 41186 31632
rect 41250 31568 41258 31632
rect 40938 30544 41258 31568
rect 40938 30480 40946 30544
rect 41010 30480 41026 30544
rect 41090 30480 41106 30544
rect 41170 30480 41186 30544
rect 41250 30480 41258 30544
rect 40938 29456 41258 30480
rect 40938 29392 40946 29456
rect 41010 29392 41026 29456
rect 41090 29392 41106 29456
rect 41170 29392 41186 29456
rect 41250 29392 41258 29456
rect 40938 28368 41258 29392
rect 40938 28304 40946 28368
rect 41010 28304 41026 28368
rect 41090 28304 41106 28368
rect 41170 28304 41186 28368
rect 41250 28304 41258 28368
rect 40938 27280 41258 28304
rect 40938 27216 40946 27280
rect 41010 27216 41026 27280
rect 41090 27216 41106 27280
rect 41170 27216 41186 27280
rect 41250 27216 41258 27280
rect 40938 26192 41258 27216
rect 43602 41968 43922 41984
rect 43602 41904 43610 41968
rect 43674 41904 43690 41968
rect 43754 41904 43770 41968
rect 43834 41904 43850 41968
rect 43914 41904 43922 41968
rect 43602 40880 43922 41904
rect 43602 40816 43610 40880
rect 43674 40816 43690 40880
rect 43754 40816 43770 40880
rect 43834 40816 43850 40880
rect 43914 40816 43922 40880
rect 43602 39792 43922 40816
rect 43602 39728 43610 39792
rect 43674 39728 43690 39792
rect 43754 39728 43770 39792
rect 43834 39728 43850 39792
rect 43914 39728 43922 39792
rect 43602 38704 43922 39728
rect 43602 38640 43610 38704
rect 43674 38640 43690 38704
rect 43754 38640 43770 38704
rect 43834 38640 43850 38704
rect 43914 38640 43922 38704
rect 43602 37616 43922 38640
rect 43602 37552 43610 37616
rect 43674 37552 43690 37616
rect 43754 37552 43770 37616
rect 43834 37552 43850 37616
rect 43914 37552 43922 37616
rect 43602 36528 43922 37552
rect 43602 36464 43610 36528
rect 43674 36464 43690 36528
rect 43754 36464 43770 36528
rect 43834 36464 43850 36528
rect 43914 36464 43922 36528
rect 43602 35440 43922 36464
rect 43602 35376 43610 35440
rect 43674 35376 43690 35440
rect 43754 35376 43770 35440
rect 43834 35376 43850 35440
rect 43914 35376 43922 35440
rect 43602 34352 43922 35376
rect 43602 34288 43610 34352
rect 43674 34288 43690 34352
rect 43754 34288 43770 34352
rect 43834 34288 43850 34352
rect 43914 34288 43922 34352
rect 43602 33264 43922 34288
rect 43602 33200 43610 33264
rect 43674 33200 43690 33264
rect 43754 33200 43770 33264
rect 43834 33200 43850 33264
rect 43914 33200 43922 33264
rect 43602 32176 43922 33200
rect 43602 32112 43610 32176
rect 43674 32112 43690 32176
rect 43754 32112 43770 32176
rect 43834 32112 43850 32176
rect 43914 32112 43922 32176
rect 43602 31088 43922 32112
rect 43602 31024 43610 31088
rect 43674 31024 43690 31088
rect 43754 31024 43770 31088
rect 43834 31024 43850 31088
rect 43914 31024 43922 31088
rect 43602 30000 43922 31024
rect 43602 29936 43610 30000
rect 43674 29936 43690 30000
rect 43754 29936 43770 30000
rect 43834 29936 43850 30000
rect 43914 29936 43922 30000
rect 43602 28912 43922 29936
rect 43602 28848 43610 28912
rect 43674 28848 43690 28912
rect 43754 28848 43770 28912
rect 43834 28848 43850 28912
rect 43914 28848 43922 28912
rect 43602 27824 43922 28848
rect 43602 27760 43610 27824
rect 43674 27760 43690 27824
rect 43754 27760 43770 27824
rect 43834 27760 43850 27824
rect 43914 27760 43922 27824
rect 43602 26736 43922 27760
rect 43602 26672 43610 26736
rect 43674 26672 43690 26736
rect 43754 26672 43770 26736
rect 43834 26672 43850 26736
rect 43914 26672 43922 26736
rect 43602 26609 43922 26672
rect 46266 41424 46586 41984
rect 46266 41360 46274 41424
rect 46338 41360 46354 41424
rect 46418 41360 46434 41424
rect 46498 41360 46514 41424
rect 46578 41360 46586 41424
rect 46266 40336 46586 41360
rect 46266 40272 46274 40336
rect 46338 40326 46354 40336
rect 46418 40326 46434 40336
rect 46498 40326 46514 40336
rect 46578 40272 46586 40336
rect 46266 40090 46308 40272
rect 46544 40090 46586 40272
rect 46266 40006 46586 40090
rect 46266 39770 46308 40006
rect 46544 39770 46586 40006
rect 46266 39248 46586 39770
rect 46266 39184 46274 39248
rect 46338 39184 46354 39248
rect 46418 39184 46434 39248
rect 46498 39184 46514 39248
rect 46578 39184 46586 39248
rect 46266 38160 46586 39184
rect 46266 38096 46274 38160
rect 46338 38096 46354 38160
rect 46418 38096 46434 38160
rect 46498 38096 46514 38160
rect 46578 38096 46586 38160
rect 46266 37072 46586 38096
rect 46266 37008 46274 37072
rect 46338 37008 46354 37072
rect 46418 37008 46434 37072
rect 46498 37008 46514 37072
rect 46578 37008 46586 37072
rect 46266 35984 46586 37008
rect 46266 35920 46274 35984
rect 46338 35920 46354 35984
rect 46418 35920 46434 35984
rect 46498 35920 46514 35984
rect 46578 35920 46586 35984
rect 46266 34896 46586 35920
rect 46266 34832 46274 34896
rect 46338 34832 46354 34896
rect 46418 34832 46434 34896
rect 46498 34832 46514 34896
rect 46578 34832 46586 34896
rect 46266 33808 46586 34832
rect 46266 33744 46274 33808
rect 46338 33744 46354 33808
rect 46418 33744 46434 33808
rect 46498 33744 46514 33808
rect 46578 33744 46586 33808
rect 46266 32720 46586 33744
rect 46266 32656 46274 32720
rect 46338 32656 46354 32720
rect 46418 32656 46434 32720
rect 46498 32656 46514 32720
rect 46578 32656 46586 32720
rect 46266 31632 46586 32656
rect 46266 31568 46274 31632
rect 46338 31568 46354 31632
rect 46418 31568 46434 31632
rect 46498 31568 46514 31632
rect 46578 31568 46586 31632
rect 46266 30544 46586 31568
rect 46266 30480 46274 30544
rect 46338 30480 46354 30544
rect 46418 30480 46434 30544
rect 46498 30480 46514 30544
rect 46578 30480 46586 30544
rect 46266 29456 46586 30480
rect 46266 29392 46274 29456
rect 46338 29392 46354 29456
rect 46418 29392 46434 29456
rect 46498 29392 46514 29456
rect 46578 29392 46586 29456
rect 46266 28368 46586 29392
rect 46266 28304 46274 28368
rect 46338 28304 46354 28368
rect 46418 28304 46434 28368
rect 46498 28304 46514 28368
rect 46578 28304 46586 28368
rect 46266 27280 46586 28304
rect 46266 27216 46274 27280
rect 46338 27216 46354 27280
rect 46418 27216 46434 27280
rect 46498 27216 46514 27280
rect 46578 27216 46586 27280
rect 46266 26609 46586 27216
rect 48930 41968 49250 41984
rect 48930 41904 48938 41968
rect 49002 41904 49018 41968
rect 49082 41904 49098 41968
rect 49162 41904 49178 41968
rect 49242 41904 49250 41968
rect 48930 40880 49250 41904
rect 48930 40816 48938 40880
rect 49002 40816 49018 40880
rect 49082 40816 49098 40880
rect 49162 40816 49178 40880
rect 49242 40816 49250 40880
rect 48930 39792 49250 40816
rect 48930 39728 48938 39792
rect 49002 39728 49018 39792
rect 49082 39728 49098 39792
rect 49162 39728 49178 39792
rect 49242 39728 49250 39792
rect 48930 38704 49250 39728
rect 48930 38640 48938 38704
rect 49002 38640 49018 38704
rect 49082 38640 49098 38704
rect 49162 38640 49178 38704
rect 49242 38640 49250 38704
rect 48930 37616 49250 38640
rect 48930 37552 48938 37616
rect 49002 37552 49018 37616
rect 49082 37552 49098 37616
rect 49162 37552 49178 37616
rect 49242 37552 49250 37616
rect 48930 36528 49250 37552
rect 48930 36464 48938 36528
rect 49002 36464 49018 36528
rect 49082 36464 49098 36528
rect 49162 36464 49178 36528
rect 49242 36464 49250 36528
rect 48930 35440 49250 36464
rect 48930 35376 48938 35440
rect 49002 35376 49018 35440
rect 49082 35376 49098 35440
rect 49162 35376 49178 35440
rect 49242 35376 49250 35440
rect 48930 34352 49250 35376
rect 48930 34288 48938 34352
rect 49002 34288 49018 34352
rect 49082 34288 49098 34352
rect 49162 34288 49178 34352
rect 49242 34288 49250 34352
rect 48930 33264 49250 34288
rect 48930 33200 48938 33264
rect 49002 33200 49018 33264
rect 49082 33200 49098 33264
rect 49162 33200 49178 33264
rect 49242 33200 49250 33264
rect 48930 32176 49250 33200
rect 48930 32112 48938 32176
rect 49002 32112 49018 32176
rect 49082 32112 49098 32176
rect 49162 32112 49178 32176
rect 49242 32112 49250 32176
rect 48930 31088 49250 32112
rect 48930 31024 48938 31088
rect 49002 31024 49018 31088
rect 49082 31024 49098 31088
rect 49162 31024 49178 31088
rect 49242 31024 49250 31088
rect 48930 30000 49250 31024
rect 48930 29936 48938 30000
rect 49002 29936 49018 30000
rect 49082 29936 49098 30000
rect 49162 29936 49178 30000
rect 49242 29936 49250 30000
rect 48930 28912 49250 29936
rect 48930 28848 48938 28912
rect 49002 28848 49018 28912
rect 49082 28848 49098 28912
rect 49162 28848 49178 28912
rect 49242 28848 49250 28912
rect 48930 27824 49250 28848
rect 48930 27760 48938 27824
rect 49002 27760 49018 27824
rect 49082 27760 49098 27824
rect 49162 27760 49178 27824
rect 49242 27760 49250 27824
rect 48930 26736 49250 27760
rect 48930 26672 48938 26736
rect 49002 26672 49018 26736
rect 49082 26672 49098 26736
rect 49162 26672 49178 26736
rect 49242 26672 49250 26736
rect 48930 26609 49250 26672
rect 51594 41424 51914 41984
rect 51594 41360 51602 41424
rect 51666 41360 51682 41424
rect 51746 41360 51762 41424
rect 51826 41360 51842 41424
rect 51906 41360 51914 41424
rect 51594 40336 51914 41360
rect 51594 40272 51602 40336
rect 51666 40326 51682 40336
rect 51746 40326 51762 40336
rect 51826 40326 51842 40336
rect 51906 40272 51914 40336
rect 51594 40090 51636 40272
rect 51872 40090 51914 40272
rect 51594 40006 51914 40090
rect 51594 39770 51636 40006
rect 51872 39770 51914 40006
rect 51594 39248 51914 39770
rect 51594 39184 51602 39248
rect 51666 39184 51682 39248
rect 51746 39184 51762 39248
rect 51826 39184 51842 39248
rect 51906 39184 51914 39248
rect 51594 38160 51914 39184
rect 51594 38096 51602 38160
rect 51666 38096 51682 38160
rect 51746 38096 51762 38160
rect 51826 38096 51842 38160
rect 51906 38096 51914 38160
rect 51594 37072 51914 38096
rect 51594 37008 51602 37072
rect 51666 37008 51682 37072
rect 51746 37008 51762 37072
rect 51826 37008 51842 37072
rect 51906 37008 51914 37072
rect 51594 35984 51914 37008
rect 51594 35920 51602 35984
rect 51666 35920 51682 35984
rect 51746 35920 51762 35984
rect 51826 35920 51842 35984
rect 51906 35920 51914 35984
rect 51594 34896 51914 35920
rect 51594 34832 51602 34896
rect 51666 34832 51682 34896
rect 51746 34832 51762 34896
rect 51826 34832 51842 34896
rect 51906 34832 51914 34896
rect 51594 33808 51914 34832
rect 51594 33744 51602 33808
rect 51666 33744 51682 33808
rect 51746 33744 51762 33808
rect 51826 33744 51842 33808
rect 51906 33744 51914 33808
rect 51594 32720 51914 33744
rect 51594 32656 51602 32720
rect 51666 32656 51682 32720
rect 51746 32656 51762 32720
rect 51826 32656 51842 32720
rect 51906 32656 51914 32720
rect 51594 31632 51914 32656
rect 51594 31568 51602 31632
rect 51666 31568 51682 31632
rect 51746 31568 51762 31632
rect 51826 31568 51842 31632
rect 51906 31568 51914 31632
rect 51594 30544 51914 31568
rect 51594 30480 51602 30544
rect 51666 30480 51682 30544
rect 51746 30480 51762 30544
rect 51826 30480 51842 30544
rect 51906 30480 51914 30544
rect 51594 29456 51914 30480
rect 51594 29392 51602 29456
rect 51666 29392 51682 29456
rect 51746 29392 51762 29456
rect 51826 29392 51842 29456
rect 51906 29392 51914 29456
rect 51594 28368 51914 29392
rect 51594 28304 51602 28368
rect 51666 28304 51682 28368
rect 51746 28304 51762 28368
rect 51826 28304 51842 28368
rect 51906 28304 51914 28368
rect 51594 27280 51914 28304
rect 51594 27216 51602 27280
rect 51666 27216 51682 27280
rect 51746 27216 51762 27280
rect 51826 27216 51842 27280
rect 51906 27216 51914 27280
rect 51594 26609 51914 27216
rect 54258 41968 54578 41984
rect 54258 41904 54266 41968
rect 54330 41904 54346 41968
rect 54410 41904 54426 41968
rect 54490 41904 54506 41968
rect 54570 41904 54578 41968
rect 54258 40880 54578 41904
rect 54258 40816 54266 40880
rect 54330 40816 54346 40880
rect 54410 40816 54426 40880
rect 54490 40816 54506 40880
rect 54570 40816 54578 40880
rect 54258 39792 54578 40816
rect 54258 39728 54266 39792
rect 54330 39728 54346 39792
rect 54410 39728 54426 39792
rect 54490 39728 54506 39792
rect 54570 39728 54578 39792
rect 54258 38704 54578 39728
rect 54258 38640 54266 38704
rect 54330 38640 54346 38704
rect 54410 38640 54426 38704
rect 54490 38640 54506 38704
rect 54570 38640 54578 38704
rect 54258 37616 54578 38640
rect 54258 37552 54266 37616
rect 54330 37552 54346 37616
rect 54410 37552 54426 37616
rect 54490 37552 54506 37616
rect 54570 37552 54578 37616
rect 54258 36528 54578 37552
rect 54258 36464 54266 36528
rect 54330 36464 54346 36528
rect 54410 36464 54426 36528
rect 54490 36464 54506 36528
rect 54570 36464 54578 36528
rect 54258 35440 54578 36464
rect 54258 35376 54266 35440
rect 54330 35376 54346 35440
rect 54410 35376 54426 35440
rect 54490 35376 54506 35440
rect 54570 35376 54578 35440
rect 54258 34352 54578 35376
rect 54258 34288 54266 34352
rect 54330 34288 54346 34352
rect 54410 34288 54426 34352
rect 54490 34288 54506 34352
rect 54570 34288 54578 34352
rect 54258 33264 54578 34288
rect 54258 33200 54266 33264
rect 54330 33200 54346 33264
rect 54410 33200 54426 33264
rect 54490 33200 54506 33264
rect 54570 33200 54578 33264
rect 54258 32176 54578 33200
rect 54258 32112 54266 32176
rect 54330 32112 54346 32176
rect 54410 32112 54426 32176
rect 54490 32112 54506 32176
rect 54570 32112 54578 32176
rect 54258 31088 54578 32112
rect 54258 31024 54266 31088
rect 54330 31024 54346 31088
rect 54410 31024 54426 31088
rect 54490 31024 54506 31088
rect 54570 31024 54578 31088
rect 54258 30000 54578 31024
rect 54258 29936 54266 30000
rect 54330 29936 54346 30000
rect 54410 29936 54426 30000
rect 54490 29936 54506 30000
rect 54570 29936 54578 30000
rect 54258 28912 54578 29936
rect 54258 28848 54266 28912
rect 54330 28848 54346 28912
rect 54410 28848 54426 28912
rect 54490 28848 54506 28912
rect 54570 28848 54578 28912
rect 54258 27824 54578 28848
rect 54258 27760 54266 27824
rect 54330 27760 54346 27824
rect 54410 27760 54426 27824
rect 54490 27760 54506 27824
rect 54570 27760 54578 27824
rect 54258 26736 54578 27760
rect 54258 26672 54266 26736
rect 54330 26672 54346 26736
rect 54410 26672 54426 26736
rect 54490 26672 54506 26736
rect 54570 26672 54578 26736
rect 54258 26609 54578 26672
rect 56922 41424 57242 41984
rect 56922 41360 56930 41424
rect 56994 41360 57010 41424
rect 57074 41360 57090 41424
rect 57154 41360 57170 41424
rect 57234 41360 57242 41424
rect 56922 40336 57242 41360
rect 56922 40272 56930 40336
rect 56994 40326 57010 40336
rect 57074 40326 57090 40336
rect 57154 40326 57170 40336
rect 57234 40272 57242 40336
rect 56922 40090 56964 40272
rect 57200 40090 57242 40272
rect 56922 40006 57242 40090
rect 56922 39770 56964 40006
rect 57200 39770 57242 40006
rect 56922 39248 57242 39770
rect 56922 39184 56930 39248
rect 56994 39184 57010 39248
rect 57074 39184 57090 39248
rect 57154 39184 57170 39248
rect 57234 39184 57242 39248
rect 56922 38160 57242 39184
rect 56922 38096 56930 38160
rect 56994 38096 57010 38160
rect 57074 38096 57090 38160
rect 57154 38096 57170 38160
rect 57234 38096 57242 38160
rect 56922 37072 57242 38096
rect 56922 37008 56930 37072
rect 56994 37008 57010 37072
rect 57074 37008 57090 37072
rect 57154 37008 57170 37072
rect 57234 37008 57242 37072
rect 56922 35984 57242 37008
rect 56922 35920 56930 35984
rect 56994 35920 57010 35984
rect 57074 35920 57090 35984
rect 57154 35920 57170 35984
rect 57234 35920 57242 35984
rect 56922 34896 57242 35920
rect 56922 34832 56930 34896
rect 56994 34832 57010 34896
rect 57074 34832 57090 34896
rect 57154 34832 57170 34896
rect 57234 34832 57242 34896
rect 56922 33808 57242 34832
rect 56922 33744 56930 33808
rect 56994 33744 57010 33808
rect 57074 33744 57090 33808
rect 57154 33744 57170 33808
rect 57234 33744 57242 33808
rect 56922 32720 57242 33744
rect 56922 32656 56930 32720
rect 56994 32656 57010 32720
rect 57074 32656 57090 32720
rect 57154 32656 57170 32720
rect 57234 32656 57242 32720
rect 56922 31632 57242 32656
rect 56922 31568 56930 31632
rect 56994 31568 57010 31632
rect 57074 31568 57090 31632
rect 57154 31568 57170 31632
rect 57234 31568 57242 31632
rect 56922 30544 57242 31568
rect 56922 30480 56930 30544
rect 56994 30480 57010 30544
rect 57074 30480 57090 30544
rect 57154 30480 57170 30544
rect 57234 30480 57242 30544
rect 56922 29456 57242 30480
rect 56922 29392 56930 29456
rect 56994 29392 57010 29456
rect 57074 29392 57090 29456
rect 57154 29392 57170 29456
rect 57234 29392 57242 29456
rect 56922 28368 57242 29392
rect 56922 28304 56930 28368
rect 56994 28304 57010 28368
rect 57074 28304 57090 28368
rect 57154 28304 57170 28368
rect 57234 28304 57242 28368
rect 56922 27280 57242 28304
rect 56922 27216 56930 27280
rect 56994 27216 57010 27280
rect 57074 27216 57090 27280
rect 57154 27216 57170 27280
rect 57234 27216 57242 27280
rect 56922 26609 57242 27216
rect 59586 41968 59906 41984
rect 59586 41904 59594 41968
rect 59658 41904 59674 41968
rect 59738 41904 59754 41968
rect 59818 41904 59834 41968
rect 59898 41904 59906 41968
rect 59586 40880 59906 41904
rect 59586 40816 59594 40880
rect 59658 40816 59674 40880
rect 59738 40816 59754 40880
rect 59818 40816 59834 40880
rect 59898 40816 59906 40880
rect 59586 39792 59906 40816
rect 59586 39728 59594 39792
rect 59658 39728 59674 39792
rect 59738 39728 59754 39792
rect 59818 39728 59834 39792
rect 59898 39728 59906 39792
rect 59586 38704 59906 39728
rect 59586 38640 59594 38704
rect 59658 38640 59674 38704
rect 59738 38640 59754 38704
rect 59818 38640 59834 38704
rect 59898 38640 59906 38704
rect 59586 37616 59906 38640
rect 59586 37552 59594 37616
rect 59658 37552 59674 37616
rect 59738 37552 59754 37616
rect 59818 37552 59834 37616
rect 59898 37552 59906 37616
rect 59586 36528 59906 37552
rect 59586 36464 59594 36528
rect 59658 36464 59674 36528
rect 59738 36464 59754 36528
rect 59818 36464 59834 36528
rect 59898 36464 59906 36528
rect 59586 35440 59906 36464
rect 59586 35376 59594 35440
rect 59658 35376 59674 35440
rect 59738 35376 59754 35440
rect 59818 35376 59834 35440
rect 59898 35376 59906 35440
rect 59586 34352 59906 35376
rect 59586 34288 59594 34352
rect 59658 34288 59674 34352
rect 59738 34288 59754 34352
rect 59818 34288 59834 34352
rect 59898 34288 59906 34352
rect 59586 33264 59906 34288
rect 59586 33200 59594 33264
rect 59658 33200 59674 33264
rect 59738 33200 59754 33264
rect 59818 33200 59834 33264
rect 59898 33200 59906 33264
rect 59586 32176 59906 33200
rect 59586 32112 59594 32176
rect 59658 32112 59674 32176
rect 59738 32112 59754 32176
rect 59818 32112 59834 32176
rect 59898 32112 59906 32176
rect 59586 31088 59906 32112
rect 59586 31024 59594 31088
rect 59658 31024 59674 31088
rect 59738 31024 59754 31088
rect 59818 31024 59834 31088
rect 59898 31024 59906 31088
rect 59586 30000 59906 31024
rect 59586 29936 59594 30000
rect 59658 29936 59674 30000
rect 59738 29936 59754 30000
rect 59818 29936 59834 30000
rect 59898 29936 59906 30000
rect 59586 28912 59906 29936
rect 59586 28848 59594 28912
rect 59658 28848 59674 28912
rect 59738 28848 59754 28912
rect 59818 28848 59834 28912
rect 59898 28848 59906 28912
rect 59586 27824 59906 28848
rect 59586 27760 59594 27824
rect 59658 27760 59674 27824
rect 59738 27760 59754 27824
rect 59818 27760 59834 27824
rect 59898 27760 59906 27824
rect 59586 26736 59906 27760
rect 59586 26672 59594 26736
rect 59658 26672 59674 26736
rect 59738 26672 59754 26736
rect 59818 26672 59834 26736
rect 59898 26672 59906 26736
rect 59586 26609 59906 26672
rect 62250 41424 62570 41984
rect 62250 41360 62258 41424
rect 62322 41360 62338 41424
rect 62402 41360 62418 41424
rect 62482 41360 62498 41424
rect 62562 41360 62570 41424
rect 62250 40336 62570 41360
rect 62250 40272 62258 40336
rect 62322 40326 62338 40336
rect 62402 40326 62418 40336
rect 62482 40326 62498 40336
rect 62562 40272 62570 40336
rect 62250 40090 62292 40272
rect 62528 40090 62570 40272
rect 62250 40006 62570 40090
rect 62250 39770 62292 40006
rect 62528 39770 62570 40006
rect 62250 39248 62570 39770
rect 62250 39184 62258 39248
rect 62322 39184 62338 39248
rect 62402 39184 62418 39248
rect 62482 39184 62498 39248
rect 62562 39184 62570 39248
rect 62250 38160 62570 39184
rect 62250 38096 62258 38160
rect 62322 38096 62338 38160
rect 62402 38096 62418 38160
rect 62482 38096 62498 38160
rect 62562 38096 62570 38160
rect 62250 37072 62570 38096
rect 62250 37008 62258 37072
rect 62322 37008 62338 37072
rect 62402 37008 62418 37072
rect 62482 37008 62498 37072
rect 62562 37008 62570 37072
rect 62250 35984 62570 37008
rect 62250 35920 62258 35984
rect 62322 35920 62338 35984
rect 62402 35920 62418 35984
rect 62482 35920 62498 35984
rect 62562 35920 62570 35984
rect 62250 34896 62570 35920
rect 62250 34832 62258 34896
rect 62322 34832 62338 34896
rect 62402 34832 62418 34896
rect 62482 34832 62498 34896
rect 62562 34832 62570 34896
rect 62250 33808 62570 34832
rect 62250 33744 62258 33808
rect 62322 33744 62338 33808
rect 62402 33744 62418 33808
rect 62482 33744 62498 33808
rect 62562 33744 62570 33808
rect 62250 32720 62570 33744
rect 62250 32656 62258 32720
rect 62322 32656 62338 32720
rect 62402 32656 62418 32720
rect 62482 32656 62498 32720
rect 62562 32656 62570 32720
rect 62250 31632 62570 32656
rect 62250 31568 62258 31632
rect 62322 31568 62338 31632
rect 62402 31568 62418 31632
rect 62482 31568 62498 31632
rect 62562 31568 62570 31632
rect 62250 30544 62570 31568
rect 62250 30480 62258 30544
rect 62322 30480 62338 30544
rect 62402 30480 62418 30544
rect 62482 30480 62498 30544
rect 62562 30480 62570 30544
rect 62250 29456 62570 30480
rect 62250 29392 62258 29456
rect 62322 29392 62338 29456
rect 62402 29392 62418 29456
rect 62482 29392 62498 29456
rect 62562 29392 62570 29456
rect 62250 28368 62570 29392
rect 62250 28304 62258 28368
rect 62322 28304 62338 28368
rect 62402 28304 62418 28368
rect 62482 28304 62498 28368
rect 62562 28304 62570 28368
rect 62250 27280 62570 28304
rect 62250 27216 62258 27280
rect 62322 27216 62338 27280
rect 62402 27216 62418 27280
rect 62482 27216 62498 27280
rect 62562 27216 62570 27280
rect 62250 26609 62570 27216
rect 64914 41968 65234 41984
rect 64914 41904 64922 41968
rect 64986 41904 65002 41968
rect 65066 41904 65082 41968
rect 65146 41904 65162 41968
rect 65226 41904 65234 41968
rect 64914 40880 65234 41904
rect 64914 40816 64922 40880
rect 64986 40816 65002 40880
rect 65066 40816 65082 40880
rect 65146 40816 65162 40880
rect 65226 40816 65234 40880
rect 64914 39792 65234 40816
rect 64914 39728 64922 39792
rect 64986 39728 65002 39792
rect 65066 39728 65082 39792
rect 65146 39728 65162 39792
rect 65226 39728 65234 39792
rect 64914 38704 65234 39728
rect 64914 38640 64922 38704
rect 64986 38640 65002 38704
rect 65066 38640 65082 38704
rect 65146 38640 65162 38704
rect 65226 38640 65234 38704
rect 64914 37616 65234 38640
rect 64914 37552 64922 37616
rect 64986 37552 65002 37616
rect 65066 37552 65082 37616
rect 65146 37552 65162 37616
rect 65226 37552 65234 37616
rect 64914 36528 65234 37552
rect 64914 36464 64922 36528
rect 64986 36464 65002 36528
rect 65066 36464 65082 36528
rect 65146 36464 65162 36528
rect 65226 36464 65234 36528
rect 64914 35440 65234 36464
rect 64914 35376 64922 35440
rect 64986 35376 65002 35440
rect 65066 35376 65082 35440
rect 65146 35376 65162 35440
rect 65226 35376 65234 35440
rect 64914 34352 65234 35376
rect 64914 34288 64922 34352
rect 64986 34288 65002 34352
rect 65066 34288 65082 34352
rect 65146 34288 65162 34352
rect 65226 34288 65234 34352
rect 64914 33264 65234 34288
rect 64914 33200 64922 33264
rect 64986 33200 65002 33264
rect 65066 33200 65082 33264
rect 65146 33200 65162 33264
rect 65226 33200 65234 33264
rect 64914 32176 65234 33200
rect 64914 32112 64922 32176
rect 64986 32112 65002 32176
rect 65066 32112 65082 32176
rect 65146 32112 65162 32176
rect 65226 32112 65234 32176
rect 64914 31088 65234 32112
rect 64914 31024 64922 31088
rect 64986 31024 65002 31088
rect 65066 31024 65082 31088
rect 65146 31024 65162 31088
rect 65226 31024 65234 31088
rect 64914 30000 65234 31024
rect 64914 29936 64922 30000
rect 64986 29936 65002 30000
rect 65066 29936 65082 30000
rect 65146 29936 65162 30000
rect 65226 29936 65234 30000
rect 64914 28912 65234 29936
rect 64914 28848 64922 28912
rect 64986 28848 65002 28912
rect 65066 28848 65082 28912
rect 65146 28848 65162 28912
rect 65226 28848 65234 28912
rect 64914 27824 65234 28848
rect 64914 27760 64922 27824
rect 64986 27760 65002 27824
rect 65066 27760 65082 27824
rect 65146 27760 65162 27824
rect 65226 27760 65234 27824
rect 64914 26736 65234 27760
rect 64914 26672 64922 26736
rect 64986 26672 65002 26736
rect 65066 26672 65082 26736
rect 65146 26672 65162 26736
rect 65226 26672 65234 26736
rect 64914 26609 65234 26672
rect 67578 41424 67898 41984
rect 67578 41360 67586 41424
rect 67650 41360 67666 41424
rect 67730 41360 67746 41424
rect 67810 41360 67826 41424
rect 67890 41360 67898 41424
rect 67578 40336 67898 41360
rect 67578 40272 67586 40336
rect 67650 40326 67666 40336
rect 67730 40326 67746 40336
rect 67810 40326 67826 40336
rect 67890 40272 67898 40336
rect 67578 40090 67620 40272
rect 67856 40090 67898 40272
rect 67578 40006 67898 40090
rect 67578 39770 67620 40006
rect 67856 39770 67898 40006
rect 67578 39248 67898 39770
rect 67578 39184 67586 39248
rect 67650 39184 67666 39248
rect 67730 39184 67746 39248
rect 67810 39184 67826 39248
rect 67890 39184 67898 39248
rect 67578 38160 67898 39184
rect 67578 38096 67586 38160
rect 67650 38096 67666 38160
rect 67730 38096 67746 38160
rect 67810 38096 67826 38160
rect 67890 38096 67898 38160
rect 67578 37072 67898 38096
rect 67578 37008 67586 37072
rect 67650 37008 67666 37072
rect 67730 37008 67746 37072
rect 67810 37008 67826 37072
rect 67890 37008 67898 37072
rect 67578 35984 67898 37008
rect 67578 35920 67586 35984
rect 67650 35920 67666 35984
rect 67730 35920 67746 35984
rect 67810 35920 67826 35984
rect 67890 35920 67898 35984
rect 67578 34896 67898 35920
rect 67578 34832 67586 34896
rect 67650 34832 67666 34896
rect 67730 34832 67746 34896
rect 67810 34832 67826 34896
rect 67890 34832 67898 34896
rect 67578 33808 67898 34832
rect 67578 33744 67586 33808
rect 67650 33744 67666 33808
rect 67730 33744 67746 33808
rect 67810 33744 67826 33808
rect 67890 33744 67898 33808
rect 67578 32720 67898 33744
rect 67578 32656 67586 32720
rect 67650 32656 67666 32720
rect 67730 32656 67746 32720
rect 67810 32656 67826 32720
rect 67890 32656 67898 32720
rect 67578 31632 67898 32656
rect 67578 31568 67586 31632
rect 67650 31568 67666 31632
rect 67730 31568 67746 31632
rect 67810 31568 67826 31632
rect 67890 31568 67898 31632
rect 67578 30544 67898 31568
rect 67578 30480 67586 30544
rect 67650 30480 67666 30544
rect 67730 30480 67746 30544
rect 67810 30480 67826 30544
rect 67890 30480 67898 30544
rect 67578 29456 67898 30480
rect 67578 29392 67586 29456
rect 67650 29392 67666 29456
rect 67730 29392 67746 29456
rect 67810 29392 67826 29456
rect 67890 29392 67898 29456
rect 67578 28368 67898 29392
rect 67578 28304 67586 28368
rect 67650 28304 67666 28368
rect 67730 28304 67746 28368
rect 67810 28304 67826 28368
rect 67890 28304 67898 28368
rect 67578 27280 67898 28304
rect 67578 27216 67586 27280
rect 67650 27216 67666 27280
rect 67730 27216 67746 27280
rect 67810 27216 67826 27280
rect 67890 27216 67898 27280
rect 67578 26609 67898 27216
rect 70242 41968 70562 41984
rect 70242 41904 70250 41968
rect 70314 41904 70330 41968
rect 70394 41904 70410 41968
rect 70474 41904 70490 41968
rect 70554 41904 70562 41968
rect 70242 40880 70562 41904
rect 70242 40816 70250 40880
rect 70314 40816 70330 40880
rect 70394 40816 70410 40880
rect 70474 40816 70490 40880
rect 70554 40816 70562 40880
rect 70242 39792 70562 40816
rect 70242 39728 70250 39792
rect 70314 39728 70330 39792
rect 70394 39728 70410 39792
rect 70474 39728 70490 39792
rect 70554 39728 70562 39792
rect 70242 38704 70562 39728
rect 70242 38640 70250 38704
rect 70314 38640 70330 38704
rect 70394 38640 70410 38704
rect 70474 38640 70490 38704
rect 70554 38640 70562 38704
rect 70242 37616 70562 38640
rect 70242 37552 70250 37616
rect 70314 37552 70330 37616
rect 70394 37552 70410 37616
rect 70474 37552 70490 37616
rect 70554 37552 70562 37616
rect 70242 36528 70562 37552
rect 70242 36464 70250 36528
rect 70314 36464 70330 36528
rect 70394 36464 70410 36528
rect 70474 36464 70490 36528
rect 70554 36464 70562 36528
rect 70242 35440 70562 36464
rect 70242 35376 70250 35440
rect 70314 35376 70330 35440
rect 70394 35376 70410 35440
rect 70474 35376 70490 35440
rect 70554 35376 70562 35440
rect 70242 34352 70562 35376
rect 70242 34288 70250 34352
rect 70314 34288 70330 34352
rect 70394 34288 70410 34352
rect 70474 34288 70490 34352
rect 70554 34288 70562 34352
rect 70242 33264 70562 34288
rect 70242 33200 70250 33264
rect 70314 33200 70330 33264
rect 70394 33200 70410 33264
rect 70474 33200 70490 33264
rect 70554 33200 70562 33264
rect 70242 32176 70562 33200
rect 70242 32112 70250 32176
rect 70314 32112 70330 32176
rect 70394 32112 70410 32176
rect 70474 32112 70490 32176
rect 70554 32112 70562 32176
rect 70242 31088 70562 32112
rect 70242 31024 70250 31088
rect 70314 31024 70330 31088
rect 70394 31024 70410 31088
rect 70474 31024 70490 31088
rect 70554 31024 70562 31088
rect 70242 30000 70562 31024
rect 70242 29936 70250 30000
rect 70314 29936 70330 30000
rect 70394 29936 70410 30000
rect 70474 29936 70490 30000
rect 70554 29936 70562 30000
rect 70242 28912 70562 29936
rect 70242 28848 70250 28912
rect 70314 28848 70330 28912
rect 70394 28848 70410 28912
rect 70474 28848 70490 28912
rect 70554 28848 70562 28912
rect 70242 27824 70562 28848
rect 70242 27760 70250 27824
rect 70314 27760 70330 27824
rect 70394 27760 70410 27824
rect 70474 27760 70490 27824
rect 70554 27760 70562 27824
rect 70242 26736 70562 27760
rect 70242 26672 70250 26736
rect 70314 26672 70330 26736
rect 70394 26672 70410 26736
rect 70474 26672 70490 26736
rect 70554 26672 70562 26736
rect 70242 26609 70562 26672
rect 72906 41424 73226 41984
rect 72906 41360 72914 41424
rect 72978 41360 72994 41424
rect 73058 41360 73074 41424
rect 73138 41360 73154 41424
rect 73218 41360 73226 41424
rect 72906 40336 73226 41360
rect 72906 40272 72914 40336
rect 72978 40326 72994 40336
rect 73058 40326 73074 40336
rect 73138 40326 73154 40336
rect 73218 40272 73226 40336
rect 72906 40090 72948 40272
rect 73184 40090 73226 40272
rect 72906 40006 73226 40090
rect 72906 39770 72948 40006
rect 73184 39770 73226 40006
rect 72906 39248 73226 39770
rect 72906 39184 72914 39248
rect 72978 39184 72994 39248
rect 73058 39184 73074 39248
rect 73138 39184 73154 39248
rect 73218 39184 73226 39248
rect 72906 38160 73226 39184
rect 72906 38096 72914 38160
rect 72978 38096 72994 38160
rect 73058 38096 73074 38160
rect 73138 38096 73154 38160
rect 73218 38096 73226 38160
rect 72906 37072 73226 38096
rect 72906 37008 72914 37072
rect 72978 37008 72994 37072
rect 73058 37008 73074 37072
rect 73138 37008 73154 37072
rect 73218 37008 73226 37072
rect 72906 35984 73226 37008
rect 72906 35920 72914 35984
rect 72978 35920 72994 35984
rect 73058 35920 73074 35984
rect 73138 35920 73154 35984
rect 73218 35920 73226 35984
rect 72906 34896 73226 35920
rect 72906 34832 72914 34896
rect 72978 34832 72994 34896
rect 73058 34832 73074 34896
rect 73138 34832 73154 34896
rect 73218 34832 73226 34896
rect 72906 33808 73226 34832
rect 72906 33744 72914 33808
rect 72978 33744 72994 33808
rect 73058 33744 73074 33808
rect 73138 33744 73154 33808
rect 73218 33744 73226 33808
rect 72906 32720 73226 33744
rect 72906 32656 72914 32720
rect 72978 32656 72994 32720
rect 73058 32656 73074 32720
rect 73138 32656 73154 32720
rect 73218 32656 73226 32720
rect 72906 31632 73226 32656
rect 72906 31568 72914 31632
rect 72978 31568 72994 31632
rect 73058 31568 73074 31632
rect 73138 31568 73154 31632
rect 73218 31568 73226 31632
rect 72906 30544 73226 31568
rect 72906 30480 72914 30544
rect 72978 30480 72994 30544
rect 73058 30480 73074 30544
rect 73138 30480 73154 30544
rect 73218 30480 73226 30544
rect 72906 29456 73226 30480
rect 72906 29392 72914 29456
rect 72978 29392 72994 29456
rect 73058 29392 73074 29456
rect 73138 29392 73154 29456
rect 73218 29392 73226 29456
rect 72906 28368 73226 29392
rect 72906 28304 72914 28368
rect 72978 28304 72994 28368
rect 73058 28304 73074 28368
rect 73138 28304 73154 28368
rect 73218 28304 73226 28368
rect 72906 27280 73226 28304
rect 72906 27216 72914 27280
rect 72978 27216 72994 27280
rect 73058 27216 73074 27280
rect 73138 27216 73154 27280
rect 73218 27216 73226 27280
rect 72906 26609 73226 27216
rect 75570 41968 75890 41984
rect 75570 41904 75578 41968
rect 75642 41904 75658 41968
rect 75722 41904 75738 41968
rect 75802 41904 75818 41968
rect 75882 41904 75890 41968
rect 75570 40880 75890 41904
rect 75570 40816 75578 40880
rect 75642 40816 75658 40880
rect 75722 40816 75738 40880
rect 75802 40816 75818 40880
rect 75882 40816 75890 40880
rect 75570 39792 75890 40816
rect 75570 39728 75578 39792
rect 75642 39728 75658 39792
rect 75722 39728 75738 39792
rect 75802 39728 75818 39792
rect 75882 39728 75890 39792
rect 75570 38704 75890 39728
rect 75570 38640 75578 38704
rect 75642 38640 75658 38704
rect 75722 38640 75738 38704
rect 75802 38640 75818 38704
rect 75882 38640 75890 38704
rect 75570 37616 75890 38640
rect 75570 37552 75578 37616
rect 75642 37552 75658 37616
rect 75722 37552 75738 37616
rect 75802 37552 75818 37616
rect 75882 37552 75890 37616
rect 75570 36528 75890 37552
rect 75570 36464 75578 36528
rect 75642 36464 75658 36528
rect 75722 36464 75738 36528
rect 75802 36464 75818 36528
rect 75882 36464 75890 36528
rect 75570 35440 75890 36464
rect 75570 35376 75578 35440
rect 75642 35376 75658 35440
rect 75722 35376 75738 35440
rect 75802 35376 75818 35440
rect 75882 35376 75890 35440
rect 75570 34352 75890 35376
rect 75570 34288 75578 34352
rect 75642 34288 75658 34352
rect 75722 34288 75738 34352
rect 75802 34288 75818 34352
rect 75882 34288 75890 34352
rect 75570 33264 75890 34288
rect 75570 33200 75578 33264
rect 75642 33200 75658 33264
rect 75722 33200 75738 33264
rect 75802 33200 75818 33264
rect 75882 33200 75890 33264
rect 75570 32176 75890 33200
rect 75570 32112 75578 32176
rect 75642 32112 75658 32176
rect 75722 32112 75738 32176
rect 75802 32112 75818 32176
rect 75882 32112 75890 32176
rect 75570 31088 75890 32112
rect 75570 31024 75578 31088
rect 75642 31024 75658 31088
rect 75722 31024 75738 31088
rect 75802 31024 75818 31088
rect 75882 31024 75890 31088
rect 75570 30000 75890 31024
rect 75570 29936 75578 30000
rect 75642 29936 75658 30000
rect 75722 29936 75738 30000
rect 75802 29936 75818 30000
rect 75882 29936 75890 30000
rect 75570 28912 75890 29936
rect 75570 28848 75578 28912
rect 75642 28848 75658 28912
rect 75722 28848 75738 28912
rect 75802 28848 75818 28912
rect 75882 28848 75890 28912
rect 75570 27824 75890 28848
rect 75570 27760 75578 27824
rect 75642 27760 75658 27824
rect 75722 27760 75738 27824
rect 75802 27760 75818 27824
rect 75882 27760 75890 27824
rect 75570 26736 75890 27760
rect 75570 26672 75578 26736
rect 75642 26672 75658 26736
rect 75722 26672 75738 26736
rect 75802 26672 75818 26736
rect 75882 26672 75890 26736
rect 75570 26609 75890 26672
rect 78234 41424 78554 41984
rect 78234 41360 78242 41424
rect 78306 41360 78322 41424
rect 78386 41360 78402 41424
rect 78466 41360 78482 41424
rect 78546 41360 78554 41424
rect 78234 40336 78554 41360
rect 78234 40272 78242 40336
rect 78306 40326 78322 40336
rect 78386 40326 78402 40336
rect 78466 40326 78482 40336
rect 78546 40272 78554 40336
rect 78234 40090 78276 40272
rect 78512 40090 78554 40272
rect 78234 40006 78554 40090
rect 78234 39770 78276 40006
rect 78512 39770 78554 40006
rect 78234 39248 78554 39770
rect 78234 39184 78242 39248
rect 78306 39184 78322 39248
rect 78386 39184 78402 39248
rect 78466 39184 78482 39248
rect 78546 39184 78554 39248
rect 78234 38160 78554 39184
rect 78234 38096 78242 38160
rect 78306 38096 78322 38160
rect 78386 38096 78402 38160
rect 78466 38096 78482 38160
rect 78546 38096 78554 38160
rect 78234 37072 78554 38096
rect 78234 37008 78242 37072
rect 78306 37008 78322 37072
rect 78386 37008 78402 37072
rect 78466 37008 78482 37072
rect 78546 37008 78554 37072
rect 78234 35984 78554 37008
rect 78234 35920 78242 35984
rect 78306 35920 78322 35984
rect 78386 35920 78402 35984
rect 78466 35920 78482 35984
rect 78546 35920 78554 35984
rect 78234 34896 78554 35920
rect 78234 34832 78242 34896
rect 78306 34832 78322 34896
rect 78386 34832 78402 34896
rect 78466 34832 78482 34896
rect 78546 34832 78554 34896
rect 78234 33808 78554 34832
rect 78234 33744 78242 33808
rect 78306 33744 78322 33808
rect 78386 33744 78402 33808
rect 78466 33744 78482 33808
rect 78546 33744 78554 33808
rect 78234 32720 78554 33744
rect 78234 32656 78242 32720
rect 78306 32656 78322 32720
rect 78386 32656 78402 32720
rect 78466 32656 78482 32720
rect 78546 32656 78554 32720
rect 78234 31632 78554 32656
rect 78234 31568 78242 31632
rect 78306 31568 78322 31632
rect 78386 31568 78402 31632
rect 78466 31568 78482 31632
rect 78546 31568 78554 31632
rect 78234 30544 78554 31568
rect 78234 30480 78242 30544
rect 78306 30480 78322 30544
rect 78386 30480 78402 30544
rect 78466 30480 78482 30544
rect 78546 30480 78554 30544
rect 78234 29456 78554 30480
rect 78234 29392 78242 29456
rect 78306 29392 78322 29456
rect 78386 29392 78402 29456
rect 78466 29392 78482 29456
rect 78546 29392 78554 29456
rect 78234 28368 78554 29392
rect 78234 28304 78242 28368
rect 78306 28304 78322 28368
rect 78386 28304 78402 28368
rect 78466 28304 78482 28368
rect 78546 28304 78554 28368
rect 78234 27280 78554 28304
rect 78234 27216 78242 27280
rect 78306 27216 78322 27280
rect 78386 27216 78402 27280
rect 78466 27216 78482 27280
rect 78546 27216 78554 27280
rect 78234 26609 78554 27216
rect 80898 41968 81218 41984
rect 80898 41904 80906 41968
rect 80970 41904 80986 41968
rect 81050 41904 81066 41968
rect 81130 41904 81146 41968
rect 81210 41904 81218 41968
rect 80898 40880 81218 41904
rect 80898 40816 80906 40880
rect 80970 40816 80986 40880
rect 81050 40816 81066 40880
rect 81130 40816 81146 40880
rect 81210 40816 81218 40880
rect 80898 39792 81218 40816
rect 80898 39728 80906 39792
rect 80970 39728 80986 39792
rect 81050 39728 81066 39792
rect 81130 39728 81146 39792
rect 81210 39728 81218 39792
rect 80898 38704 81218 39728
rect 80898 38640 80906 38704
rect 80970 38640 80986 38704
rect 81050 38640 81066 38704
rect 81130 38640 81146 38704
rect 81210 38640 81218 38704
rect 80898 37616 81218 38640
rect 80898 37552 80906 37616
rect 80970 37552 80986 37616
rect 81050 37552 81066 37616
rect 81130 37552 81146 37616
rect 81210 37552 81218 37616
rect 80898 36528 81218 37552
rect 80898 36464 80906 36528
rect 80970 36464 80986 36528
rect 81050 36464 81066 36528
rect 81130 36464 81146 36528
rect 81210 36464 81218 36528
rect 80898 35440 81218 36464
rect 80898 35376 80906 35440
rect 80970 35376 80986 35440
rect 81050 35376 81066 35440
rect 81130 35376 81146 35440
rect 81210 35376 81218 35440
rect 80898 34352 81218 35376
rect 80898 34288 80906 34352
rect 80970 34288 80986 34352
rect 81050 34288 81066 34352
rect 81130 34288 81146 34352
rect 81210 34288 81218 34352
rect 80898 33264 81218 34288
rect 80898 33200 80906 33264
rect 80970 33200 80986 33264
rect 81050 33200 81066 33264
rect 81130 33200 81146 33264
rect 81210 33200 81218 33264
rect 80898 32176 81218 33200
rect 80898 32112 80906 32176
rect 80970 32112 80986 32176
rect 81050 32112 81066 32176
rect 81130 32112 81146 32176
rect 81210 32112 81218 32176
rect 80898 31088 81218 32112
rect 80898 31024 80906 31088
rect 80970 31024 80986 31088
rect 81050 31024 81066 31088
rect 81130 31024 81146 31088
rect 81210 31024 81218 31088
rect 80898 30000 81218 31024
rect 80898 29936 80906 30000
rect 80970 29936 80986 30000
rect 81050 29936 81066 30000
rect 81130 29936 81146 30000
rect 81210 29936 81218 30000
rect 80898 28912 81218 29936
rect 80898 28848 80906 28912
rect 80970 28848 80986 28912
rect 81050 28848 81066 28912
rect 81130 28848 81146 28912
rect 81210 28848 81218 28912
rect 80898 27824 81218 28848
rect 80898 27760 80906 27824
rect 80970 27760 80986 27824
rect 81050 27760 81066 27824
rect 81130 27760 81146 27824
rect 81210 27760 81218 27824
rect 80898 26736 81218 27760
rect 80898 26672 80906 26736
rect 80970 26672 80986 26736
rect 81050 26672 81066 26736
rect 81130 26672 81146 26736
rect 81210 26672 81218 26736
rect 80898 26609 81218 26672
rect 83562 41424 83882 41984
rect 83562 41360 83570 41424
rect 83634 41360 83650 41424
rect 83714 41360 83730 41424
rect 83794 41360 83810 41424
rect 83874 41360 83882 41424
rect 83562 40336 83882 41360
rect 83562 40272 83570 40336
rect 83634 40326 83650 40336
rect 83714 40326 83730 40336
rect 83794 40326 83810 40336
rect 83874 40272 83882 40336
rect 83562 40090 83604 40272
rect 83840 40090 83882 40272
rect 83562 40006 83882 40090
rect 83562 39770 83604 40006
rect 83840 39770 83882 40006
rect 83562 39248 83882 39770
rect 83562 39184 83570 39248
rect 83634 39184 83650 39248
rect 83714 39184 83730 39248
rect 83794 39184 83810 39248
rect 83874 39184 83882 39248
rect 83562 38160 83882 39184
rect 83562 38096 83570 38160
rect 83634 38096 83650 38160
rect 83714 38096 83730 38160
rect 83794 38096 83810 38160
rect 83874 38096 83882 38160
rect 83562 37072 83882 38096
rect 83562 37008 83570 37072
rect 83634 37008 83650 37072
rect 83714 37008 83730 37072
rect 83794 37008 83810 37072
rect 83874 37008 83882 37072
rect 83562 35984 83882 37008
rect 83562 35920 83570 35984
rect 83634 35920 83650 35984
rect 83714 35920 83730 35984
rect 83794 35920 83810 35984
rect 83874 35920 83882 35984
rect 83562 34896 83882 35920
rect 83562 34832 83570 34896
rect 83634 34832 83650 34896
rect 83714 34832 83730 34896
rect 83794 34832 83810 34896
rect 83874 34832 83882 34896
rect 83562 33808 83882 34832
rect 83562 33744 83570 33808
rect 83634 33744 83650 33808
rect 83714 33744 83730 33808
rect 83794 33744 83810 33808
rect 83874 33744 83882 33808
rect 83562 32720 83882 33744
rect 83562 32656 83570 32720
rect 83634 32656 83650 32720
rect 83714 32656 83730 32720
rect 83794 32656 83810 32720
rect 83874 32656 83882 32720
rect 83562 31632 83882 32656
rect 83562 31568 83570 31632
rect 83634 31568 83650 31632
rect 83714 31568 83730 31632
rect 83794 31568 83810 31632
rect 83874 31568 83882 31632
rect 83562 30544 83882 31568
rect 83562 30480 83570 30544
rect 83634 30480 83650 30544
rect 83714 30480 83730 30544
rect 83794 30480 83810 30544
rect 83874 30480 83882 30544
rect 83562 29456 83882 30480
rect 83562 29392 83570 29456
rect 83634 29392 83650 29456
rect 83714 29392 83730 29456
rect 83794 29392 83810 29456
rect 83874 29392 83882 29456
rect 83562 28368 83882 29392
rect 83562 28304 83570 28368
rect 83634 28304 83650 28368
rect 83714 28304 83730 28368
rect 83794 28304 83810 28368
rect 83874 28304 83882 28368
rect 83562 27280 83882 28304
rect 83562 27216 83570 27280
rect 83634 27216 83650 27280
rect 83714 27216 83730 27280
rect 83794 27216 83810 27280
rect 83874 27216 83882 27280
rect 83562 26609 83882 27216
rect 86226 41968 86546 41984
rect 86226 41904 86234 41968
rect 86298 41904 86314 41968
rect 86378 41904 86394 41968
rect 86458 41904 86474 41968
rect 86538 41904 86546 41968
rect 86226 40880 86546 41904
rect 86226 40816 86234 40880
rect 86298 40816 86314 40880
rect 86378 40816 86394 40880
rect 86458 40816 86474 40880
rect 86538 40816 86546 40880
rect 86226 39792 86546 40816
rect 86226 39728 86234 39792
rect 86298 39728 86314 39792
rect 86378 39728 86394 39792
rect 86458 39728 86474 39792
rect 86538 39728 86546 39792
rect 86226 38704 86546 39728
rect 86226 38640 86234 38704
rect 86298 38640 86314 38704
rect 86378 38640 86394 38704
rect 86458 38640 86474 38704
rect 86538 38640 86546 38704
rect 86226 37616 86546 38640
rect 86226 37552 86234 37616
rect 86298 37552 86314 37616
rect 86378 37552 86394 37616
rect 86458 37552 86474 37616
rect 86538 37552 86546 37616
rect 86226 36528 86546 37552
rect 86226 36464 86234 36528
rect 86298 36464 86314 36528
rect 86378 36464 86394 36528
rect 86458 36464 86474 36528
rect 86538 36464 86546 36528
rect 86226 35440 86546 36464
rect 86226 35376 86234 35440
rect 86298 35376 86314 35440
rect 86378 35376 86394 35440
rect 86458 35376 86474 35440
rect 86538 35376 86546 35440
rect 86226 34352 86546 35376
rect 86226 34288 86234 34352
rect 86298 34288 86314 34352
rect 86378 34288 86394 34352
rect 86458 34288 86474 34352
rect 86538 34288 86546 34352
rect 86226 33264 86546 34288
rect 86226 33200 86234 33264
rect 86298 33200 86314 33264
rect 86378 33200 86394 33264
rect 86458 33200 86474 33264
rect 86538 33200 86546 33264
rect 86226 32176 86546 33200
rect 86226 32112 86234 32176
rect 86298 32112 86314 32176
rect 86378 32112 86394 32176
rect 86458 32112 86474 32176
rect 86538 32112 86546 32176
rect 86226 31088 86546 32112
rect 86226 31024 86234 31088
rect 86298 31024 86314 31088
rect 86378 31024 86394 31088
rect 86458 31024 86474 31088
rect 86538 31024 86546 31088
rect 86226 30000 86546 31024
rect 86226 29936 86234 30000
rect 86298 29936 86314 30000
rect 86378 29936 86394 30000
rect 86458 29936 86474 30000
rect 86538 29936 86546 30000
rect 86226 28912 86546 29936
rect 86226 28848 86234 28912
rect 86298 28848 86314 28912
rect 86378 28848 86394 28912
rect 86458 28848 86474 28912
rect 86538 28848 86546 28912
rect 86226 27824 86546 28848
rect 86226 27760 86234 27824
rect 86298 27760 86314 27824
rect 86378 27760 86394 27824
rect 86458 27760 86474 27824
rect 86538 27760 86546 27824
rect 86226 26736 86546 27760
rect 86226 26672 86234 26736
rect 86298 26672 86314 26736
rect 86378 26672 86394 26736
rect 86458 26672 86474 26736
rect 86538 26672 86546 26736
rect 86226 26609 86546 26672
rect 88890 41424 89210 41984
rect 88890 41360 88898 41424
rect 88962 41360 88978 41424
rect 89042 41360 89058 41424
rect 89122 41360 89138 41424
rect 89202 41360 89210 41424
rect 88890 40336 89210 41360
rect 88890 40272 88898 40336
rect 88962 40326 88978 40336
rect 89042 40326 89058 40336
rect 89122 40326 89138 40336
rect 89202 40272 89210 40336
rect 88890 40090 88932 40272
rect 89168 40090 89210 40272
rect 88890 40006 89210 40090
rect 88890 39770 88932 40006
rect 89168 39770 89210 40006
rect 88890 39248 89210 39770
rect 88890 39184 88898 39248
rect 88962 39184 88978 39248
rect 89042 39184 89058 39248
rect 89122 39184 89138 39248
rect 89202 39184 89210 39248
rect 88890 38160 89210 39184
rect 88890 38096 88898 38160
rect 88962 38096 88978 38160
rect 89042 38096 89058 38160
rect 89122 38096 89138 38160
rect 89202 38096 89210 38160
rect 88890 37072 89210 38096
rect 88890 37008 88898 37072
rect 88962 37008 88978 37072
rect 89042 37008 89058 37072
rect 89122 37008 89138 37072
rect 89202 37008 89210 37072
rect 88890 35984 89210 37008
rect 88890 35920 88898 35984
rect 88962 35920 88978 35984
rect 89042 35920 89058 35984
rect 89122 35920 89138 35984
rect 89202 35920 89210 35984
rect 88890 34896 89210 35920
rect 88890 34832 88898 34896
rect 88962 34832 88978 34896
rect 89042 34832 89058 34896
rect 89122 34832 89138 34896
rect 89202 34832 89210 34896
rect 88890 33808 89210 34832
rect 88890 33744 88898 33808
rect 88962 33744 88978 33808
rect 89042 33744 89058 33808
rect 89122 33744 89138 33808
rect 89202 33744 89210 33808
rect 88890 32720 89210 33744
rect 88890 32656 88898 32720
rect 88962 32656 88978 32720
rect 89042 32656 89058 32720
rect 89122 32656 89138 32720
rect 89202 32656 89210 32720
rect 88890 31632 89210 32656
rect 88890 31568 88898 31632
rect 88962 31568 88978 31632
rect 89042 31568 89058 31632
rect 89122 31568 89138 31632
rect 89202 31568 89210 31632
rect 88890 30544 89210 31568
rect 88890 30480 88898 30544
rect 88962 30480 88978 30544
rect 89042 30480 89058 30544
rect 89122 30480 89138 30544
rect 89202 30480 89210 30544
rect 88890 29456 89210 30480
rect 88890 29392 88898 29456
rect 88962 29392 88978 29456
rect 89042 29392 89058 29456
rect 89122 29392 89138 29456
rect 89202 29392 89210 29456
rect 88890 28368 89210 29392
rect 88890 28304 88898 28368
rect 88962 28304 88978 28368
rect 89042 28304 89058 28368
rect 89122 28304 89138 28368
rect 89202 28304 89210 28368
rect 88890 27280 89210 28304
rect 88890 27216 88898 27280
rect 88962 27216 88978 27280
rect 89042 27216 89058 27280
rect 89122 27216 89138 27280
rect 89202 27216 89210 27280
rect 88890 26609 89210 27216
rect 91554 41968 91874 41984
rect 91554 41904 91562 41968
rect 91626 41904 91642 41968
rect 91706 41904 91722 41968
rect 91786 41904 91802 41968
rect 91866 41904 91874 41968
rect 91554 40880 91874 41904
rect 91554 40816 91562 40880
rect 91626 40816 91642 40880
rect 91706 40816 91722 40880
rect 91786 40816 91802 40880
rect 91866 40816 91874 40880
rect 91554 39792 91874 40816
rect 91554 39728 91562 39792
rect 91626 39728 91642 39792
rect 91706 39728 91722 39792
rect 91786 39728 91802 39792
rect 91866 39728 91874 39792
rect 91554 38704 91874 39728
rect 91554 38640 91562 38704
rect 91626 38640 91642 38704
rect 91706 38640 91722 38704
rect 91786 38640 91802 38704
rect 91866 38640 91874 38704
rect 91554 37616 91874 38640
rect 91554 37552 91562 37616
rect 91626 37552 91642 37616
rect 91706 37552 91722 37616
rect 91786 37552 91802 37616
rect 91866 37552 91874 37616
rect 91554 36528 91874 37552
rect 91554 36464 91562 36528
rect 91626 36464 91642 36528
rect 91706 36464 91722 36528
rect 91786 36464 91802 36528
rect 91866 36464 91874 36528
rect 91554 35440 91874 36464
rect 91554 35376 91562 35440
rect 91626 35376 91642 35440
rect 91706 35376 91722 35440
rect 91786 35376 91802 35440
rect 91866 35376 91874 35440
rect 91554 34352 91874 35376
rect 91554 34288 91562 34352
rect 91626 34288 91642 34352
rect 91706 34288 91722 34352
rect 91786 34288 91802 34352
rect 91866 34288 91874 34352
rect 91554 33264 91874 34288
rect 91554 33200 91562 33264
rect 91626 33200 91642 33264
rect 91706 33200 91722 33264
rect 91786 33200 91802 33264
rect 91866 33200 91874 33264
rect 91554 32176 91874 33200
rect 91554 32112 91562 32176
rect 91626 32112 91642 32176
rect 91706 32112 91722 32176
rect 91786 32112 91802 32176
rect 91866 32112 91874 32176
rect 91554 31088 91874 32112
rect 91554 31024 91562 31088
rect 91626 31024 91642 31088
rect 91706 31024 91722 31088
rect 91786 31024 91802 31088
rect 91866 31024 91874 31088
rect 91554 30000 91874 31024
rect 91554 29936 91562 30000
rect 91626 29936 91642 30000
rect 91706 29936 91722 30000
rect 91786 29936 91802 30000
rect 91866 29936 91874 30000
rect 91554 28912 91874 29936
rect 91554 28848 91562 28912
rect 91626 28848 91642 28912
rect 91706 28848 91722 28912
rect 91786 28848 91802 28912
rect 91866 28848 91874 28912
rect 91554 27824 91874 28848
rect 91554 27760 91562 27824
rect 91626 27760 91642 27824
rect 91706 27760 91722 27824
rect 91786 27760 91802 27824
rect 91866 27760 91874 27824
rect 91554 26736 91874 27760
rect 91554 26672 91562 26736
rect 91626 26672 91642 26736
rect 91706 26672 91722 26736
rect 91786 26672 91802 26736
rect 91866 26672 91874 26736
rect 91554 26609 91874 26672
rect 40938 26128 40946 26192
rect 41010 26128 41026 26192
rect 41090 26128 41106 26192
rect 41170 26128 41186 26192
rect 41250 26128 41258 26192
rect 40938 25104 41258 26128
rect 40938 25040 40946 25104
rect 41010 25040 41026 25104
rect 41090 25040 41106 25104
rect 41170 25040 41186 25104
rect 41250 25040 41258 25104
rect 40938 24016 41258 25040
rect 40938 23952 40946 24016
rect 41010 23952 41026 24016
rect 41090 23952 41106 24016
rect 41170 23952 41186 24016
rect 41250 23952 41258 24016
rect 40938 22928 41258 23952
rect 40938 22864 40946 22928
rect 41010 22864 41026 22928
rect 41090 22864 41106 22928
rect 41170 22864 41186 22928
rect 41250 22864 41258 22928
rect 40938 21840 41258 22864
rect 40938 21776 40946 21840
rect 41010 21776 41026 21840
rect 41090 21776 41106 21840
rect 41170 21776 41186 21840
rect 41250 21776 41258 21840
rect 40938 20752 41258 21776
rect 40938 20688 40946 20752
rect 41010 20688 41026 20752
rect 41090 20688 41106 20752
rect 41170 20688 41186 20752
rect 41250 20688 41258 20752
rect 40938 19664 41258 20688
rect 40938 19600 40946 19664
rect 41010 19600 41026 19664
rect 41090 19600 41106 19664
rect 41170 19600 41186 19664
rect 41250 19600 41258 19664
rect 40938 18576 41258 19600
rect 40938 18512 40946 18576
rect 41010 18512 41026 18576
rect 41090 18512 41106 18576
rect 41170 18512 41186 18576
rect 41250 18512 41258 18576
rect 40938 17488 41258 18512
rect 40938 17424 40946 17488
rect 41010 17424 41026 17488
rect 41090 17424 41106 17488
rect 41170 17424 41186 17488
rect 41250 17424 41258 17488
rect 40938 16400 41258 17424
rect 40938 16336 40946 16400
rect 41010 16336 41026 16400
rect 41090 16336 41106 16400
rect 41170 16336 41186 16400
rect 41250 16336 41258 16400
rect 40938 15312 41258 16336
rect 40938 15248 40946 15312
rect 41010 15248 41026 15312
rect 41090 15248 41106 15312
rect 41170 15248 41186 15312
rect 41250 15248 41258 15312
rect 40938 14224 41258 15248
rect 40938 14160 40946 14224
rect 41010 14160 41026 14224
rect 41090 14160 41106 14224
rect 41170 14160 41186 14224
rect 41250 14160 41258 14224
rect 40938 13136 41258 14160
rect 40938 13072 40946 13136
rect 41010 13072 41026 13136
rect 41090 13072 41106 13136
rect 41170 13072 41186 13136
rect 41250 13072 41258 13136
rect 40938 12048 41258 13072
rect 40938 11984 40946 12048
rect 41010 11984 41026 12048
rect 41090 11984 41106 12048
rect 41170 11984 41186 12048
rect 41250 11984 41258 12048
rect 40938 10960 41258 11984
rect 40938 10896 40946 10960
rect 41010 10896 41026 10960
rect 41090 10896 41106 10960
rect 41170 10896 41186 10960
rect 41250 10896 41258 10960
rect 40938 9872 41258 10896
rect 40938 9808 40946 9872
rect 41010 9808 41026 9872
rect 41090 9808 41106 9872
rect 41170 9808 41186 9872
rect 41250 9808 41258 9872
rect 40938 8784 41258 9808
rect 40938 8720 40946 8784
rect 41010 8720 41026 8784
rect 41090 8720 41106 8784
rect 41170 8720 41186 8784
rect 41250 8720 41258 8784
rect 40938 7696 41258 8720
rect 40938 7632 40946 7696
rect 41010 7632 41026 7696
rect 41090 7632 41106 7696
rect 41170 7632 41186 7696
rect 41250 7632 41258 7696
rect 40938 6608 41258 7632
rect 40938 6544 40946 6608
rect 41010 6544 41026 6608
rect 41090 6544 41106 6608
rect 41170 6544 41186 6608
rect 41250 6544 41258 6608
rect 40938 5520 41258 6544
rect 40938 5456 40946 5520
rect 41010 5456 41026 5520
rect 41090 5456 41106 5520
rect 41170 5456 41186 5520
rect 41250 5456 41258 5520
rect 40938 4432 41258 5456
rect 40938 4368 40946 4432
rect 41010 4368 41026 4432
rect 41090 4368 41106 4432
rect 41170 4368 41186 4432
rect 41250 4368 41258 4432
rect 40938 4326 41258 4368
rect 40938 4090 40980 4326
rect 41216 4090 41258 4326
rect 40938 4006 41258 4090
rect 40938 3770 40980 4006
rect 41216 3770 41258 4006
rect 40938 3344 41258 3770
rect 40938 3280 40946 3344
rect 41010 3280 41026 3344
rect 41090 3280 41106 3344
rect 41170 3280 41186 3344
rect 41250 3280 41258 3344
rect 40938 2256 41258 3280
rect 40938 2192 40946 2256
rect 41010 2192 41026 2256
rect 41090 2192 41106 2256
rect 41170 2192 41186 2256
rect 41250 2192 41258 2256
rect 40938 1168 41258 2192
rect 40938 1104 40946 1168
rect 41010 1104 41026 1168
rect 41090 1104 41106 1168
rect 41170 1104 41186 1168
rect 41250 1104 41258 1168
rect 40938 80 41258 1104
rect 40938 16 40946 80
rect 41010 16 41026 80
rect 41090 16 41106 80
rect 41170 16 41186 80
rect 41250 16 41258 80
rect 40938 0 41258 16
<< via4 >>
rect 3684 40272 3714 40326
rect 3714 40272 3730 40326
rect 3730 40272 3794 40326
rect 3794 40272 3810 40326
rect 3810 40272 3874 40326
rect 3874 40272 3890 40326
rect 3890 40272 3920 40326
rect 3684 40090 3920 40272
rect 3684 39770 3920 40006
rect 3272 20534 3508 20770
rect 9012 40272 9042 40326
rect 9042 40272 9058 40326
rect 9058 40272 9122 40326
rect 9122 40272 9138 40326
rect 9138 40272 9202 40326
rect 9202 40272 9218 40326
rect 9218 40272 9248 40326
rect 9012 40090 9248 40272
rect 9012 39770 9248 40006
rect 14340 40272 14370 40326
rect 14370 40272 14386 40326
rect 14386 40272 14450 40326
rect 14450 40272 14466 40326
rect 14466 40272 14530 40326
rect 14530 40272 14546 40326
rect 14546 40272 14576 40326
rect 14340 40090 14576 40272
rect 14340 39770 14576 40006
rect 19668 40272 19698 40326
rect 19698 40272 19714 40326
rect 19714 40272 19778 40326
rect 19778 40272 19794 40326
rect 19794 40272 19858 40326
rect 19858 40272 19874 40326
rect 19874 40272 19904 40326
rect 19668 40090 19904 40272
rect 19668 39770 19904 40006
rect 24996 40272 25026 40326
rect 25026 40272 25042 40326
rect 25042 40272 25106 40326
rect 25106 40272 25122 40326
rect 25122 40272 25186 40326
rect 25186 40272 25202 40326
rect 25202 40272 25232 40326
rect 24996 40090 25232 40272
rect 24996 39770 25232 40006
rect 30324 40272 30354 40326
rect 30354 40272 30370 40326
rect 30370 40272 30434 40326
rect 30434 40272 30450 40326
rect 30450 40272 30514 40326
rect 30514 40272 30530 40326
rect 30530 40272 30560 40326
rect 30324 40090 30560 40272
rect 30324 39770 30560 40006
rect 35652 40272 35682 40326
rect 35682 40272 35698 40326
rect 35698 40272 35762 40326
rect 35762 40272 35778 40326
rect 35778 40272 35842 40326
rect 35842 40272 35858 40326
rect 35858 40272 35888 40326
rect 35652 40090 35888 40272
rect 35652 39770 35888 40006
rect 6348 22320 6378 22326
rect 6378 22320 6394 22326
rect 6394 22320 6458 22326
rect 6458 22320 6474 22326
rect 6474 22320 6538 22326
rect 6538 22320 6554 22326
rect 6554 22320 6584 22326
rect 6348 22090 6584 22320
rect 6348 21770 6584 22006
rect 31424 20534 31660 20770
rect 38316 22320 38346 22326
rect 38346 22320 38362 22326
rect 38362 22320 38426 22326
rect 38426 22320 38442 22326
rect 38442 22320 38506 22326
rect 38506 22320 38522 22326
rect 38522 22320 38552 22326
rect 38316 22090 38552 22320
rect 38316 21770 38552 22006
rect 4192 19324 4428 19410
rect 4192 19260 4278 19324
rect 4278 19260 4342 19324
rect 4342 19260 4428 19324
rect 4192 19174 4428 19260
rect 6768 20004 7004 20090
rect 6768 19940 6854 20004
rect 6854 19940 6918 20004
rect 6918 19940 7004 20004
rect 6768 19854 7004 19940
rect 13576 19854 13812 20090
rect 27928 19854 28164 20090
rect 31424 19854 31660 20090
rect 5112 17284 5348 17370
rect 5112 17220 5198 17284
rect 5198 17220 5262 17284
rect 5262 17220 5348 17284
rect 5112 17134 5348 17220
rect 5664 16604 5900 16690
rect 5664 16540 5750 16604
rect 5750 16540 5814 16604
rect 5814 16540 5900 16604
rect 5664 16454 5900 16540
rect 3684 4090 3920 4326
rect 3684 3770 3920 4006
rect 37864 20534 38100 20770
rect 31424 19188 31660 19410
rect 31424 19174 31510 19188
rect 31510 19174 31574 19188
rect 31574 19174 31660 19188
rect 31424 18036 31510 18050
rect 31510 18036 31574 18050
rect 31574 18036 31660 18050
rect 31424 17814 31660 18036
rect 13576 17134 13812 17370
rect 27928 17134 28164 17370
rect 36208 16604 36444 16690
rect 36208 16540 36294 16604
rect 36294 16540 36358 16604
rect 36358 16540 36444 16604
rect 36208 16454 36444 16540
rect 7320 15774 7556 16010
rect 31424 15774 31660 16010
rect 7136 15244 7372 15330
rect 7136 15180 7222 15244
rect 7222 15180 7286 15244
rect 7286 15180 7372 15244
rect 7136 15094 7372 15180
rect 31424 15094 31660 15330
rect 7320 11014 7556 11250
rect 31424 11014 31660 11250
rect 35652 4090 35888 4326
rect 35652 3770 35888 4006
rect 40980 40272 41010 40326
rect 41010 40272 41026 40326
rect 41026 40272 41090 40326
rect 41090 40272 41106 40326
rect 41106 40272 41170 40326
rect 41170 40272 41186 40326
rect 41186 40272 41216 40326
rect 40980 40090 41216 40272
rect 40980 39770 41216 40006
rect 46308 40272 46338 40326
rect 46338 40272 46354 40326
rect 46354 40272 46418 40326
rect 46418 40272 46434 40326
rect 46434 40272 46498 40326
rect 46498 40272 46514 40326
rect 46514 40272 46544 40326
rect 46308 40090 46544 40272
rect 46308 39770 46544 40006
rect 51636 40272 51666 40326
rect 51666 40272 51682 40326
rect 51682 40272 51746 40326
rect 51746 40272 51762 40326
rect 51762 40272 51826 40326
rect 51826 40272 51842 40326
rect 51842 40272 51872 40326
rect 51636 40090 51872 40272
rect 51636 39770 51872 40006
rect 56964 40272 56994 40326
rect 56994 40272 57010 40326
rect 57010 40272 57074 40326
rect 57074 40272 57090 40326
rect 57090 40272 57154 40326
rect 57154 40272 57170 40326
rect 57170 40272 57200 40326
rect 56964 40090 57200 40272
rect 56964 39770 57200 40006
rect 62292 40272 62322 40326
rect 62322 40272 62338 40326
rect 62338 40272 62402 40326
rect 62402 40272 62418 40326
rect 62418 40272 62482 40326
rect 62482 40272 62498 40326
rect 62498 40272 62528 40326
rect 62292 40090 62528 40272
rect 62292 39770 62528 40006
rect 67620 40272 67650 40326
rect 67650 40272 67666 40326
rect 67666 40272 67730 40326
rect 67730 40272 67746 40326
rect 67746 40272 67810 40326
rect 67810 40272 67826 40326
rect 67826 40272 67856 40326
rect 67620 40090 67856 40272
rect 67620 39770 67856 40006
rect 72948 40272 72978 40326
rect 72978 40272 72994 40326
rect 72994 40272 73058 40326
rect 73058 40272 73074 40326
rect 73074 40272 73138 40326
rect 73138 40272 73154 40326
rect 73154 40272 73184 40326
rect 72948 40090 73184 40272
rect 72948 39770 73184 40006
rect 78276 40272 78306 40326
rect 78306 40272 78322 40326
rect 78322 40272 78386 40326
rect 78386 40272 78402 40326
rect 78402 40272 78466 40326
rect 78466 40272 78482 40326
rect 78482 40272 78512 40326
rect 78276 40090 78512 40272
rect 78276 39770 78512 40006
rect 83604 40272 83634 40326
rect 83634 40272 83650 40326
rect 83650 40272 83714 40326
rect 83714 40272 83730 40326
rect 83730 40272 83794 40326
rect 83794 40272 83810 40326
rect 83810 40272 83840 40326
rect 83604 40090 83840 40272
rect 83604 39770 83840 40006
rect 88932 40272 88962 40326
rect 88962 40272 88978 40326
rect 88978 40272 89042 40326
rect 89042 40272 89058 40326
rect 89058 40272 89122 40326
rect 89122 40272 89138 40326
rect 89138 40272 89168 40326
rect 88932 40090 89168 40272
rect 88932 39770 89168 40006
rect 66752 20684 66988 20770
rect 66752 20620 66838 20684
rect 66838 20620 66902 20684
rect 66902 20620 66988 20684
rect 66752 20534 66988 20620
rect 41544 20004 41780 20090
rect 41544 19940 41630 20004
rect 41630 19940 41694 20004
rect 41694 19940 41780 20004
rect 41544 19854 41780 19940
rect 66936 20004 67172 20090
rect 66936 19940 67022 20004
rect 67022 19940 67086 20004
rect 67086 19940 67172 20004
rect 66936 19854 67172 19940
rect 41912 17964 42148 18050
rect 41912 17900 41998 17964
rect 41998 17900 42062 17964
rect 42062 17900 42148 17964
rect 41912 17814 42148 17900
rect 67672 17964 67908 18050
rect 67672 17900 67758 17964
rect 67758 17900 67822 17964
rect 67822 17900 67908 17964
rect 67672 17814 67908 17900
rect 41728 16604 41964 16690
rect 41728 16540 41814 16604
rect 41814 16540 41878 16604
rect 41878 16540 41964 16604
rect 41728 16454 41964 16540
rect 68224 16604 68460 16690
rect 68224 16540 68310 16604
rect 68310 16540 68374 16604
rect 68374 16540 68460 16604
rect 68224 16454 68460 16540
rect 40980 4090 41216 4326
rect 40980 3770 41216 4006
<< metal5 >>
rect 3642 40348 3962 40350
rect 8970 40348 9290 40350
rect 14298 40348 14618 40350
rect 19626 40348 19946 40350
rect 24954 40348 25274 40350
rect 30282 40348 30602 40350
rect 35610 40348 35930 40350
rect 40938 40348 41258 40350
rect 46266 40348 46586 40350
rect 51594 40348 51914 40350
rect 56922 40348 57242 40350
rect 62250 40348 62570 40350
rect 67578 40348 67898 40350
rect 72906 40348 73226 40350
rect 78234 40348 78554 40350
rect 83562 40348 83882 40350
rect 88890 40348 89210 40350
rect 538 40326 93642 40348
rect 538 40090 3684 40326
rect 3920 40090 9012 40326
rect 9248 40090 14340 40326
rect 14576 40090 19668 40326
rect 19904 40090 24996 40326
rect 25232 40090 30324 40326
rect 30560 40090 35652 40326
rect 35888 40090 40980 40326
rect 41216 40090 46308 40326
rect 46544 40090 51636 40326
rect 51872 40090 56964 40326
rect 57200 40090 62292 40326
rect 62528 40090 67620 40326
rect 67856 40090 72948 40326
rect 73184 40090 78276 40326
rect 78512 40090 83604 40326
rect 83840 40090 88932 40326
rect 89168 40090 93642 40326
rect 538 40006 93642 40090
rect 538 39770 3684 40006
rect 3920 39770 9012 40006
rect 9248 39770 14340 40006
rect 14576 39770 19668 40006
rect 19904 39770 24996 40006
rect 25232 39770 30324 40006
rect 30560 39770 35652 40006
rect 35888 39770 40980 40006
rect 41216 39770 46308 40006
rect 46544 39770 51636 40006
rect 51872 39770 56964 40006
rect 57200 39770 62292 40006
rect 62528 39770 67620 40006
rect 67856 39770 72948 40006
rect 73184 39770 78276 40006
rect 78512 39770 83604 40006
rect 83840 39770 88932 40006
rect 89168 39770 93642 40006
rect 538 39748 93642 39770
rect 3642 39746 3962 39748
rect 8970 39746 9290 39748
rect 14298 39746 14618 39748
rect 19626 39746 19946 39748
rect 24954 39746 25274 39748
rect 30282 39746 30602 39748
rect 35610 39746 35930 39748
rect 40938 39746 41258 39748
rect 46266 39746 46586 39748
rect 51594 39746 51914 39748
rect 56922 39746 57242 39748
rect 62250 39746 62570 39748
rect 67578 39746 67898 39748
rect 72906 39746 73226 39748
rect 78234 39746 78554 39748
rect 83562 39746 83882 39748
rect 88890 39746 89210 39748
rect 6306 22348 6626 22350
rect 38274 22348 38594 22350
rect 538 22326 93642 22348
rect 538 22090 6348 22326
rect 6584 22090 38316 22326
rect 38552 22090 93642 22326
rect 538 22006 93642 22090
rect 538 21770 6348 22006
rect 6584 21770 38316 22006
rect 38552 21770 93642 22006
rect 538 21748 93642 21770
rect 6306 21746 6626 21748
rect 38274 21746 38594 21748
rect 3230 20770 31702 20812
rect 3230 20534 3272 20770
rect 3508 20534 31424 20770
rect 31660 20534 31702 20770
rect 3230 20492 31702 20534
rect 37822 20770 67030 20812
rect 37822 20534 37864 20770
rect 38100 20534 66752 20770
rect 66988 20534 67030 20770
rect 37822 20492 67030 20534
rect 6726 20090 13854 20132
rect 6726 19854 6768 20090
rect 7004 19854 13576 20090
rect 13812 19854 13854 20090
rect 6726 19812 13854 19854
rect 27886 20090 31702 20132
rect 27886 19854 27928 20090
rect 28164 19854 31424 20090
rect 31660 19854 31702 20090
rect 27886 19812 31702 19854
rect 41502 20090 54886 20132
rect 41502 19854 41544 20090
rect 41780 19854 54886 20090
rect 41502 19812 54886 19854
rect 4150 19410 31702 19452
rect 4150 19174 4192 19410
rect 4428 19174 31424 19410
rect 31660 19174 31702 19410
rect 4150 19132 31702 19174
rect 54566 18772 54886 19812
rect 63950 20090 67214 20132
rect 63950 19854 66936 20090
rect 67172 19854 67214 20090
rect 63950 19812 67214 19854
rect 63950 18772 64270 19812
rect 54566 18452 64270 18772
rect 12798 18050 31702 18092
rect 12798 17814 31424 18050
rect 31660 17814 31702 18050
rect 12798 17772 31702 17814
rect 41870 18050 67950 18092
rect 41870 17814 41912 18050
rect 42148 17814 67672 18050
rect 67908 17814 67950 18050
rect 41870 17772 67950 17814
rect 12798 17412 13118 17772
rect 5070 17370 13118 17412
rect 5070 17134 5112 17370
rect 5348 17134 13118 17370
rect 5070 17092 13118 17134
rect 13534 17370 28206 17412
rect 13534 17134 13576 17370
rect 13812 17134 27928 17370
rect 28164 17134 28206 17370
rect 13534 17092 28206 17134
rect 5622 16690 36486 16732
rect 5622 16454 5664 16690
rect 5900 16454 36208 16690
rect 36444 16454 36486 16690
rect 5622 16412 36486 16454
rect 41686 16690 68502 16732
rect 41686 16454 41728 16690
rect 41964 16454 68224 16690
rect 68460 16454 68502 16690
rect 41686 16412 68502 16454
rect 7278 16010 31702 16052
rect 7278 15774 7320 16010
rect 7556 15774 31424 16010
rect 31660 15774 31702 16010
rect 7278 15732 31702 15774
rect 7094 15330 31702 15372
rect 7094 15094 7136 15330
rect 7372 15094 31424 15330
rect 31660 15094 31702 15330
rect 7094 15052 31702 15094
rect 7278 11250 31702 11292
rect 7278 11014 7320 11250
rect 7556 11014 31424 11250
rect 31660 11014 31702 11250
rect 7278 10972 31702 11014
rect 3642 4348 3962 4350
rect 35610 4348 35930 4350
rect 40938 4348 41258 4350
rect 538 4326 93642 4348
rect 538 4090 3684 4326
rect 3920 4090 35652 4326
rect 35888 4090 40980 4326
rect 41216 4090 93642 4326
rect 538 4006 93642 4090
rect 538 3770 3684 4006
rect 3920 3770 35652 4006
rect 35888 3770 40980 4006
rect 41216 3770 93642 4006
rect 538 3748 93642 3770
rect 3642 3746 3962 3748
rect 35610 3746 35930 3748
rect 40938 3746 41258 3748
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1918 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1607194113
transform 1 0 814 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607194113
transform 1 0 1918 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607194113
transform 1 0 814 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_250 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 538 0 1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1607194113
transform 1 0 538 0 -1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1607194113
transform 1 0 4126 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1607194113
transform 1 0 3022 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607194113
transform 1 0 3482 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3022 0 -1 592
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3390 0 -1 592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5966 0 1 592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5230 0 1 592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5690 0 -1 592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607194113
transform 1 0 4586 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1607194113
transform 1 0 7346 0 1 592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607194113
transform 1 0 6242 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1607194113
transform 1 0 7438 0 -1 592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1607194113
transform 1 0 6334 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1607194113
transform 1 0 6150 0 1 592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607194113
transform 1 0 6242 0 -1 592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 8082 0 1 592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1607194113
transform -1 0 8450 0 1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1607194113
transform -1 0 8450 0 -1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607194113
transform 1 0 1918 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607194113
transform 1 0 814 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607194113
transform 1 0 538 0 -1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607194113
transform 1 0 3482 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607194113
transform 1 0 3022 0 -1 1680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607194113
transform 1 0 3390 0 -1 1680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607194113
transform 1 0 5690 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607194113
transform 1 0 4586 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607194113
transform 1 0 6794 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_80
timestamp 1607194113
transform 1 0 7898 0 -1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607194113
transform -1 0 8450 0 -1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1607194113
transform 1 0 1918 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607194113
transform 1 0 814 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607194113
transform 1 0 538 0 1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1607194113
transform 1 0 4126 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1607194113
transform 1 0 3022 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1607194113
transform 1 0 5966 0 1 1680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1607194113
transform 1 0 5230 0 1 1680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_74
timestamp 1607194113
transform 1 0 7346 0 1 1680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1607194113
transform 1 0 6242 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607194113
transform 1 0 6150 0 1 1680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_82
timestamp 1607194113
transform 1 0 8082 0 1 1680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607194113
transform -1 0 8450 0 1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607194113
transform 1 0 1918 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607194113
transform 1 0 814 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607194113
transform 1 0 538 0 -1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607194113
transform 1 0 3482 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607194113
transform 1 0 3022 0 -1 2768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607194113
transform 1 0 3390 0 -1 2768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1607194113
transform 1 0 5690 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1607194113
transform 1 0 4586 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1607194113
transform 1 0 6794 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_80
timestamp 1607194113
transform 1 0 7898 0 -1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607194113
transform -1 0 8450 0 -1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1607194113
transform 1 0 1918 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607194113
transform 1 0 814 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607194113
transform 1 0 538 0 1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1607194113
transform 1 0 4126 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1607194113
transform 1 0 3022 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1607194113
transform 1 0 5966 0 1 2768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1607194113
transform 1 0 5230 0 1 2768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_74
timestamp 1607194113
transform 1 0 7346 0 1 2768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1607194113
transform 1 0 6242 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607194113
transform 1 0 6150 0 1 2768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1607194113
transform 1 0 8082 0 1 2768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607194113
transform -1 0 8450 0 1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1607194113
transform 1 0 1918 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607194113
transform 1 0 814 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1607194113
transform 1 0 1918 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607194113
transform 1 0 814 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607194113
transform 1 0 538 0 1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607194113
transform 1 0 538 0 -1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1607194113
transform 1 0 4126 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1607194113
transform 1 0 3022 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1607194113
transform 1 0 3482 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1607194113
transform 1 0 3022 0 -1 3856
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607194113
transform 1 0 3390 0 -1 3856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1607194113
transform 1 0 5966 0 1 3856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1607194113
transform 1 0 5230 0 1 3856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1607194113
transform 1 0 5690 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1607194113
transform 1 0 4586 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_74
timestamp 1607194113
transform 1 0 7346 0 1 3856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1607194113
transform 1 0 6242 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1607194113
transform 1 0 6794 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607194113
transform 1 0 6150 0 1 3856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp 1607194113
transform 1 0 8082 0 1 3856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_80
timestamp 1607194113
transform 1 0 7898 0 -1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607194113
transform -1 0 8450 0 1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607194113
transform -1 0 8450 0 -1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1607194113
transform 1 0 1918 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607194113
transform 1 0 814 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607194113
transform 1 0 538 0 -1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1607194113
transform 1 0 3482 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1607194113
transform 1 0 3022 0 -1 4944
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607194113
transform 1 0 3390 0 -1 4944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1607194113
transform 1 0 5690 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1607194113
transform 1 0 4586 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1607194113
transform 1 0 6794 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_80
timestamp 1607194113
transform 1 0 7898 0 -1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607194113
transform -1 0 8450 0 -1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1607194113
transform 1 0 1918 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607194113
transform 1 0 814 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607194113
transform 1 0 538 0 1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1607194113
transform 1 0 4126 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1607194113
transform 1 0 3022 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1607194113
transform 1 0 5966 0 1 4944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1607194113
transform 1 0 5230 0 1 4944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_74
timestamp 1607194113
transform 1 0 7346 0 1 4944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1607194113
transform 1 0 6242 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607194113
transform 1 0 6150 0 1 4944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_82
timestamp 1607194113
transform 1 0 8082 0 1 4944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607194113
transform -1 0 8450 0 1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1607194113
transform 1 0 1918 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607194113
transform 1 0 814 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607194113
transform 1 0 538 0 -1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1607194113
transform 1 0 3482 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1607194113
transform 1 0 3022 0 -1 6032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607194113
transform 1 0 3390 0 -1 6032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1607194113
transform 1 0 5690 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1607194113
transform 1 0 4586 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1607194113
transform 1 0 6794 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_80
timestamp 1607194113
transform 1 0 7898 0 -1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607194113
transform -1 0 8450 0 -1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1607194113
transform 1 0 1918 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607194113
transform 1 0 814 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607194113
transform 1 0 538 0 1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1607194113
transform 1 0 4126 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1607194113
transform 1 0 3022 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1607194113
transform 1 0 5966 0 1 6032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1607194113
transform 1 0 5230 0 1 6032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_74
timestamp 1607194113
transform 1 0 7346 0 1 6032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1607194113
transform 1 0 6242 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607194113
transform 1 0 6150 0 1 6032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_82
timestamp 1607194113
transform 1 0 8082 0 1 6032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607194113
transform -1 0 8450 0 1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1607194113
transform 1 0 1918 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607194113
transform 1 0 814 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607194113
transform 1 0 538 0 -1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1607194113
transform 1 0 3482 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1607194113
transform 1 0 3022 0 -1 7120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607194113
transform 1 0 3390 0 -1 7120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1607194113
transform 1 0 5690 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1607194113
transform 1 0 4586 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1607194113
transform 1 0 6794 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_80
timestamp 1607194113
transform 1 0 7898 0 -1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607194113
transform -1 0 8450 0 -1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607194113
transform 1 0 1918 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607194113
transform 1 0 814 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1607194113
transform 1 0 1918 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607194113
transform 1 0 814 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607194113
transform 1 0 538 0 -1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607194113
transform 1 0 538 0 1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1607194113
transform 1 0 3482 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607194113
transform 1 0 3022 0 -1 8208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1607194113
transform 1 0 4126 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1607194113
transform 1 0 3022 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607194113
transform 1 0 3390 0 -1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1607194113
transform 1 0 5690 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1607194113
transform 1 0 4586 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1607194113
transform 1 0 5966 0 1 7120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1607194113
transform 1 0 5230 0 1 7120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1607194113
transform 1 0 6794 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_74
timestamp 1607194113
transform 1 0 7346 0 1 7120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1607194113
transform 1 0 6242 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607194113
transform 1 0 6150 0 1 7120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_80
timestamp 1607194113
transform 1 0 7898 0 -1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_82
timestamp 1607194113
transform 1 0 8082 0 1 7120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607194113
transform -1 0 8450 0 -1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607194113
transform -1 0 8450 0 1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1607194113
transform 1 0 1918 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607194113
transform 1 0 814 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607194113
transform 1 0 538 0 1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1607194113
transform 1 0 4126 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1607194113
transform 1 0 3022 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1607194113
transform 1 0 5966 0 1 8208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1607194113
transform 1 0 5230 0 1 8208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_74
timestamp 1607194113
transform 1 0 7346 0 1 8208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1607194113
transform 1 0 6242 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607194113
transform 1 0 6150 0 1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_82
timestamp 1607194113
transform 1 0 8082 0 1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607194113
transform -1 0 8450 0 1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1607194113
transform 1 0 1918 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607194113
transform 1 0 814 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607194113
transform 1 0 538 0 -1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1607194113
transform 1 0 3482 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1607194113
transform 1 0 3022 0 -1 9296
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607194113
transform 1 0 3390 0 -1 9296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1607194113
transform 1 0 5690 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1607194113
transform 1 0 4586 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1607194113
transform 1 0 6794 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_80
timestamp 1607194113
transform 1 0 7898 0 -1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607194113
transform -1 0 8450 0 -1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1607194113
transform 1 0 1918 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607194113
transform 1 0 814 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607194113
transform 1 0 538 0 1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1607194113
transform 1 0 4126 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1607194113
transform 1 0 3022 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1607194113
transform 1 0 5966 0 1 9296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1607194113
transform 1 0 5230 0 1 9296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1607194113
transform 1 0 7346 0 1 9296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1607194113
transform 1 0 6242 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607194113
transform 1 0 6150 0 1 9296
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_82
timestamp 1607194113
transform 1 0 8082 0 1 9296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607194113
transform -1 0 8450 0 1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607194113
transform 1 0 1918 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607194113
transform 1 0 814 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607194113
transform 1 0 538 0 -1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1607194113
transform 1 0 3482 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607194113
transform 1 0 3022 0 -1 10384
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607194113
transform 1 0 3390 0 -1 10384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1607194113
transform 1 0 4586 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5690 0 -1 10384
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1607194113
transform 1 0 7806 0 -1 10384
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 7622 0 -1 10384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__D
timestamp 1607194113
transform 1 0 7438 0 -1 10384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607194113
transform -1 0 8450 0 -1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607194113
transform 1 0 1918 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607194113
transform 1 0 814 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1607194113
transform 1 0 1918 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607194113
transform 1 0 814 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607194113
transform 1 0 538 0 -1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607194113
transform 1 0 538 0 1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1607194113
transform 1 0 3482 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607194113
transform 1 0 3022 0 -1 11472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1607194113
transform 1 0 4126 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1607194113
transform 1 0 3022 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607194113
transform 1 0 3390 0 -1 11472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1607194113
transform 1 0 5690 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1607194113
transform 1 0 4586 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1607194113
transform 1 0 5966 0 1 10384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1607194113
transform 1 0 5230 0 1 10384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1607194113
transform 1 0 6794 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_74
timestamp 1607194113
transform 1 0 7346 0 1 10384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1607194113
transform 1 0 6242 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607194113
transform 1 0 6150 0 1 10384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_80
timestamp 1607194113
transform 1 0 7898 0 -1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_82
timestamp 1607194113
transform 1 0 8082 0 1 10384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607194113
transform -1 0 8450 0 -1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607194113
transform -1 0 8450 0 1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1607194113
transform 1 0 1918 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607194113
transform 1 0 814 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607194113
transform 1 0 538 0 1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1607194113
transform 1 0 4126 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1607194113
transform 1 0 3022 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1607194113
transform 1 0 5966 0 1 11472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1607194113
transform 1 0 5230 0 1 11472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_74
timestamp 1607194113
transform 1 0 7346 0 1 11472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1607194113
transform 1 0 6242 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607194113
transform 1 0 6150 0 1 11472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1607194113
transform 1 0 8082 0 1 11472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607194113
transform -1 0 8450 0 1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607194113
transform 1 0 1918 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607194113
transform 1 0 814 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607194113
transform 1 0 538 0 -1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607194113
transform 1 0 3482 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607194113
transform 1 0 3022 0 -1 12560
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607194113
transform 1 0 3390 0 -1 12560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1607194113
transform 1 0 5690 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1607194113
transform 1 0 4586 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1607194113
transform 1 0 6794 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_80
timestamp 1607194113
transform 1 0 7898 0 -1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607194113
transform -1 0 8450 0 -1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1607194113
transform 1 0 1918 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607194113
transform 1 0 814 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607194113
transform 1 0 538 0 1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1607194113
transform 1 0 4126 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1607194113
transform 1 0 3022 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1607194113
transform 1 0 5966 0 1 12560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1607194113
transform 1 0 5230 0 1 12560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_74
timestamp 1607194113
transform 1 0 7346 0 1 12560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1607194113
transform 1 0 6242 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607194113
transform 1 0 6150 0 1 12560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_82
timestamp 1607194113
transform 1 0 8082 0 1 12560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607194113
transform -1 0 8450 0 1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607194113
transform 1 0 1918 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607194113
transform 1 0 814 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607194113
transform 1 0 538 0 -1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1607194113
transform 1 0 3482 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607194113
transform 1 0 3022 0 -1 13648
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607194113
transform 1 0 3390 0 -1 13648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1607194113
transform 1 0 5690 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1607194113
transform 1 0 4586 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1607194113
transform 1 0 6794 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_80
timestamp 1607194113
transform 1 0 7898 0 -1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607194113
transform -1 0 8450 0 -1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1607194113
transform 1 0 1918 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607194113
transform 1 0 814 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607194113
transform 1 0 538 0 1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1607194113
transform 1 0 4126 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1607194113
transform 1 0 3022 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1607194113
transform 1 0 5966 0 1 13648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1607194113
transform 1 0 5230 0 1 13648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_74
timestamp 1607194113
transform 1 0 7346 0 1 13648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1607194113
transform 1 0 6242 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607194113
transform 1 0 6150 0 1 13648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_82
timestamp 1607194113
transform 1 0 8082 0 1 13648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607194113
transform -1 0 8450 0 1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1607194113
transform 1 0 1918 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607194113
transform 1 0 814 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1607194113
transform 1 0 1918 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607194113
transform 1 0 814 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607194113
transform 1 0 538 0 1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607194113
transform 1 0 538 0 -1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1607194113
transform 1 0 4126 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1607194113
transform 1 0 3022 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1607194113
transform 1 0 3482 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1607194113
transform 1 0 3022 0 -1 14736
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607194113
transform 1 0 3390 0 -1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1607194113
transform 1 0 5966 0 1 14736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1607194113
transform 1 0 5230 0 1 14736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1607194113
transform 1 0 4586 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1361_
timestamp 1607194113
transform 1 0 5690 0 -1 14736
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_27_76
timestamp 1607194113
transform 1 0 7530 0 1 14736
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1607194113
transform 1 0 6978 0 1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1607194113
transform 1 0 6242 0 1 14736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1607194113
transform 1 0 7622 0 -1 14736
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__CLK
timestamp 1607194113
transform 1 0 7438 0 -1 14736
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A
timestamp 1607194113
transform 1 0 7346 0 1 14736
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607194113
transform 1 0 6150 0 1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 7070 0 1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_82
timestamp 1607194113
transform 1 0 8082 0 1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607194113
transform -1 0 8450 0 1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607194113
transform -1 0 8450 0 -1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1607194113
transform 1 0 1918 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607194113
transform 1 0 814 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607194113
transform 1 0 538 0 -1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1607194113
transform 1 0 3482 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1607194113
transform 1 0 3022 0 -1 15824
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607194113
transform 1 0 3390 0 -1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_52
timestamp 1607194113
transform 1 0 5322 0 -1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_44
timestamp 1607194113
transform 1 0 4586 0 -1 15824
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1360_
timestamp 1607194113
transform 1 0 5414 0 -1 15824
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_28_74
timestamp 1607194113
transform 1 0 7346 0 -1 15824
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__CLK
timestamp 1607194113
transform 1 0 7162 0 -1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_82
timestamp 1607194113
transform 1 0 8082 0 -1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607194113
transform -1 0 8450 0 -1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1607194113
transform 1 0 1918 0 1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1607194113
transform 1 0 814 0 1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607194113
transform 1 0 538 0 1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1607194113
transform 1 0 3022 0 1 15824
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__B1
timestamp 1607194113
transform 1 0 3758 0 1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3942 0 1 15824
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1607194113
transform 1 0 5782 0 1 15824
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A2_N
timestamp 1607194113
transform 1 0 5598 0 1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__B2
timestamp 1607194113
transform 1 0 5414 0 1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1607194113
transform 1 0 6886 0 1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1607194113
transform 1 0 6242 0 1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__A
timestamp 1607194113
transform 1 0 6702 0 1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607194113
transform 1 0 6150 0 1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1307_
timestamp 1607194113
transform 1 0 6426 0 1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_81
timestamp 1607194113
transform 1 0 7990 0 1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607194113
transform -1 0 8450 0 1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1607194113
transform 1 0 1918 0 -1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607194113
transform 1 0 814 0 -1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607194113
transform 1 0 538 0 -1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1607194113
transform 1 0 3482 0 -1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1607194113
transform 1 0 3022 0 -1 16912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607194113
transform 1 0 3390 0 -1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_48
timestamp 1607194113
transform 1 0 4954 0 -1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_44
timestamp 1607194113
transform 1 0 4586 0 -1 16912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A2_N
timestamp 1607194113
transform 1 0 5046 0 -1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__B2
timestamp 1607194113
transform 1 0 5230 0 -1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__B1
timestamp 1607194113
transform 1 0 5414 0 -1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1306_
timestamp 1607194113
transform 1 0 5598 0 -1 16912
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_71
timestamp 1607194113
transform 1 0 7070 0 -1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607194113
transform -1 0 8450 0 -1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1607194113
transform 1 0 1918 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607194113
transform 1 0 814 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607194113
transform 1 0 538 0 1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1607194113
transform 1 0 4126 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1607194113
transform 1 0 3022 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1607194113
transform 1 0 5966 0 1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1607194113
transform 1 0 5230 0 1 16912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_74
timestamp 1607194113
transform 1 0 7346 0 1 16912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1607194113
transform 1 0 6242 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607194113
transform 1 0 6150 0 1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_82
timestamp 1607194113
transform 1 0 8082 0 1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607194113
transform -1 0 8450 0 1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1607194113
transform 1 0 1918 0 -1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1607194113
transform 1 0 814 0 -1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607194113
transform 1 0 538 0 -1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1607194113
transform 1 0 3482 0 -1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1607194113
transform 1 0 3022 0 -1 18000
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607194113
transform 1 0 3390 0 -1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_50
timestamp 1607194113
transform 1 0 5138 0 -1 18000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_44
timestamp 1607194113
transform 1 0 4586 0 -1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A
timestamp 1607194113
transform 1 0 4954 0 -1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1359_
timestamp 1607194113
transform 1 0 5690 0 -1 18000
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1313_
timestamp 1607194113
transform 1 0 4678 0 -1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1607194113
transform 1 0 7622 0 -1 18000
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1607194113
transform 1 0 7438 0 -1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607194113
transform -1 0 8450 0 -1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607194113
transform 1 0 1918 0 -1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607194113
transform 1 0 814 0 -1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1607194113
transform 1 0 1918 0 1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607194113
transform 1 0 814 0 1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607194113
transform 1 0 538 0 -1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607194113
transform 1 0 538 0 1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1607194113
transform 1 0 3022 0 -1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_33
timestamp 1607194113
transform 1 0 3574 0 1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_27
timestamp 1607194113
transform 1 0 3022 0 1 18000
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__B1
timestamp 1607194113
transform 1 0 3206 0 -1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607194113
transform 1 0 3390 0 -1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1358_
timestamp 1607194113
transform 1 0 3666 0 1 18000
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1314_
timestamp 1607194113
transform 1 0 3482 0 -1 19088
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_34_56
timestamp 1607194113
transform 1 0 5690 0 -1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_48
timestamp 1607194113
transform 1 0 4954 0 -1 19088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_55
timestamp 1607194113
transform 1 0 5598 0 1 18000
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__CLK
timestamp 1607194113
transform 1 0 5414 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__B1
timestamp 1607194113
transform 1 0 5782 0 -1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1312_
timestamp 1607194113
transform 1 0 5966 0 -1 19088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_34_75
timestamp 1607194113
transform 1 0 7438 0 -1 19088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_77
timestamp 1607194113
transform 1 0 7622 0 1 18000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_70
timestamp 1607194113
transform 1 0 6978 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_62
timestamp 1607194113
transform 1 0 6242 0 1 18000
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1607194113
transform 1 0 7438 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607194113
transform 1 0 6150 0 1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1309_
timestamp 1607194113
transform 1 0 7162 0 1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607194113
transform -1 0 8450 0 -1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607194113
transform -1 0 8450 0 1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_11
timestamp 1607194113
transform 1 0 1550 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1607194113
transform 1 0 814 0 1 19088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607194113
transform 1 0 538 0 1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1357_
timestamp 1607194113
transform 1 0 1642 0 1 19088
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_35_33
timestamp 1607194113
transform 1 0 3574 0 1 19088
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__CLK
timestamp 1607194113
transform 1 0 3390 0 1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1607194113
transform 1 0 3942 0 1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1607194113
transform 1 0 4126 0 1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_54
timestamp 1607194113
transform 1 0 5506 0 1 19088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1607194113
transform 1 0 4402 0 1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_74
timestamp 1607194113
transform 1 0 7346 0 1 19088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1607194113
transform 1 0 6242 0 1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1607194113
transform 1 0 6058 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607194113
transform 1 0 6150 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_82
timestamp 1607194113
transform 1 0 8082 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607194113
transform -1 0 8450 0 1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1607194113
transform 1 0 1918 0 -1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1607194113
transform 1 0 814 0 -1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607194113
transform 1 0 538 0 -1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1607194113
transform 1 0 3482 0 -1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1607194113
transform 1 0 3022 0 -1 20176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607194113
transform 1 0 3390 0 -1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_44
timestamp 1607194113
transform 1 0 4586 0 -1 20176
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1356_
timestamp 1607194113
transform 1 0 5138 0 -1 20176
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_36_71
timestamp 1607194113
transform 1 0 7070 0 -1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__CLK
timestamp 1607194113
transform 1 0 6886 0 -1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607194113
transform -1 0 8450 0 -1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_19
timestamp 1607194113
transform 1 0 2286 0 1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_15
timestamp 1607194113
transform 1 0 1918 0 1 20176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1607194113
transform 1 0 814 0 1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607194113
transform 1 0 538 0 1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_38
timestamp 1607194113
transform 1 0 4034 0 1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__B1
timestamp 1607194113
transform 1 0 2378 0 1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1317_
timestamp 1607194113
transform 1 0 2562 0 1 20176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_37_58
timestamp 1607194113
transform 1 0 5874 0 1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_50
timestamp 1607194113
transform 1 0 5138 0 1 20176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_79
timestamp 1607194113
transform 1 0 7806 0 1 20176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_67
timestamp 1607194113
transform 1 0 6702 0 1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1607194113
transform 1 0 6518 0 1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607194113
transform 1 0 6150 0 1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1318_
timestamp 1607194113
transform 1 0 6242 0 1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607194113
transform -1 0 8450 0 1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1607194113
transform 1 0 1918 0 -1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1607194113
transform 1 0 814 0 -1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607194113
transform 1 0 538 0 -1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_32
timestamp 1607194113
transform 1 0 3482 0 -1 21264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1607194113
transform 1 0 3022 0 -1 21264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607194113
transform 1 0 3390 0 -1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_40
timestamp 1607194113
transform 1 0 4218 0 -1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1355_
timestamp 1607194113
transform 1 0 4494 0 -1 21264
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_38_73
timestamp 1607194113
transform 1 0 7254 0 -1 21264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_64
timestamp 1607194113
transform 1 0 6426 0 -1 21264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__CLK
timestamp 1607194113
transform 1 0 6242 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A
timestamp 1607194113
transform 1 0 6794 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1607194113
transform 1 0 6978 0 -1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_81
timestamp 1607194113
transform 1 0 7990 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607194113
transform -1 0 8450 0 -1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_15
timestamp 1607194113
transform 1 0 1918 0 1 21264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1607194113
transform 1 0 814 0 1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607194113
transform 1 0 538 0 1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_27
timestamp 1607194113
transform 1 0 3022 0 1 21264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__B1
timestamp 1607194113
transform 1 0 3574 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1319_
timestamp 1607194113
transform 1 0 3758 0 1 21264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2654 0 1 21264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1607194113
transform 1 0 5966 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1607194113
transform 1 0 5230 0 1 21264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_74
timestamp 1607194113
transform 1 0 7346 0 1 21264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1607194113
transform 1 0 6242 0 1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607194113
transform 1 0 6150 0 1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_82
timestamp 1607194113
transform 1 0 8082 0 1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607194113
transform -1 0 8450 0 1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_15
timestamp 1607194113
transform 1 0 1918 0 -1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1607194113
transform 1 0 814 0 -1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607194113
transform 1 0 538 0 -1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1316_
timestamp 1607194113
transform 1 0 2286 0 -1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_32
timestamp 1607194113
transform 1 0 3482 0 -1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_23
timestamp 1607194113
transform 1 0 2654 0 -1 22352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__B1
timestamp 1607194113
transform 1 0 3574 0 -1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607194113
transform 1 0 3390 0 -1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1321_
timestamp 1607194113
transform 1 0 3758 0 -1 22352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_40_51
timestamp 1607194113
transform 1 0 5230 0 -1 22352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__B1
timestamp 1607194113
transform 1 0 5782 0 -1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1325_
timestamp 1607194113
transform 1 0 5966 0 -1 22352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_40_75
timestamp 1607194113
transform 1 0 7438 0 -1 22352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607194113
transform -1 0 8450 0 -1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1607194113
transform 1 0 1918 0 -1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1607194113
transform 1 0 814 0 -1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_11
timestamp 1607194113
transform 1 0 1550 0 1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1607194113
transform 1 0 814 0 1 22352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607194113
transform 1 0 538 0 -1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607194113
transform 1 0 538 0 1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1354_
timestamp 1607194113
transform 1 0 1642 0 1 22352
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_42_37
timestamp 1607194113
transform 1 0 3942 0 -1 23440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1607194113
transform 1 0 3022 0 -1 23440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_39
timestamp 1607194113
transform 1 0 4126 0 1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_33
timestamp 1607194113
transform 1 0 3574 0 1 22352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1607194113
transform 1 0 3390 0 1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1607194113
transform 1 0 3758 0 -1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607194113
transform 1 0 3390 0 -1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1322_
timestamp 1607194113
transform 1 0 3482 0 -1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_45
timestamp 1607194113
transform 1 0 4678 0 -1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_56
timestamp 1607194113
transform 1 0 5690 0 1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_44
timestamp 1607194113
transform 1 0 4586 0 1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1353_
timestamp 1607194113
transform 1 0 4770 0 -1 23440
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1310_
timestamp 1607194113
transform 1 0 4218 0 1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1607194113
transform 1 0 7806 0 -1 23440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_67
timestamp 1607194113
transform 1 0 6702 0 -1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_79
timestamp 1607194113
transform 1 0 7806 0 1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_67
timestamp 1607194113
transform 1 0 6702 0 1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_60
timestamp 1607194113
transform 1 0 6058 0 1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__CLK
timestamp 1607194113
transform 1 0 6518 0 -1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 1607194113
transform 1 0 6518 0 1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607194113
transform 1 0 6150 0 1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1324_
timestamp 1607194113
transform 1 0 6242 0 1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607194113
transform -1 0 8450 0 -1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607194113
transform -1 0 8450 0 1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1607194113
transform 1 0 814 0 1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__B1
timestamp 1607194113
transform 1 0 1918 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607194113
transform 1 0 538 0 1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1323_
timestamp 1607194113
transform 1 0 2102 0 1 23440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_43_33
timestamp 1607194113
transform 1 0 3574 0 1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1607194113
transform 1 0 5782 0 1 23440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_45
timestamp 1607194113
transform 1 0 4678 0 1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_77
timestamp 1607194113
transform 1 0 7622 0 1 23440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_70
timestamp 1607194113
transform 1 0 6978 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_62
timestamp 1607194113
transform 1 0 6242 0 1 23440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1607194113
transform 1 0 7438 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607194113
transform 1 0 6150 0 1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1607194113
transform 1 0 7162 0 1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607194113
transform -1 0 8450 0 1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1607194113
transform 1 0 1918 0 -1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1607194113
transform 1 0 814 0 -1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1607194113
transform 1 0 538 0 -1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_27
timestamp 1607194113
transform 1 0 3022 0 -1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__B1
timestamp 1607194113
transform 1 0 3206 0 -1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607194113
transform 1 0 3390 0 -1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1302_
timestamp 1607194113
transform 1 0 3482 0 -1 24528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_44_50
timestamp 1607194113
transform 1 0 5138 0 -1 24528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__B2
timestamp 1607194113
transform 1 0 4954 0 -1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1406_
timestamp 1607194113
transform 1 0 5690 0 -1 24528
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1607194113
transform 1 0 7622 0 -1 24528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__CLK
timestamp 1607194113
transform 1 0 7438 0 -1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1607194113
transform -1 0 8450 0 -1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_18
timestamp 1607194113
transform 1 0 2194 0 1 24528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_11
timestamp 1607194113
transform 1 0 1550 0 1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 1607194113
transform 1 0 814 0 1 24528
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1607194113
transform 1 0 2010 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1607194113
transform 1 0 538 0 1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1297_
timestamp 1607194113
transform 1 0 1642 0 1 24528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1363_
timestamp 1607194113
transform 1 0 2746 0 1 24528
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1607194113
transform 1 0 5782 0 1 24528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_45
timestamp 1607194113
transform 1 0 4678 0 1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__CLK
timestamp 1607194113
transform 1 0 4494 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_77
timestamp 1607194113
transform 1 0 7622 0 1 24528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_70
timestamp 1607194113
transform 1 0 6978 0 1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_62
timestamp 1607194113
transform 1 0 6242 0 1 24528
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1607194113
transform 1 0 7438 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607194113
transform 1 0 6150 0 1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1284_
timestamp 1607194113
transform 1 0 7070 0 1 24528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1607194113
transform -1 0 8450 0 1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1607194113
transform 1 0 1918 0 -1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1607194113
transform 1 0 814 0 -1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1607194113
transform 1 0 538 0 -1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_37
timestamp 1607194113
transform 1 0 3942 0 -1 25616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1607194113
transform 1 0 3022 0 -1 25616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A
timestamp 1607194113
transform 1 0 3758 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607194113
transform 1 0 3390 0 -1 25616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1607194113
transform 1 0 3482 0 -1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_59
timestamp 1607194113
transform 1 0 5966 0 -1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__B1
timestamp 1607194113
transform 1 0 4310 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1300_
timestamp 1607194113
transform 1 0 4494 0 -1 25616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_46_71
timestamp 1607194113
transform 1 0 7070 0 -1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1607194113
transform -1 0 8450 0 -1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1607194113
transform 1 0 1918 0 -1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1607194113
transform 1 0 814 0 -1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_15
timestamp 1607194113
transform 1 0 1918 0 1 25616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1607194113
transform 1 0 814 0 1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1607194113
transform 1 0 538 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1607194113
transform 1 0 538 0 1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_39
timestamp 1607194113
transform 1 0 4126 0 -1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_32
timestamp 1607194113
transform 1 0 3482 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1607194113
transform 1 0 3022 0 -1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1607194113
transform 1 0 4126 0 1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1607194113
transform 1 0 3942 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__B1
timestamp 1607194113
transform 1 0 2470 0 1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607194113
transform 1 0 3390 0 -1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1298_
timestamp 1607194113
transform 1 0 2654 0 1 25616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1296_
timestamp 1607194113
transform 1 0 3666 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_51
timestamp 1607194113
transform 1 0 5230 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1607194113
transform 1 0 5966 0 1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1607194113
transform 1 0 5230 0 1 25616
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1364_
timestamp 1607194113
transform 1 0 5506 0 -1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_48_75
timestamp 1607194113
transform 1 0 7438 0 -1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_79
timestamp 1607194113
transform 1 0 7806 0 1 25616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_67
timestamp 1607194113
transform 1 0 6702 0 1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__CLK
timestamp 1607194113
transform 1 0 7254 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1607194113
transform 1 0 6518 0 1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607194113
transform 1 0 6150 0 1 25616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1299_
timestamp 1607194113
transform 1 0 6242 0 1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1607194113
transform -1 0 8450 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1607194113
transform -1 0 8450 0 1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_15
timestamp 1607194113
transform 1 0 1918 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1607194113
transform 1 0 814 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1607194113
transform 1 0 538 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1365_
timestamp 1607194113
transform 1 0 2286 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__CLK
timestamp 1607194113
transform 1 0 4034 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_58
timestamp 1607194113
transform 1 0 5874 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_50
timestamp 1607194113
transform 1 0 5138 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_40
timestamp 1607194113
transform 1 0 4218 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1160_
timestamp 1607194113
transform 1 0 4770 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_74
timestamp 1607194113
transform 1 0 7346 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1607194113
transform 1 0 6242 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607194113
transform 1 0 6150 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_86
timestamp 1607194113
transform 1 0 8450 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B1
timestamp 1607194113
transform 1 0 9186 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1230_
timestamp 1607194113
transform 1 0 9370 0 1 26704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_49_112
timestamp 1607194113
transform 1 0 10842 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A1
timestamp 1607194113
transform 1 0 13234 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A2
timestamp 1607194113
transform 1 0 13050 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B1
timestamp 1607194113
transform 1 0 11578 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607194113
transform 1 0 11762 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0999_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 11854 0 1 26704
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_49_156
timestamp 1607194113
transform 1 0 14890 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_152
timestamp 1607194113
transform 1 0 14522 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_140
timestamp 1607194113
transform 1 0 13418 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 14982 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_168
timestamp 1607194113
transform 1 0 15994 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_160
timestamp 1607194113
transform 1 0 15258 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_i_A
timestamp 1607194113
transform 1 0 16822 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1607194113
transform 1 0 16638 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk_i
timestamp 1607194113
transform 1 0 16086 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1607194113
transform 1 0 16362 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_184
timestamp 1607194113
transform 1 0 17466 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_179
timestamp 1607194113
transform 1 0 17006 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__CLK
timestamp 1607194113
transform 1 0 17834 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607194113
transform 1 0 17374 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1404_
timestamp 1607194113
transform 1 0 18018 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_209
timestamp 1607194113
transform 1 0 19766 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1229_
timestamp 1607194113
transform 1 0 20502 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_3
timestamp 1607194113
transform 1 0 814 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1607194113
transform 1 0 538 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1607194113
transform 1 0 906 0 -1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1607194113
transform 1 0 3482 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1607194113
transform 1 0 3022 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__CLK
timestamp 1607194113
transform 1 0 2838 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__D
timestamp 1607194113
transform 1 0 2654 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607194113
transform 1 0 3390 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_56
timestamp 1607194113
transform 1 0 5690 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1607194113
transform 1 0 4586 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_62
timestamp 1607194113
transform 1 0 6242 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B1
timestamp 1607194113
transform 1 0 6334 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1216_
timestamp 1607194113
transform 1 0 6518 0 -1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_93
timestamp 1607194113
transform 1 0 9094 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 1607194113
transform 1 0 8910 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_87
timestamp 1607194113
transform 1 0 8542 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A2_N
timestamp 1607194113
transform 1 0 8358 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B2
timestamp 1607194113
transform 1 0 8174 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1_N
timestamp 1607194113
transform 1 0 7990 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607194113
transform 1 0 9002 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_105
timestamp 1607194113
transform 1 0 10198 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 1607194113
transform 1 0 10750 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0993_
timestamp 1607194113
transform 1 0 10934 0 -1 27792
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_50_138
timestamp 1607194113
transform 1 0 13234 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_128
timestamp 1607194113
transform 1 0 12314 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A2
timestamp 1607194113
transform 1 0 12130 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1607194113
transform 1 0 12682 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0951_
timestamp 1607194113
transform 1 0 12866 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_154
timestamp 1607194113
transform 1 0 14706 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_50_150
timestamp 1607194113
transform 1 0 14338 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607194113
transform 1 0 14614 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_165
timestamp 1607194113
transform 1 0 15718 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B1
timestamp 1607194113
transform 1 0 15258 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk_i
timestamp 1607194113
transform 1 0 15442 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1232_
timestamp 1607194113
transform 1 0 15810 0 -1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_184
timestamp 1607194113
transform 1 0 17466 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B2
timestamp 1607194113
transform 1 0 17282 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__B1
timestamp 1607194113
transform 1 0 17834 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1231_
timestamp 1607194113
transform 1 0 18018 0 -1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_215
timestamp 1607194113
transform 1 0 20318 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_208
timestamp 1607194113
transform 1 0 19674 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A1_N
timestamp 1607194113
transform 1 0 19490 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607194113
transform 1 0 20226 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_11
timestamp 1607194113
transform 1 0 1550 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1607194113
transform 1 0 814 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1607194113
transform 1 0 538 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1352_
timestamp 1607194113
transform 1 0 1642 0 1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_33
timestamp 1607194113
transform 1 0 3574 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__CLK
timestamp 1607194113
transform 1 0 3390 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1607194113
transform 1 0 5782 0 1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_45
timestamp 1607194113
transform 1 0 4678 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_62
timestamp 1607194113
transform 1 0 6242 0 1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607194113
transform 1 0 6150 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1415_
timestamp 1607194113
transform 1 0 6610 0 1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_96
timestamp 1607194113
transform 1 0 9370 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_87
timestamp 1607194113
transform 1 0 8542 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__CLK
timestamp 1607194113
transform 1 0 8358 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1607194113
transform 1 0 9094 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_108
timestamp 1607194113
transform 1 0 10474 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1607194113
transform 1 0 11578 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607194113
transform 1 0 11762 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 11854 0 1 27792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_51_154
timestamp 1607194113
transform 1 0 14706 0 1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_142
timestamp 1607194113
transform 1 0 13602 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B1
timestamp 1607194113
transform 1 0 15074 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A2
timestamp 1607194113
transform 1 0 13418 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_175
timestamp 1607194113
transform 1 0 16638 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A2
timestamp 1607194113
transform 1 0 15258 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1010_
timestamp 1607194113
transform 1 0 15442 0 1 27792
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_51_184
timestamp 1607194113
transform 1 0 17466 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__CLK
timestamp 1607194113
transform 1 0 17742 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607194113
transform 1 0 17374 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1414_
timestamp 1607194113
transform 1 0 17926 0 1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1607194113
transform 1 0 19674 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1607194113
transform 1 0 1918 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1607194113
transform 1 0 814 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1607194113
transform 1 0 538 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1607194113
transform 1 0 3482 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1607194113
transform 1 0 3022 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607194113
transform 1 0 3390 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_56
timestamp 1607194113
transform 1 0 5690 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1607194113
transform 1 0 4586 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_69
timestamp 1607194113
transform 1 0 6886 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_64
timestamp 1607194113
transform 1 0 6426 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0682_
timestamp 1607194113
transform 1 0 6518 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_89
timestamp 1607194113
transform 1 0 8726 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_81
timestamp 1607194113
transform 1 0 7990 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607194113
transform 1 0 9002 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0994_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 9094 0 -1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_52_114
timestamp 1607194113
transform 1 0 11026 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_102
timestamp 1607194113
transform 1 0 9922 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A1
timestamp 1607194113
transform 1 0 11302 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _1002_
timestamp 1607194113
transform 1 0 11486 0 -1 28880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_52_138
timestamp 1607194113
transform 1 0 13234 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A2
timestamp 1607194113
transform 1 0 13050 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_150
timestamp 1607194113
transform 1 0 14338 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1607194113
transform 1 0 15074 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607194113
transform 1 0 14614 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0944_
timestamp 1607194113
transform 1 0 14706 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_175
timestamp 1607194113
transform 1 0 16638 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_160
timestamp 1607194113
transform 1 0 15258 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1607194113
transform 1 0 15626 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__B
timestamp 1607194113
transform 1 0 15810 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15994 0 -1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B1
timestamp 1607194113
transform 1 0 17190 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1217_
timestamp 1607194113
transform 1 0 17374 0 -1 28880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1607194113
transform 1 0 20318 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1607194113
transform 1 0 20134 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_205
timestamp 1607194113
transform 1 0 19398 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A2_N
timestamp 1607194113
transform 1 0 19214 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B2
timestamp 1607194113
transform 1 0 19030 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1_N
timestamp 1607194113
transform 1 0 18846 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607194113
transform 1 0 20226 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_11
timestamp 1607194113
transform 1 0 1550 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1607194113
transform 1 0 814 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1607194113
transform 1 0 538 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1351_
timestamp 1607194113
transform 1 0 1642 0 1 28880
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_53_33
timestamp 1607194113
transform 1 0 3574 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__CLK
timestamp 1607194113
transform 1 0 3390 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1607194113
transform 1 0 5782 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_45
timestamp 1607194113
transform 1 0 4678 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_73
timestamp 1607194113
transform 1 0 7254 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_62
timestamp 1607194113
transform 1 0 6242 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607194113
transform 1 0 6150 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1159_
timestamp 1607194113
transform 1 0 6426 0 1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_53_88
timestamp 1607194113
transform 1 0 8634 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0942_
timestamp 1607194113
transform 1 0 7990 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_53_116
timestamp 1607194113
transform 1 0 11210 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_104
timestamp 1607194113
transform 1 0 10106 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_100
timestamp 1607194113
transform 1 0 9738 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__D
timestamp 1607194113
transform 1 0 11026 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1000_
timestamp 1607194113
transform 1 0 10198 0 1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_53_131
timestamp 1607194113
transform 1 0 12590 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_123
timestamp 1607194113
transform 1 0 11854 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1607194113
transform 1 0 13142 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607194113
transform 1 0 11762 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1607194113
transform 1 0 12866 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1607194113
transform 1 0 14430 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_139
timestamp 1607194113
transform 1 0 13326 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_175
timestamp 1607194113
transform 1 0 16638 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_163
timestamp 1607194113
transform 1 0 15534 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_187
timestamp 1607194113
transform 1 0 17742 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607194113
transform 1 0 17374 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1607194113
transform 1 0 17466 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_216
timestamp 1607194113
transform 1 0 20410 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_204
timestamp 1607194113
transform 1 0 19306 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1607194113
transform 1 0 19122 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1607194113
transform 1 0 18846 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_11
timestamp 1607194113
transform 1 0 1550 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 1607194113
transform 1 0 814 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1607194113
transform 1 0 1918 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1607194113
transform 1 0 814 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1607194113
transform 1 0 538 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1607194113
transform 1 0 538 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1350_
timestamp 1607194113
transform 1 0 1642 0 1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_55_33
timestamp 1607194113
transform 1 0 3574 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1607194113
transform 1 0 3482 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1607194113
transform 1 0 3022 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__CLK
timestamp 1607194113
transform 1 0 3390 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607194113
transform 1 0 3390 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_53
timestamp 1607194113
transform 1 0 5414 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_45
timestamp 1607194113
transform 1 0 4678 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1607194113
transform 1 0 4586 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _0943_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5690 0 -1 29968
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _0679_
timestamp 1607194113
transform 1 0 5046 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_72
timestamp 1607194113
transform 1 0 7162 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_62
timestamp 1607194113
transform 1 0 6242 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_73
timestamp 1607194113
transform 1 0 7254 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607194113
transform 1 0 6150 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1004_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6334 0 1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_55_89
timestamp 1607194113
transform 1 0 8726 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_91
timestamp 1607194113
transform 1 0 8910 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1607194113
transform 1 0 8358 0 -1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607194113
transform 1 0 9002 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1283_
timestamp 1607194113
transform 1 0 9094 0 -1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0950_
timestamp 1607194113
transform 1 0 9462 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _0908_
timestamp 1607194113
transform 1 0 7898 0 1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1607194113
transform 1 0 10934 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_101
timestamp 1607194113
transform 1 0 9830 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_114
timestamp 1607194113
transform 1 0 11026 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_102
timestamp 1607194113
transform 1 0 9922 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1220_
timestamp 1607194113
transform 1 0 11302 0 -1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_55_123
timestamp 1607194113
transform 1 0 11854 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_121
timestamp 1607194113
transform 1 0 11670 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_138
timestamp 1607194113
transform 1 0 13234 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_128
timestamp 1607194113
transform 1 0 12314 0 -1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__D
timestamp 1607194113
transform 1 0 12130 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607194113
transform 1 0 11762 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1607194113
transform 1 0 12866 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_4  _0995_
timestamp 1607194113
transform 1 0 11946 0 1 29968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_55_155
timestamp 1607194113
transform 1 0 14798 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_143
timestamp 1607194113
transform 1 0 13694 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_154
timestamp 1607194113
transform 1 0 14706 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_150
timestamp 1607194113
transform 1 0 14338 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B2
timestamp 1607194113
transform 1 0 13510 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607194113
transform 1 0 14614 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_167
timestamp 1607194113
transform 1 0 15902 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_166
timestamp 1607194113
transform 1 0 15810 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__CLK
timestamp 1607194113
transform 1 0 15902 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1374_
timestamp 1607194113
transform 1 0 16086 0 -1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_55_184
timestamp 1607194113
transform 1 0 17466 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_179
timestamp 1607194113
transform 1 0 17006 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_196
timestamp 1607194113
transform 1 0 18570 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1607194113
transform 1 0 17834 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__CLK
timestamp 1607194113
transform 1 0 17742 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607194113
transform 1 0 17374 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1373_
timestamp 1607194113
transform 1 0 17926 0 1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1607194113
transform 1 0 18662 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1607194113
transform 1 0 19674 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_215
timestamp 1607194113
transform 1 0 20318 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_202
timestamp 1607194113
transform 1 0 19122 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1607194113
transform 1 0 18938 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607194113
transform 1 0 20226 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1607194113
transform 1 0 1918 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1607194113
transform 1 0 814 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1607194113
transform 1 0 538 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_38
timestamp 1607194113
transform 1 0 4034 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_32
timestamp 1607194113
transform 1 0 3482 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1607194113
transform 1 0 3022 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1607194113
transform 1 0 4126 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607194113
transform 1 0 3390 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_57
timestamp 1607194113
transform 1 0 5782 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_45
timestamp 1607194113
transform 1 0 4678 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1607194113
transform 1 0 5230 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1607194113
transform 1 0 4310 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0680_
timestamp 1607194113
transform 1 0 5414 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_74
timestamp 1607194113
transform 1 0 7346 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _0949_
timestamp 1607194113
transform 1 0 6518 0 -1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_93
timestamp 1607194113
transform 1 0 9094 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_56_86
timestamp 1607194113
transform 1 0 8450 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607194113
transform 1 0 9002 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_113
timestamp 1607194113
transform 1 0 10934 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_101
timestamp 1607194113
transform 1 0 9830 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__D
timestamp 1607194113
transform 1 0 9922 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0683_
timestamp 1607194113
transform 1 0 10106 0 -1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B2
timestamp 1607194113
transform 1 0 13234 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1001_
timestamp 1607194113
transform 1 0 11670 0 -1 31056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_56_154
timestamp 1607194113
transform 1 0 14706 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_150
timestamp 1607194113
transform 1 0 14338 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_142
timestamp 1607194113
transform 1 0 13602 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B1
timestamp 1607194113
transform 1 0 13418 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607194113
transform 1 0 14614 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__B1
timestamp 1607194113
transform 1 0 15810 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1278_
timestamp 1607194113
transform 1 0 15994 0 -1 31056
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_56_194
timestamp 1607194113
transform 1 0 18386 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1607194113
transform 1 0 17650 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A1_N
timestamp 1607194113
transform 1 0 17466 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1607194113
transform 1 0 18478 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_215
timestamp 1607194113
transform 1 0 20318 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_211
timestamp 1607194113
transform 1 0 19950 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_199
timestamp 1607194113
transform 1 0 18846 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607194113
transform 1 0 20226 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_11
timestamp 1607194113
transform 1 0 1550 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_3
timestamp 1607194113
transform 1 0 814 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1607194113
transform 1 0 538 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1339_
timestamp 1607194113
transform 1 0 1642 0 1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_35
timestamp 1607194113
transform 1 0 3758 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__CLK
timestamp 1607194113
transform 1 0 3574 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__D
timestamp 1607194113
transform 1 0 3390 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_53
timestamp 1607194113
transform 1 0 5414 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B
timestamp 1607194113
transform 1 0 5966 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1607194113
transform 1 0 4862 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0668_
timestamp 1607194113
transform 1 0 5046 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_72
timestamp 1607194113
transform 1 0 7162 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_62
timestamp 1607194113
transform 1 0 6242 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607194113
transform 1 0 6150 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0670_
timestamp 1607194113
transform 1 0 6334 0 1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_96
timestamp 1607194113
transform 1 0 9370 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_84
timestamp 1607194113
transform 1 0 8266 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1607194113
transform 1 0 7898 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_112
timestamp 1607194113
transform 1 0 10842 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0909_
timestamp 1607194113
transform 1 0 10474 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_136
timestamp 1607194113
transform 1 0 13050 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_123
timestamp 1607194113
transform 1 0 11854 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_120
timestamp 1607194113
transform 1 0 11578 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607194113
transform 1 0 11762 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0958_
timestamp 1607194113
transform 1 0 12406 0 1 31056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_57_148
timestamp 1607194113
transform 1 0 14154 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_178
timestamp 1607194113
transform 1 0 16914 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_166
timestamp 1607194113
transform 1 0 15810 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_160
timestamp 1607194113
transform 1 0 15258 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1607194113
transform 1 0 15442 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B1
timestamp 1607194113
transform 1 0 17190 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607194113
transform 1 0 17374 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1279_
timestamp 1607194113
transform 1 0 17466 0 1 31056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_212
timestamp 1607194113
transform 1 0 20042 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_202
timestamp 1607194113
transform 1 0 19122 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1_N
timestamp 1607194113
transform 1 0 18938 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0962_
timestamp 1607194113
transform 1 0 19674 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1607194113
transform 1 0 1918 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1607194113
transform 1 0 814 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1607194113
transform 1 0 538 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1607194113
transform 1 0 3482 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1607194113
transform 1 0 3022 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607194113
transform 1 0 3390 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_55
timestamp 1607194113
transform 1 0 5598 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_44
timestamp 1607194113
transform 1 0 4586 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A
timestamp 1607194113
transform 1 0 5138 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__C
timestamp 1607194113
transform 1 0 5966 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1607194113
transform 1 0 5322 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_72
timestamp 1607194113
transform 1 0 7162 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1607194113
transform 1 0 7714 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1607194113
transform 1 0 6150 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0867_
timestamp 1607194113
transform 1 0 6334 0 -1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1607194113
transform 1 0 9094 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_91
timestamp 1607194113
transform 1 0 8910 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_83
timestamp 1607194113
transform 1 0 8174 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607194113
transform 1 0 9002 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1607194113
transform 1 0 7898 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_113
timestamp 1607194113
transform 1 0 10934 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_105
timestamp 1607194113
transform 1 0 10198 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 11210 0 -1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_136
timestamp 1607194113
transform 1 0 13050 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_127
timestamp 1607194113
transform 1 0 12222 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A
timestamp 1607194113
transform 1 0 12038 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1607194113
transform 1 0 12590 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1607194113
transform 1 0 12774 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_158
timestamp 1607194113
transform 1 0 15074 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_152
timestamp 1607194113
transform 1 0 14522 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_148
timestamp 1607194113
transform 1 0 14154 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607194113
transform 1 0 14614 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0959_
timestamp 1607194113
transform 1 0 14706 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_170
timestamp 1607194113
transform 1 0 16178 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B1
timestamp 1607194113
transform 1 0 16730 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1218_
timestamp 1607194113
transform 1 0 16914 0 -1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_58_196
timestamp 1607194113
transform 1 0 18570 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1_N
timestamp 1607194113
transform 1 0 18386 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_215
timestamp 1607194113
transform 1 0 20318 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_206
timestamp 1607194113
transform 1 0 19490 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607194113
transform 1 0 20226 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0672_
timestamp 1607194113
transform 1 0 19122 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_15
timestamp 1607194113
transform 1 0 1918 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1607194113
transform 1 0 814 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1607194113
transform 1 0 538 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1331_
timestamp 1607194113
transform 1 0 2470 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_59_53
timestamp 1607194113
transform 1 0 5414 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_42
timestamp 1607194113
transform 1 0 4402 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__CLK
timestamp 1607194113
transform 1 0 4218 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1607194113
transform 1 0 4954 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1607194113
transform 1 0 5138 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_74
timestamp 1607194113
transform 1 0 7346 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_62
timestamp 1607194113
transform 1 0 6242 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607194113
transform 1 0 6150 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0907_
timestamp 1607194113
transform 1 0 6978 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_98
timestamp 1607194113
transform 1 0 9554 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_86
timestamp 1607194113
transform 1 0 8450 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_110
timestamp 1607194113
transform 1 0 10658 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_123
timestamp 1607194113
transform 1 0 11854 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607194113
transform 1 0 11762 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1021_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 12130 0 1 32144
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_59_155
timestamp 1607194113
transform 1 0 14798 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_140
timestamp 1607194113
transform 1 0 13418 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1006_
timestamp 1607194113
transform 1 0 14154 0 1 32144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_59_175
timestamp 1607194113
transform 1 0 16638 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_59_163
timestamp 1607194113
transform 1 0 15534 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15810 0 1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__CLK
timestamp 1607194113
transform 1 0 17190 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607194113
transform 1 0 17374 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1413_
timestamp 1607194113
transform 1 0 17466 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_59_215
timestamp 1607194113
transform 1 0 20318 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_203
timestamp 1607194113
transform 1 0 19214 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1607194113
transform 1 0 1918 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1607194113
transform 1 0 814 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1607194113
transform 1 0 538 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1607194113
transform 1 0 3482 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1607194113
transform 1 0 3022 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607194113
transform 1 0 3390 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_44
timestamp 1607194113
transform 1 0 4586 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1444_
timestamp 1607194113
transform 1 0 4678 0 -1 33232
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_60_78
timestamp 1607194113
transform 1 0 7714 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1607194113
transform 1 0 6610 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__CLK
timestamp 1607194113
transform 1 0 6426 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_93
timestamp 1607194113
transform 1 0 9094 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_90
timestamp 1607194113
transform 1 0 8818 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607194113
transform 1 0 9002 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_101
timestamp 1607194113
transform 1 0 9830 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1520_
timestamp 1607194113
transform 1 0 10014 0 -1 33232
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1607194113
transform 1 0 12774 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_124
timestamp 1607194113
transform 1 0 11946 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__CLK
timestamp 1607194113
transform 1 0 11762 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1607194113
transform 1 0 12498 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_154
timestamp 1607194113
transform 1 0 14706 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_152
timestamp 1607194113
transform 1 0 14522 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_144
timestamp 1607194113
transform 1 0 13786 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1607194113
transform 1 0 13326 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607194113
transform 1 0 14614 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1607194113
transform 1 0 13510 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_178
timestamp 1607194113
transform 1 0 16914 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_166
timestamp 1607194113
transform 1 0 15810 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A2_N
timestamp 1607194113
transform 1 0 18662 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1007_
timestamp 1607194113
transform 1 0 17190 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1607194113
transform 1 0 20318 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_213
timestamp 1607194113
transform 1 0 20134 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_201
timestamp 1607194113
transform 1 0 19030 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1_N
timestamp 1607194113
transform 1 0 18846 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607194113
transform 1 0 20226 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1607194113
transform 1 0 1918 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1607194113
transform 1 0 814 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_15
timestamp 1607194113
transform 1 0 1918 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1607194113
transform 1 0 814 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1607194113
transform 1 0 538 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1607194113
transform 1 0 538 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2102 0 1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1607194113
transform 1 0 3482 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1607194113
transform 1 0 3022 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_36
timestamp 1607194113
transform 1 0 3850 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_28
timestamp 1607194113
transform 1 0 3114 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__B1
timestamp 1607194113
transform 1 0 3942 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly_A
timestamp 1607194113
transform 1 0 2930 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1607194113
transform 1 0 3390 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 4126 0 1 33232
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_62_48
timestamp 1607194113
transform 1 0 4954 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_44
timestamp 1607194113
transform 1 0 4586 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_53
timestamp 1607194113
transform 1 0 5414 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1332_
timestamp 1607194113
transform 1 0 5046 0 -1 34320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_70
timestamp 1607194113
transform 1 0 6978 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1607194113
transform 1 0 7346 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1607194113
transform 1 0 6242 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__CLK
timestamp 1607194113
transform 1 0 6794 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607194113
transform 1 0 6150 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_82
timestamp 1607194113
transform 1 0 8082 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_86
timestamp 1607194113
transform 1 0 8450 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__B1
timestamp 1607194113
transform 1 0 8818 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1607194113
transform 1 0 9002 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1445_
timestamp 1607194113
transform 1 0 8726 0 1 33232
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _1170_
timestamp 1607194113
transform 1 0 9094 0 -1 34320
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_119
timestamp 1607194113
transform 1 0 11486 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_107
timestamp 1607194113
transform 1 0 10382 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_110
timestamp 1607194113
transform 1 0 10658 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__CLK
timestamp 1607194113
transform 1 0 10474 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_131
timestamp 1607194113
transform 1 0 12590 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B1
timestamp 1607194113
transform 1 0 13142 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607194113
transform 1 0 11762 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0685_
timestamp 1607194113
transform 1 0 11854 0 1 33232
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1607194113
transform 1 0 14706 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_151
timestamp 1607194113
transform 1 0 14430 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_143
timestamp 1607194113
transform 1 0 13694 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_148
timestamp 1607194113
transform 1 0 14154 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_139
timestamp 1607194113
transform 1 0 13326 0 1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1607194113
transform 1 0 13694 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1607194113
transform 1 0 14614 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1607194113
transform 1 0 13878 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_166
timestamp 1607194113
transform 1 0 15810 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_172
timestamp 1607194113
transform 1 0 16362 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_160
timestamp 1607194113
transform 1 0 15258 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B1
timestamp 1607194113
transform 1 0 15902 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1280_
timestamp 1607194113
transform 1 0 16086 0 -1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_189
timestamp 1607194113
transform 1 0 17926 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_195
timestamp 1607194113
transform 1 0 18478 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_187
timestamp 1607194113
transform 1 0 17742 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_180
timestamp 1607194113
transform 1 0 17098 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B2
timestamp 1607194113
transform 1 0 17742 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1_N
timestamp 1607194113
transform 1 0 17558 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607194113
transform 1 0 17374 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1607194113
transform 1 0 17466 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1607194113
transform 1 0 18754 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_215
timestamp 1607194113
transform 1 0 20318 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_213
timestamp 1607194113
transform 1 0 20134 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1607194113
transform 1 0 19030 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_213
timestamp 1607194113
transform 1 0 20134 0 1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_201
timestamp 1607194113
transform 1 0 19030 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1607194113
transform 1 0 20226 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1607194113
transform 1 0 1918 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1607194113
transform 1 0 814 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1607194113
transform 1 0 538 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1340_
timestamp 1607194113
transform 1 0 2286 0 1 34320
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1607194113
transform 1 0 4034 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_52
timestamp 1607194113
transform 1 0 5322 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1607194113
transform 1 0 4218 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_79
timestamp 1607194113
transform 1 0 7806 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_67
timestamp 1607194113
transform 1 0 6702 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_60
timestamp 1607194113
transform 1 0 6058 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A
timestamp 1607194113
transform 1 0 6242 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1607194113
transform 1 0 6150 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1607194113
transform 1 0 6426 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_91
timestamp 1607194113
transform 1 0 8910 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_115
timestamp 1607194113
transform 1 0 11118 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_103
timestamp 1607194113
transform 1 0 10014 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_138
timestamp 1607194113
transform 1 0 13234 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_131
timestamp 1607194113
transform 1 0 12590 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_123
timestamp 1607194113
transform 1 0 11854 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_121
timestamp 1607194113
transform 1 0 11670 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1607194113
transform 1 0 12682 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1607194113
transform 1 0 11762 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0666_
timestamp 1607194113
transform 1 0 12866 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_150
timestamp 1607194113
transform 1 0 14338 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_178
timestamp 1607194113
transform 1 0 16914 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_174
timestamp 1607194113
transform 1 0 16546 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_162
timestamp 1607194113
transform 1 0 15442 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_198
timestamp 1607194113
transform 1 0 18754 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_186
timestamp 1607194113
transform 1 0 17650 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_182
timestamp 1607194113
transform 1 0 17282 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_i_A
timestamp 1607194113
transform 1 0 17466 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A
timestamp 1607194113
transform 1 0 18570 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk_i
timestamp 1607194113
transform 1 0 17006 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1607194113
transform 1 0 17374 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1277_
timestamp 1607194113
transform 1 0 18202 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_214
timestamp 1607194113
transform 1 0 20226 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_210
timestamp 1607194113
transform 1 0 19858 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A
timestamp 1607194113
transform 1 0 20318 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1329_
timestamp 1607194113
transform 1 0 20502 0 1 34320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_64_11
timestamp 1607194113
transform 1 0 1550 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_3
timestamp 1607194113
transform 1 0 814 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1607194113
transform 1 0 538 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:1.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 1826 0 -1 35408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1607194113
transform 1 0 3482 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_23
timestamp 1607194113
transform 1 0 2654 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1607194113
transform 1 0 3390 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_50
timestamp 1607194113
transform 1 0 5138 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_44
timestamp 1607194113
transform 1 0 4586 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1333_
timestamp 1607194113
transform 1 0 5230 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_72
timestamp 1607194113
transform 1 0 7162 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__CLK
timestamp 1607194113
transform 1 0 6978 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_93
timestamp 1607194113
transform 1 0 9094 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_84
timestamp 1607194113
transform 1 0 8266 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1607194113
transform 1 0 9002 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1446_
timestamp 1607194113
transform 1 0 9830 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_64_134
timestamp 1607194113
transform 1 0 12866 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_122
timestamp 1607194113
transform 1 0 11762 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__CLK
timestamp 1607194113
transform 1 0 11578 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1607194113
transform 1 0 13050 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1024_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13234 0 -1 35408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_64_145
timestamp 1607194113
transform 1 0 13878 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1607194113
transform 1 0 14982 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1607194113
transform 1 0 14614 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1607194113
transform 1 0 14706 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1607194113
transform 1 0 15166 0 -1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__CLK
timestamp 1607194113
transform 1 0 15534 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1372_
timestamp 1607194113
transform 1 0 15718 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_64_184
timestamp 1607194113
transform 1 0 17466 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0674_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 18202 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_215
timestamp 1607194113
transform 1 0 20318 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_206
timestamp 1607194113
transform 1 0 19490 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A2
timestamp 1607194113
transform 1 0 19306 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1607194113
transform 1 0 20226 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_19
timestamp 1607194113
transform 1 0 2286 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_15
timestamp 1607194113
transform 1 0 1918 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1607194113
transform 1 0 814 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1607194113
transform 1 0 538 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__CLK
timestamp 1607194113
transform 1 0 4126 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1341_
timestamp 1607194113
transform 1 0 2378 0 1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_53
timestamp 1607194113
transform 1 0 5414 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_41
timestamp 1607194113
transform 1 0 4310 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_74
timestamp 1607194113
transform 1 0 7346 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_62
timestamp 1607194113
transform 1 0 6242 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1607194113
transform 1 0 6150 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_98
timestamp 1607194113
transform 1 0 9554 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_86
timestamp 1607194113
transform 1 0 8450 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1169_
timestamp 1607194113
transform 1 0 9646 0 1 35408
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_65_113
timestamp 1607194113
transform 1 0 10934 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_121
timestamp 1607194113
transform 1 0 11670 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1607194113
transform 1 0 11762 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1447_
timestamp 1607194113
transform 1 0 11854 0 1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_156
timestamp 1607194113
transform 1 0 14890 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_152
timestamp 1607194113
transform 1 0 14522 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_144
timestamp 1607194113
transform 1 0 13786 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__CLK
timestamp 1607194113
transform 1 0 13602 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk_i
timestamp 1607194113
transform 1 0 14614 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_175
timestamp 1607194113
transform 1 0 16638 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_168
timestamp 1607194113
transform 1 0 15994 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1607194113
transform 1 0 16362 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_196
timestamp 1607194113
transform 1 0 18570 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_184
timestamp 1607194113
transform 1 0 17466 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1607194113
transform 1 0 18386 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1607194113
transform 1 0 17190 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1607194113
transform 1 0 17374 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0675_
timestamp 1607194113
transform 1 0 17558 0 1 35408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_65_208
timestamp 1607194113
transform 1 0 19674 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1328_
timestamp 1607194113
transform 1 0 20042 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_11
timestamp 1607194113
transform 1 0 1550 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_3
timestamp 1607194113
transform 1 0 814 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1607194113
transform 1 0 538 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:2.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 1826 0 -1 36496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1607194113
transform 1 0 3482 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_23
timestamp 1607194113
transform 1 0 2654 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1607194113
transform 1 0 3390 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_52
timestamp 1607194113
transform 1 0 5322 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_44
timestamp 1607194113
transform 1 0 4586 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1334_
timestamp 1607194113
transform 1 0 5506 0 -1 36496
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_75
timestamp 1607194113
transform 1 0 7438 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__CLK
timestamp 1607194113
transform 1 0 7254 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_97
timestamp 1607194113
transform 1 0 9462 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_93
timestamp 1607194113
transform 1 0 9094 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_91
timestamp 1607194113
transform 1 0 8910 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_87
timestamp 1607194113
transform 1 0 8542 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1607194113
transform 1 0 9002 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1162_
timestamp 1607194113
transform 1 0 9554 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_114
timestamp 1607194113
transform 1 0 11026 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_102
timestamp 1607194113
transform 1 0 9922 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1168_
timestamp 1607194113
transform 1 0 11118 0 -1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_66_129
timestamp 1607194113
transform 1 0 12406 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_154
timestamp 1607194113
transform 1 0 14706 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1607194113
transform 1 0 13510 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1607194113
transform 1 0 14614 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_165
timestamp 1607194113
transform 1 0 15718 0 -1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__CLK
timestamp 1607194113
transform 1 0 16270 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk_i
timestamp 1607194113
transform 1 0 15442 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1521_
timestamp 1607194113
transform 1 0 16454 0 -1 36496
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_66_192
timestamp 1607194113
transform 1 0 18202 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_215
timestamp 1607194113
transform 1 0 20318 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_211
timestamp 1607194113
transform 1 0 19950 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_203
timestamp 1607194113
transform 1 0 19214 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1607194113
transform 1 0 20226 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1607194113
transform 1 0 18938 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1607194113
transform 1 0 1918 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1607194113
transform 1 0 814 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_3
timestamp 1607194113
transform 1 0 814 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1607194113
transform 1 0 538 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1607194113
transform 1 0 538 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:3.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 1550 0 1 36496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_68_38
timestamp 1607194113
transform 1 0 4034 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_32
timestamp 1607194113
transform 1 0 3482 0 -1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1607194113
transform 1 0 3022 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_20
timestamp 1607194113
transform 1 0 2378 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1607194113
transform 1 0 3390 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1342_
timestamp 1607194113
transform 1 0 3114 0 1 36496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1335_
timestamp 1607194113
transform 1 0 4126 0 -1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_67_49
timestamp 1607194113
transform 1 0 5046 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__CLK
timestamp 1607194113
transform 1 0 4862 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__CLK
timestamp 1607194113
transform 1 0 5874 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_72
timestamp 1607194113
transform 1 0 7162 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_60
timestamp 1607194113
transform 1 0 6058 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_74
timestamp 1607194113
transform 1 0 7346 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1607194113
transform 1 0 6242 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1607194113
transform 1 0 6150 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_93
timestamp 1607194113
transform 1 0 9094 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_84
timestamp 1607194113
transform 1 0 8266 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_94
timestamp 1607194113
transform 1 0 9186 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_86
timestamp 1607194113
transform 1 0 8450 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A
timestamp 1607194113
transform 1 0 9462 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1607194113
transform 1 0 9002 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1164_
timestamp 1607194113
transform 1 0 9646 0 1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_118
timestamp 1607194113
transform 1 0 11394 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_101
timestamp 1607194113
transform 1 0 9830 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_115
timestamp 1607194113
transform 1 0 11118 0 1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_103
timestamp 1607194113
transform 1 0 10014 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1166_
timestamp 1607194113
transform 1 0 10106 0 -1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_67_135
timestamp 1607194113
transform 1 0 12958 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_123
timestamp 1607194113
transform 1 0 11854 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_121
timestamp 1607194113
transform 1 0 11670 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1607194113
transform 1 0 11762 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1167_
timestamp 1607194113
transform 1 0 12130 0 -1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_68_154
timestamp 1607194113
transform 1 0 14706 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_152
timestamp 1607194113
transform 1 0 14522 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_140
timestamp 1607194113
transform 1 0 13418 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_147
timestamp 1607194113
transform 1 0 14062 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1607194113
transform 1 0 14614 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_171
timestamp 1607194113
transform 1 0 16270 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_162
timestamp 1607194113
transform 1 0 15442 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_173
timestamp 1607194113
transform 1 0 16454 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1607194113
transform 1 0 15902 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_159
timestamp 1607194113
transform 1 0 15166 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1607194113
transform 1 0 15994 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0984_
timestamp 1607194113
transform 1 0 15626 0 -1 37584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1607194113
transform 1 0 16178 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_188
timestamp 1607194113
transform 1 0 17834 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1607194113
transform 1 0 18294 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_181
timestamp 1607194113
transform 1 0 17190 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B
timestamp 1607194113
transform 1 0 18110 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1607194113
transform 1 0 17374 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 17006 0 -1 37584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1005_
timestamp 1607194113
transform 1 0 17466 0 1 36496
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_68_200
timestamp 1607194113
transform 1 0 18938 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_205
timestamp 1607194113
transform 1 0 19398 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__CLK
timestamp 1607194113
transform 1 0 20042 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1607194113
transform 1 0 20502 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B
timestamp 1607194113
transform 1 0 19674 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1607194113
transform 1 0 20226 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1522_
timestamp 1607194113
transform 1 0 20318 0 -1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1013_
timestamp 1607194113
transform 1 0 19858 0 1 36496
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_69_15
timestamp 1607194113
transform 1 0 1918 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1607194113
transform 1 0 814 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1607194113
transform 1 0 538 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1343_
timestamp 1607194113
transform 1 0 2102 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_38
timestamp 1607194113
transform 1 0 4034 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__CLK
timestamp 1607194113
transform 1 0 3850 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_58
timestamp 1607194113
transform 1 0 5874 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_50
timestamp 1607194113
transform 1 0 5138 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_74
timestamp 1607194113
transform 1 0 7346 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_62
timestamp 1607194113
transform 1 0 6242 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1607194113
transform 1 0 6150 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1451_
timestamp 1607194113
transform 1 0 7438 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_96
timestamp 1607194113
transform 1 0 9370 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__CLK
timestamp 1607194113
transform 1 0 9186 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_108
timestamp 1607194113
transform 1 0 10474 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_129
timestamp 1607194113
transform 1 0 12406 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_123
timestamp 1607194113
transform 1 0 11854 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_69_120
timestamp 1607194113
transform 1 0 11578 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1607194113
transform 1 0 11762 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1448_
timestamp 1607194113
transform 1 0 12498 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_151
timestamp 1607194113
transform 1 0 14430 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__CLK
timestamp 1607194113
transform 1 0 14246 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_175
timestamp 1607194113
transform 1 0 16638 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1607194113
transform 1 0 15902 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_163
timestamp 1607194113
transform 1 0 15534 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0977_
timestamp 1607194113
transform 1 0 15994 0 1 37584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_69_195
timestamp 1607194113
transform 1 0 18478 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__C
timestamp 1607194113
transform 1 0 18294 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1607194113
transform 1 0 17374 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0991_
timestamp 1607194113
transform 1 0 17466 0 1 37584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_69_207
timestamp 1607194113
transform 1 0 19582 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1023_
timestamp 1607194113
transform 1 0 20134 0 1 37584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_70_11
timestamp 1607194113
transform 1 0 1550 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_3
timestamp 1607194113
transform 1 0 814 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1607194113
transform 1 0 538 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:4.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 1826 0 -1 38672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_70_32
timestamp 1607194113
transform 1 0 3482 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_23
timestamp 1607194113
transform 1 0 2654 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1607194113
transform 1 0 3390 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1336_
timestamp 1607194113
transform 1 0 4034 0 -1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_59
timestamp 1607194113
transform 1 0 5966 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__CLK
timestamp 1607194113
transform 1 0 5782 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_71
timestamp 1607194113
transform 1 0 7070 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_93
timestamp 1607194113
transform 1 0 9094 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1607194113
transform 1 0 8910 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_83
timestamp 1607194113
transform 1 0 8174 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1607194113
transform 1 0 9002 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_101
timestamp 1607194113
transform 1 0 9830 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1449_
timestamp 1607194113
transform 1 0 10014 0 -1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_136
timestamp 1607194113
transform 1 0 13050 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_124
timestamp 1607194113
transform 1 0 11946 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__CLK
timestamp 1607194113
transform 1 0 11762 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_154
timestamp 1607194113
transform 1 0 14706 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_152
timestamp 1607194113
transform 1 0 14522 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_148
timestamp 1607194113
transform 1 0 14154 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1607194113
transform 1 0 14614 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_177
timestamp 1607194113
transform 1 0 16822 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_166
timestamp 1607194113
transform 1 0 15810 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0961_
timestamp 1607194113
transform 1 0 16178 0 -1 38672
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_70_196
timestamp 1607194113
transform 1 0 18570 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__C
timestamp 1607194113
transform 1 0 18386 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0983_
timestamp 1607194113
transform 1 0 17558 0 -1 38672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_215
timestamp 1607194113
transform 1 0 20318 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_208
timestamp 1607194113
transform 1 0 19674 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1607194113
transform 1 0 20226 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_15
timestamp 1607194113
transform 1 0 1918 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1607194113
transform 1 0 814 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1607194113
transform 1 0 538 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1344_
timestamp 1607194113
transform 1 0 2194 0 1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1607194113
transform 1 0 4126 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__CLK
timestamp 1607194113
transform 1 0 3942 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_59
timestamp 1607194113
transform 1 0 5966 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_51
timestamp 1607194113
transform 1 0 5230 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_74
timestamp 1607194113
transform 1 0 7346 0 1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_62
timestamp 1607194113
transform 1 0 6242 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1607194113
transform 1 0 6150 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_96
timestamp 1607194113
transform 1 0 9370 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A2
timestamp 1607194113
transform 1 0 7898 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1163_
timestamp 1607194113
transform 1 0 8082 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_71_108
timestamp 1607194113
transform 1 0 10474 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_123
timestamp 1607194113
transform 1 0 11854 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_120
timestamp 1607194113
transform 1 0 11578 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1607194113
transform 1 0 11762 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1450_
timestamp 1607194113
transform 1 0 11946 0 1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_71_157
timestamp 1607194113
transform 1 0 14982 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_145
timestamp 1607194113
transform 1 0 13878 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__CLK
timestamp 1607194113
transform 1 0 13694 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_175
timestamp 1607194113
transform 1 0 16638 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_165
timestamp 1607194113
transform 1 0 15718 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0970_
timestamp 1607194113
transform 1 0 15994 0 1 38672
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_71_196
timestamp 1607194113
transform 1 0 18570 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1607194113
transform 1 0 17466 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1607194113
transform 1 0 17374 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0969_
timestamp 1607194113
transform 1 0 18662 0 1 38672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_71_208
timestamp 1607194113
transform 1 0 19674 0 1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__C
timestamp 1607194113
transform 1 0 19490 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0941_
timestamp 1607194113
transform 1 0 20226 0 1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1607194113
transform 1 0 1918 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1607194113
transform 1 0 814 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1607194113
transform 1 0 538 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1607194113
transform 1 0 3022 0 -1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1607194113
transform 1 0 3390 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:5.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 3482 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1607194113
transform 1 0 5414 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1607194113
transform 1 0 4310 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_77
timestamp 1607194113
transform 1 0 7622 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1607194113
transform 1 0 6518 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_93
timestamp 1607194113
transform 1 0 9094 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_89
timestamp 1607194113
transform 1 0 8726 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1607194113
transform 1 0 9002 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_117
timestamp 1607194113
transform 1 0 11302 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_105
timestamp 1607194113
transform 1 0 10198 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1165_
timestamp 1607194113
transform 1 0 11486 0 -1 39760
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_72_133
timestamp 1607194113
transform 1 0 12774 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_154
timestamp 1607194113
transform 1 0 14706 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_145
timestamp 1607194113
transform 1 0 13878 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1607194113
transform 1 0 14614 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_178
timestamp 1607194113
transform 1 0 16914 0 -1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_166
timestamp 1607194113
transform 1 0 15810 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_193
timestamp 1607194113
transform 1 0 18294 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__C
timestamp 1607194113
transform 1 0 18110 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0976_
timestamp 1607194113
transform 1 0 17282 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_72_215
timestamp 1607194113
transform 1 0 20318 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_213
timestamp 1607194113
transform 1 0 20134 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_205
timestamp 1607194113
transform 1 0 19398 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1607194113
transform 1 0 20226 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1607194113
transform 1 0 1918 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1607194113
transform 1 0 814 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1607194113
transform 1 0 538 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1607194113
transform 1 0 4126 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1607194113
transform 1 0 3022 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_59
timestamp 1607194113
transform 1 0 5966 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_51
timestamp 1607194113
transform 1 0 5230 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_62
timestamp 1607194113
transform 1 0 6242 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1607194113
transform 1 0 6150 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1338_
timestamp 1607194113
transform 1 0 6334 0 1 39760
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_73_84
timestamp 1607194113
transform 1 0 8266 0 1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__CLK
timestamp 1607194113
transform 1 0 8082 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1337_
timestamp 1607194113
transform 1 0 8818 0 1 39760
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_73_119
timestamp 1607194113
transform 1 0 11486 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_111
timestamp 1607194113
transform 1 0 10750 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__CLK
timestamp 1607194113
transform 1 0 10566 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_137
timestamp 1607194113
transform 1 0 13142 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_129
timestamp 1607194113
transform 1 0 12406 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_123
timestamp 1607194113
transform 1 0 11854 0 1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1607194113
transform 1 0 11762 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0997_
timestamp 1607194113
transform 1 0 12498 0 1 39760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_73_152
timestamp 1607194113
transform 1 0 14522 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1003_
timestamp 1607194113
transform 1 0 13878 0 1 39760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_73_176
timestamp 1607194113
transform 1 0 16730 0 1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_164
timestamp 1607194113
transform 1 0 15626 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_184
timestamp 1607194113
transform 1 0 17466 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_182
timestamp 1607194113
transform 1 0 17282 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__CLK
timestamp 1607194113
transform 1 0 18570 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1607194113
transform 1 0 17374 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1493_
timestamp 1607194113
transform 1 0 18754 0 1 39760
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_73_217
timestamp 1607194113
transform 1 0 20502 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_11
timestamp 1607194113
transform 1 0 1550 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_3
timestamp 1607194113
transform 1 0 814 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_19
timestamp 1607194113
transform 1 0 2286 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_15
timestamp 1607194113
transform 1 0 1918 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1607194113
transform 1 0 814 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1607194113
transform 1 0 538 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1607194113
transform 1 0 538 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1486_
timestamp 1607194113
transform 1 0 1642 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_75_35
timestamp 1607194113
transform 1 0 3758 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_23
timestamp 1607194113
transform 1 0 2654 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__CLK
timestamp 1607194113
transform 1 0 3574 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__D
timestamp 1607194113
transform 1 0 3390 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1607194113
transform 1 0 3390 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1487_
timestamp 1607194113
transform 1 0 3482 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1607194113
transform 1 0 2378 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_53
timestamp 1607194113
transform 1 0 5414 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_43
timestamp 1607194113
transform 1 0 4494 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_55
timestamp 1607194113
transform 1 0 5598 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__CLK
timestamp 1607194113
transform 1 0 5414 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__D
timestamp 1607194113
transform 1 0 5230 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:6.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 4586 0 1 40848
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_74_63
timestamp 1607194113
transform 1 0 6334 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1607194113
transform 1 0 6150 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1346_
timestamp 1607194113
transform 1 0 6242 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1345_
timestamp 1607194113
transform 1 0 6426 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_95
timestamp 1607194113
transform 1 0 9278 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_83
timestamp 1607194113
transform 1 0 8174 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_93
timestamp 1607194113
transform 1 0 9094 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1607194113
transform 1 0 8910 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1607194113
transform 1 0 8358 0 -1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__CLK
timestamp 1607194113
transform 1 0 7990 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__CLK
timestamp 1607194113
transform 1 0 8174 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1607194113
transform 1 0 9002 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_119
timestamp 1607194113
transform 1 0 11486 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_107
timestamp 1607194113
transform 1 0 10382 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_113
timestamp 1607194113
transform 1 0 10934 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_105
timestamp 1607194113
transform 1 0 10198 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1488_
timestamp 1607194113
transform 1 0 11026 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_75_123
timestamp 1607194113
transform 1 0 11854 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_135
timestamp 1607194113
transform 1 0 12958 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__CLK
timestamp 1607194113
transform 1 0 12774 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1607194113
transform 1 0 11762 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1489_
timestamp 1607194113
transform 1 0 12038 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_158
timestamp 1607194113
transform 1 0 15074 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_146
timestamp 1607194113
transform 1 0 13970 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_154
timestamp 1607194113
transform 1 0 14706 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_147
timestamp 1607194113
transform 1 0 14062 0 -1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__CLK
timestamp 1607194113
transform 1 0 13786 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1607194113
transform 1 0 14614 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1490_
timestamp 1607194113
transform 1 0 14890 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_75_178
timestamp 1607194113
transform 1 0 16914 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_170
timestamp 1607194113
transform 1 0 16178 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_177
timestamp 1607194113
transform 1 0 16822 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__CLK
timestamp 1607194113
transform 1 0 16638 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__CLK
timestamp 1607194113
transform 1 0 17190 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__CLK
timestamp 1607194113
transform 1 0 17190 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1607194113
transform 1 0 17374 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1492_
timestamp 1607194113
transform 1 0 17466 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1491_
timestamp 1607194113
transform 1 0 17374 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_215
timestamp 1607194113
transform 1 0 20318 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_203
timestamp 1607194113
transform 1 0 19214 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_215
timestamp 1607194113
transform 1 0 20318 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_202
timestamp 1607194113
transform 1 0 19122 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1607194113
transform 1 0 20226 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1607194113
transform 1 0 1918 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1607194113
transform 1 0 814 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1607194113
transform 1 0 538 0 -1 41936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1607194113
transform 1 0 3482 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1607194113
transform 1 0 3022 0 -1 41936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1607194113
transform 1 0 3390 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_56
timestamp 1607194113
transform 1 0 5690 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1607194113
transform 1 0 4586 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_75
timestamp 1607194113
transform 1 0 7438 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_63
timestamp 1607194113
transform 1 0 6334 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1607194113
transform 1 0 6242 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_94
timestamp 1607194113
transform 1 0 9186 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_87
timestamp 1607194113
transform 1 0 8542 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1607194113
transform 1 0 9094 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_118
timestamp 1607194113
transform 1 0 11394 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_106
timestamp 1607194113
transform 1 0 10290 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_137
timestamp 1607194113
transform 1 0 13142 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_125
timestamp 1607194113
transform 1 0 12038 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1607194113
transform 1 0 11946 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_156
timestamp 1607194113
transform 1 0 14890 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_149
timestamp 1607194113
transform 1 0 14246 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1607194113
transform 1 0 14798 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_168
timestamp 1607194113
transform 1 0 15994 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_187
timestamp 1607194113
transform 1 0 17742 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_180
timestamp 1607194113
transform 1 0 17098 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1607194113
transform 1 0 17650 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_211
timestamp 1607194113
transform 1 0 19950 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_199
timestamp 1607194113
transform 1 0 18846 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1607194113
transform 1 0 20502 0 -1 41936
box -38 -48 130 592
use delayline_9_hd_25_1  inst_tdelay_line
timestamp 1607276668
transform -1 0 32076 0 1 1472
box 800 800 20764 22385
use sky130_fd_sc_hd__decap_12  FILLER_1_368
timestamp 1607194113
transform 1 0 34394 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_368
timestamp 1607194113
transform 1 0 34394 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1607194113
transform 1 0 34118 0 1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1607194113
transform 1 0 34118 0 -1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_392
timestamp 1607194113
transform 1 0 36602 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_380
timestamp 1607194113
transform 1 0 35498 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_392
timestamp 1607194113
transform 1 0 36602 0 -1 592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_380
timestamp 1607194113
transform 1 0 35498 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_404
timestamp 1607194113
transform 1 0 37706 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_409
timestamp 1607194113
transform 1 0 38166 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_397
timestamp 1607194113
transform 1 0 37062 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607194113
transform 1 0 36970 0 -1 592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_427
timestamp 1607194113
transform 1 0 39822 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_424
timestamp 1607194113
transform 1 0 39546 0 1 592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_416
timestamp 1607194113
transform 1 0 38810 0 1 592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_428
timestamp 1607194113
transform 1 0 39914 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_421
timestamp 1607194113
transform 1 0 39270 0 -1 592
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1607194113
transform 1 0 39730 0 1 592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607194113
transform 1 0 39822 0 -1 592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_368
timestamp 1607194113
transform 1 0 34394 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1607194113
transform 1 0 34118 0 -1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_392
timestamp 1607194113
transform 1 0 36602 0 -1 1680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_380
timestamp 1607194113
transform 1 0 35498 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_409
timestamp 1607194113
transform 1 0 38166 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_397
timestamp 1607194113
transform 1 0 37062 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1607194113
transform 1 0 36970 0 -1 1680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1607194113
transform 1 0 40374 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1607194113
transform 1 0 39270 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_368
timestamp 1607194113
transform 1 0 34394 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1607194113
transform 1 0 34118 0 1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_392
timestamp 1607194113
transform 1 0 36602 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_380
timestamp 1607194113
transform 1 0 35498 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_404
timestamp 1607194113
transform 1 0 37706 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_427
timestamp 1607194113
transform 1 0 39822 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_424
timestamp 1607194113
transform 1 0 39546 0 1 1680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_416
timestamp 1607194113
transform 1 0 38810 0 1 1680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1607194113
transform 1 0 39730 0 1 1680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_370
timestamp 1607194113
transform 1 0 34578 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_inp_i
timestamp 1607194113
transform 1 0 34394 0 -1 2768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1607194113
transform 1 0 34118 0 -1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_394
timestamp 1607194113
transform 1 0 36786 0 -1 2768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_382
timestamp 1607194113
transform 1 0 35682 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_409
timestamp 1607194113
transform 1 0 38166 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_397
timestamp 1607194113
transform 1 0 37062 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1607194113
transform 1 0 36970 0 -1 2768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1607194113
transform 1 0 40374 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1607194113
transform 1 0 39270 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_368
timestamp 1607194113
transform 1 0 34394 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1607194113
transform 1 0 34118 0 1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_392
timestamp 1607194113
transform 1 0 36602 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_380
timestamp 1607194113
transform 1 0 35498 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_404
timestamp 1607194113
transform 1 0 37706 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_427
timestamp 1607194113
transform 1 0 39822 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_424
timestamp 1607194113
transform 1 0 39546 0 1 2768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_416
timestamp 1607194113
transform 1 0 38810 0 1 2768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1607194113
transform 1 0 39730 0 1 2768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_368
timestamp 1607194113
transform 1 0 34394 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_368
timestamp 1607194113
transform 1 0 34394 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1607194113
transform 1 0 34118 0 -1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1607194113
transform 1 0 34118 0 1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_392
timestamp 1607194113
transform 1 0 36602 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_380
timestamp 1607194113
transform 1 0 35498 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_392
timestamp 1607194113
transform 1 0 36602 0 -1 3856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_380
timestamp 1607194113
transform 1 0 35498 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_404
timestamp 1607194113
transform 1 0 37706 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_409
timestamp 1607194113
transform 1 0 38166 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_397
timestamp 1607194113
transform 1 0 37062 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1607194113
transform 1 0 36970 0 -1 3856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_427
timestamp 1607194113
transform 1 0 39822 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_424
timestamp 1607194113
transform 1 0 39546 0 1 3856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_416
timestamp 1607194113
transform 1 0 38810 0 1 3856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1607194113
transform 1 0 40374 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1607194113
transform 1 0 39270 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1607194113
transform 1 0 39730 0 1 3856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_368
timestamp 1607194113
transform 1 0 34394 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1607194113
transform 1 0 34118 0 -1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_392
timestamp 1607194113
transform 1 0 36602 0 -1 4944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_380
timestamp 1607194113
transform 1 0 35498 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_409
timestamp 1607194113
transform 1 0 38166 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_397
timestamp 1607194113
transform 1 0 37062 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1607194113
transform 1 0 36970 0 -1 4944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1607194113
transform 1 0 40374 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1607194113
transform 1 0 39270 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_368
timestamp 1607194113
transform 1 0 34394 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1607194113
transform 1 0 34118 0 1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_392
timestamp 1607194113
transform 1 0 36602 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_380
timestamp 1607194113
transform 1 0 35498 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_404
timestamp 1607194113
transform 1 0 37706 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_427
timestamp 1607194113
transform 1 0 39822 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_424
timestamp 1607194113
transform 1 0 39546 0 1 4944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_416
timestamp 1607194113
transform 1 0 38810 0 1 4944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1607194113
transform 1 0 39730 0 1 4944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_368
timestamp 1607194113
transform 1 0 34394 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1607194113
transform 1 0 34118 0 -1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_392
timestamp 1607194113
transform 1 0 36602 0 -1 6032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_380
timestamp 1607194113
transform 1 0 35498 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_409
timestamp 1607194113
transform 1 0 38166 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_397
timestamp 1607194113
transform 1 0 37062 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1607194113
transform 1 0 36970 0 -1 6032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1607194113
transform 1 0 40374 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1607194113
transform 1 0 39270 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_368
timestamp 1607194113
transform 1 0 34394 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1607194113
transform 1 0 34118 0 1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_392
timestamp 1607194113
transform 1 0 36602 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_380
timestamp 1607194113
transform 1 0 35498 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_404
timestamp 1607194113
transform 1 0 37706 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_427
timestamp 1607194113
transform 1 0 39822 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_424
timestamp 1607194113
transform 1 0 39546 0 1 6032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_416
timestamp 1607194113
transform 1 0 38810 0 1 6032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1607194113
transform 1 0 39730 0 1 6032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_368
timestamp 1607194113
transform 1 0 34394 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1607194113
transform 1 0 34118 0 -1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_392
timestamp 1607194113
transform 1 0 36602 0 -1 7120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_380
timestamp 1607194113
transform 1 0 35498 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_409
timestamp 1607194113
transform 1 0 38166 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_397
timestamp 1607194113
transform 1 0 37062 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1607194113
transform 1 0 36970 0 -1 7120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1607194113
transform 1 0 40374 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1607194113
transform 1 0 39270 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_368
timestamp 1607194113
transform 1 0 34394 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_368
timestamp 1607194113
transform 1 0 34394 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1607194113
transform 1 0 34118 0 1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1607194113
transform 1 0 34118 0 -1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_392
timestamp 1607194113
transform 1 0 36602 0 -1 8208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_380
timestamp 1607194113
transform 1 0 35498 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_392
timestamp 1607194113
transform 1 0 36602 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_380
timestamp 1607194113
transform 1 0 35498 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_409
timestamp 1607194113
transform 1 0 38166 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_397
timestamp 1607194113
transform 1 0 37062 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_404
timestamp 1607194113
transform 1 0 37706 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1607194113
transform 1 0 36970 0 -1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1607194113
transform 1 0 40374 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1607194113
transform 1 0 39270 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_427
timestamp 1607194113
transform 1 0 39822 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_424
timestamp 1607194113
transform 1 0 39546 0 1 7120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_416
timestamp 1607194113
transform 1 0 38810 0 1 7120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1607194113
transform 1 0 39730 0 1 7120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_368
timestamp 1607194113
transform 1 0 34394 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1607194113
transform 1 0 34118 0 1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_392
timestamp 1607194113
transform 1 0 36602 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_380
timestamp 1607194113
transform 1 0 35498 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_404
timestamp 1607194113
transform 1 0 37706 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_427
timestamp 1607194113
transform 1 0 39822 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_424
timestamp 1607194113
transform 1 0 39546 0 1 8208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_416
timestamp 1607194113
transform 1 0 38810 0 1 8208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1607194113
transform 1 0 39730 0 1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_368
timestamp 1607194113
transform 1 0 34394 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1607194113
transform 1 0 34118 0 -1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_392
timestamp 1607194113
transform 1 0 36602 0 -1 9296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_380
timestamp 1607194113
transform 1 0 35498 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_409
timestamp 1607194113
transform 1 0 38166 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_397
timestamp 1607194113
transform 1 0 37062 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1607194113
transform 1 0 36970 0 -1 9296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1607194113
transform 1 0 40374 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1607194113
transform 1 0 39270 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_368
timestamp 1607194113
transform 1 0 34394 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1607194113
transform 1 0 34118 0 1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_392
timestamp 1607194113
transform 1 0 36602 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_380
timestamp 1607194113
transform 1 0 35498 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_404
timestamp 1607194113
transform 1 0 37706 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_427
timestamp 1607194113
transform 1 0 39822 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_424
timestamp 1607194113
transform 1 0 39546 0 1 9296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_416
timestamp 1607194113
transform 1 0 38810 0 1 9296
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1607194113
transform 1 0 39730 0 1 9296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_368
timestamp 1607194113
transform 1 0 34394 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1607194113
transform 1 0 34118 0 -1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_392
timestamp 1607194113
transform 1 0 36602 0 -1 10384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_380
timestamp 1607194113
transform 1 0 35498 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_409
timestamp 1607194113
transform 1 0 38166 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_397
timestamp 1607194113
transform 1 0 37062 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1607194113
transform 1 0 36970 0 -1 10384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1607194113
transform 1 0 40374 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1607194113
transform 1 0 39270 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_368
timestamp 1607194113
transform 1 0 34394 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_370
timestamp 1607194113
transform 1 0 34578 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[8]
timestamp 1607194113
transform 1 0 34394 0 1 10384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1607194113
transform 1 0 34118 0 1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1607194113
transform 1 0 34118 0 -1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_392
timestamp 1607194113
transform 1 0 36602 0 -1 11472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_380
timestamp 1607194113
transform 1 0 35498 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_394
timestamp 1607194113
transform 1 0 36786 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_382
timestamp 1607194113
transform 1 0 35682 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_409
timestamp 1607194113
transform 1 0 38166 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_397
timestamp 1607194113
transform 1 0 37062 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_406
timestamp 1607194113
transform 1 0 37890 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1607194113
transform 1 0 36970 0 -1 11472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1607194113
transform 1 0 40374 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1607194113
transform 1 0 39270 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_427
timestamp 1607194113
transform 1 0 39822 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_418
timestamp 1607194113
transform 1 0 38994 0 1 10384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1607194113
transform 1 0 39730 0 1 10384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_368
timestamp 1607194113
transform 1 0 34394 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1607194113
transform 1 0 34118 0 1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_392
timestamp 1607194113
transform 1 0 36602 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_380
timestamp 1607194113
transform 1 0 35498 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_404
timestamp 1607194113
transform 1 0 37706 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_427
timestamp 1607194113
transform 1 0 39822 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_424
timestamp 1607194113
transform 1 0 39546 0 1 11472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_416
timestamp 1607194113
transform 1 0 38810 0 1 11472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1607194113
transform 1 0 39730 0 1 11472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_368
timestamp 1607194113
transform 1 0 34394 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1607194113
transform 1 0 34118 0 -1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_392
timestamp 1607194113
transform 1 0 36602 0 -1 12560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_380
timestamp 1607194113
transform 1 0 35498 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_409
timestamp 1607194113
transform 1 0 38166 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_397
timestamp 1607194113
transform 1 0 37062 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1607194113
transform 1 0 36970 0 -1 12560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1607194113
transform 1 0 40374 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1607194113
transform 1 0 39270 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_368
timestamp 1607194113
transform 1 0 34394 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1607194113
transform 1 0 34118 0 1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_392
timestamp 1607194113
transform 1 0 36602 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_380
timestamp 1607194113
transform 1 0 35498 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_404
timestamp 1607194113
transform 1 0 37706 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_427
timestamp 1607194113
transform 1 0 39822 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_424
timestamp 1607194113
transform 1 0 39546 0 1 12560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_416
timestamp 1607194113
transform 1 0 38810 0 1 12560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1607194113
transform 1 0 39730 0 1 12560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_368
timestamp 1607194113
transform 1 0 34394 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1607194113
transform 1 0 34118 0 -1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_392
timestamp 1607194113
transform 1 0 36602 0 -1 13648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_380
timestamp 1607194113
transform 1 0 35498 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_409
timestamp 1607194113
transform 1 0 38166 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_397
timestamp 1607194113
transform 1 0 37062 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1607194113
transform 1 0 36970 0 -1 13648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1607194113
transform 1 0 40374 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1607194113
transform 1 0 39270 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_368
timestamp 1607194113
transform 1 0 34394 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1607194113
transform 1 0 34118 0 1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_392
timestamp 1607194113
transform 1 0 36602 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_380
timestamp 1607194113
transform 1 0 35498 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_404
timestamp 1607194113
transform 1 0 37706 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_427
timestamp 1607194113
transform 1 0 39822 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_424
timestamp 1607194113
transform 1 0 39546 0 1 13648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_416
timestamp 1607194113
transform 1 0 38810 0 1 13648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1607194113
transform 1 0 39730 0 1 13648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_370
timestamp 1607194113
transform 1 0 34578 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_368
timestamp 1607194113
transform 1 0 34394 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[7]
timestamp 1607194113
transform 1 0 34394 0 1 14736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1607194113
transform 1 0 34118 0 -1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1607194113
transform 1 0 34118 0 1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_394
timestamp 1607194113
transform 1 0 36786 0 1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_382
timestamp 1607194113
transform 1 0 35682 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_392
timestamp 1607194113
transform 1 0 36602 0 -1 14736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_380
timestamp 1607194113
transform 1 0 35498 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_409
timestamp 1607194113
transform 1 0 38166 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_397
timestamp 1607194113
transform 1 0 37062 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__CLK
timestamp 1607194113
transform 1 0 37062 0 1 14736
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1607194113
transform 1 0 36970 0 -1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1411_
timestamp 1607194113
transform 1 0 37246 0 1 14736
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_27_427
timestamp 1607194113
transform 1 0 39822 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_418
timestamp 1607194113
transform 1 0 38994 0 1 14736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1607194113
transform 1 0 40374 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1607194113
transform 1 0 39270 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1607194113
transform 1 0 39730 0 1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_368
timestamp 1607194113
transform 1 0 34394 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1607194113
transform 1 0 34118 0 -1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_392
timestamp 1607194113
transform 1 0 36602 0 -1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_380
timestamp 1607194113
transform 1 0 35498 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__CLK
timestamp 1607194113
transform 1 0 36786 0 -1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1607194113
transform 1 0 36970 0 -1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1410_
timestamp 1607194113
transform 1 0 37062 0 -1 15824
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_28_428
timestamp 1607194113
transform 1 0 39914 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_416
timestamp 1607194113
transform 1 0 38810 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_368
timestamp 1607194113
transform 1 0 34394 0 1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1607194113
transform 1 0 34118 0 1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_388
timestamp 1607194113
transform 1 0 36234 0 1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_380
timestamp 1607194113
transform 1 0 35498 0 1 15824
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B1
timestamp 1607194113
transform 1 0 36326 0 1 15824
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1223_
timestamp 1607194113
transform 1 0 36510 0 1 15824
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_407
timestamp 1607194113
transform 1 0 37982 0 1 15824
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1607194113
transform 1 0 38718 0 1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_427
timestamp 1607194113
transform 1 0 39822 0 1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_418
timestamp 1607194113
transform 1 0 38994 0 1 15824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1607194113
transform 1 0 39730 0 1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_368
timestamp 1607194113
transform 1 0 34394 0 -1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1607194113
transform 1 0 34118 0 -1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_392
timestamp 1607194113
transform 1 0 36602 0 -1 16912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_380
timestamp 1607194113
transform 1 0 35498 0 -1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_405
timestamp 1607194113
transform 1 0 37798 0 -1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_401
timestamp 1607194113
transform 1 0 37430 0 -1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_397
timestamp 1607194113
transform 1 0 37062 0 -1 16912
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1607194113
transform 1 0 36970 0 -1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1607194113
transform 1 0 37522 0 -1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_425
timestamp 1607194113
transform 1 0 39638 0 -1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_417
timestamp 1607194113
transform 1 0 38902 0 -1 16912
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__CLK
timestamp 1607194113
transform 1 0 39822 0 -1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1369_
timestamp 1607194113
transform 1 0 40006 0 -1 16912
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_31_370
timestamp 1607194113
transform 1 0 34578 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[6]
timestamp 1607194113
transform 1 0 34394 0 1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1607194113
transform 1 0 34118 0 1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_382
timestamp 1607194113
transform 1 0 35682 0 1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B1
timestamp 1607194113
transform 1 0 35774 0 1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1224_
timestamp 1607194113
transform 1 0 35958 0 1 16912
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_413
timestamp 1607194113
transform 1 0 38534 0 1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_401
timestamp 1607194113
transform 1 0 37430 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1607194113
transform 1 0 38718 0 1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1607194113
transform 1 0 39178 0 1 16912
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A
timestamp 1607194113
transform 1 0 38994 0 1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__B1
timestamp 1607194113
transform 1 0 39546 0 1 16912
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1607194113
transform 1 0 39730 0 1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1288_
timestamp 1607194113
transform 1 0 39822 0 1 16912
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_368
timestamp 1607194113
transform 1 0 34394 0 -1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1607194113
transform 1 0 34118 0 -1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_392
timestamp 1607194113
transform 1 0 36602 0 -1 18000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_380
timestamp 1607194113
transform 1 0 35498 0 -1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_409
timestamp 1607194113
transform 1 0 38166 0 -1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_397
timestamp 1607194113
transform 1 0 37062 0 -1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__B1
timestamp 1607194113
transform 1 0 38258 0 -1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1607194113
transform 1 0 36970 0 -1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1286_
timestamp 1607194113
transform 1 0 38442 0 -1 18000
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_32_428
timestamp 1607194113
transform 1 0 39914 0 -1 18000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_370
timestamp 1607194113
transform 1 0 34578 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[5]
timestamp 1607194113
transform 1 0 34394 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1607194113
transform 1 0 34118 0 1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1607194113
transform 1 0 34118 0 -1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1408_
timestamp 1607194113
transform 1 0 34762 0 1 18000
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1227_
timestamp 1607194113
transform 1 0 34394 0 -1 19088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_34_384
timestamp 1607194113
transform 1 0 35866 0 -1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1607194113
transform 1 0 36694 0 1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__CLK
timestamp 1607194113
transform 1 0 36510 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_409
timestamp 1607194113
transform 1 0 38166 0 -1 19088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_397
timestamp 1607194113
transform 1 0 37062 0 -1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1607194113
transform 1 0 37798 0 1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1607194113
transform 1 0 36970 0 -1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_431
timestamp 1607194113
transform 1 0 40190 0 1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_427
timestamp 1607194113
transform 1 0 39822 0 1 18000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_425
timestamp 1607194113
transform 1 0 39638 0 1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_417
timestamp 1607194113
transform 1 0 38902 0 1 18000
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__CLK
timestamp 1607194113
transform 1 0 38902 0 -1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__CLK
timestamp 1607194113
transform 1 0 40282 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1607194113
transform 1 0 39730 0 1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1409_
timestamp 1607194113
transform 1 0 39086 0 -1 19088
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1370_
timestamp 1607194113
transform 1 0 40466 0 1 18000
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_35_372
timestamp 1607194113
transform 1 0 34762 0 1 19088
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[4]
timestamp 1607194113
transform 1 0 34394 0 1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B1
timestamp 1607194113
transform 1 0 34578 0 1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1607194113
transform 1 0 34118 0 1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_394
timestamp 1607194113
transform 1 0 36786 0 1 19088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_382
timestamp 1607194113
transform 1 0 35682 0 1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_378
timestamp 1607194113
transform 1 0 35314 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1607194113
transform 1 0 35406 0 1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_398
timestamp 1607194113
transform 1 0 37154 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B1
timestamp 1607194113
transform 1 0 37246 0 1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1226_
timestamp 1607194113
transform 1 0 37430 0 1 19088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_430
timestamp 1607194113
transform 1 0 40098 0 1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_425
timestamp 1607194113
transform 1 0 39638 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_419
timestamp 1607194113
transform 1 0 39086 0 1 19088
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A1_N
timestamp 1607194113
transform 1 0 38902 0 1 19088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1607194113
transform 1 0 39730 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1607194113
transform 1 0 39822 0 1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_368
timestamp 1607194113
transform 1 0 34394 0 -1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1607194113
transform 1 0 34118 0 -1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_392
timestamp 1607194113
transform 1 0 36602 0 -1 20176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_380
timestamp 1607194113
transform 1 0 35498 0 -1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_409
timestamp 1607194113
transform 1 0 38166 0 -1 20176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_397
timestamp 1607194113
transform 1 0 37062 0 -1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1607194113
transform 1 0 36970 0 -1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_417
timestamp 1607194113
transform 1 0 38902 0 -1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__B1
timestamp 1607194113
transform 1 0 38994 0 -1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1228_
timestamp 1607194113
transform 1 0 39178 0 -1 20176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_37_370
timestamp 1607194113
transform 1 0 34578 0 1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[3]
timestamp 1607194113
transform 1 0 34394 0 1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1607194113
transform 1 0 34118 0 1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_392
timestamp 1607194113
transform 1 0 36602 0 1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_382
timestamp 1607194113
transform 1 0 35682 0 1 20176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A
timestamp 1607194113
transform 1 0 36050 0 1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1222_
timestamp 1607194113
transform 1 0 36234 0 1 20176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_404
timestamp 1607194113
transform 1 0 37706 0 1 20176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_433
timestamp 1607194113
transform 1 0 40374 0 1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_427
timestamp 1607194113
transform 1 0 39822 0 1 20176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_424
timestamp 1607194113
transform 1 0 39546 0 1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_416
timestamp 1607194113
transform 1 0 38810 0 1 20176
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__CLK
timestamp 1607194113
transform 1 0 40466 0 1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1607194113
transform 1 0 39730 0 1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__B1
timestamp 1607194113
transform 1 0 34394 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1607194113
transform 1 0 34118 0 -1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1293_
timestamp 1607194113
transform 1 0 34578 0 -1 21264
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_38_394
timestamp 1607194113
transform 1 0 36786 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_386
timestamp 1607194113
transform 1 0 36050 0 -1 21264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_401
timestamp 1607194113
transform 1 0 37430 0 -1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_397
timestamp 1607194113
transform 1 0 37062 0 -1 21264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__B1
timestamp 1607194113
transform 1 0 37522 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1607194113
transform 1 0 36970 0 -1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1291_
timestamp 1607194113
transform 1 0 37706 0 -1 21264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_38_420
timestamp 1607194113
transform 1 0 39178 0 -1 21264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__CLK
timestamp 1607194113
transform 1 0 39730 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1368_
timestamp 1607194113
transform 1 0 39914 0 -1 21264
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_40_368
timestamp 1607194113
transform 1 0 34394 0 -1 22352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[2]
timestamp 1607194113
transform 1 0 34762 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1607194113
transform 1 0 34946 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1607194113
transform 1 0 34118 0 1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1607194113
transform 1 0 34118 0 -1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1225_
timestamp 1607194113
transform 1 0 34394 0 1 21264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_395
timestamp 1607194113
transform 1 0 36878 0 -1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_383
timestamp 1607194113
transform 1 0 35774 0 -1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_376
timestamp 1607194113
transform 1 0 35130 0 -1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_376
timestamp 1607194113
transform 1 0 35130 0 1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__CLK
timestamp 1607194113
transform 1 0 35406 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A
timestamp 1607194113
transform 1 0 35590 0 -1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1367_
timestamp 1607194113
transform 1 0 35590 0 1 21264
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1292_
timestamp 1607194113
transform 1 0 35314 0 -1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_409
timestamp 1607194113
transform 1 0 38166 0 -1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_397
timestamp 1607194113
transform 1 0 37062 0 -1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_412
timestamp 1607194113
transform 1 0 38442 0 1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_400
timestamp 1607194113
transform 1 0 37338 0 1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1607194113
transform 1 0 36970 0 -1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_421
timestamp 1607194113
transform 1 0 39270 0 -1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_432
timestamp 1607194113
transform 1 0 40282 0 1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_424
timestamp 1607194113
transform 1 0 39546 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A
timestamp 1607194113
transform 1 0 40098 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__B1
timestamp 1607194113
transform 1 0 39546 0 -1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1607194113
transform 1 0 39730 0 1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1295_
timestamp 1607194113
transform 1 0 39730 0 -1 22352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 1607194113
transform 1 0 39822 0 1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[1]
timestamp 1607194113
transform 1 0 34762 0 1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A
timestamp 1607194113
transform 1 0 34946 0 1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1607194113
transform 1 0 34118 0 1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1221_
timestamp 1607194113
transform 1 0 34394 0 1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_388
timestamp 1607194113
transform 1 0 36234 0 1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_376
timestamp 1607194113
transform 1 0 35130 0 1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_406
timestamp 1607194113
transform 1 0 37890 0 1 22352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1607194113
transform 1 0 37338 0 1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1285_
timestamp 1607194113
transform 1 0 37522 0 1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1607194113
transform 1 0 38626 0 1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_433
timestamp 1607194113
transform 1 0 40374 0 1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_427
timestamp 1607194113
transform 1 0 39822 0 1 22352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_425
timestamp 1607194113
transform 1 0 39638 0 1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_417
timestamp 1607194113
transform 1 0 38902 0 1 22352
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__CLK
timestamp 1607194113
transform 1 0 40466 0 1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1607194113
transform 1 0 39730 0 1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_tdelay_line_en_i[0]
timestamp 1607194113
transform 1 0 34762 0 -1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A
timestamp 1607194113
transform 1 0 34946 0 -1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1607194113
transform 1 0 34118 0 -1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1290_
timestamp 1607194113
transform 1 0 34394 0 -1 23440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_388
timestamp 1607194113
transform 1 0 36234 0 -1 23440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_376
timestamp 1607194113
transform 1 0 35130 0 -1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_403
timestamp 1607194113
transform 1 0 37614 0 -1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_397
timestamp 1607194113
transform 1 0 37062 0 -1 23440
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__CLK
timestamp 1607194113
transform 1 0 37706 0 -1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1607194113
transform 1 0 36970 0 -1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1362_
timestamp 1607194113
transform 1 0 37890 0 -1 23440
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_433
timestamp 1607194113
transform 1 0 40374 0 -1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_425
timestamp 1607194113
transform 1 0 39638 0 -1 23440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1607194113
transform 1 0 40466 0 -1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_368
timestamp 1607194113
transform 1 0 34394 0 1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A2_N
timestamp 1607194113
transform 1 0 34486 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__B2
timestamp 1607194113
transform 1 0 34670 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__B1
timestamp 1607194113
transform 1 0 34854 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1607194113
transform 1 0 34118 0 1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1233_
timestamp 1607194113
transform 1 0 35038 0 1 23440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_393
timestamp 1607194113
transform 1 0 36694 0 1 23440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1_N
timestamp 1607194113
transform 1 0 36510 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__CLK
timestamp 1607194113
transform 1 0 37062 0 1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1403_
timestamp 1607194113
transform 1 0 37246 0 1 23440
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_43_427
timestamp 1607194113
transform 1 0 39822 0 1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_418
timestamp 1607194113
transform 1 0 38994 0 1 23440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1607194113
transform 1 0 39730 0 1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_368
timestamp 1607194113
transform 1 0 34394 0 -1 24528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1607194113
transform 1 0 34118 0 -1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_395
timestamp 1607194113
transform 1 0 36878 0 -1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_391
timestamp 1607194113
transform 1 0 36510 0 -1 24528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_379
timestamp 1607194113
transform 1 0 35406 0 -1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk_i
timestamp 1607194113
transform 1 0 35130 0 -1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_414
timestamp 1607194113
transform 1 0 38626 0 -1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_402
timestamp 1607194113
transform 1 0 37522 0 -1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A
timestamp 1607194113
transform 1 0 37338 0 -1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1607194113
transform 1 0 36970 0 -1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1607194113
transform 1 0 37062 0 -1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_426
timestamp 1607194113
transform 1 0 39730 0 -1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_368
timestamp 1607194113
transform 1 0 34394 0 1 24528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_i_A
timestamp 1607194113
transform 1 0 34946 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1607194113
transform 1 0 34118 0 1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_379
timestamp 1607194113
transform 1 0 35406 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A2_N
timestamp 1607194113
transform 1 0 35590 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__B2
timestamp 1607194113
transform 1 0 35774 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__B1
timestamp 1607194113
transform 1 0 35958 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk_i
timestamp 1607194113
transform 1 0 35130 0 1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1304_
timestamp 1607194113
transform 1 0 36142 0 1 24528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_45_415
timestamp 1607194113
transform 1 0 38718 0 1 24528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_403
timestamp 1607194113
transform 1 0 37614 0 1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_433
timestamp 1607194113
transform 1 0 40374 0 1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_427
timestamp 1607194113
transform 1 0 39822 0 1 24528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_45_423
timestamp 1607194113
transform 1 0 39454 0 1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__CLK
timestamp 1607194113
transform 1 0 40466 0 1 24528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1607194113
transform 1 0 39730 0 1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_370
timestamp 1607194113
transform 1 0 34578 0 -1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__CLK
timestamp 1607194113
transform 1 0 34394 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1607194113
transform 1 0 34118 0 -1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1607194113
transform 1 0 34118 0 1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1417_
timestamp 1607194113
transform 1 0 34394 0 1 25616
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_47_387
timestamp 1607194113
transform 1 0 36142 0 1 25616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_394
timestamp 1607194113
transform 1 0 36786 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_382
timestamp 1607194113
transform 1 0 35682 0 -1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__B2
timestamp 1607194113
transform 1 0 36510 0 1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A2
timestamp 1607194113
transform 1 0 36694 0 1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0954_
timestamp 1607194113
transform 1 0 36878 0 1 25616
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_47_409
timestamp 1607194113
transform 1 0 38166 0 1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_397
timestamp 1607194113
transform 1 0 37062 0 -1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A2_N
timestamp 1607194113
transform 1 0 37338 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B2
timestamp 1607194113
transform 1 0 37522 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B1
timestamp 1607194113
transform 1 0 37706 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1607194113
transform 1 0 36970 0 -1 25616
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1209_
timestamp 1607194113
transform 1 0 37890 0 -1 25616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_427
timestamp 1607194113
transform 1 0 39822 0 1 25616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_425
timestamp 1607194113
transform 1 0 39638 0 1 25616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_421
timestamp 1607194113
transform 1 0 39270 0 1 25616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_422
timestamp 1607194113
transform 1 0 39362 0 -1 25616
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__CLK
timestamp 1607194113
transform 1 0 39914 0 -1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1607194113
transform 1 0 39730 0 1 25616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1420_
timestamp 1607194113
transform 1 0 40098 0 -1 25616
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1607194113
transform 1 0 34118 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1213_
timestamp 1607194113
transform 1 0 34394 0 -1 26704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_48_394
timestamp 1607194113
transform 1 0 36786 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_386
timestamp 1607194113
transform 1 0 36050 0 -1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A1_N
timestamp 1607194113
transform 1 0 35866 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_400
timestamp 1607194113
transform 1 0 37338 0 -1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A2_N
timestamp 1607194113
transform 1 0 38074 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B2
timestamp 1607194113
transform 1 0 38258 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B1
timestamp 1607194113
transform 1 0 38442 0 -1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1607194113
transform 1 0 36970 0 -1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1210_
timestamp 1607194113
transform 1 0 38626 0 -1 26704
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1607194113
transform 1 0 37062 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_430
timestamp 1607194113
transform 1 0 40098 0 -1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_235
timestamp 1607194113
transform 1 0 22158 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_223
timestamp 1607194113
transform 1 0 21054 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A
timestamp 1607194113
transform 1 0 20870 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_245
timestamp 1607194113
transform 1 0 23078 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_241
timestamp 1607194113
transform 1 0 22710 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B2
timestamp 1607194113
transform 1 0 22802 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607194113
transform 1 0 22986 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0988_
timestamp 1607194113
transform 1 0 23170 0 1 26704
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_49_273
timestamp 1607194113
transform 1 0 25654 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_262
timestamp 1607194113
transform 1 0 24642 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1607194113
transform 1 0 25470 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B1
timestamp 1607194113
transform 1 0 24458 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1607194113
transform 1 0 25194 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_293
timestamp 1607194113
transform 1 0 27494 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_285
timestamp 1607194113
transform 1 0 26758 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1607194113
transform 1 0 27586 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_306
timestamp 1607194113
transform 1 0 28690 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_299
timestamp 1607194113
transform 1 0 28046 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1607194113
transform 1 0 27862 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A2
timestamp 1607194113
transform 1 0 29058 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B2
timestamp 1607194113
transform 1 0 29242 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607194113
transform 1 0 28598 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0980_
timestamp 1607194113
transform 1 0 29426 0 1 26704
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_49_330
timestamp 1607194113
transform 1 0 30898 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1607194113
transform 1 0 30714 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1607194113
transform 1 0 31450 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_351
timestamp 1607194113
transform 1 0 32830 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_339
timestamp 1607194113
transform 1 0 31726 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk_i
timestamp 1607194113
transform 1 0 33014 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_369
timestamp 1607194113
transform 1 0 34486 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_356
timestamp 1607194113
transform 1 0 33290 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A2_N
timestamp 1607194113
transform 1 0 33842 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__B2
timestamp 1607194113
transform 1 0 34026 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__B1
timestamp 1607194113
transform 1 0 34302 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607194113
transform 1 0 34210 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_377
timestamp 1607194113
transform 1 0 35222 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A2
timestamp 1607194113
transform 1 0 35498 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__B2
timestamp 1607194113
transform 1 0 35682 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0966_
timestamp 1607194113
transform 1 0 35866 0 1 26704
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_49_410
timestamp 1607194113
transform 1 0 38258 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_398
timestamp 1607194113
transform 1 0 37154 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_428
timestamp 1607194113
transform 1 0 39914 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_426
timestamp 1607194113
transform 1 0 39730 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_422
timestamp 1607194113
transform 1 0 39362 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607194113
transform 1 0 39822 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1607194113
transform 1 0 21422 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_242
timestamp 1607194113
transform 1 0 22802 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B1
timestamp 1607194113
transform 1 0 23354 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1215_
timestamp 1607194113
transform 1 0 23538 0 -1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1607194113
transform 1 0 22526 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_276
timestamp 1607194113
transform 1 0 25930 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_274
timestamp 1607194113
transform 1 0 25746 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_270
timestamp 1607194113
transform 1 0 25378 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B2
timestamp 1607194113
transform 1 0 25194 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A2_N
timestamp 1607194113
transform 1 0 25010 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607194113
transform 1 0 25838 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1405_
timestamp 1607194113
transform 1 0 27034 0 -1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1607194113
transform 1 0 28966 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__CLK
timestamp 1607194113
transform 1 0 28782 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_328
timestamp 1607194113
transform 1 0 30714 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_321
timestamp 1607194113
transform 1 0 30070 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607194113
transform 1 0 31450 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1607194113
transform 1 0 30438 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_337
timestamp 1607194113
transform 1 0 31542 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A2
timestamp 1607194113
transform 1 0 31634 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B2
timestamp 1607194113
transform 1 0 31818 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0973_
timestamp 1607194113
transform 1 0 32002 0 -1 27792
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_50_370
timestamp 1607194113
transform 1 0 34578 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_358
timestamp 1607194113
transform 1 0 33474 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B1
timestamp 1607194113
transform 1 0 33290 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_388
timestamp 1607194113
transform 1 0 36234 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_382
timestamp 1607194113
transform 1 0 35682 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_i_A
timestamp 1607194113
transform 1 0 36050 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk_i
timestamp 1607194113
transform 1 0 35774 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_398
timestamp 1607194113
transform 1 0 37154 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_396
timestamp 1607194113
transform 1 0 36970 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__CLK
timestamp 1607194113
transform 1 0 37706 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607194113
transform 1 0 37062 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1459_
timestamp 1607194113
transform 1 0 37890 0 -1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_427
timestamp 1607194113
transform 1 0 39822 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__D
timestamp 1607194113
transform 1 0 39638 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_232
timestamp 1607194113
transform 1 0 21882 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_220
timestamp 1607194113
transform 1 0 20778 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1607194113
transform 1 0 21698 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__B
timestamp 1607194113
transform 1 0 20870 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1018_
timestamp 1607194113
transform 1 0 21054 0 1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_51_249
timestamp 1607194113
transform 1 0 23446 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__CLK
timestamp 1607194113
transform 1 0 23998 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607194113
transform 1 0 22986 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0953_
timestamp 1607194113
transform 1 0 23078 0 1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_276
timestamp 1607194113
transform 1 0 25930 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1416_
timestamp 1607194113
transform 1 0 24182 0 1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_51_288
timestamp 1607194113
transform 1 0 27034 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1607194113
transform 1 0 27586 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_314
timestamp 1607194113
transform 1 0 29426 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_306
timestamp 1607194113
transform 1 0 28690 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_297
timestamp 1607194113
transform 1 0 27862 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B1
timestamp 1607194113
transform 1 0 29518 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607194113
transform 1 0 28598 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1607194113
transform 1 0 31450 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A2
timestamp 1607194113
transform 1 0 29702 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _0968_
timestamp 1607194113
transform 1 0 29886 0 1 27792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_51_350
timestamp 1607194113
transform 1 0 32738 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_338
timestamp 1607194113
transform 1 0 31634 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_365
timestamp 1607194113
transform 1 0 34118 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_358
timestamp 1607194113
transform 1 0 33474 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A2_N
timestamp 1607194113
transform 1 0 33750 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B2
timestamp 1607194113
transform 1 0 33934 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607194113
transform 1 0 34210 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1212_
timestamp 1607194113
transform 1 0 34302 0 1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_51_394
timestamp 1607194113
transform 1 0 36786 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_383
timestamp 1607194113
transform 1 0 35774 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1607194113
transform 1 0 36510 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_406
timestamp 1607194113
transform 1 0 37890 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_428
timestamp 1607194113
transform 1 0 39914 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_426
timestamp 1607194113
transform 1 0 39730 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_418
timestamp 1607194113
transform 1 0 38994 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B1
timestamp 1607194113
transform 1 0 40190 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1_N
timestamp 1607194113
transform 1 0 40374 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607194113
transform 1 0 39822 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_228
timestamp 1607194113
transform 1 0 21514 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1607194113
transform 1 0 21422 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_245
timestamp 1607194113
transform 1 0 23078 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_240
timestamp 1607194113
transform 1 0 22618 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_239
timestamp 1607194113
transform 1 0 22526 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B
timestamp 1607194113
transform 1 0 22802 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B1
timestamp 1607194113
transform 1 0 22710 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1607194113
transform 1 0 22894 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607194113
transform 1 0 22986 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0985_
timestamp 1607194113
transform 1 0 23170 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_53_255
timestamp 1607194113
transform 1 0 23998 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1607194113
transform 1 0 23814 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _0990_
timestamp 1607194113
transform 1 0 23078 0 -1 28880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1607194113
transform 1 0 24918 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_276
timestamp 1607194113
transform 1 0 25930 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_264
timestamp 1607194113
transform 1 0 24826 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_i_A
timestamp 1607194113
transform 1 0 25654 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1607194113
transform 1 0 24642 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A
timestamp 1607194113
transform 1 0 24366 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk_i
timestamp 1607194113
transform 1 0 25378 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607194113
transform 1 0 25838 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1214_
timestamp 1607194113
transform 1 0 24550 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_289
timestamp 1607194113
transform 1 0 27126 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_277
timestamp 1607194113
transform 1 0 26022 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B1
timestamp 1607194113
transform 1 0 26298 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A2
timestamp 1607194113
transform 1 0 26482 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _0982_
timestamp 1607194113
transform 1 0 26666 0 -1 28880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_53_301
timestamp 1607194113
transform 1 0 28230 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_303
timestamp 1607194113
transform 1 0 28414 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1
timestamp 1607194113
transform 1 0 28230 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1607194113
transform 1 0 28690 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B
timestamp 1607194113
transform 1 0 28874 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A2
timestamp 1607194113
transform 1 0 28966 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607194113
transform 1 0 28598 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0963_
timestamp 1607194113
transform 1 0 29058 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0956_
timestamp 1607194113
transform 1 0 29150 0 -1 28880
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_53_317
timestamp 1607194113
transform 1 0 29702 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_335
timestamp 1607194113
transform 1 0 31358 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_327
timestamp 1607194113
transform 1 0 30622 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A1
timestamp 1607194113
transform 1 0 30438 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B1
timestamp 1607194113
transform 1 0 30070 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A2
timestamp 1607194113
transform 1 0 30254 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607194113
transform 1 0 31450 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0975_
timestamp 1607194113
transform 1 0 30438 0 1 28880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_53_344
timestamp 1607194113
transform 1 0 32186 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_352
timestamp 1607194113
transform 1 0 32922 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_340
timestamp 1607194113
transform 1 0 31818 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1607194113
transform 1 0 32002 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1607194113
transform 1 0 31542 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1607194113
transform 1 0 34302 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_364
timestamp 1607194113
transform 1 0 34026 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_356
timestamp 1607194113
transform 1 0 33290 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_364
timestamp 1607194113
transform 1 0 34026 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__CLK
timestamp 1607194113
transform 1 0 34302 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B1
timestamp 1607194113
transform 1 0 34118 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607194113
transform 1 0 34210 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1418_
timestamp 1607194113
transform 1 0 34486 0 -1 28880
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_53_387
timestamp 1607194113
transform 1 0 36142 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_379
timestamp 1607194113
transform 1 0 35406 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_388
timestamp 1607194113
transform 1 0 36234 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1_N
timestamp 1607194113
transform 1 0 36326 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0784_
timestamp 1607194113
transform 1 0 36510 0 1 28880
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_52_396
timestamp 1607194113
transform 1 0 36970 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607194113
transform 1 0 37062 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_411
timestamp 1607194113
transform 1 0 38350 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_410
timestamp 1607194113
transform 1 0 38258 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A1_N
timestamp 1607194113
transform 1 0 38350 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2_N
timestamp 1607194113
transform 1 0 38166 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B2
timestamp 1607194113
transform 1 0 37982 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1607194113
transform 1 0 38718 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_398
timestamp 1607194113
transform 1 0 37154 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _0741_
timestamp 1607194113
transform 1 0 38534 0 -1 28880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_428
timestamp 1607194113
transform 1 0 39914 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_426
timestamp 1607194113
transform 1 0 39730 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_418
timestamp 1607194113
transform 1 0 38994 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_429
timestamp 1607194113
transform 1 0 40006 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607194113
transform 1 0 39822 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_227
timestamp 1607194113
transform 1 0 21422 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_255
timestamp 1607194113
transform 1 0 23998 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_239
timestamp 1607194113
transform 1 0 22526 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__B
timestamp 1607194113
transform 1 0 22802 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1607194113
transform 1 0 23814 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1172_
timestamp 1607194113
transform 1 0 22986 0 -1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_54_276
timestamp 1607194113
transform 1 0 25930 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_267
timestamp 1607194113
transform 1 0 25102 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607194113
transform 1 0 25838 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_284
timestamp 1607194113
transform 1 0 26666 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A1
timestamp 1607194113
transform 1 0 26942 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A2
timestamp 1607194113
transform 1 0 27126 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A3
timestamp 1607194113
transform 1 0 27310 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1273_
timestamp 1607194113
transform 1 0 27494 0 -1 29968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_54_312
timestamp 1607194113
transform 1 0 29242 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B1
timestamp 1607194113
transform 1 0 29058 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__B
timestamp 1607194113
transform 1 0 29610 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_335
timestamp 1607194113
transform 1 0 31358 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_327
timestamp 1607194113
transform 1 0 30622 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1607194113
transform 1 0 30438 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607194113
transform 1 0 31450 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0947_
timestamp 1607194113
transform 1 0 29794 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_54_346
timestamp 1607194113
transform 1 0 32370 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__B
timestamp 1607194113
transform 1 0 32186 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0971_
timestamp 1607194113
transform 1 0 31542 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_54_367
timestamp 1607194113
transform 1 0 34302 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_358
timestamp 1607194113
transform 1 0 33474 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A
timestamp 1607194113
transform 1 0 34118 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1211_
timestamp 1607194113
transform 1 0 33750 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_391
timestamp 1607194113
transform 1 0 36510 0 -1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_379
timestamp 1607194113
transform 1 0 35406 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_410
timestamp 1607194113
transform 1 0 38258 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_402
timestamp 1607194113
transform 1 0 37522 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_398
timestamp 1607194113
transform 1 0 37154 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A1_N
timestamp 1607194113
transform 1 0 38350 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607194113
transform 1 0 37062 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0826_
timestamp 1607194113
transform 1 0 38534 0 -1 29968
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1607194113
transform 1 0 37246 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_429
timestamp 1607194113
transform 1 0 40006 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_236
timestamp 1607194113
transform 1 0 22250 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1607194113
transform 1 0 21882 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_220
timestamp 1607194113
transform 1 0 20778 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_243
timestamp 1607194113
transform 1 0 22894 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1607194113
transform 1 0 22342 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A2
timestamp 1607194113
transform 1 0 22710 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A3
timestamp 1607194113
transform 1 0 22526 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607194113
transform 1 0 22986 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1276_
timestamp 1607194113
transform 1 0 23078 0 1 29968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_55_276
timestamp 1607194113
transform 1 0 25930 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_264
timestamp 1607194113
transform 1 0 24826 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__B1
timestamp 1607194113
transform 1 0 24642 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_296
timestamp 1607194113
transform 1 0 27770 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_284
timestamp 1607194113
transform 1 0 26666 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B
timestamp 1607194113
transform 1 0 26942 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0978_
timestamp 1607194113
transform 1 0 27126 0 1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_55_306
timestamp 1607194113
transform 1 0 28690 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_304
timestamp 1607194113
transform 1 0 28506 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607194113
transform 1 0 28598 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_330
timestamp 1607194113
transform 1 0 30898 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_318
timestamp 1607194113
transform 1 0 29794 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_354
timestamp 1607194113
transform 1 0 33106 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_342
timestamp 1607194113
transform 1 0 32002 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_370
timestamp 1607194113
transform 1 0 34578 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607194113
transform 1 0 34210 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1607194113
transform 1 0 34302 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_390
timestamp 1607194113
transform 1 0 36418 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1607194113
transform 1 0 35682 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1_N
timestamp 1607194113
transform 1 0 36694 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0855_
timestamp 1607194113
transform 1 0 36878 0 1 29968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_415
timestamp 1607194113
transform 1 0 38718 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2_N
timestamp 1607194113
transform 1 0 38534 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B2
timestamp 1607194113
transform 1 0 38350 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_428
timestamp 1607194113
transform 1 0 39914 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607194113
transform 1 0 39822 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_231
timestamp 1607194113
transform 1 0 21790 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_227
timestamp 1607194113
transform 1 0 21422 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__CLK
timestamp 1607194113
transform 1 0 21882 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1375_
timestamp 1607194113
transform 1 0 22066 0 -1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1607194113
transform 1 0 23814 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_276
timestamp 1607194113
transform 1 0 25930 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_273
timestamp 1607194113
transform 1 0 25654 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_265
timestamp 1607194113
transform 1 0 24918 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607194113
transform 1 0 25838 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_288
timestamp 1607194113
transform 1 0 27034 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1378_
timestamp 1607194113
transform 1 0 27310 0 -1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_312
timestamp 1607194113
transform 1 0 29242 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__CLK
timestamp 1607194113
transform 1 0 29058 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_324
timestamp 1607194113
transform 1 0 30346 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607194113
transform 1 0 31450 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_337
timestamp 1607194113
transform 1 0 31542 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1376_
timestamp 1607194113
transform 1 0 32646 0 -1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_370
timestamp 1607194113
transform 1 0 34578 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__CLK
timestamp 1607194113
transform 1 0 34394 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 1607194113
transform 1 0 34946 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_392
timestamp 1607194113
transform 1 0 36602 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_380
timestamp 1607194113
transform 1 0 35498 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__CLK
timestamp 1607194113
transform 1 0 36878 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1182_
timestamp 1607194113
transform 1 0 35130 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607194113
transform 1 0 37062 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1377_
timestamp 1607194113
transform 1 0 37154 0 -1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_429
timestamp 1607194113
transform 1 0 40006 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_417
timestamp 1607194113
transform 1 0 38902 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_236
timestamp 1607194113
transform 1 0 22250 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_232
timestamp 1607194113
transform 1 0 21882 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_224
timestamp 1607194113
transform 1 0 21146 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1607194113
transform 1 0 21974 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_245
timestamp 1607194113
transform 1 0 23078 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 1607194113
transform 1 0 22802 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607194113
transform 1 0 22986 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1016_
timestamp 1607194113
transform 1 0 23170 0 1 31056
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_57_274
timestamp 1607194113
transform 1 0 25746 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_262
timestamp 1607194113
transform 1 0 24642 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A1
timestamp 1607194113
transform 1 0 24458 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_287
timestamp 1607194113
transform 1 0 26942 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A
timestamp 1607194113
transform 1 0 26758 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1607194113
transform 1 0 26482 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_299
timestamp 1607194113
transform 1 0 28046 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607194113
transform 1 0 28598 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1379_
timestamp 1607194113
transform 1 0 28690 0 1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_327
timestamp 1607194113
transform 1 0 30622 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__CLK
timestamp 1607194113
transform 1 0 30438 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_339
timestamp 1607194113
transform 1 0 31726 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B1
timestamp 1607194113
transform 1 0 31818 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1275_
timestamp 1607194113
transform 1 0 32002 0 1 31056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1607194113
transform 1 0 34302 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_360
timestamp 1607194113
transform 1 0 33658 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A1_N
timestamp 1607194113
transform 1 0 33474 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607194113
transform 1 0 34210 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_379
timestamp 1607194113
transform 1 0 35406 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B1
timestamp 1607194113
transform 1 0 35498 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1274_
timestamp 1607194113
transform 1 0 35682 0 1 31056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_410
timestamp 1607194113
transform 1 0 38258 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_398
timestamp 1607194113
transform 1 0 37154 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_431
timestamp 1607194113
transform 1 0 40190 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_426
timestamp 1607194113
transform 1 0 39730 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_422
timestamp 1607194113
transform 1 0 39362 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607194113
transform 1 0 39822 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1607194113
transform 1 0 39914 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__B
timestamp 1607194113
transform 1 0 21422 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A
timestamp 1607194113
transform 1 0 21606 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1234_
timestamp 1607194113
transform 1 0 21790 0 -1 32144
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_58_250
timestamp 1607194113
transform 1 0 23538 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_238
timestamp 1607194113
transform 1 0 22434 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A
timestamp 1607194113
transform 1 0 23630 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1173_
timestamp 1607194113
transform 1 0 23814 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_276
timestamp 1607194113
transform 1 0 25930 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_269
timestamp 1607194113
transform 1 0 25286 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_257
timestamp 1607194113
transform 1 0 24182 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607194113
transform 1 0 25838 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_289
timestamp 1607194113
transform 1 0 27126 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_281
timestamp 1607194113
transform 1 0 26390 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A1
timestamp 1607194113
transform 1 0 27402 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A2
timestamp 1607194113
transform 1 0 27586 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A3
timestamp 1607194113
transform 1 0 27770 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1607194113
transform 1 0 26114 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__B1
timestamp 1607194113
transform 1 0 29518 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1272_
timestamp 1607194113
transform 1 0 27954 0 -1 32144
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_58_335
timestamp 1607194113
transform 1 0 31358 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_329
timestamp 1607194113
transform 1 0 30806 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_317
timestamp 1607194113
transform 1 0 29702 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607194113
transform 1 0 31450 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1607194113
transform 1 0 32646 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_337
timestamp 1607194113
transform 1 0 31542 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_373
timestamp 1607194113
transform 1 0 34854 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_361
timestamp 1607194113
transform 1 0 33750 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_385
timestamp 1607194113
transform 1 0 35958 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_410
timestamp 1607194113
transform 1 0 38258 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_398
timestamp 1607194113
transform 1 0 37154 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607194113
transform 1 0 37062 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_432
timestamp 1607194113
transform 1 0 40282 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_418
timestamp 1607194113
transform 1 0 38994 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1607194113
transform 1 0 40098 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1128_
timestamp 1607194113
transform 1 0 39270 0 -1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_60_227
timestamp 1607194113
transform 1 0 21422 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_219
timestamp 1607194113
transform 1 0 20686 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_228
timestamp 1607194113
transform 1 0 21514 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1607194113
transform 1 0 21974 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1022_
timestamp 1607194113
transform 1 0 20686 0 1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1014_
timestamp 1607194113
transform 1 0 20778 0 -1 33232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1607194113
transform 1 0 22158 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_250
timestamp 1607194113
transform 1 0 23538 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_238
timestamp 1607194113
transform 1 0 22434 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_245
timestamp 1607194113
transform 1 0 23078 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_240
timestamp 1607194113
transform 1 0 22618 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607194113
transform 1 0 22986 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_262
timestamp 1607194113
transform 1 0 24642 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_265
timestamp 1607194113
transform 1 0 24918 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_257
timestamp 1607194113
transform 1 0 24182 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__CLK
timestamp 1607194113
transform 1 0 25010 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk_i
timestamp 1607194113
transform 1 0 25010 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_271
timestamp 1607194113
transform 1 0 25470 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_i_A
timestamp 1607194113
transform 1 0 25286 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607194113
transform 1 0 25838 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1412_
timestamp 1607194113
transform 1 0 25194 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _0707_
timestamp 1607194113
transform 1 0 25930 0 -1 33232
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1607194113
transform 1 0 27586 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_287
timestamp 1607194113
transform 1 0 26942 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A2
timestamp 1607194113
transform 1 0 27402 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B2
timestamp 1607194113
transform 1 0 27218 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_311
timestamp 1607194113
transform 1 0 29150 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1607194113
transform 1 0 28690 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_306
timestamp 1607194113
transform 1 0 28690 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_299
timestamp 1607194113
transform 1 0 28046 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607194113
transform 1 0 28598 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1607194113
transform 1 0 28874 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_335
timestamp 1607194113
transform 1 0 31358 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_323
timestamp 1607194113
transform 1 0 30254 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_330
timestamp 1607194113
transform 1 0 30898 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_318
timestamp 1607194113
transform 1 0 29794 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607194113
transform 1 0 31450 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_350
timestamp 1607194113
transform 1 0 32738 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_342
timestamp 1607194113
transform 1 0 32002 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1380_
timestamp 1607194113
transform 1 0 31542 0 -1 33232
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1607194113
transform 1 0 33014 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_358
timestamp 1607194113
transform 1 0 33474 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_364
timestamp 1607194113
transform 1 0 34026 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_356
timestamp 1607194113
transform 1 0 33290 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__CLK
timestamp 1607194113
transform 1 0 33842 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__CLK
timestamp 1607194113
transform 1 0 33290 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_373
timestamp 1607194113
transform 1 0 34854 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1607194113
transform 1 0 34670 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607194113
transform 1 0 34210 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1177_
timestamp 1607194113
transform 1 0 34302 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1421_
timestamp 1607194113
transform 1 0 34026 0 -1 33232
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_60_395
timestamp 1607194113
transform 1 0 36878 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_383
timestamp 1607194113
transform 1 0 35774 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_395
timestamp 1607194113
transform 1 0 36878 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_383
timestamp 1607194113
transform 1 0 35774 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A
timestamp 1607194113
transform 1 0 35222 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1207_
timestamp 1607194113
transform 1 0 35406 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_398
timestamp 1607194113
transform 1 0 37154 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_411
timestamp 1607194113
transform 1 0 38350 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_407
timestamp 1607194113
transform 1 0 37982 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__CLK
timestamp 1607194113
transform 1 0 37706 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607194113
transform 1 0 37062 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1464_
timestamp 1607194113
transform 1 0 37890 0 -1 33232
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1126_
timestamp 1607194113
transform 1 0 38442 0 1 32144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_60_425
timestamp 1607194113
transform 1 0 39638 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_428
timestamp 1607194113
transform 1 0 39914 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_419
timestamp 1607194113
transform 1 0 39086 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607194113
transform 1 0 39822 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1129_
timestamp 1607194113
transform 1 0 40374 0 -1 33232
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _1124_
timestamp 1607194113
transform 1 0 40006 0 1 32144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_61_226
timestamp 1607194113
transform 1 0 21330 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_219
timestamp 1607194113
transform 1 0 20686 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1607194113
transform 1 0 20778 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0868_
timestamp 1607194113
transform 1 0 20962 0 1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_249
timestamp 1607194113
transform 1 0 23446 0 1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_245
timestamp 1607194113
transform 1 0 23078 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_238
timestamp 1607194113
transform 1 0 22434 0 1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__B1
timestamp 1607194113
transform 1 0 23998 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607194113
transform 1 0 22986 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1607194113
transform 1 0 23170 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_273
timestamp 1607194113
transform 1 0 25654 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1219_
timestamp 1607194113
transform 1 0 24182 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_61_287
timestamp 1607194113
transform 1 0 26942 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1607194113
transform 1 0 26390 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1174_
timestamp 1607194113
transform 1 0 26574 0 1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_315
timestamp 1607194113
transform 1 0 29518 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_310
timestamp 1607194113
transform 1 0 29058 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_306
timestamp 1607194113
transform 1 0 28690 0 1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_299
timestamp 1607194113
transform 1 0 28046 0 1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1607194113
transform 1 0 28598 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1236_
timestamp 1607194113
transform 1 0 29150 0 1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_326
timestamp 1607194113
transform 1 0 30530 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1271_
timestamp 1607194113
transform 1 0 31266 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1607194113
transform 1 0 30254 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_352
timestamp 1607194113
transform 1 0 32922 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A1_N
timestamp 1607194113
transform 1 0 32738 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1607194113
transform 1 0 34302 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_364
timestamp 1607194113
transform 1 0 34026 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1607194113
transform 1 0 34210 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_394
timestamp 1607194113
transform 1 0 36786 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_382
timestamp 1607194113
transform 1 0 35682 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1607194113
transform 1 0 35406 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_406
timestamp 1607194113
transform 1 0 37890 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_426
timestamp 1607194113
transform 1 0 39730 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_418
timestamp 1607194113
transform 1 0 38994 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1607194113
transform 1 0 39822 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1127_
timestamp 1607194113
transform 1 0 39914 0 1 33232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1607194113
transform 1 0 21422 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__CLK
timestamp 1607194113
transform 1 0 21790 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1371_
timestamp 1607194113
transform 1 0 21974 0 -1 34320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_252
timestamp 1607194113
transform 1 0 23722 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_272
timestamp 1607194113
transform 1 0 25562 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_264
timestamp 1607194113
transform 1 0 24826 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B
timestamp 1607194113
transform 1 0 25654 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1607194113
transform 1 0 25838 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0708_
timestamp 1607194113
transform 1 0 25930 0 -1 34320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_287
timestamp 1607194113
transform 1 0 26942 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__C
timestamp 1607194113
transform 1 0 26758 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_312
timestamp 1607194113
transform 1 0 29242 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1607194113
transform 1 0 28782 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_299
timestamp 1607194113
transform 1 0 28046 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1241_
timestamp 1607194113
transform 1 0 28874 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1607194113
transform 1 0 30346 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1607194113
transform 1 0 31450 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_344
timestamp 1607194113
transform 1 0 32186 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_337
timestamp 1607194113
transform 1 0 31542 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A
timestamp 1607194113
transform 1 0 32002 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1270_
timestamp 1607194113
transform 1 0 31634 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B2
timestamp 1607194113
transform 1 0 34946 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A1_N
timestamp 1607194113
transform 1 0 34762 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1208_
timestamp 1607194113
transform 1 0 33290 0 -1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_388
timestamp 1607194113
transform 1 0 36234 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_376
timestamp 1607194113
transform 1 0 35130 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_410
timestamp 1607194113
transform 1 0 38258 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_398
timestamp 1607194113
transform 1 0 37154 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_396
timestamp 1607194113
transform 1 0 36970 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1607194113
transform 1 0 37062 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_422
timestamp 1607194113
transform 1 0 39362 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0747_
timestamp 1607194113
transform 1 0 39638 0 -1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_228
timestamp 1607194113
transform 1 0 21514 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__B
timestamp 1607194113
transform 1 0 21330 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1607194113
transform 1 0 23078 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_240
timestamp 1607194113
transform 1 0 22618 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1607194113
transform 1 0 22986 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_257
timestamp 1607194113
transform 1 0 24182 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A2
timestamp 1607194113
transform 1 0 25838 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B2
timestamp 1607194113
transform 1 0 25654 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0805_
timestamp 1607194113
transform 1 0 24366 0 1 34320
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_63_292
timestamp 1607194113
transform 1 0 27402 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_277
timestamp 1607194113
transform 1 0 26022 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__C
timestamp 1607194113
transform 1 0 27218 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__B
timestamp 1607194113
transform 1 0 26206 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0806_
timestamp 1607194113
transform 1 0 26390 0 1 34320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_314
timestamp 1607194113
transform 1 0 29426 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_306
timestamp 1607194113
transform 1 0 28690 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_304
timestamp 1607194113
transform 1 0 28506 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A
timestamp 1607194113
transform 1 0 29518 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1607194113
transform 1 0 28598 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_333
timestamp 1607194113
transform 1 0 31174 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_321
timestamp 1607194113
transform 1 0 30070 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1237_
timestamp 1607194113
transform 1 0 29702 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_345
timestamp 1607194113
transform 1 0 32278 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_367
timestamp 1607194113
transform 1 0 34302 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_357
timestamp 1607194113
transform 1 0 33382 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__CLK
timestamp 1607194113
transform 1 0 34578 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk_i
timestamp 1607194113
transform 1 0 33934 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1607194113
transform 1 0 34210 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1422_
timestamp 1607194113
transform 1 0 34762 0 1 34320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1607194113
transform 1 0 36510 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_412
timestamp 1607194113
transform 1 0 38442 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_403
timestamp 1607194113
transform 1 0 37614 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1607194113
transform 1 0 38166 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_424
timestamp 1607194113
transform 1 0 39546 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1607194113
transform 1 0 39822 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0829_
timestamp 1607194113
transform 1 0 39914 0 1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__B1
timestamp 1607194113
transform 1 0 21422 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1281_
timestamp 1607194113
transform 1 0 21606 0 -1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_249
timestamp 1607194113
transform 1 0 23446 0 -1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A2_N
timestamp 1607194113
transform 1 0 23262 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__B2
timestamp 1607194113
transform 1 0 23078 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1267_
timestamp 1607194113
transform 1 0 23814 0 -1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_276
timestamp 1607194113
transform 1 0 25930 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1607194113
transform 1 0 25470 0 -1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_259
timestamp 1607194113
transform 1 0 24366 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A
timestamp 1607194113
transform 1 0 24182 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1607194113
transform 1 0 25838 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_284
timestamp 1607194113
transform 1 0 26666 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B1
timestamp 1607194113
transform 1 0 26850 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1205_
timestamp 1607194113
transform 1 0 27034 0 -1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_304
timestamp 1607194113
transform 1 0 28506 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0695_
timestamp 1607194113
transform 1 0 29242 0 -1 35408
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1607194113
transform 1 0 30714 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__B2
timestamp 1607194113
transform 1 0 30530 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1607194113
transform 1 0 31450 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_353
timestamp 1607194113
transform 1 0 33014 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_349
timestamp 1607194113
transform 1 0 32646 0 -1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1607194113
transform 1 0 31542 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1381_
timestamp 1607194113
transform 1 0 33106 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_64_375
timestamp 1607194113
transform 1 0 35038 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__CLK
timestamp 1607194113
transform 1 0 34854 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_384
timestamp 1607194113
transform 1 0 35866 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1607194113
transform 1 0 35590 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_398
timestamp 1607194113
transform 1 0 37154 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_396
timestamp 1607194113
transform 1 0 36970 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__CLK
timestamp 1607194113
transform 1 0 37338 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1607194113
transform 1 0 37062 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1385_
timestamp 1607194113
transform 1 0 37522 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_432
timestamp 1607194113
transform 1 0 40282 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_421
timestamp 1607194113
transform 1 0 39270 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1607194113
transform 1 0 40006 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_226
timestamp 1607194113
transform 1 0 21330 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__A2
timestamp 1607194113
transform 1 0 21146 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_238
timestamp 1607194113
transform 1 0 22434 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1607194113
transform 1 0 22986 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1382_
timestamp 1607194113
transform 1 0 23078 0 1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_275
timestamp 1607194113
transform 1 0 25838 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_266
timestamp 1607194113
transform 1 0 25010 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__CLK
timestamp 1607194113
transform 1 0 24826 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1607194113
transform 1 0 25562 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_287
timestamp 1607194113
transform 1 0 26942 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_299
timestamp 1607194113
transform 1 0 28046 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1607194113
transform 1 0 28598 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0795_
timestamp 1607194113
transform 1 0 28690 0 1 35408
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_65_334
timestamp 1607194113
transform 1 0 31266 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_322
timestamp 1607194113
transform 1 0 30162 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B2
timestamp 1607194113
transform 1 0 29978 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_340
timestamp 1607194113
transform 1 0 31818 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1269_
timestamp 1607194113
transform 1 0 31910 0 1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1607194113
transform 1 0 34854 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_365
timestamp 1607194113
transform 1 0 34118 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_359
timestamp 1607194113
transform 1 0 33566 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A
timestamp 1607194113
transform 1 0 34670 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A1_N
timestamp 1607194113
transform 1 0 33382 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1607194113
transform 1 0 34210 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1204_
timestamp 1607194113
transform 1 0 34302 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_385
timestamp 1607194113
transform 1 0 35958 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_397
timestamp 1607194113
transform 1 0 37062 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__CLK
timestamp 1607194113
transform 1 0 37154 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1426_
timestamp 1607194113
transform 1 0 37338 0 1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_431
timestamp 1607194113
transform 1 0 40190 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_419
timestamp 1607194113
transform 1 0 39086 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1607194113
transform 1 0 39822 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1607194113
transform 1 0 39914 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_228
timestamp 1607194113
transform 1 0 21514 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_219
timestamp 1607194113
transform 1 0 20686 0 1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_231
timestamp 1607194113
transform 1 0 21790 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_223
timestamp 1607194113
transform 1 0 21054 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1607194113
transform 1 0 21606 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1330_
timestamp 1607194113
transform 1 0 21238 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1607194113
transform 1 0 21330 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_245
timestamp 1607194113
transform 1 0 23078 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_240
timestamp 1607194113
transform 1 0 22618 0 1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_243
timestamp 1607194113
transform 1 0 22894 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B1
timestamp 1607194113
transform 1 0 23078 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1607194113
transform 1 0 22986 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1268_
timestamp 1607194113
transform 1 0 23262 0 -1 36496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_269
timestamp 1607194113
transform 1 0 25286 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_257
timestamp 1607194113
transform 1 0 24182 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_276
timestamp 1607194113
transform 1 0 25930 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_263
timestamp 1607194113
transform 1 0 24734 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1607194113
transform 1 0 25838 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1607194113
transform 1 0 27494 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1607194113
transform 1 0 26390 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_288
timestamp 1607194113
transform 1 0 27034 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1423_
timestamp 1607194113
transform 1 0 27402 0 -1 36496
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_67_309
timestamp 1607194113
transform 1 0 28966 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_313
timestamp 1607194113
transform 1 0 29334 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__CLK
timestamp 1607194113
transform 1 0 29150 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1607194113
transform 1 0 28598 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1607194113
transform 1 0 28690 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_333
timestamp 1607194113
transform 1 0 31174 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_321
timestamp 1607194113
transform 1 0 30070 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_333
timestamp 1607194113
transform 1 0 31174 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_325
timestamp 1607194113
transform 1 0 30438 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1607194113
transform 1 0 31450 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0936_
timestamp 1607194113
transform 1 0 31358 0 1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_67_353
timestamp 1607194113
transform 1 0 33014 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_349
timestamp 1607194113
transform 1 0 32646 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_343
timestamp 1607194113
transform 1 0 32094 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_337
timestamp 1607194113
transform 1 0 31542 0 -1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_i_A
timestamp 1607194113
transform 1 0 32186 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B1
timestamp 1607194113
transform 1 0 32830 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A1
timestamp 1607194113
transform 1 0 32646 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk_i
timestamp 1607194113
transform 1 0 32370 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1206_
timestamp 1607194113
transform 1 0 32738 0 -1 36496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1607194113
transform 1 0 34302 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_365
timestamp 1607194113
transform 1 0 34118 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_368
timestamp 1607194113
transform 1 0 34394 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1_N
timestamp 1607194113
transform 1 0 34210 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1607194113
transform 1 0 34210 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_391
timestamp 1607194113
transform 1 0 36510 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_379
timestamp 1607194113
transform 1 0 35406 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_392
timestamp 1607194113
transform 1 0 36602 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_380
timestamp 1607194113
transform 1 0 35498 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_399
timestamp 1607194113
transform 1 0 37246 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_398
timestamp 1607194113
transform 1 0 37154 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_396
timestamp 1607194113
transform 1 0 36970 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1607194113
transform 1 0 37430 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A
timestamp 1607194113
transform 1 0 37430 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1607194113
transform 1 0 37062 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1260_
timestamp 1607194113
transform 1 0 37614 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1197_
timestamp 1607194113
transform 1 0 37614 0 1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_415
timestamp 1607194113
transform 1 0 38718 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_407
timestamp 1607194113
transform 1 0 37982 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_407
timestamp 1607194113
transform 1 0 37982 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_428
timestamp 1607194113
transform 1 0 39914 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_419
timestamp 1607194113
transform 1 0 39086 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A2
timestamp 1607194113
transform 1 0 40466 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B1
timestamp 1607194113
transform 1 0 38810 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1607194113
transform 1 0 38994 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1607194113
transform 1 0 40098 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1607194113
transform 1 0 39822 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0938_
timestamp 1607194113
transform 1 0 39178 0 -1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0864_
timestamp 1607194113
transform 1 0 40282 0 1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_234
timestamp 1607194113
transform 1 0 22066 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_246
timestamp 1607194113
transform 1 0 23170 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_276
timestamp 1607194113
transform 1 0 25930 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_274
timestamp 1607194113
transform 1 0 25746 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_270
timestamp 1607194113
transform 1 0 25378 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_258
timestamp 1607194113
transform 1 0 24274 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1607194113
transform 1 0 25838 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_284
timestamp 1607194113
transform 1 0 26666 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0934_
timestamp 1607194113
transform 1 0 26942 0 -1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_68_309
timestamp 1607194113
transform 1 0 28966 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_301
timestamp 1607194113
transform 1 0 28230 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A
timestamp 1607194113
transform 1 0 29242 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1263_
timestamp 1607194113
transform 1 0 29426 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_330
timestamp 1607194113
transform 1 0 30898 0 -1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_318
timestamp 1607194113
transform 1 0 29794 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1607194113
transform 1 0 31450 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_341
timestamp 1607194113
transform 1 0 31910 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_337
timestamp 1607194113
transform 1 0 31542 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _0926_
timestamp 1607194113
transform 1 0 32002 0 -1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_68_372
timestamp 1607194113
transform 1 0 34762 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_360
timestamp 1607194113
transform 1 0 33658 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B1
timestamp 1607194113
transform 1 0 33474 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A1
timestamp 1607194113
transform 1 0 33290 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_384
timestamp 1607194113
transform 1 0 35866 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_396
timestamp 1607194113
transform 1 0 36970 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A1_N
timestamp 1607194113
transform 1 0 38626 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1607194113
transform 1 0 37062 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1201_
timestamp 1607194113
transform 1 0 37154 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_427
timestamp 1607194113
transform 1 0 39822 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_420
timestamp 1607194113
transform 1 0 39178 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_416
timestamp 1607194113
transform 1 0 38810 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B1
timestamp 1607194113
transform 1 0 40190 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1607194113
transform 1 0 39270 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A2
timestamp 1607194113
transform 1 0 40374 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0869_
timestamp 1607194113
transform 1 0 39454 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_234
timestamp 1607194113
transform 1 0 22066 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_222
timestamp 1607194113
transform 1 0 20962 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__CLK
timestamp 1607194113
transform 1 0 22802 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1607194113
transform 1 0 22986 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1383_
timestamp 1607194113
transform 1 0 23078 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_275
timestamp 1607194113
transform 1 0 25838 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_264
timestamp 1607194113
transform 1 0 24826 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1607194113
transform 1 0 25378 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1607194113
transform 1 0 25562 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_296
timestamp 1607194113
transform 1 0 27770 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_287
timestamp 1607194113
transform 1 0 26942 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1607194113
transform 1 0 27218 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0925_
timestamp 1607194113
transform 1 0 27402 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_312
timestamp 1607194113
transform 1 0 29242 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_304
timestamp 1607194113
transform 1 0 28506 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1607194113
transform 1 0 29610 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1607194113
transform 1 0 29058 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1607194113
transform 1 0 28598 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0924_
timestamp 1607194113
transform 1 0 28690 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_333
timestamp 1607194113
transform 1 0 31174 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_321
timestamp 1607194113
transform 1 0 30070 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1607194113
transform 1 0 29794 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_337
timestamp 1607194113
transform 1 0 31542 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A2_N
timestamp 1607194113
transform 1 0 31634 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B2
timestamp 1607194113
transform 1 0 31818 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1265_
timestamp 1607194113
transform 1 0 32002 0 1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_69_367
timestamp 1607194113
transform 1 0 34302 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_360
timestamp 1607194113
transform 1 0 33658 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A
timestamp 1607194113
transform 1 0 34578 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A1_N
timestamp 1607194113
transform 1 0 33474 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1607194113
transform 1 0 34210 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1200_
timestamp 1607194113
transform 1 0 34762 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_388
timestamp 1607194113
transform 1 0 36234 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_376
timestamp 1607194113
transform 1 0 35130 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B2
timestamp 1607194113
transform 1 0 36326 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1264_
timestamp 1607194113
transform 1 0 36510 0 1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_409
timestamp 1607194113
transform 1 0 38166 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A1_N
timestamp 1607194113
transform 1 0 37982 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_432
timestamp 1607194113
transform 1 0 40282 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_428
timestamp 1607194113
transform 1 0 39914 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_421
timestamp 1607194113
transform 1 0 39270 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B
timestamp 1607194113
transform 1 0 40374 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1607194113
transform 1 0 39822 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_227
timestamp 1607194113
transform 1 0 21422 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_247
timestamp 1607194113
transform 1 0 23262 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_239
timestamp 1607194113
transform 1 0 22526 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__B1
timestamp 1607194113
transform 1 0 23354 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1266_
timestamp 1607194113
transform 1 0 23538 0 -1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_276
timestamp 1607194113
transform 1 0 25930 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_274
timestamp 1607194113
transform 1 0 25746 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_270
timestamp 1607194113
transform 1 0 25378 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A2_N
timestamp 1607194113
transform 1 0 25194 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__B2
timestamp 1607194113
transform 1 0 25010 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1607194113
transform 1 0 25838 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_292
timestamp 1607194113
transform 1 0 27402 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_288
timestamp 1607194113
transform 1 0 27034 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1424_
timestamp 1607194113
transform 1 0 27494 0 -1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_314
timestamp 1607194113
transform 1 0 29426 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__CLK
timestamp 1607194113
transform 1 0 29242 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_334
timestamp 1607194113
transform 1 0 31266 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_326
timestamp 1607194113
transform 1 0 30530 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1607194113
transform 1 0 31450 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_349
timestamp 1607194113
transform 1 0 32646 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_337
timestamp 1607194113
transform 1 0 31542 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__CLK
timestamp 1607194113
transform 1 0 33106 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk_i
timestamp 1607194113
transform 1 0 32830 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_375
timestamp 1607194113
transform 1 0 35038 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1384_
timestamp 1607194113
transform 1 0 33290 0 -1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_70_395
timestamp 1607194113
transform 1 0 36878 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_387
timestamp 1607194113
transform 1 0 36142 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_410
timestamp 1607194113
transform 1 0 38258 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_398
timestamp 1607194113
transform 1 0 37154 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1607194113
transform 1 0 37062 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_434
timestamp 1607194113
transform 1 0 40466 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_418
timestamp 1607194113
transform 1 0 38994 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__B1
timestamp 1607194113
transform 1 0 39086 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 39270 0 -1 38672
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_71_230
timestamp 1607194113
transform 1 0 21698 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_218
timestamp 1607194113
transform 1 0 20594 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_245
timestamp 1607194113
transform 1 0 23078 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_242
timestamp 1607194113
transform 1 0 22802 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1607194113
transform 1 0 22986 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_269
timestamp 1607194113
transform 1 0 25286 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_257
timestamp 1607194113
transform 1 0 24182 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_281
timestamp 1607194113
transform 1 0 26390 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0932_
timestamp 1607194113
transform 1 0 26574 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_71_306
timestamp 1607194113
transform 1 0 28690 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_297
timestamp 1607194113
transform 1 0 27862 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1607194113
transform 1 0 28598 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_330
timestamp 1607194113
transform 1 0 30898 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_318
timestamp 1607194113
transform 1 0 29794 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_338
timestamp 1607194113
transform 1 0 31634 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A1
timestamp 1607194113
transform 1 0 33106 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0928_
timestamp 1607194113
transform 1 0 31818 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_71_367
timestamp 1607194113
transform 1 0 34302 0 1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_358
timestamp 1607194113
transform 1 0 33474 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__CLK
timestamp 1607194113
transform 1 0 34670 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B1
timestamp 1607194113
transform 1 0 33290 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1607194113
transform 1 0 34210 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1425_
timestamp 1607194113
transform 1 0 34854 0 1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_392
timestamp 1607194113
transform 1 0 36602 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_404
timestamp 1607194113
transform 1 0 37706 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_428
timestamp 1607194113
transform 1 0 39914 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_424
timestamp 1607194113
transform 1 0 39546 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_416
timestamp 1607194113
transform 1 0 38810 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1607194113
transform 1 0 39822 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_233
timestamp 1607194113
transform 1 0 21974 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1607194113
transform 1 0 21238 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_232
timestamp 1607194113
transform 1 0 21882 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__B
timestamp 1607194113
transform 1 0 21698 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1607194113
transform 1 0 21422 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0957_
timestamp 1607194113
transform 1 0 21054 0 -1 39760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1607194113
transform 1 0 21606 0 1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_245
timestamp 1607194113
transform 1 0 23078 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_241
timestamp 1607194113
transform 1 0 22710 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_256
timestamp 1607194113
transform 1 0 24090 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_244
timestamp 1607194113
transform 1 0 22986 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1607194113
transform 1 0 22986 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_269
timestamp 1607194113
transform 1 0 25286 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_257
timestamp 1607194113
transform 1 0 24182 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_276
timestamp 1607194113
transform 1 0 25930 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_274
timestamp 1607194113
transform 1 0 25746 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_268
timestamp 1607194113
transform 1 0 25194 0 -1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1607194113
transform 1 0 25838 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0935_
timestamp 1607194113
transform 1 0 25378 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_73_296
timestamp 1607194113
transform 1 0 27770 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_279
timestamp 1607194113
transform 1 0 26206 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_284
timestamp 1607194113
transform 1 0 26666 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__B1
timestamp 1607194113
transform 1 0 26942 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1203_
timestamp 1607194113
transform 1 0 27126 0 -1 39760
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _0933_
timestamp 1607194113
transform 1 0 26942 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_73_315
timestamp 1607194113
transform 1 0 29518 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_304
timestamp 1607194113
transform 1 0 28506 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_305
timestamp 1607194113
transform 1 0 28598 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1607194113
transform 1 0 28598 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0937_
timestamp 1607194113
transform 1 0 28690 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_73_335
timestamp 1607194113
transform 1 0 31358 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_327
timestamp 1607194113
transform 1 0 30622 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_335
timestamp 1607194113
transform 1 0 31358 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_329
timestamp 1607194113
transform 1 0 30806 0 -1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_317
timestamp 1607194113
transform 1 0 29702 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1607194113
transform 1 0 31450 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_347
timestamp 1607194113
transform 1 0 32462 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_354
timestamp 1607194113
transform 1 0 33106 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_346
timestamp 1607194113
transform 1 0 32370 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0929_
timestamp 1607194113
transform 1 0 31542 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0927_
timestamp 1607194113
transform 1 0 31634 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1607194113
transform 1 0 34302 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_365
timestamp 1607194113
transform 1 0 34118 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_359
timestamp 1607194113
transform 1 0 33566 0 1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_374
timestamp 1607194113
transform 1 0 34946 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A1_N
timestamp 1607194113
transform 1 0 34762 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1607194113
transform 1 0 34210 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1202_
timestamp 1607194113
transform 1 0 33290 0 -1 39760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_73_395
timestamp 1607194113
transform 1 0 36878 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_391
timestamp 1607194113
transform 1 0 36510 0 1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_379
timestamp 1607194113
transform 1 0 35406 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_394
timestamp 1607194113
transform 1 0 36786 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_386
timestamp 1607194113
transform 1 0 36050 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_407
timestamp 1607194113
transform 1 0 37982 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_414
timestamp 1607194113
transform 1 0 38626 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_402
timestamp 1607194113
transform 1 0 37522 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1607194113
transform 1 0 37798 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1607194113
transform 1 0 37062 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0939_
timestamp 1607194113
transform 1 0 36970 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0862_
timestamp 1607194113
transform 1 0 37154 0 -1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_428
timestamp 1607194113
transform 1 0 39914 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_419
timestamp 1607194113
transform 1 0 39086 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_426
timestamp 1607194113
transform 1 0 39730 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1607194113
transform 1 0 39822 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1262_
timestamp 1607194113
transform 1 0 40466 0 -1 39760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_74_219
timestamp 1607194113
transform 1 0 20686 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__CLK
timestamp 1607194113
transform 1 0 20778 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1494_
timestamp 1607194113
transform 1 0 20962 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1607194113
transform 1 0 23814 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_241
timestamp 1607194113
transform 1 0 22710 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_276
timestamp 1607194113
transform 1 0 25930 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_273
timestamp 1607194113
transform 1 0 25654 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_265
timestamp 1607194113
transform 1 0 24918 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1607194113
transform 1 0 25838 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_284
timestamp 1607194113
transform 1 0 26666 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1497_
timestamp 1607194113
transform 1 0 26758 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_306
timestamp 1607194113
transform 1 0 28690 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__CLK
timestamp 1607194113
transform 1 0 28506 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_330
timestamp 1607194113
transform 1 0 30898 0 -1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_318
timestamp 1607194113
transform 1 0 29794 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1607194113
transform 1 0 31450 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_337
timestamp 1607194113
transform 1 0 31542 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1499_
timestamp 1607194113
transform 1 0 31818 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_74_361
timestamp 1607194113
transform 1 0 33750 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__CLK
timestamp 1607194113
transform 1 0 34118 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__CLK
timestamp 1607194113
transform 1 0 33566 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1500_
timestamp 1607194113
transform 1 0 34302 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_74_394
timestamp 1607194113
transform 1 0 36786 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_386
timestamp 1607194113
transform 1 0 36050 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__CLK
timestamp 1607194113
transform 1 0 36878 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1607194113
transform 1 0 37062 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1501_
timestamp 1607194113
transform 1 0 37154 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_74_417
timestamp 1607194113
transform 1 0 38902 0 -1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__CLK
timestamp 1607194113
transform 1 0 39454 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1502_
timestamp 1607194113
transform 1 0 39638 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_227
timestamp 1607194113
transform 1 0 21422 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_239
timestamp 1607194113
transform 1 0 22526 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__CLK
timestamp 1607194113
transform 1 0 22802 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1607194113
transform 1 0 22986 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1495_
timestamp 1607194113
transform 1 0 23078 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_75_266
timestamp 1607194113
transform 1 0 25010 0 1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__D
timestamp 1607194113
transform 1 0 24826 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1496_
timestamp 1607194113
transform 1 0 25562 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1607194113
transform 1 0 27494 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__CLK
timestamp 1607194113
transform 1 0 27310 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1607194113
transform 1 0 28598 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1498_
timestamp 1607194113
transform 1 0 28690 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_327
timestamp 1607194113
transform 1 0 30622 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__CLK
timestamp 1607194113
transform 1 0 30438 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_346
timestamp 1607194113
transform 1 0 32370 0 1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_75_339
timestamp 1607194113
transform 1 0 31726 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1607194113
transform 1 0 32922 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0923_
timestamp 1607194113
transform 1 0 32002 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1607194113
transform 1 0 33106 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1607194113
transform 1 0 34302 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_365
timestamp 1607194113
transform 1 0 34118 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_357
timestamp 1607194113
transform 1 0 33382 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1607194113
transform 1 0 34210 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_393
timestamp 1607194113
transform 1 0 36694 0 1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_387
timestamp 1607194113
transform 1 0 36142 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_379
timestamp 1607194113
transform 1 0 35406 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0896_
timestamp 1607194113
transform 1 0 36326 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_410
timestamp 1607194113
transform 1 0 38258 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1607194113
transform 1 0 37246 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0922_
timestamp 1607194113
transform 1 0 37430 0 1 40848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_428
timestamp 1607194113
transform 1 0 39914 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_426
timestamp 1607194113
transform 1 0 39730 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_422
timestamp 1607194113
transform 1 0 39362 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1607194113
transform 1 0 39822 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_230
timestamp 1607194113
transform 1 0 21698 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_218
timestamp 1607194113
transform 1 0 20594 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_249
timestamp 1607194113
transform 1 0 23446 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_242
timestamp 1607194113
transform 1 0 22802 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1607194113
transform 1 0 23354 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_273
timestamp 1607194113
transform 1 0 25654 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_261
timestamp 1607194113
transform 1 0 24550 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_292
timestamp 1607194113
transform 1 0 27402 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_280
timestamp 1607194113
transform 1 0 26298 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1607194113
transform 1 0 26206 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_311
timestamp 1607194113
transform 1 0 29150 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_304
timestamp 1607194113
transform 1 0 28506 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1607194113
transform 1 0 29058 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_335
timestamp 1607194113
transform 1 0 31358 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_323
timestamp 1607194113
transform 1 0 30254 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_354
timestamp 1607194113
transform 1 0 33106 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_342
timestamp 1607194113
transform 1 0 32002 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1607194113
transform 1 0 31910 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_373
timestamp 1607194113
transform 1 0 34854 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_366
timestamp 1607194113
transform 1 0 34210 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1607194113
transform 1 0 34762 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_385
timestamp 1607194113
transform 1 0 35958 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_404
timestamp 1607194113
transform 1 0 37706 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_397
timestamp 1607194113
transform 1 0 37062 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1607194113
transform 1 0 37614 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_428
timestamp 1607194113
transform 1 0 39914 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_416
timestamp 1607194113
transform 1 0 38810 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1607194113
transform 1 0 40466 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1607194113
transform 1 0 41478 0 -1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_451
timestamp 1607194113
transform 1 0 42030 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_439
timestamp 1607194113
transform 1 0 40926 0 1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_452
timestamp 1607194113
transform 1 0 42122 0 -1 592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_440
timestamp 1607194113
transform 1 0 41018 0 -1 592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_462
timestamp 1607194113
transform 1 0 43042 0 -1 1680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_458
timestamp 1607194113
transform 1 0 42674 0 -1 1680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1607194113
transform 1 0 42766 0 -1 592
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1607194113
transform 1 0 42582 0 -1 1680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607194113
transform 1 0 42674 0 -1 592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1607194113
transform -1 0 43410 0 1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1607194113
transform -1 0 43410 0 -1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1607194113
transform -1 0 43410 0 -1 592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_451
timestamp 1607194113
transform 1 0 42030 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_439
timestamp 1607194113
transform 1 0 40926 0 1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1607194113
transform 1 0 41478 0 -1 2768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_451
timestamp 1607194113
transform 1 0 42030 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_439
timestamp 1607194113
transform 1 0 40926 0 1 1680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_458
timestamp 1607194113
transform 1 0 42674 0 -1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_inp_i
timestamp 1607194113
transform 1 0 42950 0 -1 2768
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1607194113
transform 1 0 42582 0 -1 2768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1607194113
transform -1 0 43410 0 1 1680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1607194113
transform -1 0 43410 0 -1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1607194113
transform -1 0 43410 0 1 2768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_451
timestamp 1607194113
transform 1 0 42030 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_439
timestamp 1607194113
transform 1 0 40926 0 1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1607194113
transform 1 0 41478 0 -1 3856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_462
timestamp 1607194113
transform 1 0 43042 0 -1 3856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_458
timestamp 1607194113
transform 1 0 42674 0 -1 3856
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1607194113
transform 1 0 42582 0 -1 3856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1607194113
transform -1 0 43410 0 -1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1607194113
transform -1 0 43410 0 1 3856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1607194113
transform 1 0 41478 0 -1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_451
timestamp 1607194113
transform 1 0 42030 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_439
timestamp 1607194113
transform 1 0 40926 0 1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1607194113
transform 1 0 41478 0 -1 4944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_462
timestamp 1607194113
transform 1 0 43042 0 -1 6032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_458
timestamp 1607194113
transform 1 0 42674 0 -1 6032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_462
timestamp 1607194113
transform 1 0 43042 0 -1 4944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_458
timestamp 1607194113
transform 1 0 42674 0 -1 4944
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1607194113
transform 1 0 42582 0 -1 4944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1607194113
transform 1 0 42582 0 -1 6032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1607194113
transform -1 0 43410 0 -1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1607194113
transform -1 0 43410 0 1 4944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1607194113
transform -1 0 43410 0 -1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1607194113
transform 1 0 41478 0 -1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_451
timestamp 1607194113
transform 1 0 42030 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_439
timestamp 1607194113
transform 1 0 40926 0 1 6032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_462
timestamp 1607194113
transform 1 0 43042 0 -1 7120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_458
timestamp 1607194113
transform 1 0 42674 0 -1 7120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1607194113
transform 1 0 42582 0 -1 7120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1607194113
transform -1 0 43410 0 1 6032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1607194113
transform -1 0 43410 0 -1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_451
timestamp 1607194113
transform 1 0 42030 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_439
timestamp 1607194113
transform 1 0 40926 0 1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1607194113
transform 1 0 41478 0 -1 8208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_451
timestamp 1607194113
transform 1 0 42030 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_439
timestamp 1607194113
transform 1 0 40926 0 1 7120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_462
timestamp 1607194113
transform 1 0 43042 0 -1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_458
timestamp 1607194113
transform 1 0 42674 0 -1 8208
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1607194113
transform 1 0 42582 0 -1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1607194113
transform -1 0 43410 0 1 7120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1607194113
transform -1 0 43410 0 -1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1607194113
transform -1 0 43410 0 1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1607194113
transform 1 0 41478 0 -1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_451
timestamp 1607194113
transform 1 0 42030 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_439
timestamp 1607194113
transform 1 0 40926 0 1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1607194113
transform 1 0 41478 0 -1 9296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_462
timestamp 1607194113
transform 1 0 43042 0 -1 10384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_458
timestamp 1607194113
transform 1 0 42674 0 -1 10384
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_462
timestamp 1607194113
transform 1 0 43042 0 -1 9296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_458
timestamp 1607194113
transform 1 0 42674 0 -1 9296
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1607194113
transform 1 0 42582 0 -1 9296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1607194113
transform 1 0 42582 0 -1 10384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1607194113
transform -1 0 43410 0 -1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1607194113
transform -1 0 43410 0 1 9296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1607194113
transform -1 0 43410 0 -1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1607194113
transform 1 0 41478 0 -1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_451
timestamp 1607194113
transform 1 0 42030 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_439
timestamp 1607194113
transform 1 0 40926 0 1 10384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_462
timestamp 1607194113
transform 1 0 43042 0 -1 11472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_458
timestamp 1607194113
transform 1 0 42674 0 -1 11472
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1607194113
transform 1 0 42582 0 -1 11472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1607194113
transform -1 0 43410 0 1 10384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1607194113
transform -1 0 43410 0 -1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_451
timestamp 1607194113
transform 1 0 42030 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_439
timestamp 1607194113
transform 1 0 40926 0 1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1607194113
transform 1 0 41478 0 -1 12560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_451
timestamp 1607194113
transform 1 0 42030 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_439
timestamp 1607194113
transform 1 0 40926 0 1 11472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_462
timestamp 1607194113
transform 1 0 43042 0 -1 12560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_458
timestamp 1607194113
transform 1 0 42674 0 -1 12560
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1607194113
transform 1 0 42582 0 -1 12560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1607194113
transform -1 0 43410 0 1 11472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1607194113
transform -1 0 43410 0 -1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1607194113
transform -1 0 43410 0 1 12560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_451
timestamp 1607194113
transform 1 0 42030 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_439
timestamp 1607194113
transform 1 0 40926 0 1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1607194113
transform 1 0 41478 0 -1 13648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_462
timestamp 1607194113
transform 1 0 43042 0 -1 13648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_458
timestamp 1607194113
transform 1 0 42674 0 -1 13648
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1607194113
transform 1 0 42582 0 -1 13648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1607194113
transform -1 0 43410 0 -1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1607194113
transform -1 0 43410 0 1 13648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_452
timestamp 1607194113
transform 1 0 42122 0 -1 15824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_440
timestamp 1607194113
transform 1 0 41018 0 -1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_451
timestamp 1607194113
transform 1 0 42030 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_439
timestamp 1607194113
transform 1 0 40926 0 1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1607194113
transform 1 0 41478 0 -1 14736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_458
timestamp 1607194113
transform 1 0 42674 0 -1 14736
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1607194113
transform 1 0 42582 0 -1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_462
timestamp 1607194113
transform 1 0 43042 0 -1 14736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1607194113
transform -1 0 43410 0 -1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_458
timestamp 1607194113
transform 1 0 42674 0 -1 15824
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_456
timestamp 1607194113
transform 1 0 42490 0 -1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1607194113
transform 1 0 42582 0 -1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_462
timestamp 1607194113
transform 1 0 43042 0 -1 15824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1607194113
transform -1 0 43410 0 1 14736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1607194113
transform -1 0 43410 0 -1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_448
timestamp 1607194113
transform 1 0 41754 0 -1 16912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_451
timestamp 1607194113
transform 1 0 42030 0 1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_439
timestamp 1607194113
transform 1 0 40926 0 1 15824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_462
timestamp 1607194113
transform 1 0 43042 0 -1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_458
timestamp 1607194113
transform 1 0 42674 0 -1 16912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_456
timestamp 1607194113
transform 1 0 42490 0 -1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1607194113
transform 1 0 42582 0 -1 16912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1607194113
transform -1 0 43410 0 1 15824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1607194113
transform -1 0 43410 0 -1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_453
timestamp 1607194113
transform 1 0 42214 0 1 18000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_453
timestamp 1607194113
transform 1 0 42214 0 -1 18000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_441
timestamp 1607194113
transform 1 0 41110 0 -1 18000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_443
timestamp 1607194113
transform 1 0 41294 0 1 16912
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A
timestamp 1607194113
transform 1 0 40926 0 -1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1607194113
transform 1 0 40650 0 -1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_461
timestamp 1607194113
transform 1 0 42950 0 1 18000
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_462
timestamp 1607194113
transform 1 0 43042 0 -1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_458
timestamp 1607194113
transform 1 0 42674 0 -1 18000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_455
timestamp 1607194113
transform 1 0 42398 0 1 16912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1607194113
transform 1 0 42582 0 -1 18000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1607194113
transform -1 0 43410 0 1 16912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1607194113
transform -1 0 43410 0 -1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1607194113
transform -1 0 43410 0 1 18000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_449
timestamp 1607194113
transform 1 0 41846 0 -1 20176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_438
timestamp 1607194113
transform 1 0 40834 0 -1 20176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_442
timestamp 1607194113
transform 1 0 41202 0 1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_450
timestamp 1607194113
transform 1 0 41938 0 -1 19088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_438
timestamp 1607194113
transform 1 0 40834 0 -1 19088
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A1_N
timestamp 1607194113
transform 1 0 40650 0 -1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1607194113
transform 1 0 41570 0 -1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_462
timestamp 1607194113
transform 1 0 43042 0 -1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_458
timestamp 1607194113
transform 1 0 42674 0 -1 19088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_456
timestamp 1607194113
transform 1 0 42490 0 -1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1607194113
transform 1 0 42582 0 -1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1607194113
transform -1 0 43410 0 -1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_462
timestamp 1607194113
transform 1 0 43042 0 1 19088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_454
timestamp 1607194113
transform 1 0 42306 0 1 19088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1607194113
transform -1 0 43410 0 1 19088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_462
timestamp 1607194113
transform 1 0 43042 0 -1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_458
timestamp 1607194113
transform 1 0 42674 0 -1 20176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1607194113
transform 1 0 42582 0 -1 20176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1607194113
transform -1 0 43410 0 -1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_447
timestamp 1607194113
transform 1 0 41662 0 -1 21264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1407_
timestamp 1607194113
transform 1 0 40650 0 1 20176
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_38_462
timestamp 1607194113
transform 1 0 43042 0 -1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_458
timestamp 1607194113
transform 1 0 42674 0 -1 21264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_455
timestamp 1607194113
transform 1 0 42398 0 -1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_455
timestamp 1607194113
transform 1 0 42398 0 1 20176
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[3]
timestamp 1607194113
transform 1 0 42950 0 1 20176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1607194113
transform 1 0 42582 0 -1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1607194113
transform -1 0 43410 0 1 20176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1607194113
transform -1 0 43410 0 -1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_444
timestamp 1607194113
transform 1 0 41386 0 1 21264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_460
timestamp 1607194113
transform 1 0 42858 0 1 21264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_456
timestamp 1607194113
transform 1 0 42490 0 1 21264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[2]
timestamp 1607194113
transform 1 0 42950 0 1 21264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1607194113
transform -1 0 43410 0 1 21264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_454
timestamp 1607194113
transform 1 0 42306 0 -1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_442
timestamp 1607194113
transform 1 0 41202 0 -1 22352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_462
timestamp 1607194113
transform 1 0 43042 0 -1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_458
timestamp 1607194113
transform 1 0 42674 0 -1 22352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1607194113
transform 1 0 42582 0 -1 22352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1607194113
transform -1 0 43410 0 -1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_451
timestamp 1607194113
transform 1 0 42030 0 -1 23440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_439
timestamp 1607194113
transform 1 0 40926 0 -1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A
timestamp 1607194113
transform 1 0 40742 0 -1 23440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1366_
timestamp 1607194113
transform 1 0 40650 0 1 22352
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_462
timestamp 1607194113
transform 1 0 43042 0 -1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_458
timestamp 1607194113
transform 1 0 42674 0 -1 23440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_455
timestamp 1607194113
transform 1 0 42398 0 1 22352
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[1]
timestamp 1607194113
transform 1 0 42950 0 1 22352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1607194113
transform 1 0 42582 0 -1 23440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1607194113
transform -1 0 43410 0 1 22352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1607194113
transform -1 0 43410 0 -1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_451
timestamp 1607194113
transform 1 0 42030 0 1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_439
timestamp 1607194113
transform 1 0 40926 0 1 23440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1607194113
transform -1 0 43410 0 1 23440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_450
timestamp 1607194113
transform 1 0 41938 0 -1 24528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_438
timestamp 1607194113
transform 1 0 40834 0 -1 24528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_462
timestamp 1607194113
transform 1 0 43042 0 -1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_458
timestamp 1607194113
transform 1 0 42674 0 -1 24528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_456
timestamp 1607194113
transform 1 0 42490 0 -1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1607194113
transform 1 0 42582 0 -1 24528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1607194113
transform -1 0 43410 0 -1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1419_
timestamp 1607194113
transform 1 0 40650 0 1 24528
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_45_455
timestamp 1607194113
transform 1 0 42398 0 1 24528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1607194113
transform -1 0 43410 0 1 24528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_449
timestamp 1607194113
transform 1 0 41846 0 -1 25616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_462
timestamp 1607194113
transform 1 0 43042 0 -1 25616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_458
timestamp 1607194113
transform 1 0 42674 0 -1 25616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1607194113
transform 1 0 42582 0 -1 25616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1607194113
transform -1 0 43410 0 -1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_454
timestamp 1607194113
transform 1 0 42306 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_442
timestamp 1607194113
transform 1 0 41202 0 -1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_453
timestamp 1607194113
transform 1 0 42214 0 1 25616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_442
timestamp 1607194113
transform 1 0 41202 0 1 25616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1607194113
transform 1 0 41938 0 1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1607194113
transform 1 0 40926 0 1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_462
timestamp 1607194113
transform 1 0 43042 0 -1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_458
timestamp 1607194113
transform 1 0 42674 0 -1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_461
timestamp 1607194113
transform 1 0 42950 0 1 25616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1607194113
transform 1 0 42582 0 -1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1607194113
transform -1 0 43410 0 1 25616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1607194113
transform -1 0 43410 0 -1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_452
timestamp 1607194113
transform 1 0 42122 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_440
timestamp 1607194113
transform 1 0 41018 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _0728_
timestamp 1607194113
transform 1 0 42214 0 1 26704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1607194113
transform 1 0 44054 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A2_N
timestamp 1607194113
transform 1 0 43870 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B2
timestamp 1607194113
transform 1 0 43686 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_489
timestamp 1607194113
transform 1 0 45526 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_485
timestamp 1607194113
transform 1 0 45158 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607194113
transform 1 0 45434 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_513
timestamp 1607194113
transform 1 0 47734 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_501
timestamp 1607194113
transform 1 0 46630 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_526
timestamp 1607194113
transform 1 0 48930 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1146_
timestamp 1607194113
transform 1 0 48286 0 1 26704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1142_
timestamp 1607194113
transform 1 0 49666 0 1 26704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_49_541
timestamp 1607194113
transform 1 0 50310 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607194113
transform 1 0 51046 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1458_
timestamp 1607194113
transform 1 0 51138 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_49_571
timestamp 1607194113
transform 1 0 53070 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__CLK
timestamp 1607194113
transform 1 0 52886 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1607194113
transform 1 0 53622 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_592
timestamp 1607194113
transform 1 0 55002 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_580
timestamp 1607194113
transform 1 0 53898 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_604
timestamp 1607194113
transform 1 0 56106 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__CLK
timestamp 1607194113
transform 1 0 56474 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607194113
transform 1 0 56658 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1460_
timestamp 1607194113
transform 1 0 56750 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_49_642
timestamp 1607194113
transform 1 0 59602 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_630
timestamp 1607194113
transform 1 0 58498 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_451
timestamp 1607194113
transform 1 0 42030 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_439
timestamp 1607194113
transform 1 0 40926 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_455
timestamp 1607194113
transform 1 0 42398 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B1
timestamp 1607194113
transform 1 0 42490 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A2_N
timestamp 1607194113
transform 1 0 44238 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607194113
transform 1 0 42674 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0737_
timestamp 1607194113
transform 1 0 42766 0 -1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_492
timestamp 1607194113
transform 1 0 45802 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_479
timestamp 1607194113
transform 1 0 44606 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B2
timestamp 1607194113
transform 1 0 44422 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0742_
timestamp 1607194113
transform 1 0 44974 0 -1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_50_511
timestamp 1607194113
transform 1 0 47550 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_504
timestamp 1607194113
transform 1 0 46906 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1149_
timestamp 1607194113
transform 1 0 47274 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_535
timestamp 1607194113
transform 1 0 49758 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_523
timestamp 1607194113
transform 1 0 48654 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607194113
transform 1 0 48286 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1147_
timestamp 1607194113
transform 1 0 49942 0 -1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1607194113
transform 1 0 48378 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_548
timestamp 1607194113
transform 1 0 50954 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1607194113
transform 1 0 50770 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1607194113
transform 1 0 51322 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 51506 0 -1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_50_579
timestamp 1607194113
transform 1 0 53806 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_575
timestamp 1607194113
transform 1 0 53438 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_563
timestamp 1607194113
transform 1 0 52334 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_600
timestamp 1607194113
transform 1 0 55738 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_588
timestamp 1607194113
transform 1 0 54634 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607194113
transform 1 0 53898 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1139_
timestamp 1607194113
transform 1 0 53990 0 -1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_50_612
timestamp 1607194113
transform 1 0 56842 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1140_
timestamp 1607194113
transform 1 0 57210 0 -1 27792
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_50_642
timestamp 1607194113
transform 1 0 59602 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_633
timestamp 1607194113
transform 1 0 58774 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__B1
timestamp 1607194113
transform 1 0 58590 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1607194113
transform 1 0 58406 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607194113
transform 1 0 59510 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_453
timestamp 1607194113
transform 1 0 42214 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A2_N
timestamp 1607194113
transform 1 0 42030 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0761_
timestamp 1607194113
transform 1 0 40558 0 1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_51_459
timestamp 1607194113
transform 1 0 42766 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1_N
timestamp 1607194113
transform 1 0 42858 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0760_
timestamp 1607194113
transform 1 0 43042 0 1 27792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_51_489
timestamp 1607194113
transform 1 0 45526 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_480
timestamp 1607194113
transform 1 0 44698 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B2
timestamp 1607194113
transform 1 0 44514 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1607194113
transform 1 0 46078 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607194113
transform 1 0 45434 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 46262 0 1 27792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_4  _1457_
timestamp 1607194113
transform 1 0 48102 0 1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1138_
timestamp 1607194113
transform 1 0 49850 0 1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_51_558
timestamp 1607194113
transform 1 0 51874 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_550
timestamp 1607194113
transform 1 0 51138 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_547
timestamp 1607194113
transform 1 0 50862 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__CLK
timestamp 1607194113
transform 1 0 50494 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__B
timestamp 1607194113
transform 1 0 50678 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607194113
transform 1 0 51046 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1144_
timestamp 1607194113
transform 1 0 51966 0 1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_570
timestamp 1607194113
transform 1 0 52978 0 1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1607194113
transform 1 0 52794 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B
timestamp 1607194113
transform 1 0 53346 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1044_
timestamp 1607194113
transform 1 0 53530 0 1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_51_595
timestamp 1607194113
transform 1 0 55278 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_583
timestamp 1607194113
transform 1 0 54174 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_611
timestamp 1607194113
transform 1 0 56750 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_603
timestamp 1607194113
transform 1 0 56014 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_i_A
timestamp 1607194113
transform 1 0 56198 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk_i
timestamp 1607194113
transform 1 0 56382 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607194113
transform 1 0 56658 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1141_
timestamp 1607194113
transform 1 0 56842 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_635
timestamp 1607194113
transform 1 0 58958 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_626
timestamp 1607194113
transform 1 0 58130 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A1
timestamp 1607194113
transform 1 0 57946 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1607194113
transform 1 0 58682 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_647
timestamp 1607194113
transform 1 0 60062 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_453
timestamp 1607194113
transform 1 0 42214 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_441
timestamp 1607194113
transform 1 0 41110 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B1
timestamp 1607194113
transform 1 0 42490 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A1_N
timestamp 1607194113
transform 1 0 42766 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607194113
transform 1 0 42674 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0733_
timestamp 1607194113
transform 1 0 42950 0 -1 28880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1607194113
transform 1 0 45526 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1607194113
transform 1 0 44422 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_513
timestamp 1607194113
transform 1 0 47734 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1607194113
transform 1 0 46630 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_520
timestamp 1607194113
transform 1 0 48378 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A2
timestamp 1607194113
transform 1 0 49942 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607194113
transform 1 0 48286 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1148_
timestamp 1607194113
transform 1 0 48654 0 -1 28880
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_52_557
timestamp 1607194113
transform 1 0 51782 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_549
timestamp 1607194113
transform 1 0 51046 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_541
timestamp 1607194113
transform 1 0 50310 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__B1
timestamp 1607194113
transform 1 0 50126 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0732_
timestamp 1607194113
transform 1 0 50678 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_579
timestamp 1607194113
transform 1 0 53806 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_571
timestamp 1607194113
transform 1 0 53070 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__D
timestamp 1607194113
transform 1 0 52886 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1048_
timestamp 1607194113
transform 1 0 52058 0 -1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_52_584
timestamp 1607194113
transform 1 0 54266 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607194113
transform 1 0 53898 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1461_
timestamp 1607194113
transform 1 0 55002 0 -1 28880
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1607194113
transform 1 0 53990 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_613
timestamp 1607194113
transform 1 0 56934 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__CLK
timestamp 1607194113
transform 1 0 56750 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0735_
timestamp 1607194113
transform 1 0 57486 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_635
timestamp 1607194113
transform 1 0 58958 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_623
timestamp 1607194113
transform 1 0 57854 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607194113
transform 1 0 59510 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1607194113
transform 1 0 59602 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_646
timestamp 1607194113
transform 1 0 59970 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_440
timestamp 1607194113
transform 1 0 41018 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A1_N
timestamp 1607194113
transform 1 0 41202 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B1
timestamp 1607194113
transform 1 0 41386 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0824_
timestamp 1607194113
transform 1 0 41570 0 1 28880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_466
timestamp 1607194113
transform 1 0 43410 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B2
timestamp 1607194113
transform 1 0 43226 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A2_N
timestamp 1607194113
transform 1 0 43042 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_486
timestamp 1607194113
transform 1 0 45250 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_478
timestamp 1607194113
transform 1 0 44514 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607194113
transform 1 0 45434 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0765_
timestamp 1607194113
transform 1 0 45526 0 1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_498
timestamp 1607194113
transform 1 0 46354 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B1
timestamp 1607194113
transform 1 0 46722 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A1_N
timestamp 1607194113
transform 1 0 46906 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0839_
timestamp 1607194113
transform 1 0 47090 0 1 28880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_53_534
timestamp 1607194113
transform 1 0 49666 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_524
timestamp 1607194113
transform 1 0 48746 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A2_N
timestamp 1607194113
transform 1 0 48562 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0739_
timestamp 1607194113
transform 1 0 49298 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_553
timestamp 1607194113
transform 1 0 51414 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_546
timestamp 1607194113
transform 1 0 50770 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607194113
transform 1 0 51046 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1607194113
transform 1 0 51138 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_565
timestamp 1607194113
transform 1 0 52518 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1607194113
transform 1 0 52794 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1136_
timestamp 1607194113
transform 1 0 52978 0 1 28880
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_53_595
timestamp 1607194113
transform 1 0 55278 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_586
timestamp 1607194113
transform 1 0 54450 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B1
timestamp 1607194113
transform 1 0 54266 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1607194113
transform 1 0 55002 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_611
timestamp 1607194113
transform 1 0 56750 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_607
timestamp 1607194113
transform 1 0 56382 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607194113
transform 1 0 56658 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1607194113
transform 1 0 57854 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A1_N
timestamp 1607194113
transform 1 0 58038 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0764_
timestamp 1607194113
transform 1 0 58222 0 1 28880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_53_647
timestamp 1607194113
transform 1 0 60062 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B2
timestamp 1607194113
transform 1 0 59878 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B1
timestamp 1607194113
transform 1 0 59694 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1607194113
transform 1 0 60430 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_440
timestamp 1607194113
transform 1 0 41018 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_453
timestamp 1607194113
transform 1 0 42214 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_441
timestamp 1607194113
transform 1 0 41110 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A1_N
timestamp 1607194113
transform 1 0 41110 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B1
timestamp 1607194113
transform 1 0 41294 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B1
timestamp 1607194113
transform 1 0 42306 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0819_
timestamp 1607194113
transform 1 0 41478 0 1 29968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_465
timestamp 1607194113
transform 1 0 43318 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_475
timestamp 1607194113
transform 1 0 44238 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A1_N
timestamp 1607194113
transform 1 0 42490 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A2_N
timestamp 1607194113
transform 1 0 43134 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B2
timestamp 1607194113
transform 1 0 42950 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607194113
transform 1 0 42674 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0827_
timestamp 1607194113
transform 1 0 43686 0 1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_4  _0822_
timestamp 1607194113
transform 1 0 42766 0 -1 29968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_489
timestamp 1607194113
transform 1 0 45526 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_486
timestamp 1607194113
transform 1 0 45250 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_478
timestamp 1607194113
transform 1 0 44514 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_487
timestamp 1607194113
transform 1 0 45342 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607194113
transform 1 0 45434 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_501
timestamp 1607194113
transform 1 0 46630 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_511
timestamp 1607194113
transform 1 0 47550 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_499
timestamp 1607194113
transform 1 0 46446 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1
timestamp 1607194113
transform 1 0 46722 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1_N
timestamp 1607194113
transform 1 0 46906 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0838_
timestamp 1607194113
transform 1 0 47090 0 1 29968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_534
timestamp 1607194113
transform 1 0 49666 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_522
timestamp 1607194113
transform 1 0 48562 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_528
timestamp 1607194113
transform 1 0 49114 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_520
timestamp 1607194113
transform 1 0 48378 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1607194113
transform 1 0 48930 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607194113
transform 1 0 48286 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0727_
timestamp 1607194113
transform 1 0 48562 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_550
timestamp 1607194113
transform 1 0 51138 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_546
timestamp 1607194113
transform 1 0 50770 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_555
timestamp 1607194113
transform 1 0 51598 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_540
timestamp 1607194113
transform 1 0 50218 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607194113
transform 1 0 51046 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1133_
timestamp 1607194113
transform 1 0 50954 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_54_574
timestamp 1607194113
transform 1 0 53346 0 -1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1607194113
transform 1 0 53162 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1462_
timestamp 1607194113
transform 1 0 52242 0 1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1135_
timestamp 1607194113
transform 1 0 52334 0 -1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_55_583
timestamp 1607194113
transform 1 0 54174 0 1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_590
timestamp 1607194113
transform 1 0 54818 0 -1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__CLK
timestamp 1607194113
transform 1 0 53990 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1607194113
transform 1 0 54634 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607194113
transform 1 0 53898 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1134_
timestamp 1607194113
transform 1 0 54726 0 1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1131_
timestamp 1607194113
transform 1 0 53990 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_54_599
timestamp 1607194113
transform 1 0 55646 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk_i
timestamp 1607194113
transform 1 0 55370 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1607194113
transform 1 0 55738 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_596
timestamp 1607194113
transform 1 0 55370 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_611
timestamp 1607194113
transform 1 0 56750 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_608
timestamp 1607194113
transform 1 0 56474 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_615
timestamp 1607194113
transform 1 0 57118 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_603
timestamp 1607194113
transform 1 0 56014 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk_i
timestamp 1607194113
transform 1 0 57486 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607194113
transform 1 0 56658 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_623
timestamp 1607194113
transform 1 0 57854 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_642
timestamp 1607194113
transform 1 0 59602 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_640
timestamp 1607194113
transform 1 0 59418 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_636
timestamp 1607194113
transform 1 0 59050 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_624
timestamp 1607194113
transform 1 0 57946 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_i_A
timestamp 1607194113
transform 1 0 57762 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A1_N
timestamp 1607194113
transform 1 0 58222 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607194113
transform 1 0 59510 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0841_
timestamp 1607194113
transform 1 0 58406 0 1 29968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_55_649
timestamp 1607194113
transform 1 0 60246 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B2
timestamp 1607194113
transform 1 0 60062 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B1
timestamp 1607194113
transform 1 0 59878 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk_i
timestamp 1607194113
transform 1 0 60338 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_453
timestamp 1607194113
transform 1 0 42214 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_441
timestamp 1607194113
transform 1 0 41110 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_471
timestamp 1607194113
transform 1 0 43870 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_459
timestamp 1607194113
transform 1 0 42766 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_457
timestamp 1607194113
transform 1 0 42582 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1607194113
transform 1 0 44054 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607194113
transform 1 0 42674 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0759_
timestamp 1607194113
transform 1 0 44238 0 -1 31056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_493
timestamp 1607194113
transform 1 0 45894 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2_N
timestamp 1607194113
transform 1 0 45710 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_517
timestamp 1607194113
transform 1 0 48102 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_505
timestamp 1607194113
transform 1 0 46998 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_529
timestamp 1607194113
transform 1 0 49206 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607194113
transform 1 0 48286 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0842_
timestamp 1607194113
transform 1 0 48378 0 -1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_553
timestamp 1607194113
transform 1 0 51414 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_541
timestamp 1607194113
transform 1 0 50310 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_574
timestamp 1607194113
transform 1 0 53346 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_561
timestamp 1607194113
transform 1 0 52150 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1607194113
transform 1 0 53162 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1109_
timestamp 1607194113
transform 1 0 52334 0 -1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_56_593
timestamp 1607194113
transform 1 0 55094 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_581
timestamp 1607194113
transform 1 0 53990 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607194113
transform 1 0 53898 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1049_
timestamp 1607194113
transform 1 0 54266 0 -1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_56_617
timestamp 1607194113
transform 1 0 57302 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_605
timestamp 1607194113
transform 1 0 56198 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1113_
timestamp 1607194113
transform 1 0 57578 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_642
timestamp 1607194113
transform 1 0 59602 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_640
timestamp 1607194113
transform 1 0 59418 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_632
timestamp 1607194113
transform 1 0 58682 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607194113
transform 1 0 59510 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_443
timestamp 1607194113
transform 1 0 41294 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_467
timestamp 1607194113
transform 1 0 43502 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_455
timestamp 1607194113
transform 1 0 42398 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_489
timestamp 1607194113
transform 1 0 45526 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_487
timestamp 1607194113
transform 1 0 45342 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_479
timestamp 1607194113
transform 1 0 44606 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607194113
transform 1 0 45434 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_507
timestamp 1607194113
transform 1 0 47182 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_501
timestamp 1607194113
transform 1 0 46630 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1607194113
transform 1 0 46906 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_531
timestamp 1607194113
transform 1 0 49390 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_519
timestamp 1607194113
transform 1 0 48286 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_543
timestamp 1607194113
transform 1 0 50494 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1607194113
transform 1 0 51966 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607194113
transform 1 0 51046 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1117_
timestamp 1607194113
transform 1 0 51138 0 1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_57_574
timestamp 1607194113
transform 1 0 53346 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_569
timestamp 1607194113
transform 1 0 52886 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_561
timestamp 1607194113
transform 1 0 52150 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1607194113
transform 1 0 52978 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_594
timestamp 1607194113
transform 1 0 55186 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_582
timestamp 1607194113
transform 1 0 54082 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1607194113
transform 1 0 55002 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1041_
timestamp 1607194113
transform 1 0 54174 0 1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_57_619
timestamp 1607194113
transform 1 0 57486 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_611
timestamp 1607194113
transform 1 0 56750 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_606
timestamp 1607194113
transform 1 0 56290 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607194113
transform 1 0 56658 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1468_
timestamp 1607194113
transform 1 0 57578 0 1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_639
timestamp 1607194113
transform 1 0 59326 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_650
timestamp 1607194113
transform 1 0 60338 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1607194113
transform 1 0 60062 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_454
timestamp 1607194113
transform 1 0 42306 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_442
timestamp 1607194113
transform 1 0 41202 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_438
timestamp 1607194113
transform 1 0 40834 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1607194113
transform 1 0 40926 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1607194113
transform 1 0 44238 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_471
timestamp 1607194113
transform 1 0 43870 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_459
timestamp 1607194113
transform 1 0 42766 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607194113
transform 1 0 42674 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_496
timestamp 1607194113
transform 1 0 46170 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B1
timestamp 1607194113
transform 1 0 44330 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A2_N
timestamp 1607194113
transform 1 0 45986 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0837_
timestamp 1607194113
transform 1 0 44514 0 -1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_58_511
timestamp 1607194113
transform 1 0 47550 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1607194113
transform 1 0 47366 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1114_
timestamp 1607194113
transform 1 0 46722 0 -1 32144
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_58_535
timestamp 1607194113
transform 1 0 49758 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_523
timestamp 1607194113
transform 1 0 48654 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607194113
transform 1 0 48286 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1465_
timestamp 1607194113
transform 1 0 49850 0 -1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1607194113
transform 1 0 48378 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1607194113
transform 1 0 51782 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__CLK
timestamp 1607194113
transform 1 0 51598 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_572
timestamp 1607194113
transform 1 0 53162 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1607194113
transform 1 0 52886 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_596
timestamp 1607194113
transform 1 0 55370 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_584
timestamp 1607194113
transform 1 0 54266 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607194113
transform 1 0 53898 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1607194113
transform 1 0 53990 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_608
timestamp 1607194113
transform 1 0 56474 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _1112_
timestamp 1607194113
transform 1 0 57578 0 -1 32144
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_58_635
timestamp 1607194113
transform 1 0 58958 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__B1
timestamp 1607194113
transform 1 0 58774 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607194113
transform 1 0 59510 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0710_
timestamp 1607194113
transform 1 0 59602 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_646
timestamp 1607194113
transform 1 0 59970 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_438
timestamp 1607194113
transform 1 0 40834 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__CLK
timestamp 1607194113
transform 1 0 41202 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B
timestamp 1607194113
transform 1 0 40650 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1463_
timestamp 1607194113
transform 1 0 41386 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_59_463
timestamp 1607194113
transform 1 0 43134 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1607194113
transform 1 0 43686 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1110_
timestamp 1607194113
transform 1 0 43870 0 1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_59_489
timestamp 1607194113
transform 1 0 45526 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_482
timestamp 1607194113
transform 1 0 44882 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__C
timestamp 1607194113
transform 1 0 44698 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607194113
transform 1 0 45434 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_517
timestamp 1607194113
transform 1 0 48102 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_497
timestamp 1607194113
transform 1 0 46262 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B1
timestamp 1607194113
transform 1 0 47918 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A1
timestamp 1607194113
transform 1 0 47734 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1122_
timestamp 1607194113
transform 1 0 46446 0 1 32144
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_59_532
timestamp 1607194113
transform 1 0 49482 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__C
timestamp 1607194113
transform 1 0 49298 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1111_
timestamp 1607194113
transform 1 0 48470 0 1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_59_550
timestamp 1607194113
transform 1 0 51138 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_548
timestamp 1607194113
transform 1 0 50954 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_544
timestamp 1607194113
transform 1 0 50586 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607194113
transform 1 0 51046 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1467_
timestamp 1607194113
transform 1 0 51230 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_572
timestamp 1607194113
transform 1 0 53162 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__CLK
timestamp 1607194113
transform 1 0 52978 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_596
timestamp 1607194113
transform 1 0 55370 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_584
timestamp 1607194113
transform 1 0 54266 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_611
timestamp 1607194113
transform 1 0 56750 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_608
timestamp 1607194113
transform 1 0 56474 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607194113
transform 1 0 56658 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_623
timestamp 1607194113
transform 1 0 57854 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B1
timestamp 1607194113
transform 1 0 58406 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0717_
timestamp 1607194113
transform 1 0 58590 0 1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_651
timestamp 1607194113
transform 1 0 60430 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A2_N
timestamp 1607194113
transform 1 0 60246 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A1_N
timestamp 1607194113
transform 1 0 60062 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_451
timestamp 1607194113
transform 1 0 42030 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A2
timestamp 1607194113
transform 1 0 41846 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B1
timestamp 1607194113
transform 1 0 41662 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_471
timestamp 1607194113
transform 1 0 43870 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_459
timestamp 1607194113
transform 1 0 42766 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_457
timestamp 1607194113
transform 1 0 42582 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607194113
transform 1 0 42674 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0745_
timestamp 1607194113
transform 1 0 43502 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_488
timestamp 1607194113
transform 1 0 45434 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__D
timestamp 1607194113
transform 1 0 44422 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1042_
timestamp 1607194113
transform 1 0 44606 0 -1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_60_513
timestamp 1607194113
transform 1 0 47734 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_500
timestamp 1607194113
transform 1 0 46538 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1607194113
transform 1 0 47550 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1121_
timestamp 1607194113
transform 1 0 46722 0 -1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_535
timestamp 1607194113
transform 1 0 49758 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_520
timestamp 1607194113
transform 1 0 48378 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607194113
transform 1 0 48286 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1116_
timestamp 1607194113
transform 1 0 48930 0 -1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_559
timestamp 1607194113
transform 1 0 51966 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_547
timestamp 1607194113
transform 1 0 50862 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_579
timestamp 1607194113
transform 1 0 53806 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_571
timestamp 1607194113
transform 1 0 53070 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_593
timestamp 1607194113
transform 1 0 55094 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_581
timestamp 1607194113
transform 1 0 53990 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607194113
transform 1 0 53898 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1607194113
transform 1 0 54726 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_613
timestamp 1607194113
transform 1 0 56934 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_605
timestamp 1607194113
transform 1 0 56198 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1_N
timestamp 1607194113
transform 1 0 57118 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0808_
timestamp 1607194113
transform 1 0 57302 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_60_637
timestamp 1607194113
transform 1 0 59142 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B2
timestamp 1607194113
transform 1 0 58958 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B1
timestamp 1607194113
transform 1 0 59326 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B1
timestamp 1607194113
transform 1 0 58774 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607194113
transform 1 0 59510 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0812_
timestamp 1607194113
transform 1 0 59602 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_62_453
timestamp 1607194113
transform 1 0 42214 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_441
timestamp 1607194113
transform 1 0 41110 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1607194113
transform 1 0 41846 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_437
timestamp 1607194113
transform 1 0 40742 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1607194113
transform 1 0 40558 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_471
timestamp 1607194113
transform 1 0 43870 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_459
timestamp 1607194113
transform 1 0 42766 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_457
timestamp 1607194113
transform 1 0 42582 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_469
timestamp 1607194113
transform 1 0 43686 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_461
timestamp 1607194113
transform 1 0 42950 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1607194113
transform 1 0 43870 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1607194113
transform 1 0 42674 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1607194113
transform 1 0 44054 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_486
timestamp 1607194113
transform 1 0 45250 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_489
timestamp 1607194113
transform 1 0 45526 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_476
timestamp 1607194113
transform 1 0 44330 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1607194113
transform 1 0 45434 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1607194113
transform 1 0 44974 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_517
timestamp 1607194113
transform 1 0 48102 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_509
timestamp 1607194113
transform 1 0 47366 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_498
timestamp 1607194113
transform 1 0 46354 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_511
timestamp 1607194113
transform 1 0 47550 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_501
timestamp 1607194113
transform 1 0 46630 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1120_
timestamp 1607194113
transform 1 0 46722 0 -1 34320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1115_
timestamp 1607194113
transform 1 0 46906 0 1 33232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_532
timestamp 1607194113
transform 1 0 49482 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_520
timestamp 1607194113
transform 1 0 48378 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_535
timestamp 1607194113
transform 1 0 49758 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_523
timestamp 1607194113
transform 1 0 48654 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1607194113
transform 1 0 48286 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_550
timestamp 1607194113
transform 1 0 51138 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_544
timestamp 1607194113
transform 1 0 50586 0 -1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_553
timestamp 1607194113
transform 1 0 51414 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_547
timestamp 1607194113
transform 1 0 50862 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A1_N
timestamp 1607194113
transform 1 0 51230 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1607194113
transform 1 0 51414 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1607194113
transform 1 0 51046 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0800_
timestamp 1607194113
transform 1 0 51598 0 -1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1607194113
transform 1 0 51138 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_579
timestamp 1607194113
transform 1 0 53806 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_575
timestamp 1607194113
transform 1 0 53438 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_561
timestamp 1607194113
transform 1 0 52150 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A2_N
timestamp 1607194113
transform 1 0 53254 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B2
timestamp 1607194113
transform 1 0 53070 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A1_N
timestamp 1607194113
transform 1 0 52334 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B1
timestamp 1607194113
transform 1 0 52518 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0702_
timestamp 1607194113
transform 1 0 52702 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_594
timestamp 1607194113
transform 1 0 55186 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_581
timestamp 1607194113
transform 1 0 53990 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_599
timestamp 1607194113
transform 1 0 55646 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_587
timestamp 1607194113
transform 1 0 54542 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__C
timestamp 1607194113
transform 1 0 54174 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A2_N
timestamp 1607194113
transform 1 0 54358 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B2
timestamp 1607194113
transform 1 0 54174 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1607194113
transform 1 0 53898 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0721_
timestamp 1607194113
transform 1 0 54358 0 -1 34320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_618
timestamp 1607194113
transform 1 0 57394 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_606
timestamp 1607194113
transform 1 0 56290 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_619
timestamp 1607194113
transform 1 0 57486 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_611
timestamp 1607194113
transform 1 0 56750 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_607
timestamp 1607194113
transform 1 0 56382 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A1_N
timestamp 1607194113
transform 1 0 57578 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1607194113
transform 1 0 56658 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_638
timestamp 1607194113
transform 1 0 59234 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_630
timestamp 1607194113
transform 1 0 58498 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_642
timestamp 1607194113
transform 1 0 59602 0 1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B2
timestamp 1607194113
transform 1 0 59418 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B1
timestamp 1607194113
transform 1 0 59234 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1607194113
transform 1 0 59510 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0720_
timestamp 1607194113
transform 1 0 59602 0 -1 34320
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_4  _0712_
timestamp 1607194113
transform 1 0 57762 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__D
timestamp 1607194113
transform 1 0 60430 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0815_
timestamp 1607194113
transform 1 0 59970 0 1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_63_444
timestamp 1607194113
transform 1 0 41386 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_468
timestamp 1607194113
transform 1 0 43594 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_456
timestamp 1607194113
transform 1 0 42490 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_489
timestamp 1607194113
transform 1 0 45526 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_480
timestamp 1607194113
transform 1 0 44698 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1607194113
transform 1 0 45434 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__CLK
timestamp 1607194113
transform 1 0 48010 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1466_
timestamp 1607194113
transform 1 0 46262 0 1 34320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_527
timestamp 1607194113
transform 1 0 49022 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_518
timestamp 1607194113
transform 1 0 48194 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1607194113
transform 1 0 48746 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_550
timestamp 1607194113
transform 1 0 51138 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_547
timestamp 1607194113
transform 1 0 50862 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_539
timestamp 1607194113
transform 1 0 50126 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__C
timestamp 1607194113
transform 1 0 51506 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1607194113
transform 1 0 51046 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0816_
timestamp 1607194113
transform 1 0 51690 0 1 34320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_63_565
timestamp 1607194113
transform 1 0 52518 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B1
timestamp 1607194113
transform 1 0 53070 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0699_
timestamp 1607194113
transform 1 0 53254 0 1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_593
timestamp 1607194113
transform 1 0 55094 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A1_N
timestamp 1607194113
transform 1 0 54910 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A2_N
timestamp 1607194113
transform 1 0 54726 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_611
timestamp 1607194113
transform 1 0 56750 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_609
timestamp 1607194113
transform 1 0 56566 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_605
timestamp 1607194113
transform 1 0 56198 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1607194113
transform 1 0 56658 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_623
timestamp 1607194113
transform 1 0 57854 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1607194113
transform 1 0 57946 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1_N
timestamp 1607194113
transform 1 0 59602 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0715_
timestamp 1607194113
transform 1 0 58130 0 1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_646
timestamp 1607194113
transform 1 0 59970 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A2_N
timestamp 1607194113
transform 1 0 59786 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_444
timestamp 1607194113
transform 1 0 41386 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_459
timestamp 1607194113
transform 1 0 42766 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_456
timestamp 1607194113
transform 1 0 42490 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__CLK
timestamp 1607194113
transform 1 0 43042 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1607194113
transform 1 0 42674 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1387_
timestamp 1607194113
transform 1 0 43226 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_64_483
timestamp 1607194113
transform 1 0 44974 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1518_
timestamp 1607194113
transform 1 0 45710 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_64_512
timestamp 1607194113
transform 1 0 47642 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__CLK
timestamp 1607194113
transform 1 0 47458 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_528
timestamp 1607194113
transform 1 0 49114 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_520
timestamp 1607194113
transform 1 0 48378 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_518
timestamp 1607194113
transform 1 0 48194 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__C
timestamp 1607194113
transform 1 0 49298 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1607194113
transform 1 0 48286 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0796_
timestamp 1607194113
transform 1 0 49482 0 -1 35408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_64_549
timestamp 1607194113
transform 1 0 51046 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_541
timestamp 1607194113
transform 1 0 50310 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0791_
timestamp 1607194113
transform 1 0 51230 0 -1 35408
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_64_577
timestamp 1607194113
transform 1 0 53622 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_569
timestamp 1607194113
transform 1 0 52886 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A2
timestamp 1607194113
transform 1 0 52702 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B2
timestamp 1607194113
transform 1 0 52518 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_592
timestamp 1607194113
transform 1 0 55002 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__C
timestamp 1607194113
transform 1 0 54818 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1607194113
transform 1 0 53898 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0859_
timestamp 1607194113
transform 1 0 53990 0 -1 35408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_616
timestamp 1607194113
transform 1 0 57210 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_604
timestamp 1607194113
transform 1 0 56106 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_642
timestamp 1607194113
transform 1 0 59602 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_640
timestamp 1607194113
transform 1 0 59418 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_628
timestamp 1607194113
transform 1 0 58314 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1607194113
transform 1 0 59510 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_443
timestamp 1607194113
transform 1 0 41294 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_455
timestamp 1607194113
transform 1 0 42398 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1607194113
transform 1 0 42766 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1428_
timestamp 1607194113
transform 1 0 42950 0 1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_492
timestamp 1607194113
transform 1 0 45802 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_480
timestamp 1607194113
transform 1 0 44698 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1607194113
transform 1 0 45434 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1607194113
transform 1 0 45526 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_507
timestamp 1607194113
transform 1 0 47182 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1607194113
transform 1 0 46906 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_531
timestamp 1607194113
transform 1 0 49390 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_519
timestamp 1607194113
transform 1 0 48286 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__C
timestamp 1607194113
transform 1 0 48378 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0696_
timestamp 1607194113
transform 1 0 48562 0 1 35408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_550
timestamp 1607194113
transform 1 0 51138 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_543
timestamp 1607194113
transform 1 0 50494 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1607194113
transform 1 0 51046 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_562
timestamp 1607194113
transform 1 0 52242 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B1
timestamp 1607194113
transform 1 0 52426 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0798_
timestamp 1607194113
transform 1 0 52610 0 1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_598
timestamp 1607194113
transform 1 0 55554 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_586
timestamp 1607194113
transform 1 0 54450 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1_N
timestamp 1607194113
transform 1 0 54266 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A2_N
timestamp 1607194113
transform 1 0 54082 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_617
timestamp 1607194113
transform 1 0 57302 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A
timestamp 1607194113
transform 1 0 57118 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1607194113
transform 1 0 56658 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1253_
timestamp 1607194113
transform 1 0 56750 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_623
timestamp 1607194113
transform 1 0 57854 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2_N
timestamp 1607194113
transform 1 0 59602 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1607194113
transform 1 0 57946 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0810_
timestamp 1607194113
transform 1 0 58130 0 1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_644
timestamp 1607194113
transform 1 0 59786 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_450
timestamp 1607194113
transform 1 0 41938 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_438
timestamp 1607194113
transform 1 0 40834 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B2
timestamp 1607194113
transform 1 0 40650 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_471
timestamp 1607194113
transform 1 0 43870 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_459
timestamp 1607194113
transform 1 0 42766 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1607194113
transform 1 0 42674 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_492
timestamp 1607194113
transform 1 0 45802 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_483
timestamp 1607194113
transform 1 0 44974 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1607194113
transform 1 0 45342 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1607194113
transform 1 0 45526 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_516
timestamp 1607194113
transform 1 0 48010 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_504
timestamp 1607194113
transform 1 0 46906 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_532
timestamp 1607194113
transform 1 0 49482 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_520
timestamp 1607194113
transform 1 0 48378 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1607194113
transform 1 0 48286 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_544
timestamp 1607194113
transform 1 0 50586 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _0689_
timestamp 1607194113
transform 1 0 50954 0 -1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_66_578
timestamp 1607194113
transform 1 0 53714 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_566
timestamp 1607194113
transform 1 0 52610 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A2
timestamp 1607194113
transform 1 0 52426 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B2
timestamp 1607194113
transform 1 0 52242 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_596
timestamp 1607194113
transform 1 0 55370 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_584
timestamp 1607194113
transform 1 0 54266 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1607194113
transform 1 0 53898 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1607194113
transform 1 0 53990 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_604
timestamp 1607194113
transform 1 0 56106 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__CLK
timestamp 1607194113
transform 1 0 56290 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1390_
timestamp 1607194113
transform 1 0 56474 0 -1 36496
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_642
timestamp 1607194113
transform 1 0 59602 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_639
timestamp 1607194113
transform 1 0 59326 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_627
timestamp 1607194113
transform 1 0 58222 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1607194113
transform 1 0 59510 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_449
timestamp 1607194113
transform 1 0 41846 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_448
timestamp 1607194113
transform 1 0 41754 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_436
timestamp 1607194113
transform 1 0 40650 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1607194113
transform 1 0 41662 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0917_
timestamp 1607194113
transform 1 0 40558 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_457
timestamp 1607194113
transform 1 0 42582 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_474
timestamp 1607194113
transform 1 0 44146 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A1_N
timestamp 1607194113
transform 1 0 44238 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A1_N
timestamp 1607194113
transform 1 0 43962 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1607194113
transform 1 0 42674 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1261_
timestamp 1607194113
transform 1 0 42766 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1198_
timestamp 1607194113
transform 1 0 42490 0 1 36496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_68_485
timestamp 1607194113
transform 1 0 45158 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_477
timestamp 1607194113
transform 1 0 44422 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_486
timestamp 1607194113
transform 1 0 45250 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A1
timestamp 1607194113
transform 1 0 45342 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B1
timestamp 1607194113
transform 1 0 45526 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__B1
timestamp 1607194113
transform 1 0 45526 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1607194113
transform 1 0 45434 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0793_
timestamp 1607194113
transform 1 0 45710 0 -1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _0692_
timestamp 1607194113
transform 1 0 45710 0 1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_68_517
timestamp 1607194113
transform 1 0 48102 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_505
timestamp 1607194113
transform 1 0 46998 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1607194113
transform 1 0 48102 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1607194113
transform 1 0 46998 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_532
timestamp 1607194113
transform 1 0 49482 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_520
timestamp 1607194113
transform 1 0 48378 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_537
timestamp 1607194113
transform 1 0 49942 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_529
timestamp 1607194113
transform 1 0 49206 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1607194113
transform 1 0 48286 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1607194113
transform 1 0 50034 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_550
timestamp 1607194113
transform 1 0 51138 0 1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_541
timestamp 1607194113
transform 1 0 50310 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1607194113
transform 1 0 51046 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1433_
timestamp 1607194113
transform 1 0 50586 0 -1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1392_
timestamp 1607194113
transform 1 0 51690 0 1 36496
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_68_577
timestamp 1607194113
transform 1 0 53622 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_565
timestamp 1607194113
transform 1 0 52518 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_577
timestamp 1607194113
transform 1 0 53622 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__CLK
timestamp 1607194113
transform 1 0 52334 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__CLK
timestamp 1607194113
transform 1 0 53438 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_589
timestamp 1607194113
transform 1 0 54726 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_581
timestamp 1607194113
transform 1 0 53990 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_589
timestamp 1607194113
transform 1 0 54726 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1607194113
transform 1 0 53898 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1257_
timestamp 1607194113
transform 1 0 54818 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_68_606
timestamp 1607194113
transform 1 0 56290 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_618
timestamp 1607194113
transform 1 0 57394 0 1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_611
timestamp 1607194113
transform 1 0 56750 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_609
timestamp 1607194113
transform 1 0 56566 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_601
timestamp 1607194113
transform 1 0 55830 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1607194113
transform 1 0 56842 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1607194113
transform 1 0 56658 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1255_
timestamp 1607194113
transform 1 0 57026 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1190_
timestamp 1607194113
transform 1 0 57026 0 1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_640
timestamp 1607194113
transform 1 0 59418 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_632
timestamp 1607194113
transform 1 0 58682 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_641
timestamp 1607194113
transform 1 0 59510 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_629
timestamp 1607194113
transform 1 0 58406 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1607194113
transform 1 0 57946 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1_N
timestamp 1607194113
transform 1 0 58498 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1607194113
transform 1 0 59510 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1194_
timestamp 1607194113
transform 1 0 59602 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1607194113
transform 1 0 58130 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_454
timestamp 1607194113
transform 1 0 42306 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_444
timestamp 1607194113
transform 1 0 41386 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A
timestamp 1607194113
transform 1 0 41754 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1607194113
transform 1 0 41202 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0916_
timestamp 1607194113
transform 1 0 40558 0 1 37584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1607194113
transform 1 0 41938 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_466
timestamp 1607194113
transform 1 0 43410 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_492
timestamp 1607194113
transform 1 0 45802 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_486
timestamp 1607194113
transform 1 0 45250 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_478
timestamp 1607194113
transform 1 0 44514 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1607194113
transform 1 0 45434 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1607194113
transform 1 0 45526 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_504
timestamp 1607194113
transform 1 0 46906 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B1
timestamp 1607194113
transform 1 0 47090 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A2
timestamp 1607194113
transform 1 0 47274 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0910_
timestamp 1607194113
transform 1 0 47458 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_534
timestamp 1607194113
transform 1 0 49666 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_522
timestamp 1607194113
transform 1 0 48562 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_546
timestamp 1607194113
transform 1 0 50770 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1607194113
transform 1 0 50862 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1607194113
transform 1 0 51046 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1191_
timestamp 1607194113
transform 1 0 51138 0 1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_578
timestamp 1607194113
transform 1 0 53714 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_566
timestamp 1607194113
transform 1 0 52610 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_596
timestamp 1607194113
transform 1 0 55370 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A
timestamp 1607194113
transform 1 0 54818 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1256_
timestamp 1607194113
transform 1 0 55002 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_619
timestamp 1607194113
transform 1 0 57486 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_611
timestamp 1607194113
transform 1 0 56750 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_607
timestamp 1607194113
transform 1 0 56382 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk_i
timestamp 1607194113
transform 1 0 56106 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk_i
timestamp 1607194113
transform 1 0 57670 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1607194113
transform 1 0 56658 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_626
timestamp 1607194113
transform 1 0 58130 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_i_A
timestamp 1607194113
transform 1 0 57946 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1192_
timestamp 1607194113
transform 1 0 58222 0 1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_645
timestamp 1607194113
transform 1 0 59878 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A1_N
timestamp 1607194113
transform 1 0 59694 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_446
timestamp 1607194113
transform 1 0 41570 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1607194113
transform 1 0 41018 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0897_
timestamp 1607194113
transform 1 0 41202 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_471
timestamp 1607194113
transform 1 0 43870 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_459
timestamp 1607194113
transform 1 0 42766 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1607194113
transform 1 0 42674 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__CLK
timestamp 1607194113
transform 1 0 46170 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1427_
timestamp 1607194113
transform 1 0 44422 0 -1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_70_516
timestamp 1607194113
transform 1 0 48010 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_510
timestamp 1607194113
transform 1 0 47458 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_498
timestamp 1607194113
transform 1 0 46354 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B
timestamp 1607194113
transform 1 0 48102 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_529
timestamp 1607194113
transform 1 0 49206 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1607194113
transform 1 0 49022 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1607194113
transform 1 0 48286 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0904_
timestamp 1607194113
transform 1 0 48378 0 -1 38672
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_70_549
timestamp 1607194113
transform 1 0 51046 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_541
timestamp 1607194113
transform 1 0 50310 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__B1
timestamp 1607194113
transform 1 0 51138 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1254_
timestamp 1607194113
transform 1 0 51322 0 -1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_568
timestamp 1607194113
transform 1 0 52794 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_581
timestamp 1607194113
transform 1 0 53990 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B2
timestamp 1607194113
transform 1 0 54266 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A2
timestamp 1607194113
transform 1 0 54450 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1607194113
transform 1 0 53898 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0901_
timestamp 1607194113
transform 1 0 54634 0 -1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_70_618
timestamp 1607194113
transform 1 0 57394 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_606
timestamp 1607194113
transform 1 0 56290 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B1
timestamp 1607194113
transform 1 0 56106 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A1
timestamp 1607194113
transform 1 0 55922 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_642
timestamp 1607194113
transform 1 0 59602 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_70_638
timestamp 1607194113
transform 1 0 59234 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_630
timestamp 1607194113
transform 1 0 58498 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1607194113
transform 1 0 59510 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1607194113
transform 1 0 60154 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1432_
timestamp 1607194113
transform 1 0 60338 0 -1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_71_436
timestamp 1607194113
transform 1 0 40650 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B2
timestamp 1607194113
transform 1 0 42214 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A2
timestamp 1607194113
transform 1 0 42030 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0921_
timestamp 1607194113
transform 1 0 40742 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_71_455
timestamp 1607194113
transform 1 0 42398 0 1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _1199_
timestamp 1607194113
transform 1 0 42950 0 1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_494
timestamp 1607194113
transform 1 0 45986 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_485
timestamp 1607194113
transform 1 0 45158 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_477
timestamp 1607194113
transform 1 0 44422 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1607194113
transform 1 0 45802 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1607194113
transform 1 0 45434 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1607194113
transform 1 0 45526 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1
timestamp 1607194113
transform 1 0 47090 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0911_
timestamp 1607194113
transform 1 0 47274 0 1 38672
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_71_533
timestamp 1607194113
transform 1 0 49574 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_521
timestamp 1607194113
transform 1 0 48470 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B2
timestamp 1607194113
transform 1 0 50678 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A2
timestamp 1607194113
transform 1 0 50862 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1607194113
transform 1 0 51046 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0899_
timestamp 1607194113
transform 1 0 51138 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_71_576
timestamp 1607194113
transform 1 0 53530 0 1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_564
timestamp 1607194113
transform 1 0 52426 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_598
timestamp 1607194113
transform 1 0 55554 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B2
timestamp 1607194113
transform 1 0 53898 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A2
timestamp 1607194113
transform 1 0 54082 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0914_
timestamp 1607194113
transform 1 0 54266 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_71_611
timestamp 1607194113
transform 1 0 56750 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1607194113
transform 1 0 56658 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_635
timestamp 1607194113
transform 1 0 58958 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_623
timestamp 1607194113
transform 1 0 57854 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_647
timestamp 1607194113
transform 1 0 60062 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A
timestamp 1607194113
transform 1 0 60154 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1193_
timestamp 1607194113
transform 1 0 60338 0 1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_450
timestamp 1607194113
transform 1 0 41938 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_464
timestamp 1607194113
transform 1 0 43226 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1607194113
transform 1 0 43042 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1607194113
transform 1 0 42674 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1607194113
transform 1 0 42766 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_488
timestamp 1607194113
transform 1 0 45434 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_476
timestamp 1607194113
transform 1 0 44330 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_512
timestamp 1607194113
transform 1 0 47642 0 -1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_500
timestamp 1607194113
transform 1 0 46538 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_520
timestamp 1607194113
transform 1 0 48378 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_518
timestamp 1607194113
transform 1 0 48194 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1607194113
transform 1 0 49482 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1607194113
transform 1 0 48286 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0902_
timestamp 1607194113
transform 1 0 49666 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_555
timestamp 1607194113
transform 1 0 51598 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_543
timestamp 1607194113
transform 1 0 50494 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_579
timestamp 1607194113
transform 1 0 53806 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_567
timestamp 1607194113
transform 1 0 52702 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B2
timestamp 1607194113
transform 1 0 53990 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A2
timestamp 1607194113
transform 1 0 54174 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A1
timestamp 1607194113
transform 1 0 55646 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1607194113
transform 1 0 53898 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0912_
timestamp 1607194113
transform 1 0 54358 0 -1 39760
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_72_615
timestamp 1607194113
transform 1 0 57118 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_611
timestamp 1607194113
transform 1 0 56750 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_603
timestamp 1607194113
transform 1 0 56014 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B1
timestamp 1607194113
transform 1 0 55830 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk_i
timestamp 1607194113
transform 1 0 56842 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_642
timestamp 1607194113
transform 1 0 59602 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_639
timestamp 1607194113
transform 1 0 59326 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_627
timestamp 1607194113
transform 1 0 58222 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1607194113
transform 1 0 59510 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_444
timestamp 1607194113
transform 1 0 41386 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_440
timestamp 1607194113
transform 1 0 41018 0 1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__CLK
timestamp 1607194113
transform 1 0 41478 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1386_
timestamp 1607194113
transform 1 0 41662 0 1 39760
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_73_466
timestamp 1607194113
transform 1 0 43410 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_489
timestamp 1607194113
transform 1 0 45526 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_486
timestamp 1607194113
transform 1 0 45250 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_478
timestamp 1607194113
transform 1 0 44514 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1607194113
transform 1 0 45434 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_510
timestamp 1607194113
transform 1 0 47458 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_497
timestamp 1607194113
transform 1 0 46262 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1607194113
transform 1 0 46446 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0913_
timestamp 1607194113
transform 1 0 46630 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_73_522
timestamp 1607194113
transform 1 0 48562 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1607194113
transform 1 0 49298 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0900_
timestamp 1607194113
transform 1 0 49482 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_73_550
timestamp 1607194113
transform 1 0 51138 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_541
timestamp 1607194113
transform 1 0 50310 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1607194113
transform 1 0 51046 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_574
timestamp 1607194113
transform 1 0 53346 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_562
timestamp 1607194113
transform 1 0 52242 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1259_
timestamp 1607194113
transform 1 0 54450 0 1 39760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_618
timestamp 1607194113
transform 1 0 57394 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_611
timestamp 1607194113
transform 1 0 56750 0 1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_602
timestamp 1607194113
transform 1 0 55922 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1607194113
transform 1 0 56658 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1607194113
transform 1 0 57118 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_642
timestamp 1607194113
transform 1 0 59602 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_630
timestamp 1607194113
transform 1 0 58498 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1196_
timestamp 1607194113
transform 1 0 59878 0 1 39760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_75_452
timestamp 1607194113
transform 1 0 42122 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_440
timestamp 1607194113
transform 1 0 41018 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_444
timestamp 1607194113
transform 1 0 41386 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1607194113
transform 1 0 44054 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_460
timestamp 1607194113
transform 1 0 42858 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__CLK
timestamp 1607194113
transform 1 0 42490 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1607194113
transform 1 0 43042 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1607194113
transform 1 0 42674 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1503_
timestamp 1607194113
transform 1 0 42766 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _0915_
timestamp 1607194113
transform 1 0 43226 0 1 40848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_489
timestamp 1607194113
transform 1 0 45526 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_485
timestamp 1607194113
transform 1 0 45158 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_486
timestamp 1607194113
transform 1 0 45250 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_478
timestamp 1607194113
transform 1 0 44514 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1607194113
transform 1 0 45434 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1504_
timestamp 1607194113
transform 1 0 45434 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_75_505
timestamp 1607194113
transform 1 0 46998 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_501
timestamp 1607194113
transform 1 0 46630 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_517
timestamp 1607194113
transform 1 0 48102 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_509
timestamp 1607194113
transform 1 0 47366 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__CLK
timestamp 1607194113
transform 1 0 47182 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1505_
timestamp 1607194113
transform 1 0 47090 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_527
timestamp 1607194113
transform 1 0 49022 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_520
timestamp 1607194113
transform 1 0 48378 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__CLK
timestamp 1607194113
transform 1 0 48838 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1607194113
transform 1 0 48286 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1506_
timestamp 1607194113
transform 1 0 49482 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_75_547
timestamp 1607194113
transform 1 0 50862 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_539
timestamp 1607194113
transform 1 0 50126 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_553
timestamp 1607194113
transform 1 0 51414 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__CLK
timestamp 1607194113
transform 1 0 51230 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1607194113
transform 1 0 51046 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1507_
timestamp 1607194113
transform 1 0 51138 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_571
timestamp 1607194113
transform 1 0 53070 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_577
timestamp 1607194113
transform 1 0 53622 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_565
timestamp 1607194113
transform 1 0 52518 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__CLK
timestamp 1607194113
transform 1 0 52886 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_583
timestamp 1607194113
transform 1 0 54174 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_597
timestamp 1607194113
transform 1 0 55462 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_593
timestamp 1607194113
transform 1 0 55094 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_581
timestamp 1607194113
transform 1 0 53990 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1607194113
transform 1 0 53898 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1388_
timestamp 1607194113
transform 1 0 55554 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1258_
timestamp 1607194113
transform 1 0 54450 0 1 40848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_75_604
timestamp 1607194113
transform 1 0 56106 0 1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_619
timestamp 1607194113
transform 1 0 57486 0 -1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__CLK
timestamp 1607194113
transform 1 0 57302 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A1_N
timestamp 1607194113
transform 1 0 55922 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1607194113
transform 1 0 56658 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1389_
timestamp 1607194113
transform 1 0 56750 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_632
timestamp 1607194113
transform 1 0 58682 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_642
timestamp 1607194113
transform 1 0 59602 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_640
timestamp 1607194113
transform 1 0 59418 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_628
timestamp 1607194113
transform 1 0 58314 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__CLK
timestamp 1607194113
transform 1 0 58498 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1607194113
transform 1 0 59510 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1607194113
transform 1 0 58038 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_644
timestamp 1607194113
transform 1 0 59786 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1195_
timestamp 1607194113
transform 1 0 60062 0 1 40848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_447
timestamp 1607194113
transform 1 0 41662 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_435
timestamp 1607194113
transform 1 0 40558 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_466
timestamp 1607194113
transform 1 0 43410 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_459
timestamp 1607194113
transform 1 0 42766 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1607194113
transform 1 0 43318 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_490
timestamp 1607194113
transform 1 0 45618 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_478
timestamp 1607194113
transform 1 0 44514 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1607194113
transform 1 0 46170 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_509
timestamp 1607194113
transform 1 0 47366 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_497
timestamp 1607194113
transform 1 0 46262 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_528
timestamp 1607194113
transform 1 0 49114 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_521
timestamp 1607194113
transform 1 0 48470 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1607194113
transform 1 0 49022 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_559
timestamp 1607194113
transform 1 0 51966 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_552
timestamp 1607194113
transform 1 0 51322 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_540
timestamp 1607194113
transform 1 0 50218 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1607194113
transform 1 0 51874 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_571
timestamp 1607194113
transform 1 0 53070 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_590
timestamp 1607194113
transform 1 0 54818 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_583
timestamp 1607194113
transform 1 0 54174 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1607194113
transform 1 0 54726 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_621
timestamp 1607194113
transform 1 0 57670 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_614
timestamp 1607194113
transform 1 0 57026 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_602
timestamp 1607194113
transform 1 0 55922 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1607194113
transform 1 0 57578 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_633
timestamp 1607194113
transform 1 0 58774 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_645
timestamp 1607194113
transform 1 0 59878 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1607194113
transform 1 0 60430 0 -1 41936
box -38 -48 130 592
use delayline_9_hd_25_1  inst_idelay_line
timestamp 1607276668
transform 1 0 45434 0 1 1472
box 800 800 20764 22385
use sky130_fd_sc_hd__fill_1  FILLER_49_670
timestamp 1607194113
transform 1 0 62178 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_666
timestamp 1607194113
transform 1 0 61810 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_654
timestamp 1607194113
transform 1 0 60706 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607194113
transform 1 0 62270 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1456_
timestamp 1607194113
transform 1 0 62362 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_691
timestamp 1607194113
transform 1 0 64110 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1152_
timestamp 1607194113
transform 1 0 64846 0 1 26704
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_49_726
timestamp 1607194113
transform 1 0 67330 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_714
timestamp 1607194113
transform 1 0 66226 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__B1
timestamp 1607194113
transform 1 0 66042 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607194113
transform 1 0 67882 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1470_
timestamp 1607194113
transform 1 0 67974 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[8]
timestamp 1607194113
transform 1 0 70458 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[6]
timestamp 1607194113
transform 1 0 71286 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[5]
timestamp 1607194113
transform 1 0 71102 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[4]
timestamp 1607194113
transform 1 0 70918 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[3]
timestamp 1607194113
transform 1 0 69722 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[2]
timestamp 1607194113
transform 1 0 69906 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[1]
timestamp 1607194113
transform 1 0 70090 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[0]
timestamp 1607194113
transform 1 0 70274 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1326_
timestamp 1607194113
transform 1 0 70642 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_785
timestamp 1607194113
transform 1 0 72758 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[7]
timestamp 1607194113
transform 1 0 71470 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1607194113
transform 1 0 73034 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1100_
timestamp 1607194113
transform 1 0 71654 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_807
timestamp 1607194113
transform 1 0 74782 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_792
timestamp 1607194113
transform 1 0 73402 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B1
timestamp 1607194113
transform 1 0 73218 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607194113
transform 1 0 73494 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1099_
timestamp 1607194113
transform 1 0 73586 0 1 26704
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_49_818
timestamp 1607194113
transform 1 0 75794 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1607194113
transform 1 0 75518 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_846
timestamp 1607194113
transform 1 0 78370 0 1 26704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_842
timestamp 1607194113
transform 1 0 78002 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_830
timestamp 1607194113
transform 1 0 76898 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1607194113
transform 1 0 78094 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__CLK
timestamp 1607194113
transform 1 0 78922 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607194113
transform 1 0 79106 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1477_
timestamp 1607194113
transform 1 0 79198 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_654
timestamp 1607194113
transform 1 0 60706 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1607194113
transform 1 0 62086 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1607194113
transform 1 0 61810 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_689
timestamp 1607194113
transform 1 0 63926 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_671
timestamp 1607194113
transform 1 0 62270 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1153_
timestamp 1607194113
transform 1 0 62822 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_703
timestamp 1607194113
transform 1 0 65214 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_701
timestamp 1607194113
transform 1 0 65030 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607194113
transform 1 0 65122 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_727
timestamp 1607194113
transform 1 0 67422 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_715
timestamp 1607194113
transform 1 0 66318 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_750
timestamp 1607194113
transform 1 0 69538 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_742
timestamp 1607194113
transform 1 0 68802 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1607194113
transform 1 0 67790 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1105_
timestamp 1607194113
transform 1 0 67974 0 -1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_50_764
timestamp 1607194113
transform 1 0 70826 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_762
timestamp 1607194113
transform 1 0 70642 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_754
timestamp 1607194113
transform 1 0 69906 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__CLK
timestamp 1607194113
transform 1 0 69722 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_inp_i
timestamp 1607194113
transform 1 0 71286 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607194113
transform 1 0 70734 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0780_
timestamp 1607194113
transform 1 0 70918 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_773
timestamp 1607194113
transform 1 0 71654 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A1
timestamp 1607194113
transform 1 0 71470 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1472_
timestamp 1607194113
transform 1 0 72022 0 -1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_50_798
timestamp 1607194113
transform 1 0 73954 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__CLK
timestamp 1607194113
transform 1 0 73770 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1098_
timestamp 1607194113
transform 1 0 74506 0 -1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_50_825
timestamp 1607194113
transform 1 0 76438 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_823
timestamp 1607194113
transform 1 0 76254 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_811
timestamp 1607194113
transform 1 0 75150 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607194113
transform 1 0 76346 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_846
timestamp 1607194113
transform 1 0 78370 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_837
timestamp 1607194113
transform 1 0 77542 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1607194113
transform 1 0 78094 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_868
timestamp 1607194113
transform 1 0 80394 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B1
timestamp 1607194113
transform 1 0 78922 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1080_
timestamp 1607194113
transform 1 0 79106 0 -1 27792
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_51_659
timestamp 1607194113
transform 1 0 61166 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_681
timestamp 1607194113
transform 1 0 63190 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607194113
transform 1 0 62270 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1155_
timestamp 1607194113
transform 1 0 63926 0 1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1154_
timestamp 1607194113
transform 1 0 62362 0 1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_51_710
timestamp 1607194113
transform 1 0 65858 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_698
timestamp 1607194113
transform 1 0 64754 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_730
timestamp 1607194113
transform 1 0 67698 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_722
timestamp 1607194113
transform 1 0 66962 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_748
timestamp 1607194113
transform 1 0 69354 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_740
timestamp 1607194113
transform 1 0 68618 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607194113
transform 1 0 67882 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1104_
timestamp 1607194113
transform 1 0 67974 0 1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1097_
timestamp 1607194113
transform 1 0 69538 0 1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_51_769
timestamp 1607194113
transform 1 0 71286 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_757
timestamp 1607194113
transform 1 0 70182 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_785
timestamp 1607194113
transform 1 0 72758 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_775
timestamp 1607194113
transform 1 0 71838 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1101_
timestamp 1607194113
transform 1 0 71930 0 1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_51_794
timestamp 1607194113
transform 1 0 73586 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607194113
transform 1 0 73494 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1471_
timestamp 1607194113
transform 1 0 73862 0 1 27792
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_51_818
timestamp 1607194113
transform 1 0 75794 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__CLK
timestamp 1607194113
transform 1 0 75610 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_842
timestamp 1607194113
transform 1 0 78002 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_830
timestamp 1607194113
transform 1 0 76898 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_855
timestamp 1607194113
transform 1 0 79198 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1607194113
transform 1 0 79750 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607194113
transform 1 0 79106 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1079_
timestamp 1607194113
transform 1 0 79934 0 1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_52_658
timestamp 1607194113
transform 1 0 61074 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1607194113
transform 1 0 61258 0 -1 28880
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_52_679
timestamp 1607194113
transform 1 0 63006 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1151_
timestamp 1607194113
transform 1 0 63742 0 -1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_52_703
timestamp 1607194113
transform 1 0 65214 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_694
timestamp 1607194113
transform 1 0 64386 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607194113
transform 1 0 65122 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_728
timestamp 1607194113
transform 1 0 67514 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_723
timestamp 1607194113
transform 1 0 67054 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_715
timestamp 1607194113
transform 1 0 66318 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1088_
timestamp 1607194113
transform 1 0 67146 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_740
timestamp 1607194113
transform 1 0 68618 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1607194113
transform 1 0 69354 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0749_
timestamp 1607194113
transform 1 0 68250 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_764
timestamp 1607194113
transform 1 0 70826 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_751
timestamp 1607194113
transform 1 0 69630 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607194113
transform 1 0 70734 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_783
timestamp 1607194113
transform 1 0 72574 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A
timestamp 1607194113
transform 1 0 73126 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1607194113
transform 1 0 71562 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1036_
timestamp 1607194113
transform 1 0 71746 0 -1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_52_800
timestamp 1607194113
transform 1 0 74138 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _1102_
timestamp 1607194113
transform 1 0 73310 0 -1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_52_825
timestamp 1607194113
transform 1 0 76438 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_812
timestamp 1607194113
transform 1 0 75242 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607194113
transform 1 0 76346 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_849
timestamp 1607194113
transform 1 0 78646 0 -1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_837
timestamp 1607194113
transform 1 0 77542 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_855
timestamp 1607194113
transform 1 0 79198 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__CLK
timestamp 1607194113
transform 1 0 79290 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1478_
timestamp 1607194113
transform 1 0 79474 0 -1 28880
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_53_668
timestamp 1607194113
transform 1 0 61994 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_656
timestamp 1607194113
transform 1 0 60890 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1607194113
transform 1 0 60706 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_683
timestamp 1607194113
transform 1 0 63374 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1607194113
transform 1 0 62362 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1607194113
transform 1 0 63926 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607194113
transform 1 0 62270 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1047_
timestamp 1607194113
transform 1 0 62546 0 1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_53_710
timestamp 1607194113
transform 1 0 65858 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_698
timestamp 1607194113
transform 1 0 64754 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1150_
timestamp 1607194113
transform 1 0 64110 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_53_722
timestamp 1607194113
transform 1 0 66962 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A2
timestamp 1607194113
transform 1 0 67514 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A1
timestamp 1607194113
transform 1 0 67698 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_749
timestamp 1607194113
transform 1 0 69446 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__B1
timestamp 1607194113
transform 1 0 69262 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607194113
transform 1 0 67882 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1107_
timestamp 1607194113
transform 1 0 67974 0 1 28880
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_53_758
timestamp 1607194113
transform 1 0 70274 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1607194113
transform 1 0 70826 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1327_
timestamp 1607194113
transform 1 0 71010 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1607194113
transform 1 0 69998 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_785
timestamp 1607194113
transform 1 0 72758 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_773
timestamp 1607194113
transform 1 0 71654 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_799
timestamp 1607194113
transform 1 0 74046 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1607194113
transform 1 0 73862 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1607194113
transform 1 0 74414 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607194113
transform 1 0 73494 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1082_
timestamp 1607194113
transform 1 0 74598 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1607194113
transform 1 0 73586 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_829
timestamp 1607194113
transform 1 0 76806 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_812
timestamp 1607194113
transform 1 0 75242 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__C
timestamp 1607194113
transform 1 0 75794 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1050_
timestamp 1607194113
transform 1 0 75978 0 1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_53_840
timestamp 1607194113
transform 1 0 77818 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk_i
timestamp 1607194113
transform 1 0 77542 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_867
timestamp 1607194113
transform 1 0 80302 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_859
timestamp 1607194113
transform 1 0 79566 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_855
timestamp 1607194113
transform 1 0 79198 0 1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_852
timestamp 1607194113
transform 1 0 78922 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607194113
transform 1 0 79106 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1069_
timestamp 1607194113
transform 1 0 79658 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_55_669
timestamp 1607194113
transform 1 0 62086 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_661
timestamp 1607194113
transform 1 0 61350 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_664
timestamp 1607194113
transform 1 0 61626 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_653
timestamp 1607194113
transform 1 0 60614 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1607194113
transform 1 0 61350 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_681
timestamp 1607194113
transform 1 0 63190 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607194113
transform 1 0 62270 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1607194113
transform 1 0 62362 0 -1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1157_
timestamp 1607194113
transform 1 0 62362 0 1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_55_693
timestamp 1607194113
transform 1 0 64294 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_699
timestamp 1607194113
transform 1 0 64846 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_691
timestamp 1607194113
transform 1 0 64110 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__B
timestamp 1607194113
transform 1 0 65858 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607194113
transform 1 0 65122 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1607194113
transform 1 0 64386 0 1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1158_
timestamp 1607194113
transform 1 0 65214 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_55_724
timestamp 1607194113
transform 1 0 67146 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_713
timestamp 1607194113
transform 1 0 66134 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_722
timestamp 1607194113
transform 1 0 66962 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_718
timestamp 1607194113
transform 1 0 66594 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_714
timestamp 1607194113
transform 1 0 66226 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__A
timestamp 1607194113
transform 1 0 66042 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1607194113
transform 1 0 66686 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1028_
timestamp 1607194113
transform 1 0 67698 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1607194113
transform 1 0 66870 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_739
timestamp 1607194113
transform 1 0 68526 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_733
timestamp 1607194113
transform 1 0 67974 0 1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_734
timestamp 1607194113
transform 1 0 68066 0 -1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607194113
transform 1 0 67882 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_746
timestamp 1607194113
transform 1 0 69170 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_740
timestamp 1607194113
transform 1 0 68618 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B
timestamp 1607194113
transform 1 0 68710 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A
timestamp 1607194113
transform 1 0 68894 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1607194113
transform 1 0 68618 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1096_
timestamp 1607194113
transform 1 0 69078 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1607194113
transform 1 0 68802 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_758
timestamp 1607194113
transform 1 0 70274 0 1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_54_760
timestamp 1607194113
transform 1 0 70458 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_752
timestamp 1607194113
transform 1 0 69722 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1059_
timestamp 1607194113
transform 1 0 69906 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_769
timestamp 1607194113
transform 1 0 71286 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A
timestamp 1607194113
transform 1 0 70826 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607194113
transform 1 0 70734 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1072_
timestamp 1607194113
transform 1 0 70826 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1607194113
transform 1 0 71010 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_768
timestamp 1607194113
transform 1 0 71194 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_787
timestamp 1607194113
transform 1 0 72942 0 1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_777
timestamp 1607194113
transform 1 0 72022 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1607194113
transform 1 0 72758 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A
timestamp 1607194113
transform 1 0 72298 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1093_
timestamp 1607194113
transform 1 0 72482 0 -1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1092_
timestamp 1607194113
transform 1 0 72114 0 1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_55_794
timestamp 1607194113
transform 1 0 73586 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A
timestamp 1607194113
transform 1 0 73862 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607194113
transform 1 0 73494 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1084_
timestamp 1607194113
transform 1 0 74046 0 1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_55_806
timestamp 1607194113
transform 1 0 74690 0 1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_803
timestamp 1607194113
transform 1 0 74414 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_i_A
timestamp 1607194113
transform 1 0 74506 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk_i
timestamp 1607194113
transform 1 0 74690 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1083_
timestamp 1607194113
transform 1 0 74966 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_54_791
timestamp 1607194113
transform 1 0 73310 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_828
timestamp 1607194113
transform 1 0 76714 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_816
timestamp 1607194113
transform 1 0 75610 0 -1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__B1
timestamp 1607194113
transform 1 0 75242 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 1607194113
transform 1 0 76162 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607194113
transform 1 0 76346 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1094_
timestamp 1607194113
transform 1 0 75426 0 1 29968
box -38 -48 1326 592
use sky130_fd_sc_hd__or4_4  _1039_
timestamp 1607194113
transform 1 0 76438 0 -1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_55_839
timestamp 1607194113
transform 1 0 77726 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_845
timestamp 1607194113
transform 1 0 78278 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_834
timestamp 1607194113
transform 1 0 77266 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1607194113
transform 1 0 78002 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1607194113
transform 1 0 77450 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_867
timestamp 1607194113
transform 1 0 80302 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_855
timestamp 1607194113
transform 1 0 79198 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_851
timestamp 1607194113
transform 1 0 78830 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_858
timestamp 1607194113
transform 1 0 79474 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1607194113
transform 1 0 79290 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1607194113
transform 1 0 79842 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607194113
transform 1 0 79106 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1070_
timestamp 1607194113
transform 1 0 80026 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1607194113
transform 1 0 79014 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_670
timestamp 1607194113
transform 1 0 62178 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_666
timestamp 1607194113
transform 1 0 61810 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_654
timestamp 1607194113
transform 1 0 60706 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_682
timestamp 1607194113
transform 1 0 63282 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A
timestamp 1607194113
transform 1 0 63098 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__B
timestamp 1607194113
transform 1 0 62914 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1156_
timestamp 1607194113
transform 1 0 62270 0 -1 31056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_56_703
timestamp 1607194113
transform 1 0 65214 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_694
timestamp 1607194113
transform 1 0 64386 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607194113
transform 1 0 65122 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_715
timestamp 1607194113
transform 1 0 66318 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1469_
timestamp 1607194113
transform 1 0 66502 0 -1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_748
timestamp 1607194113
transform 1 0 69354 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_736
timestamp 1607194113
transform 1 0 68250 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1106_
timestamp 1607194113
transform 1 0 68986 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_764
timestamp 1607194113
transform 1 0 70826 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_760
timestamp 1607194113
transform 1 0 70458 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607194113
transform 1 0 70734 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1474_
timestamp 1607194113
transform 1 0 71102 0 -1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_56_788
timestamp 1607194113
transform 1 0 73034 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__CLK
timestamp 1607194113
transform 1 0 72850 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_805
timestamp 1607194113
transform 1 0 74598 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1089_
timestamp 1607194113
transform 1 0 73770 0 -1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_56_825
timestamp 1607194113
transform 1 0 76438 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_816
timestamp 1607194113
transform 1 0 75610 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607194113
transform 1 0 76346 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1607194113
transform 1 0 75334 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_831
timestamp 1607194113
transform 1 0 76990 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1473_
timestamp 1607194113
transform 1 0 77082 0 -1 31056
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_853
timestamp 1607194113
transform 1 0 79014 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__CLK
timestamp 1607194113
transform 1 0 78830 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1087_
timestamp 1607194113
transform 1 0 80118 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_670
timestamp 1607194113
transform 1 0 62178 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_662
timestamp 1607194113
transform 1 0 61442 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_679
timestamp 1607194113
transform 1 0 63006 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_672
timestamp 1607194113
transform 1 0 62362 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607194113
transform 1 0 62270 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0701_
timestamp 1607194113
transform 1 0 62638 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_709
timestamp 1607194113
transform 1 0 65766 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_703
timestamp 1607194113
transform 1 0 65214 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_691
timestamp 1607194113
transform 1 0 64110 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_i_A
timestamp 1607194113
transform 1 0 65858 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_727
timestamp 1607194113
transform 1 0 67422 0 1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_715
timestamp 1607194113
transform 1 0 66318 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk_i
timestamp 1607194113
transform 1 0 66042 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_746
timestamp 1607194113
transform 1 0 69170 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_733
timestamp 1607194113
transform 1 0 67974 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_731
timestamp 1607194113
transform 1 0 67790 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__C
timestamp 1607194113
transform 1 0 68158 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607194113
transform 1 0 67882 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0857_
timestamp 1607194113
transform 1 0 68342 0 1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_770
timestamp 1607194113
transform 1 0 71378 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_758
timestamp 1607194113
transform 1 0 70274 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_782
timestamp 1607194113
transform 1 0 72482 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_803
timestamp 1607194113
transform 1 0 74414 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_790
timestamp 1607194113
transform 1 0 73218 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1607194113
transform 1 0 73310 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607194113
transform 1 0 73494 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1090_
timestamp 1607194113
transform 1 0 73586 0 1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_818
timestamp 1607194113
transform 1 0 75794 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1085_
timestamp 1607194113
transform 1 0 75150 0 1 31056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_57_842
timestamp 1607194113
transform 1 0 78002 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_830
timestamp 1607194113
transform 1 0 76898 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_867
timestamp 1607194113
transform 1 0 80302 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_855
timestamp 1607194113
transform 1 0 79198 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607194113
transform 1 0 79106 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_670
timestamp 1607194113
transform 1 0 62178 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_658
timestamp 1607194113
transform 1 0 61074 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_682
timestamp 1607194113
transform 1 0 63282 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1607194113
transform 1 0 63374 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0858_
timestamp 1607194113
transform 1 0 63558 0 -1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_703
timestamp 1607194113
transform 1 0 65214 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_696
timestamp 1607194113
transform 1 0 64570 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__C
timestamp 1607194113
transform 1 0 64386 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607194113
transform 1 0 65122 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_727
timestamp 1607194113
transform 1 0 67422 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_715
timestamp 1607194113
transform 1 0 66318 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_735
timestamp 1607194113
transform 1 0 68158 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A1_N
timestamp 1607194113
transform 1 0 68250 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0853_
timestamp 1607194113
transform 1 0 68434 0 -1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_58_764
timestamp 1607194113
transform 1 0 70826 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_762
timestamp 1607194113
transform 1 0 70642 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_758
timestamp 1607194113
transform 1 0 70274 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B2
timestamp 1607194113
transform 1 0 70090 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B1
timestamp 1607194113
transform 1 0 69906 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607194113
transform 1 0 70734 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_779
timestamp 1607194113
transform 1 0 72206 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_772
timestamp 1607194113
transform 1 0 71562 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1607194113
transform 1 0 72022 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1607194113
transform 1 0 71746 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_806
timestamp 1607194113
transform 1 0 74690 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_799
timestamp 1607194113
transform 1 0 74046 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_791
timestamp 1607194113
transform 1 0 73310 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1607194113
transform 1 0 74506 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1607194113
transform 1 0 74230 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_825
timestamp 1607194113
transform 1 0 76438 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_818
timestamp 1607194113
transform 1 0 75794 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607194113
transform 1 0 76346 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__B1
timestamp 1607194113
transform 1 0 76990 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk_i
timestamp 1607194113
transform 1 0 77174 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0846_
timestamp 1607194113
transform 1 0 77450 0 -1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_864
timestamp 1607194113
transform 1 0 80026 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_852
timestamp 1607194113
transform 1 0 78922 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0752_
timestamp 1607194113
transform 1 0 80394 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_663
timestamp 1607194113
transform 1 0 61534 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_672
timestamp 1607194113
transform 1 0 62362 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607194113
transform 1 0 62270 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0781_
timestamp 1607194113
transform 1 0 63098 0 1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B2
timestamp 1607194113
transform 1 0 64938 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__C
timestamp 1607194113
transform 1 0 65122 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A2_N
timestamp 1607194113
transform 1 0 64754 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B1
timestamp 1607194113
transform 1 0 64570 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0786_
timestamp 1607194113
transform 1 0 65306 0 1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_59_725
timestamp 1607194113
transform 1 0 67238 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_713
timestamp 1607194113
transform 1 0 66134 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_745
timestamp 1607194113
transform 1 0 69078 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_733
timestamp 1607194113
transform 1 0 67974 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_731
timestamp 1607194113
transform 1 0 67790 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607194113
transform 1 0 67882 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1519_
timestamp 1607194113
transform 1 0 69446 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_770
timestamp 1607194113
transform 1 0 71378 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__CLK
timestamp 1607194113
transform 1 0 71194 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_782
timestamp 1607194113
transform 1 0 72482 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_790
timestamp 1607194113
transform 1 0 73218 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607194113
transform 1 0 73494 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1475_
timestamp 1607194113
transform 1 0 73586 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_59_815
timestamp 1607194113
transform 1 0 75518 0 1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__CLK
timestamp 1607194113
transform 1 0 75334 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A1_N
timestamp 1607194113
transform 1 0 75886 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0778_
timestamp 1607194113
transform 1 0 76070 0 1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_839
timestamp 1607194113
transform 1 0 77726 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B2
timestamp 1607194113
transform 1 0 77542 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_867
timestamp 1607194113
transform 1 0 80302 0 1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_855
timestamp 1607194113
transform 1 0 79198 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_851
timestamp 1607194113
transform 1 0 78830 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607194113
transform 1 0 79106 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_662
timestamp 1607194113
transform 1 0 61442 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2_N
timestamp 1607194113
transform 1 0 61258 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1_N
timestamp 1607194113
transform 1 0 61074 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_674
timestamp 1607194113
transform 1 0 62546 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _0785_
timestamp 1607194113
transform 1 0 62914 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A2_N
timestamp 1607194113
transform 1 0 64754 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__B2
timestamp 1607194113
transform 1 0 64570 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B
timestamp 1607194113
transform 1 0 64938 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A1_N
timestamp 1607194113
transform 1 0 64386 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607194113
transform 1 0 65122 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0787_
timestamp 1607194113
transform 1 0 65214 0 -1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_60_714
timestamp 1607194113
transform 1 0 66226 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B1
timestamp 1607194113
transform 1 0 66502 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A1_N
timestamp 1607194113
transform 1 0 66686 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__C
timestamp 1607194113
transform 1 0 66042 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0856_
timestamp 1607194113
transform 1 0 66870 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_748
timestamp 1607194113
transform 1 0 69354 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_741
timestamp 1607194113
transform 1 0 68710 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A2_N
timestamp 1607194113
transform 1 0 68526 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B2
timestamp 1607194113
transform 1 0 68342 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1607194113
transform 1 0 69078 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_764
timestamp 1607194113
transform 1 0 70826 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_760
timestamp 1607194113
transform 1 0 70458 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607194113
transform 1 0 70734 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_788
timestamp 1607194113
transform 1 0 73034 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_776
timestamp 1607194113
transform 1 0 71930 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_796
timestamp 1607194113
transform 1 0 73770 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A1_N
timestamp 1607194113
transform 1 0 73954 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0852_
timestamp 1607194113
transform 1 0 74138 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_60_825
timestamp 1607194113
transform 1 0 76438 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_818
timestamp 1607194113
transform 1 0 75794 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B2
timestamp 1607194113
transform 1 0 75610 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607194113
transform 1 0 76346 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_831
timestamp 1607194113
transform 1 0 76990 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1607194113
transform 1 0 77082 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0770_
timestamp 1607194113
transform 1 0 77266 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_862
timestamp 1607194113
transform 1 0 79842 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_850
timestamp 1607194113
transform 1 0 78738 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_665
timestamp 1607194113
transform 1 0 61718 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_653
timestamp 1607194113
transform 1 0 60614 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_669
timestamp 1607194113
transform 1 0 62086 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_657
timestamp 1607194113
transform 1 0 60982 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__D
timestamp 1607194113
transform 1 0 60798 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_677
timestamp 1607194113
transform 1 0 62822 0 -1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_678
timestamp 1607194113
transform 1 0 62914 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_672
timestamp 1607194113
transform 1 0 62362 0 1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__C
timestamp 1607194113
transform 1 0 64018 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1607194113
transform 1 0 63006 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1607194113
transform 1 0 63374 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1607194113
transform 1 0 62270 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0836_
timestamp 1607194113
transform 1 0 63190 0 1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0757_
timestamp 1607194113
transform 1 0 63558 0 -1 34320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_703
timestamp 1607194113
transform 1 0 65214 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_696
timestamp 1607194113
transform 1 0 64570 0 -1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_704
timestamp 1607194113
transform 1 0 65306 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_692
timestamp 1607194113
transform 1 0 64202 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__C
timestamp 1607194113
transform 1 0 64386 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A
timestamp 1607194113
transform 1 0 65398 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1607194113
transform 1 0 65122 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0788_
timestamp 1607194113
transform 1 0 65582 0 1 33232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_62_727
timestamp 1607194113
transform 1 0 67422 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_715
timestamp 1607194113
transform 1 0 66318 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_728
timestamp 1607194113
transform 1 0 67514 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_716
timestamp 1607194113
transform 1 0 66410 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A1_N
timestamp 1607194113
transform 1 0 67514 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__C1
timestamp 1607194113
transform 1 0 67698 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A2_N
timestamp 1607194113
transform 1 0 67698 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_750
timestamp 1607194113
transform 1 0 69538 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_749
timestamp 1607194113
transform 1 0 69446 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B2
timestamp 1607194113
transform 1 0 69354 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A2
timestamp 1607194113
transform 1 0 69262 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1607194113
transform 1 0 67882 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0743_
timestamp 1607194113
transform 1 0 67974 0 1 33232
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _0725_
timestamp 1607194113
transform 1 0 67882 0 -1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_764
timestamp 1607194113
transform 1 0 70826 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_762
timestamp 1607194113
transform 1 0 70642 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_761
timestamp 1607194113
transform 1 0 70550 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1607194113
transform 1 0 70734 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_788
timestamp 1607194113
transform 1 0 73034 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_776
timestamp 1607194113
transform 1 0 71930 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_785
timestamp 1607194113
transform 1 0 72758 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_773
timestamp 1607194113
transform 1 0 71654 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_792
timestamp 1607194113
transform 1 0 73402 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1607194113
transform 1 0 73494 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0803_
timestamp 1607194113
transform 1 0 73586 0 1 33232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0704_
timestamp 1607194113
transform 1 0 73494 0 -1 34320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_62_802
timestamp 1607194113
transform 1 0 74322 0 -1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_803
timestamp 1607194113
transform 1 0 74414 0 1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B
timestamp 1607194113
transform 1 0 74138 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B
timestamp 1607194113
transform 1 0 74230 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1607194113
transform 1 0 74966 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1607194113
transform 1 0 74874 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_825
timestamp 1607194113
transform 1 0 76438 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_823
timestamp 1607194113
transform 1 0 76254 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_811
timestamp 1607194113
transform 1 0 75150 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_824
timestamp 1607194113
transform 1 0 76346 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_812
timestamp 1607194113
transform 1 0 75242 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1607194113
transform 1 0 76346 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_837
timestamp 1607194113
transform 1 0 77542 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_848
timestamp 1607194113
transform 1 0 78554 0 1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_836
timestamp 1607194113
transform 1 0 77450 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _0754_
timestamp 1607194113
transform 1 0 77910 0 -1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_857
timestamp 1607194113
transform 1 0 79382 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1607194113
transform 1 0 79106 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0833_
timestamp 1607194113
transform 1 0 79198 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_63_670
timestamp 1607194113
transform 1 0 62178 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_658
timestamp 1607194113
transform 1 0 61074 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_688
timestamp 1607194113
transform 1 0 63834 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1607194113
transform 1 0 62270 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0831_
timestamp 1607194113
transform 1 0 62362 0 1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_700
timestamp 1607194113
transform 1 0 64938 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_724
timestamp 1607194113
transform 1 0 67146 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_712
timestamp 1607194113
transform 1 0 66042 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2_N
timestamp 1607194113
transform 1 0 67698 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1_N
timestamp 1607194113
transform 1 0 67974 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1607194113
transform 1 0 67882 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0818_
timestamp 1607194113
transform 1 0 68158 0 1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_765
timestamp 1607194113
transform 1 0 70918 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_753
timestamp 1607194113
transform 1 0 69814 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B2
timestamp 1607194113
transform 1 0 69630 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_789
timestamp 1607194113
transform 1 0 73126 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_777
timestamp 1607194113
transform 1 0 72022 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_800
timestamp 1607194113
transform 1 0 74138 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_794
timestamp 1607194113
transform 1 0 73586 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1607194113
transform 1 0 73494 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1397_
timestamp 1607194113
transform 1 0 74230 0 1 34320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_822
timestamp 1607194113
transform 1 0 76162 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__CLK
timestamp 1607194113
transform 1 0 75978 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_846
timestamp 1607194113
transform 1 0 78370 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_834
timestamp 1607194113
transform 1 0 77266 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_863
timestamp 1607194113
transform 1 0 79934 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_855
timestamp 1607194113
transform 1 0 79198 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1607194113
transform 1 0 79106 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1240_
timestamp 1607194113
transform 1 0 80026 0 1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_666
timestamp 1607194113
transform 1 0 61810 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_654
timestamp 1607194113
transform 1 0 60706 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_689
timestamp 1607194113
transform 1 0 63926 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_672
timestamp 1607194113
transform 1 0 62362 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0750_
timestamp 1607194113
transform 1 0 62454 0 -1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_703
timestamp 1607194113
transform 1 0 65214 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_701
timestamp 1607194113
transform 1 0 65030 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_i_A
timestamp 1607194113
transform 1 0 65766 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1607194113
transform 1 0 65122 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_726
timestamp 1607194113
transform 1 0 67330 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_714
timestamp 1607194113
transform 1 0 66226 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk_i
timestamp 1607194113
transform 1 0 65950 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_734
timestamp 1607194113
transform 1 0 68066 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__C1
timestamp 1607194113
transform 1 0 68342 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0828_
timestamp 1607194113
transform 1 0 68526 0 -1 35408
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_64_767
timestamp 1607194113
transform 1 0 71102 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_755
timestamp 1607194113
transform 1 0 69998 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A2
timestamp 1607194113
transform 1 0 69814 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1607194113
transform 1 0 70734 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1607194113
transform 1 0 70826 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_779
timestamp 1607194113
transform 1 0 72206 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_791
timestamp 1607194113
transform 1 0 73310 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1438_
timestamp 1607194113
transform 1 0 73862 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_825
timestamp 1607194113
transform 1 0 76438 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_818
timestamp 1607194113
transform 1 0 75794 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__CLK
timestamp 1607194113
transform 1 0 75610 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1607194113
transform 1 0 76346 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_849
timestamp 1607194113
transform 1 0 78646 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_837
timestamp 1607194113
transform 1 0 77542 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__CLK
timestamp 1607194113
transform 1 0 79198 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1401_
timestamp 1607194113
transform 1 0 79382 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_65_668
timestamp 1607194113
transform 1 0 61994 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_656
timestamp 1607194113
transform 1 0 60890 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A1_N
timestamp 1607194113
transform 1 0 62086 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B2
timestamp 1607194113
transform 1 0 64018 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1607194113
transform 1 0 63834 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1607194113
transform 1 0 62270 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0756_
timestamp 1607194113
transform 1 0 62362 0 1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_704
timestamp 1607194113
transform 1 0 65306 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_692
timestamp 1607194113
transform 1 0 64202 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_728
timestamp 1607194113
transform 1 0 67514 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_716
timestamp 1607194113
transform 1 0 66410 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_736
timestamp 1607194113
transform 1 0 68250 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1607194113
transform 1 0 67882 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1396_
timestamp 1607194113
transform 1 0 68986 0 1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1607194113
transform 1 0 67974 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_765
timestamp 1607194113
transform 1 0 70918 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__CLK
timestamp 1607194113
transform 1 0 70734 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_789
timestamp 1607194113
transform 1 0 73126 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_777
timestamp 1607194113
transform 1 0 72022 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1607194113
transform 1 0 73494 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1184_
timestamp 1607194113
transform 1 0 73586 0 1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_822
timestamp 1607194113
transform 1 0 76162 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_810
timestamp 1607194113
transform 1 0 75058 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A
timestamp 1607194113
transform 1 0 75610 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1246_
timestamp 1607194113
transform 1 0 75794 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_846
timestamp 1607194113
transform 1 0 78370 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_834
timestamp 1607194113
transform 1 0 77266 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_861
timestamp 1607194113
transform 1 0 79750 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A
timestamp 1607194113
transform 1 0 79566 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1607194113
transform 1 0 79106 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1238_
timestamp 1607194113
transform 1 0 79198 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_654
timestamp 1607194113
transform 1 0 60706 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A1_N
timestamp 1607194113
transform 1 0 61442 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0835_
timestamp 1607194113
transform 1 0 61626 0 -1 36496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_682
timestamp 1607194113
transform 1 0 63282 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B2
timestamp 1607194113
transform 1 0 63098 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_707
timestamp 1607194113
transform 1 0 65582 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_703
timestamp 1607194113
transform 1 0 65214 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_694
timestamp 1607194113
transform 1 0 64386 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A
timestamp 1607194113
transform 1 0 65674 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1607194113
transform 1 0 65122 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1183_
timestamp 1607194113
transform 1 0 65858 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_726
timestamp 1607194113
transform 1 0 67330 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_714
timestamp 1607194113
transform 1 0 66226 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1437_
timestamp 1607194113
transform 1 0 67422 0 -1 36496
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_748
timestamp 1607194113
transform 1 0 69354 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__CLK
timestamp 1607194113
transform 1 0 69170 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_764
timestamp 1607194113
transform 1 0 70826 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_760
timestamp 1607194113
transform 1 0 70458 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1607194113
transform 1 0 70734 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_788
timestamp 1607194113
transform 1 0 73034 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_776
timestamp 1607194113
transform 1 0 71930 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_807
timestamp 1607194113
transform 1 0 74782 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1247_
timestamp 1607194113
transform 1 0 73310 0 -1 36496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_825
timestamp 1607194113
transform 1 0 76438 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_823
timestamp 1607194113
transform 1 0 76254 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_819
timestamp 1607194113
transform 1 0 75886 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1607194113
transform 1 0 76346 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_849
timestamp 1607194113
transform 1 0 78646 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_837
timestamp 1607194113
transform 1 0 77542 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_861
timestamp 1607194113
transform 1 0 79750 0 -1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A
timestamp 1607194113
transform 1 0 80302 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_668
timestamp 1607194113
transform 1 0 61994 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_660
timestamp 1607194113
transform 1 0 61258 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1607194113
transform 1 0 61718 0 1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_653
timestamp 1607194113
transform 1 0 60614 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A1_N
timestamp 1607194113
transform 1 0 61074 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_688
timestamp 1607194113
transform 1 0 63834 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_676
timestamp 1607194113
transform 1 0 62730 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_672
timestamp 1607194113
transform 1 0 62362 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__CLK
timestamp 1607194113
transform 1 0 62270 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1607194113
transform 1 0 62270 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1391_
timestamp 1607194113
transform 1 0 62454 0 -1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1607194113
transform 1 0 62454 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1607194113
transform 1 0 64018 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_703
timestamp 1607194113
transform 1 0 65214 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_700
timestamp 1607194113
transform 1 0 64938 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_692
timestamp 1607194113
transform 1 0 64202 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_705
timestamp 1607194113
transform 1 0 65398 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_693
timestamp 1607194113
transform 1 0 64294 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1607194113
transform 1 0 65122 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_730
timestamp 1607194113
transform 1 0 67698 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_715
timestamp 1607194113
transform 1 0 66318 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_729
timestamp 1607194113
transform 1 0 67606 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_717
timestamp 1607194113
transform 1 0 66502 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0886_
timestamp 1607194113
transform 1 0 66410 0 -1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_67_749
timestamp 1607194113
transform 1 0 69446 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1607194113
transform 1 0 67882 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1248_
timestamp 1607194113
transform 1 0 68434 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1185_
timestamp 1607194113
transform 1 0 67974 0 1 36496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_764
timestamp 1607194113
transform 1 0 70826 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_762
timestamp 1607194113
transform 1 0 70642 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_754
timestamp 1607194113
transform 1 0 69906 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_761
timestamp 1607194113
transform 1 0 70550 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1607194113
transform 1 0 70734 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_776
timestamp 1607194113
transform 1 0 71930 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_785
timestamp 1607194113
transform 1 0 72758 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_773
timestamp 1607194113
transform 1 0 71654 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_i_A
timestamp 1607194113
transform 1 0 73034 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0884_
timestamp 1607194113
transform 1 0 72022 0 -1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_68_791
timestamp 1607194113
transform 1 0 73310 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_800
timestamp 1607194113
transform 1 0 74138 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1607194113
transform 1 0 73954 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk_i
timestamp 1607194113
transform 1 0 73218 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1607194113
transform 1 0 73494 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1187_
timestamp 1607194113
transform 1 0 74046 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _0883_
timestamp 1607194113
transform 1 0 73586 0 1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_825
timestamp 1607194113
transform 1 0 76438 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_823
timestamp 1607194113
transform 1 0 76254 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_815
timestamp 1607194113
transform 1 0 75518 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_824
timestamp 1607194113
transform 1 0 76346 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_820
timestamp 1607194113
transform 1 0 75978 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_812
timestamp 1607194113
transform 1 0 75242 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk_i
timestamp 1607194113
transform 1 0 76070 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1607194113
transform 1 0 76346 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_833
timestamp 1607194113
transform 1 0 77174 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_848
timestamp 1607194113
transform 1 0 78554 0 1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_836
timestamp 1607194113
transform 1 0 77450 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__CLK
timestamp 1607194113
transform 1 0 77450 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1395_
timestamp 1607194113
transform 1 0 77634 0 -1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_68_865
timestamp 1607194113
transform 1 0 80118 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_857
timestamp 1607194113
transform 1 0 79382 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_858
timestamp 1607194113
transform 1 0 79474 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1607194113
transform 1 0 80302 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1607194113
transform 1 0 79106 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1607194113
transform 1 0 79198 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_663
timestamp 1607194113
transform 1 0 61534 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_69_657
timestamp 1607194113
transform 1 0 60982 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__CLK
timestamp 1607194113
transform 1 0 62086 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1607194113
transform 1 0 61258 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1607194113
transform 1 0 62270 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1431_
timestamp 1607194113
transform 1 0 62362 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_703
timestamp 1607194113
transform 1 0 65214 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_691
timestamp 1607194113
transform 1 0 64110 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_727
timestamp 1607194113
transform 1 0 67422 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_715
timestamp 1607194113
transform 1 0 66318 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_731
timestamp 1607194113
transform 1 0 67790 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1607194113
transform 1 0 67882 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1434_
timestamp 1607194113
transform 1 0 67974 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_766
timestamp 1607194113
transform 1 0 71010 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_754
timestamp 1607194113
transform 1 0 69906 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__CLK
timestamp 1607194113
transform 1 0 69722 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_785
timestamp 1607194113
transform 1 0 72758 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_778
timestamp 1607194113
transform 1 0 72114 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1607194113
transform 1 0 72206 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0882_
timestamp 1607194113
transform 1 0 72390 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_794
timestamp 1607194113
transform 1 0 73586 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B2
timestamp 1607194113
transform 1 0 73862 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1607194113
transform 1 0 73494 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1250_
timestamp 1607194113
transform 1 0 74046 0 1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_826
timestamp 1607194113
transform 1 0 76530 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_815
timestamp 1607194113
transform 1 0 75518 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk_i
timestamp 1607194113
transform 1 0 76254 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_838
timestamp 1607194113
transform 1 0 77634 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_858
timestamp 1607194113
transform 1 0 79474 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_850
timestamp 1607194113
transform 1 0 78738 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1607194113
transform 1 0 79106 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1607194113
transform 1 0 79198 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_669
timestamp 1607194113
transform 1 0 62086 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_688
timestamp 1607194113
transform 1 0 63834 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_681
timestamp 1607194113
transform 1 0 63190 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A
timestamp 1607194113
transform 1 0 63282 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1249_
timestamp 1607194113
transform 1 0 63466 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_703
timestamp 1607194113
transform 1 0 65214 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_700
timestamp 1607194113
transform 1 0 64938 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1607194113
transform 1 0 65122 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_715
timestamp 1607194113
transform 1 0 66318 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _1189_
timestamp 1607194113
transform 1 0 66870 0 -1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_748
timestamp 1607194113
transform 1 0 69354 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_739
timestamp 1607194113
transform 1 0 68526 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A1_N
timestamp 1607194113
transform 1 0 68342 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1607194113
transform 1 0 69078 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_764
timestamp 1607194113
transform 1 0 70826 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_760
timestamp 1607194113
transform 1 0 70458 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1607194113
transform 1 0 70734 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_784
timestamp 1607194113
transform 1 0 72666 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_776
timestamp 1607194113
transform 1 0 71930 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A
timestamp 1607194113
transform 1 0 72114 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1186_
timestamp 1607194113
transform 1 0 72298 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_806
timestamp 1607194113
transform 1 0 74690 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0888_
timestamp 1607194113
transform 1 0 73402 0 -1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_70_825
timestamp 1607194113
transform 1 0 76438 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_818
timestamp 1607194113
transform 1 0 75794 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1607194113
transform 1 0 76346 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_833
timestamp 1607194113
transform 1 0 77174 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__CLK
timestamp 1607194113
transform 1 0 77266 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1436_
timestamp 1607194113
transform 1 0 77450 0 -1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_866
timestamp 1607194113
transform 1 0 80210 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_855
timestamp 1607194113
transform 1 0 79198 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1607194113
transform 1 0 79934 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_670
timestamp 1607194113
transform 1 0 62178 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_666
timestamp 1607194113
transform 1 0 61810 0 1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_654
timestamp 1607194113
transform 1 0 60706 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_684
timestamp 1607194113
transform 1 0 63466 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_672
timestamp 1607194113
transform 1 0 62362 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A2_N
timestamp 1607194113
transform 1 0 63742 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__B2
timestamp 1607194113
transform 1 0 63926 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1607194113
transform 1 0 62270 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_707
timestamp 1607194113
transform 1 0 65582 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1252_
timestamp 1607194113
transform 1 0 64110 0 1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_71_723
timestamp 1607194113
transform 1 0 67054 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_719
timestamp 1607194113
transform 1 0 66686 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1607194113
transform 1 0 66778 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_749
timestamp 1607194113
transform 1 0 69446 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_731
timestamp 1607194113
transform 1 0 67790 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1
timestamp 1607194113
transform 1 0 69262 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1607194113
transform 1 0 67882 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0894_
timestamp 1607194113
transform 1 0 67974 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_71_761
timestamp 1607194113
transform 1 0 70550 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_785
timestamp 1607194113
transform 1 0 72758 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_773
timestamp 1607194113
transform 1 0 71654 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_794
timestamp 1607194113
transform 1 0 73586 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1607194113
transform 1 0 73494 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0892_
timestamp 1607194113
transform 1 0 73770 0 1 38672
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_71_818
timestamp 1607194113
transform 1 0 75794 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_810
timestamp 1607194113
transform 1 0 75058 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B1
timestamp 1607194113
transform 1 0 75978 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1188_
timestamp 1607194113
transform 1 0 76162 0 1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_71_838
timestamp 1607194113
transform 1 0 77634 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_850
timestamp 1607194113
transform 1 0 78738 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__CLK
timestamp 1607194113
transform 1 0 78922 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1607194113
transform 1 0 79106 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1435_
timestamp 1607194113
transform 1 0 79198 0 1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_72_666
timestamp 1607194113
transform 1 0 61810 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_654
timestamp 1607194113
transform 1 0 60706 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_690
timestamp 1607194113
transform 1 0 64018 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_678
timestamp 1607194113
transform 1 0 62914 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_698
timestamp 1607194113
transform 1 0 64754 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__CLK
timestamp 1607194113
transform 1 0 64938 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1607194113
transform 1 0 65122 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1393_
timestamp 1607194113
transform 1 0 65214 0 -1 39760
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_72_722
timestamp 1607194113
transform 1 0 66962 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0895_
timestamp 1607194113
transform 1 0 67698 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_739
timestamp 1607194113
transform 1 0 68526 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_770
timestamp 1607194113
transform 1 0 71378 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_751
timestamp 1607194113
transform 1 0 69630 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1607194113
transform 1 0 71194 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1607194113
transform 1 0 70734 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1607194113
transform 1 0 70826 0 -1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_782
timestamp 1607194113
transform 1 0 72482 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0889_
timestamp 1607194113
transform 1 0 72574 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_804
timestamp 1607194113
transform 1 0 74506 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_792
timestamp 1607194113
transform 1 0 73402 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_825
timestamp 1607194113
transform 1 0 76438 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_816
timestamp 1607194113
transform 1 0 75610 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1607194113
transform 1 0 76346 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__CLK
timestamp 1607194113
transform 1 0 77174 0 -1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1394_
timestamp 1607194113
transform 1 0 77358 0 -1 39760
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_72_866
timestamp 1607194113
transform 1 0 80210 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_854
timestamp 1607194113
transform 1 0 79106 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_669
timestamp 1607194113
transform 1 0 62086 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_661
timestamp 1607194113
transform 1 0 61350 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_688
timestamp 1607194113
transform 1 0 63834 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_676
timestamp 1607194113
transform 1 0 62730 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_672
timestamp 1607194113
transform 1 0 62362 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1607194113
transform 1 0 62270 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1607194113
transform 1 0 62454 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_700
timestamp 1607194113
transform 1 0 64938 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_724
timestamp 1607194113
transform 1 0 67146 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_712
timestamp 1607194113
transform 1 0 66042 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_742
timestamp 1607194113
transform 1 0 68802 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1607194113
transform 1 0 67882 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0887_
timestamp 1607194113
transform 1 0 67974 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_73_754
timestamp 1607194113
transform 1 0 69906 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _0885_
timestamp 1607194113
transform 1 0 71010 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_73_787
timestamp 1607194113
transform 1 0 72942 0 1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_775
timestamp 1607194113
transform 1 0 71838 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_803
timestamp 1607194113
transform 1 0 74414 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1607194113
transform 1 0 73494 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0893_
timestamp 1607194113
transform 1 0 73586 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A2_N
timestamp 1607194113
transform 1 0 75150 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B2
timestamp 1607194113
transform 1 0 75334 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B1
timestamp 1607194113
transform 1 0 75518 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1251_
timestamp 1607194113
transform 1 0 75702 0 1 39760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_73_844
timestamp 1607194113
transform 1 0 78186 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_833
timestamp 1607194113
transform 1 0 77174 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1607194113
transform 1 0 77910 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_867
timestamp 1607194113
transform 1 0 80302 0 1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_855
timestamp 1607194113
transform 1 0 79198 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_852
timestamp 1607194113
transform 1 0 78922 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1607194113
transform 1 0 79106 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_665
timestamp 1607194113
transform 1 0 61718 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_654
timestamp 1607194113
transform 1 0 60706 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__CLK
timestamp 1607194113
transform 1 0 62086 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1607194113
transform 1 0 60890 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A1_N
timestamp 1607194113
transform 1 0 61534 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1429_
timestamp 1607194113
transform 1 0 61074 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_688
timestamp 1607194113
transform 1 0 63834 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_677
timestamp 1607194113
transform 1 0 62822 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1607194113
transform 1 0 62270 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1430_
timestamp 1607194113
transform 1 0 62362 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1607194113
transform 1 0 63558 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_703
timestamp 1607194113
transform 1 0 65214 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_691
timestamp 1607194113
transform 1 0 64110 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_703
timestamp 1607194113
transform 1 0 65214 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_700
timestamp 1607194113
transform 1 0 64938 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1607194113
transform 1 0 65122 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_727
timestamp 1607194113
transform 1 0 67422 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_715
timestamp 1607194113
transform 1 0 66318 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_715
timestamp 1607194113
transform 1 0 66318 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1508_
timestamp 1607194113
transform 1 0 66502 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_745
timestamp 1607194113
transform 1 0 69078 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_733
timestamp 1607194113
transform 1 0 67974 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_731
timestamp 1607194113
transform 1 0 67790 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_750
timestamp 1607194113
transform 1 0 69538 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_738
timestamp 1607194113
transform 1 0 68434 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__CLK
timestamp 1607194113
transform 1 0 68250 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1607194113
transform 1 0 67882 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_769
timestamp 1607194113
transform 1 0 71286 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_757
timestamp 1607194113
transform 1 0 70182 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_762
timestamp 1607194113
transform 1 0 70642 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1607194113
transform 1 0 70734 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1512_
timestamp 1607194113
transform 1 0 70826 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_781
timestamp 1607194113
transform 1 0 72390 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_785
timestamp 1607194113
transform 1 0 72758 0 -1 40848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__CLK
timestamp 1607194113
transform 1 0 72574 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1607194113
transform 1 0 73494 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1510_
timestamp 1607194113
transform 1 0 73586 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1509_
timestamp 1607194113
transform 1 0 73310 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_827
timestamp 1607194113
transform 1 0 76622 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_815
timestamp 1607194113
transform 1 0 75518 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_825
timestamp 1607194113
transform 1 0 76438 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_812
timestamp 1607194113
transform 1 0 75242 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__CLK
timestamp 1607194113
transform 1 0 75334 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__CLK
timestamp 1607194113
transform 1 0 75058 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1607194113
transform 1 0 76346 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_839
timestamp 1607194113
transform 1 0 77726 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_837
timestamp 1607194113
transform 1 0 77542 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__CLK
timestamp 1607194113
transform 1 0 77818 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__D
timestamp 1607194113
transform 1 0 78002 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1347_
timestamp 1607194113
transform 1 0 78186 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_75_867
timestamp 1607194113
transform 1 0 80302 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_855
timestamp 1607194113
transform 1 0 79198 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_851
timestamp 1607194113
transform 1 0 78830 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_863
timestamp 1607194113
transform 1 0 79934 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1607194113
transform 1 0 79106 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_664
timestamp 1607194113
transform 1 0 61626 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_652
timestamp 1607194113
transform 1 0 60522 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_683
timestamp 1607194113
transform 1 0 63374 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_676
timestamp 1607194113
transform 1 0 62730 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1607194113
transform 1 0 63282 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_707
timestamp 1607194113
transform 1 0 65582 0 -1 41936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_695
timestamp 1607194113
transform 1 0 64478 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__CLK
timestamp 1607194113
transform 1 0 65950 0 -1 41936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1607194113
transform 1 0 66134 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1511_
timestamp 1607194113
transform 1 0 66226 0 -1 41936
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_76_745
timestamp 1607194113
transform 1 0 69078 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_741
timestamp 1607194113
transform 1 0 68710 0 -1 41936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_733
timestamp 1607194113
transform 1 0 67974 0 -1 41936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1607194113
transform 1 0 68986 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_769
timestamp 1607194113
transform 1 0 71286 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_757
timestamp 1607194113
transform 1 0 70182 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_788
timestamp 1607194113
transform 1 0 73034 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_776
timestamp 1607194113
transform 1 0 71930 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1607194113
transform 1 0 71838 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_807
timestamp 1607194113
transform 1 0 74782 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_800
timestamp 1607194113
transform 1 0 74138 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1607194113
transform 1 0 74690 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_819
timestamp 1607194113
transform 1 0 75886 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_838
timestamp 1607194113
transform 1 0 77634 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_831
timestamp 1607194113
transform 1 0 76990 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1607194113
transform 1 0 77542 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_862
timestamp 1607194113
transform 1 0 79842 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_850
timestamp 1607194113
transform 1 0 78738 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1607194113
transform 1 0 80394 0 -1 41936
box -38 -48 130 592
use delayline_9_hd_25_1  inst_rdelay_line
timestamp 1607276668
transform 1 0 69814 0 1 1472
box 800 800 20764 22385
use sky130_fd_sc_hd__decap_12  FILLER_49_886
timestamp 1607194113
transform 1 0 82050 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_874
timestamp 1607194113
transform 1 0 80946 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_898
timestamp 1607194113
transform 1 0 83154 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_925
timestamp 1607194113
transform 1 0 85638 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_914
timestamp 1607194113
transform 1 0 84626 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_910
timestamp 1607194113
transform 1 0 84258 0 1 26704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1607194113
transform 1 0 85454 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607194113
transform 1 0 84718 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1071_
timestamp 1607194113
transform 1 0 84810 0 1 26704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_49_929
timestamp 1607194113
transform 1 0 86006 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__CLK
timestamp 1607194113
transform 1 0 86098 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1480_
timestamp 1607194113
transform 1 0 86282 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_963
timestamp 1607194113
transform 1 0 89134 0 1 26704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_951
timestamp 1607194113
transform 1 0 88030 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_971
timestamp 1607194113
transform 1 0 89870 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__CLK
timestamp 1607194113
transform 1 0 90146 0 1 26704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607194113
transform 1 0 90330 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1481_
timestamp 1607194113
transform 1 0 90422 0 1 26704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_49_996
timestamp 1607194113
transform 1 0 92170 0 1 26704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1008
timestamp 1607194113
transform 1 0 93274 0 1 26704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1607194113
transform -1 0 93642 0 1 26704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_884
timestamp 1607194113
transform 1 0 81866 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_880
timestamp 1607194113
transform 1 0 81498 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607194113
transform 1 0 81958 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1607194113
transform 1 0 82050 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_897
timestamp 1607194113
transform 1 0 83062 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_889
timestamp 1607194113
transform 1 0 82326 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1607194113
transform 1 0 83982 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1051_
timestamp 1607194113
transform 1 0 83154 0 -1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_909
timestamp 1607194113
transform 1 0 84166 0 -1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B1
timestamp 1607194113
transform 1 0 84534 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1073_
timestamp 1607194113
transform 1 0 84718 0 -1 27792
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_50_940
timestamp 1607194113
transform 1 0 87018 0 -1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_928
timestamp 1607194113
transform 1 0 85914 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607194113
transform 1 0 87570 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1607194113
transform 1 0 87662 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_967
timestamp 1607194113
transform 1 0 89502 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_962
timestamp 1607194113
transform 1 0 89042 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_950
timestamp 1607194113
transform 1 0 87938 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1607194113
transform 1 0 89226 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_982
timestamp 1607194113
transform 1 0 90882 0 -1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1062_
timestamp 1607194113
transform 1 0 90238 0 -1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_50_1005
timestamp 1607194113
transform 1 0 92998 0 -1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_993
timestamp 1607194113
transform 1 0 91894 0 -1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1607194113
transform 1 0 91618 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1008
timestamp 1607194113
transform 1 0 93274 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607194113
transform 1 0 93182 0 -1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1607194113
transform -1 0 93642 0 -1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_886
timestamp 1607194113
transform 1 0 82050 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_877
timestamp 1607194113
transform 1 0 81222 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_887
timestamp 1607194113
transform 1 0 82142 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_872
timestamp 1607194113
transform 1 0 80762 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B
timestamp 1607194113
transform 1 0 81314 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607194113
transform 1 0 81958 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1033_
timestamp 1607194113
transform 1 0 81498 0 1 27792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_52_906
timestamp 1607194113
transform 1 0 83890 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_898
timestamp 1607194113
transform 1 0 83154 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_907
timestamp 1607194113
transform 1 0 83982 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_895
timestamp 1607194113
transform 1 0 82878 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1607194113
transform 1 0 82970 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1076_
timestamp 1607194113
transform 1 0 83154 0 1 27792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_51_916
timestamp 1607194113
transform 1 0 84810 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__CLK
timestamp 1607194113
transform 1 0 84074 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607194113
transform 1 0 84718 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1479_
timestamp 1607194113
transform 1 0 84258 0 -1 28880
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1074_
timestamp 1607194113
transform 1 0 85086 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_947
timestamp 1607194113
transform 1 0 87662 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_945
timestamp 1607194113
transform 1 0 87478 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_941
timestamp 1607194113
transform 1 0 87110 0 -1 28880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_929
timestamp 1607194113
transform 1 0 86006 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_943
timestamp 1607194113
transform 1 0 87294 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_931
timestamp 1607194113
transform 1 0 86190 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607194113
transform 1 0 87570 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_959
timestamp 1607194113
transform 1 0 88766 0 -1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_963
timestamp 1607194113
transform 1 0 89134 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_955
timestamp 1607194113
transform 1 0 88398 0 1 27792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1607194113
transform 1 0 89318 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_982
timestamp 1607194113
transform 1 0 90882 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_971
timestamp 1607194113
transform 1 0 89870 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_970
timestamp 1607194113
transform 1 0 89778 0 1 27792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1607194113
transform 1 0 89594 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B1
timestamp 1607194113
transform 1 0 90146 0 1 27792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607194113
transform 1 0 90330 0 1 27792
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1067_
timestamp 1607194113
transform 1 0 90422 0 1 27792
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_4  _1052_
timestamp 1607194113
transform 1 0 90054 0 -1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_52_1005
timestamp 1607194113
transform 1 0 92998 0 -1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_997
timestamp 1607194113
transform 1 0 92262 0 -1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1003
timestamp 1607194113
transform 1 0 92814 0 1 27792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_991
timestamp 1607194113
transform 1 0 91710 0 1 27792
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1064_
timestamp 1607194113
transform 1 0 91618 0 -1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1008
timestamp 1607194113
transform 1 0 93274 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607194113
transform 1 0 93182 0 -1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1607194113
transform -1 0 93642 0 -1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1607194113
transform -1 0 93642 0 1 27792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_882
timestamp 1607194113
transform 1 0 81682 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1607194113
transform 1 0 80854 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1078_
timestamp 1607194113
transform 1 0 81038 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_53_906
timestamp 1607194113
transform 1 0 83890 0 1 28880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_894
timestamp 1607194113
transform 1 0 82786 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_925
timestamp 1607194113
transform 1 0 85638 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_912
timestamp 1607194113
transform 1 0 84442 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1607194113
transform 1 0 84534 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607194113
transform 1 0 84718 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1075_
timestamp 1607194113
transform 1 0 84810 0 1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_53_942
timestamp 1607194113
transform 1 0 87202 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A
timestamp 1607194113
transform 1 0 87018 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1055_
timestamp 1607194113
transform 1 0 86374 0 1 28880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_53_966
timestamp 1607194113
transform 1 0 89410 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_954
timestamp 1607194113
transform 1 0 88306 0 1 28880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_987
timestamp 1607194113
transform 1 0 91342 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_977
timestamp 1607194113
transform 1 0 90422 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1607194113
transform 1 0 90146 0 1 28880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607194113
transform 1 0 90330 0 1 28880
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1066_
timestamp 1607194113
transform 1 0 90514 0 1 28880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_53_1006
timestamp 1607194113
transform 1 0 93090 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_998
timestamp 1607194113
transform 1 0 92354 0 1 28880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1607194113
transform 1 0 92078 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1607194113
transform -1 0 93642 0 1 28880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_886
timestamp 1607194113
transform 1 0 82050 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_883
timestamp 1607194113
transform 1 0 81774 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_871
timestamp 1607194113
transform 1 0 80670 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__CLK
timestamp 1607194113
transform 1 0 80578 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607194113
transform 1 0 81958 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1476_
timestamp 1607194113
transform 1 0 80762 0 1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_55_903
timestamp 1607194113
transform 1 0 83614 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_891
timestamp 1607194113
transform 1 0 82510 0 1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_906
timestamp 1607194113
transform 1 0 83890 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_898
timestamp 1607194113
transform 1 0 83154 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_916
timestamp 1607194113
transform 1 0 84810 0 1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_914
timestamp 1607194113
transform 1 0 84626 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A
timestamp 1607194113
transform 1 0 84442 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607194113
transform 1 0 84718 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1607194113
transform 1 0 84166 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_922
timestamp 1607194113
transform 1 0 85362 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__CLK
timestamp 1607194113
transform 1 0 85178 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1607194113
transform 1 0 85638 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1057_
timestamp 1607194113
transform 1 0 85822 0 -1 29968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1484_
timestamp 1607194113
transform 1 0 85362 0 1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_55_941
timestamp 1607194113
transform 1 0 87110 0 1 29968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_944
timestamp 1607194113
transform 1 0 87386 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_936
timestamp 1607194113
transform 1 0 86650 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 1607194113
transform 1 0 87662 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607194113
transform 1 0 87570 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1607194113
transform 1 0 87662 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_965
timestamp 1607194113
transform 1 0 89318 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_962
timestamp 1607194113
transform 1 0 89042 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_950
timestamp 1607194113
transform 1 0 87938 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1607194113
transform 1 0 89134 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1060_
timestamp 1607194113
transform 1 0 87846 0 1 29968
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_55_977
timestamp 1607194113
transform 1 0 90422 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_973
timestamp 1607194113
transform 1 0 90054 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_985
timestamp 1607194113
transform 1 0 91158 0 -1 29968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_974
timestamp 1607194113
transform 1 0 90146 0 -1 29968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__CLK
timestamp 1607194113
transform 1 0 90514 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607194113
transform 1 0 90330 0 1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1482_
timestamp 1607194113
transform 1 0 90698 0 1 29968
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1065_
timestamp 1607194113
transform 1 0 90514 0 -1 29968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_55_999
timestamp 1607194113
transform 1 0 92446 0 1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_1005
timestamp 1607194113
transform 1 0 92998 0 -1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_997
timestamp 1607194113
transform 1 0 92262 0 -1 29968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1007
timestamp 1607194113
transform 1 0 93182 0 1 29968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1008
timestamp 1607194113
transform 1 0 93274 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607194113
transform 1 0 93182 0 -1 29968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1607194113
transform -1 0 93642 0 1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1607194113
transform -1 0 93642 0 -1 29968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_877
timestamp 1607194113
transform 1 0 81222 0 -1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607194113
transform 1 0 81958 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1607194113
transform 1 0 82050 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_901
timestamp 1607194113
transform 1 0 83430 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_889
timestamp 1607194113
transform 1 0 82326 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_920
timestamp 1607194113
transform 1 0 85178 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_913
timestamp 1607194113
transform 1 0 84534 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A
timestamp 1607194113
transform 1 0 84994 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1056_
timestamp 1607194113
transform 1 0 85730 0 -1 31056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1607194113
transform 1 0 84718 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_947
timestamp 1607194113
transform 1 0 87662 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_945
timestamp 1607194113
transform 1 0 87478 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_933
timestamp 1607194113
transform 1 0 86374 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607194113
transform 1 0 87570 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_962
timestamp 1607194113
transform 1 0 89042 0 -1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1607194113
transform 1 0 88858 0 -1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1053_
timestamp 1607194113
transform 1 0 88214 0 -1 31056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_56_983
timestamp 1607194113
transform 1 0 90974 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_971
timestamp 1607194113
transform 1 0 89870 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1607194113
transform 1 0 89594 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0767_
timestamp 1607194113
transform 1 0 91342 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_1003
timestamp 1607194113
transform 1 0 92814 0 -1 31056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_991
timestamp 1607194113
transform 1 0 91710 0 -1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1008
timestamp 1607194113
transform 1 0 93274 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607194113
transform 1 0 93182 0 -1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1607194113
transform -1 0 93642 0 -1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_884
timestamp 1607194113
transform 1 0 81866 0 1 31056
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__B1
timestamp 1607194113
transform 1 0 80486 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1086_
timestamp 1607194113
transform 1 0 80670 0 1 31056
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_57_901
timestamp 1607194113
transform 1 0 83430 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0851_
timestamp 1607194113
transform 1 0 82602 0 1 31056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_916
timestamp 1607194113
transform 1 0 84810 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_913
timestamp 1607194113
transform 1 0 84534 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607194113
transform 1 0 84718 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_940
timestamp 1607194113
transform 1 0 87018 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_928
timestamp 1607194113
transform 1 0 85914 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_957
timestamp 1607194113
transform 1 0 88582 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_952
timestamp 1607194113
transform 1 0 88122 0 1 31056
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1607194113
transform 1 0 88306 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_977
timestamp 1607194113
transform 1 0 90422 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_975
timestamp 1607194113
transform 1 0 90238 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_969
timestamp 1607194113
transform 1 0 89686 0 1 31056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607194113
transform 1 0 90330 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0844_
timestamp 1607194113
transform 1 0 90698 0 1 31056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_996
timestamp 1607194113
transform 1 0 92170 0 1 31056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1008
timestamp 1607194113
transform 1 0 93274 0 1 31056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1607194113
transform -1 0 93642 0 1 31056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_886
timestamp 1607194113
transform 1 0 82050 0 -1 32144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_884
timestamp 1607194113
transform 1 0 81866 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_872
timestamp 1607194113
transform 1 0 80762 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607194113
transform 1 0 81958 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0850_
timestamp 1607194113
transform 1 0 80854 0 1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_59_906
timestamp 1607194113
transform 1 0 83890 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_889
timestamp 1607194113
transform 1 0 82326 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_892
timestamp 1607194113
transform 1 0 82602 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A2_N
timestamp 1607194113
transform 1 0 82694 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A1_N
timestamp 1607194113
transform 1 0 82878 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0848_
timestamp 1607194113
transform 1 0 83062 0 -1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _0776_
timestamp 1607194113
transform 1 0 83062 0 1 32144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_59_916
timestamp 1607194113
transform 1 0 84810 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_914
timestamp 1607194113
transform 1 0 84626 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_925
timestamp 1607194113
transform 1 0 85638 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_913
timestamp 1607194113
transform 1 0 84534 0 -1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607194113
transform 1 0 84718 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_933
timestamp 1607194113
transform 1 0 86374 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_928
timestamp 1607194113
transform 1 0 85914 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_937
timestamp 1607194113
transform 1 0 86742 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1607194113
transform 1 0 86098 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_941
timestamp 1607194113
transform 1 0 87110 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_947
timestamp 1607194113
transform 1 0 87662 0 -1 32144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_945
timestamp 1607194113
transform 1 0 87478 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__CLK
timestamp 1607194113
transform 1 0 87294 0 1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607194113
transform 1 0 87570 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1443_
timestamp 1607194113
transform 1 0 87478 0 1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_964
timestamp 1607194113
transform 1 0 89226 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_951
timestamp 1607194113
transform 1 0 88030 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__CLK
timestamp 1607194113
transform 1 0 88122 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1483_
timestamp 1607194113
transform 1 0 88306 0 -1 32144
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_977
timestamp 1607194113
transform 1 0 90422 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_973
timestamp 1607194113
transform 1 0 90054 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607194113
transform 1 0 90330 0 1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0768_
timestamp 1607194113
transform 1 0 90790 0 -1 32144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1001
timestamp 1607194113
transform 1 0 92630 0 1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_989
timestamp 1607194113
transform 1 0 91526 0 1 32144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_1005
timestamp 1607194113
transform 1 0 92998 0 -1 32144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_997
timestamp 1607194113
transform 1 0 92262 0 -1 32144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1008
timestamp 1607194113
transform 1 0 93274 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607194113
transform 1 0 93182 0 -1 32144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1607194113
transform -1 0 93642 0 1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1607194113
transform -1 0 93642 0 -1 32144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_886
timestamp 1607194113
transform 1 0 82050 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_882
timestamp 1607194113
transform 1 0 81682 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_874
timestamp 1607194113
transform 1 0 80946 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607194113
transform 1 0 81958 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_892
timestamp 1607194113
transform 1 0 82602 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A2_N
timestamp 1607194113
transform 1 0 82694 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1_N
timestamp 1607194113
transform 1 0 82878 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0773_
timestamp 1607194113
transform 1 0 83062 0 -1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_925
timestamp 1607194113
transform 1 0 85638 0 -1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_913
timestamp 1607194113
transform 1 0 84534 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_938
timestamp 1607194113
transform 1 0 86834 0 -1 33232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_933
timestamp 1607194113
transform 1 0 86374 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__CLK
timestamp 1607194113
transform 1 0 87386 0 -1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607194113
transform 1 0 87570 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1402_
timestamp 1607194113
transform 1 0 87662 0 -1 33232
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1607194113
transform 1 0 86558 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_966
timestamp 1607194113
transform 1 0 89410 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_978
timestamp 1607194113
transform 1 0 90514 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1006
timestamp 1607194113
transform 1 0 93090 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1002
timestamp 1607194113
transform 1 0 92722 0 -1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_990
timestamp 1607194113
transform 1 0 91618 0 -1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1008
timestamp 1607194113
transform 1 0 93274 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607194113
transform 1 0 93182 0 -1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1607194113
transform -1 0 93642 0 -1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_871
timestamp 1607194113
transform 1 0 80670 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _0775_
timestamp 1607194113
transform 1 0 81406 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_61_907
timestamp 1607194113
transform 1 0 83982 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_895
timestamp 1607194113
transform 1 0 82878 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_924
timestamp 1607194113
transform 1 0 85546 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_916
timestamp 1607194113
transform 1 0 84810 0 1 33232
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A2_N
timestamp 1607194113
transform 1 0 85638 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B2
timestamp 1607194113
transform 1 0 85822 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1607194113
transform 1 0 84718 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1_N
timestamp 1607194113
transform 1 0 87662 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B1
timestamp 1607194113
transform 1 0 86006 0 1 33232
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1175_
timestamp 1607194113
transform 1 0 86190 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_61_961
timestamp 1607194113
transform 1 0 88950 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_949
timestamp 1607194113
transform 1 0 87846 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_973
timestamp 1607194113
transform 1 0 90054 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1607194113
transform 1 0 90330 0 1 33232
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0719_
timestamp 1607194113
transform 1 0 90422 0 1 33232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_1005
timestamp 1607194113
transform 1 0 92998 0 1 33232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_993
timestamp 1607194113
transform 1 0 91894 0 1 33232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1607194113
transform -1 0 93642 0 1 33232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_880
timestamp 1607194113
transform 1 0 81498 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_886
timestamp 1607194113
transform 1 0 82050 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_877
timestamp 1607194113
transform 1 0 81222 0 -1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_869
timestamp 1607194113
transform 1 0 80486 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A
timestamp 1607194113
transform 1 0 81038 0 -1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1607194113
transform 1 0 81958 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1607194113
transform 1 0 80762 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_898
timestamp 1607194113
transform 1 0 83154 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_892
timestamp 1607194113
transform 1 0 82602 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_898
timestamp 1607194113
transform 1 0 83154 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1607194113
transform 1 0 82970 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1607194113
transform 1 0 82694 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_924
timestamp 1607194113
transform 1 0 85546 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_916
timestamp 1607194113
transform 1 0 84810 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_914
timestamp 1607194113
transform 1 0 84626 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_910
timestamp 1607194113
transform 1 0 84258 0 1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_922
timestamp 1607194113
transform 1 0 85362 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_910
timestamp 1607194113
transform 1 0 84258 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B1
timestamp 1607194113
transform 1 0 85730 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1607194113
transform 1 0 84718 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_946
timestamp 1607194113
transform 1 0 87570 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_947
timestamp 1607194113
transform 1 0 87662 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_934
timestamp 1607194113
transform 1 0 86466 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1_N
timestamp 1607194113
transform 1 0 87386 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1607194113
transform 1 0 87570 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1239_
timestamp 1607194113
transform 1 0 85914 0 1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_958
timestamp 1607194113
transform 1 0 88674 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_959
timestamp 1607194113
transform 1 0 88766 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_987
timestamp 1607194113
transform 1 0 91342 0 1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_983
timestamp 1607194113
transform 1 0 90974 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_977
timestamp 1607194113
transform 1 0 90422 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_970
timestamp 1607194113
transform 1 0 89778 0 1 34320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_971
timestamp 1607194113
transform 1 0 89870 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1607194113
transform 1 0 90330 0 1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1607194113
transform 1 0 91066 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0814_
timestamp 1607194113
transform 1 0 90238 0 -1 34320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_63_999
timestamp 1607194113
transform 1 0 92446 0 1 34320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1003
timestamp 1607194113
transform 1 0 92814 0 -1 34320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_991
timestamp 1607194113
transform 1 0 91710 0 -1 34320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1007
timestamp 1607194113
transform 1 0 93182 0 1 34320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1008
timestamp 1607194113
transform 1 0 93274 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1607194113
transform 1 0 93182 0 -1 34320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1607194113
transform -1 0 93642 0 1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1607194113
transform -1 0 93642 0 -1 34320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_886
timestamp 1607194113
transform 1 0 82050 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_884
timestamp 1607194113
transform 1 0 81866 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_876
timestamp 1607194113
transform 1 0 81130 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1607194113
transform 1 0 81958 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_894
timestamp 1607194113
transform 1 0 82786 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__CLK
timestamp 1607194113
transform 1 0 83062 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1442_
timestamp 1607194113
transform 1 0 83246 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_918
timestamp 1607194113
transform 1 0 84994 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_947
timestamp 1607194113
transform 1 0 87662 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_942
timestamp 1607194113
transform 1 0 87202 0 -1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_930
timestamp 1607194113
transform 1 0 86098 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1607194113
transform 1 0 87570 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_959
timestamp 1607194113
transform 1 0 88766 0 -1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__CLK
timestamp 1607194113
transform 1 0 89502 0 -1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1400_
timestamp 1607194113
transform 1 0 89686 0 -1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1006
timestamp 1607194113
transform 1 0 93090 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1000
timestamp 1607194113
transform 1 0 92538 0 -1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_988
timestamp 1607194113
transform 1 0 91434 0 -1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1008
timestamp 1607194113
transform 1 0 93274 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1607194113
transform 1 0 93182 0 -1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1607194113
transform -1 0 93642 0 -1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_873
timestamp 1607194113
transform 1 0 80854 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_881
timestamp 1607194113
transform 1 0 81590 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_873
timestamp 1607194113
transform 1 0 80854 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A2_N
timestamp 1607194113
transform 1 0 81682 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B2
timestamp 1607194113
transform 1 0 81866 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1607194113
transform 1 0 81958 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1242_
timestamp 1607194113
transform 1 0 80486 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _1176_
timestamp 1607194113
transform 1 0 82050 0 1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0873_
timestamp 1607194113
transform 1 0 82050 0 -1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_66_900
timestamp 1607194113
transform 1 0 83338 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_902
timestamp 1607194113
transform 1 0 83522 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_924
timestamp 1607194113
transform 1 0 85546 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_912
timestamp 1607194113
transform 1 0 84442 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_920
timestamp 1607194113
transform 1 0 85178 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_916
timestamp 1607194113
transform 1 0 84810 0 1 35408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_914
timestamp 1607194113
transform 1 0 84626 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1607194113
transform 1 0 84718 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0871_
timestamp 1607194113
transform 1 0 85270 0 1 35408
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_66_947
timestamp 1607194113
transform 1 0 87662 0 -1 36496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_944
timestamp 1607194113
transform 1 0 87386 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_936
timestamp 1607194113
transform 1 0 86650 0 -1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_947
timestamp 1607194113
transform 1 0 87662 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_939
timestamp 1607194113
transform 1 0 86926 0 1 35408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B1
timestamp 1607194113
transform 1 0 86742 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1607194113
transform 1 0 86558 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1607194113
transform 1 0 87570 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A2_N
timestamp 1607194113
transform 1 0 88214 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B1
timestamp 1607194113
transform 1 0 88398 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B1
timestamp 1607194113
transform 1 0 87938 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1243_
timestamp 1607194113
transform 1 0 88122 0 1 35408
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1179_
timestamp 1607194113
transform 1 0 88582 0 -1 36496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_66_985
timestamp 1607194113
transform 1 0 91158 0 -1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_973
timestamp 1607194113
transform 1 0 90054 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_968
timestamp 1607194113
transform 1 0 89594 0 1 35408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__CLK
timestamp 1607194113
transform 1 0 90146 0 1 35408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1607194113
transform 1 0 90330 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1441_
timestamp 1607194113
transform 1 0 90422 0 1 35408
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1607194113
transform 1 0 91342 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1006
timestamp 1607194113
transform 1 0 93090 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_1002
timestamp 1607194113
transform 1 0 92722 0 -1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_990
timestamp 1607194113
transform 1 0 91618 0 -1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_996
timestamp 1607194113
transform 1 0 92170 0 1 35408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1008
timestamp 1607194113
transform 1 0 93274 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1008
timestamp 1607194113
transform 1 0 93274 0 1 35408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1607194113
transform 1 0 93182 0 -1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1607194113
transform -1 0 93642 0 -1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1607194113
transform -1 0 93642 0 1 35408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_878
timestamp 1607194113
transform 1 0 81314 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_870
timestamp 1607194113
transform 1 0 80578 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1607194113
transform 1 0 80762 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0865_
timestamp 1607194113
transform 1 0 80946 0 1 36496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_902
timestamp 1607194113
transform 1 0 83522 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_890
timestamp 1607194113
transform 1 0 82418 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_914
timestamp 1607194113
transform 1 0 84626 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1607194113
transform 1 0 84718 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0877_
timestamp 1607194113
transform 1 0 84810 0 1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_67_946
timestamp 1607194113
transform 1 0 87570 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_934
timestamp 1607194113
transform 1 0 86466 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B1
timestamp 1607194113
transform 1 0 86282 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A1
timestamp 1607194113
transform 1 0 86098 0 1 36496
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0875_
timestamp 1607194113
transform 1 0 88306 0 1 36496
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_67_977
timestamp 1607194113
transform 1 0 90422 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_968
timestamp 1607194113
transform 1 0 89594 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1607194113
transform 1 0 90330 0 1 36496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1001
timestamp 1607194113
transform 1 0 92630 0 1 36496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_989
timestamp 1607194113
transform 1 0 91526 0 1 36496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1607194113
transform -1 0 93642 0 1 36496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_873
timestamp 1607194113
transform 1 0 80854 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1607194113
transform 1 0 81958 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1178_
timestamp 1607194113
transform 1 0 82050 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0870_
timestamp 1607194113
transform 1 0 80486 0 -1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_904
timestamp 1607194113
transform 1 0 83706 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_892
timestamp 1607194113
transform 1 0 82602 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__CLK
timestamp 1607194113
transform 1 0 83798 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A
timestamp 1607194113
transform 1 0 82418 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1399_
timestamp 1607194113
transform 1 0 83982 0 -1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_68_926
timestamp 1607194113
transform 1 0 85730 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_947
timestamp 1607194113
transform 1 0 87662 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_945
timestamp 1607194113
transform 1 0 87478 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_937
timestamp 1607194113
transform 1 0 86742 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1607194113
transform 1 0 87570 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1607194113
transform 1 0 86466 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_955
timestamp 1607194113
transform 1 0 88398 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__B1
timestamp 1607194113
transform 1 0 88674 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1245_
timestamp 1607194113
transform 1 0 88858 0 -1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_68_984
timestamp 1607194113
transform 1 0 91066 0 -1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_976
timestamp 1607194113
transform 1 0 90330 0 -1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1607194113
transform 1 0 91250 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_1001
timestamp 1607194113
transform 1 0 92630 0 -1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_989
timestamp 1607194113
transform 1 0 91526 0 -1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1008
timestamp 1607194113
transform 1 0 93274 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1607194113
transform 1 0 93182 0 -1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1607194113
transform -1 0 93642 0 -1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_886
timestamp 1607194113
transform 1 0 82050 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_884
timestamp 1607194113
transform 1 0 81866 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_878
timestamp 1607194113
transform 1 0 81314 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_882
timestamp 1607194113
transform 1 0 81682 0 1 37584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_870
timestamp 1607194113
transform 1 0 80578 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1607194113
transform 1 0 81958 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_894
timestamp 1607194113
transform 1 0 82786 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_890
timestamp 1607194113
transform 1 0 82418 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A1_N
timestamp 1607194113
transform 1 0 83982 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1244_
timestamp 1607194113
transform 1 0 82510 0 1 37584
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1180_
timestamp 1607194113
transform 1 0 83062 0 -1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_924
timestamp 1607194113
transform 1 0 85546 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_915
timestamp 1607194113
transform 1 0 84718 0 -1 38672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_909
timestamp 1607194113
transform 1 0 84166 0 1 37584
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__CLK
timestamp 1607194113
transform 1 0 84534 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A1_N
timestamp 1607194113
transform 1 0 84534 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1607194113
transform 1 0 84718 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1440_
timestamp 1607194113
transform 1 0 84810 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1607194113
transform 1 0 85270 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_947
timestamp 1607194113
transform 1 0 87662 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_944
timestamp 1607194113
transform 1 0 87386 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_936
timestamp 1607194113
transform 1 0 86650 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_947
timestamp 1607194113
transform 1 0 87662 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_935
timestamp 1607194113
transform 1 0 86558 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1607194113
transform 1 0 87570 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_953
timestamp 1607194113
transform 1 0 88214 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__B1
timestamp 1607194113
transform 1 0 88766 0 -1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1181_
timestamp 1607194113
transform 1 0 88950 0 -1 38672
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0879_
timestamp 1607194113
transform 1 0 88306 0 1 37584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_70_985
timestamp 1607194113
transform 1 0 91158 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_977
timestamp 1607194113
transform 1 0 90422 0 -1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_968
timestamp 1607194113
transform 1 0 89594 0 1 37584
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__CLK
timestamp 1607194113
transform 1 0 90146 0 1 37584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1607194113
transform 1 0 90330 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1398_
timestamp 1607194113
transform 1 0 90422 0 1 37584
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_70_1003
timestamp 1607194113
transform 1 0 92814 0 -1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_991
timestamp 1607194113
transform 1 0 91710 0 -1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_996
timestamp 1607194113
transform 1 0 92170 0 1 37584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1607194113
transform 1 0 91434 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1008
timestamp 1607194113
transform 1 0 93274 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_1008
timestamp 1607194113
transform 1 0 93274 0 1 37584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1607194113
transform 1 0 93182 0 -1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1607194113
transform -1 0 93642 0 -1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1607194113
transform -1 0 93642 0 1 37584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_886
timestamp 1607194113
transform 1 0 82050 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_874
timestamp 1607194113
transform 1 0 80946 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_898
timestamp 1607194113
transform 1 0 83154 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_916
timestamp 1607194113
transform 1 0 84810 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_914
timestamp 1607194113
transform 1 0 84626 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_910
timestamp 1607194113
transform 1 0 84258 0 1 38672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1607194113
transform 1 0 84718 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_940
timestamp 1607194113
transform 1 0 87018 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_928
timestamp 1607194113
transform 1 0 85914 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_964
timestamp 1607194113
transform 1 0 89226 0 1 38672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_952
timestamp 1607194113
transform 1 0 88122 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_972
timestamp 1607194113
transform 1 0 89962 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__CLK
timestamp 1607194113
transform 1 0 90146 0 1 38672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1607194113
transform 1 0 90330 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1439_
timestamp 1607194113
transform 1 0 90422 0 1 38672
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_996
timestamp 1607194113
transform 1 0 92170 0 1 38672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_1008
timestamp 1607194113
transform 1 0 93274 0 1 38672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1607194113
transform -1 0 93642 0 1 38672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_886
timestamp 1607194113
transform 1 0 82050 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_884
timestamp 1607194113
transform 1 0 81866 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_878
timestamp 1607194113
transform 1 0 81314 0 -1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1607194113
transform 1 0 81958 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_898
timestamp 1607194113
transform 1 0 83154 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0878_
timestamp 1607194113
transform 1 0 83890 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_927
timestamp 1607194113
transform 1 0 85822 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_915
timestamp 1607194113
transform 1 0 84718 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_947
timestamp 1607194113
transform 1 0 87662 0 -1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_945
timestamp 1607194113
transform 1 0 87478 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_939
timestamp 1607194113
transform 1 0 86926 0 -1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1607194113
transform 1 0 87570 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_967
timestamp 1607194113
transform 1 0 89502 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_955
timestamp 1607194113
transform 1 0 88398 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0880_
timestamp 1607194113
transform 1 0 88674 0 -1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_979
timestamp 1607194113
transform 1 0 90606 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_1003
timestamp 1607194113
transform 1 0 92814 0 -1 39760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_991
timestamp 1607194113
transform 1 0 91710 0 -1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1008
timestamp 1607194113
transform 1 0 93274 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1607194113
transform 1 0 93182 0 -1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1607194113
transform -1 0 93642 0 -1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_877
timestamp 1607194113
transform 1 0 81222 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_873
timestamp 1607194113
transform 1 0 80854 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__CLK
timestamp 1607194113
transform 1 0 80946 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1607194113
transform 1 0 80670 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1607194113
transform 1 0 81958 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1516_
timestamp 1607194113
transform 1 0 81130 0 1 39760
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _0874_
timestamp 1607194113
transform 1 0 82050 0 -1 40848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1607194113
transform 1 0 80854 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_903
timestamp 1607194113
transform 1 0 83614 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_895
timestamp 1607194113
transform 1 0 82878 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_907
timestamp 1607194113
transform 1 0 83982 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_895
timestamp 1607194113
transform 1 0 82878 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__CLK
timestamp 1607194113
transform 1 0 83706 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1514_
timestamp 1607194113
transform 1 0 83890 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_925
timestamp 1607194113
transform 1 0 85638 0 -1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_916
timestamp 1607194113
transform 1 0 84810 0 1 39760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1607194113
transform 1 0 84718 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0872_
timestamp 1607194113
transform 1 0 85362 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_74_947
timestamp 1607194113
transform 1 0 87662 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_945
timestamp 1607194113
transform 1 0 87478 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_937
timestamp 1607194113
transform 1 0 86742 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_943
timestamp 1607194113
transform 1 0 87294 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_931
timestamp 1607194113
transform 1 0 86190 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1607194113
transform 1 0 87570 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_966
timestamp 1607194113
transform 1 0 89410 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_955
timestamp 1607194113
transform 1 0 88398 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__CLK
timestamp 1607194113
transform 1 0 88030 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1513_
timestamp 1607194113
transform 1 0 88214 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _0876_
timestamp 1607194113
transform 1 0 88582 0 1 39760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_74_972
timestamp 1607194113
transform 1 0 89962 0 -1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_977
timestamp 1607194113
transform 1 0 90422 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_974
timestamp 1607194113
transform 1 0 90146 0 1 39760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__CLK
timestamp 1607194113
transform 1 0 90330 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__D
timestamp 1607194113
transform 1 0 90514 0 -1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1607194113
transform 1 0 90330 0 1 39760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1348_
timestamp 1607194113
transform 1 0 90698 0 -1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_74_999
timestamp 1607194113
transform 1 0 92446 0 -1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_1001
timestamp 1607194113
transform 1 0 92630 0 1 39760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_989
timestamp 1607194113
transform 1 0 91526 0 1 39760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1008
timestamp 1607194113
transform 1 0 93274 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1607194113
transform 1 0 93182 0 -1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1607194113
transform -1 0 93642 0 -1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1607194113
transform -1 0 93642 0 1 39760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__CLK
timestamp 1607194113
transform 1 0 80670 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__D
timestamp 1607194113
transform 1 0 80854 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1485_
timestamp 1607194113
transform 1 0 81038 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_75_906
timestamp 1607194113
transform 1 0 83890 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_894
timestamp 1607194113
transform 1 0 82786 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_916
timestamp 1607194113
transform 1 0 84810 0 1 40848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_914
timestamp 1607194113
transform 1 0 84626 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__CLK
timestamp 1607194113
transform 1 0 85178 0 1 40848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1607194113
transform 1 0 84718 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1517_
timestamp 1607194113
transform 1 0 85362 0 1 40848
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_941
timestamp 1607194113
transform 1 0 87110 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_965
timestamp 1607194113
transform 1 0 89318 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_953
timestamp 1607194113
transform 1 0 88214 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_977
timestamp 1607194113
transform 1 0 90422 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_973
timestamp 1607194113
transform 1 0 90054 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1607194113
transform 1 0 90330 0 1 40848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1001
timestamp 1607194113
transform 1 0 92630 0 1 40848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_989
timestamp 1607194113
transform 1 0 91526 0 1 40848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1607194113
transform -1 0 93642 0 1 40848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_881
timestamp 1607194113
transform 1 0 81590 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_869
timestamp 1607194113
transform 1 0 80486 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_900
timestamp 1607194113
transform 1 0 83338 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_893
timestamp 1607194113
transform 1 0 82694 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1607194113
transform 1 0 83246 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_924
timestamp 1607194113
transform 1 0 85546 0 -1 41936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_912
timestamp 1607194113
transform 1 0 84442 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_943
timestamp 1607194113
transform 1 0 87294 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_931
timestamp 1607194113
transform 1 0 86190 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1607194113
transform 1 0 86098 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_955
timestamp 1607194113
transform 1 0 88398 0 -1 41936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__CLK
timestamp 1607194113
transform 1 0 88766 0 -1 41936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1607194113
transform 1 0 88950 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1515_
timestamp 1607194113
transform 1 0 89042 0 -1 41936
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_76_981
timestamp 1607194113
transform 1 0 90790 0 -1 41936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_1005
timestamp 1607194113
transform 1 0 92998 0 -1 41936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_993
timestamp 1607194113
transform 1 0 91894 0 -1 41936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_989
timestamp 1607194113
transform 1 0 91526 0 -1 41936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1607194113
transform 1 0 91802 0 -1 41936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1607194113
transform -1 0 93642 0 -1 41936
box -38 -48 314 592
<< labels >>
rlabel metal2 s 1200 43312 1256 44112 6 bus_in[0]
port 0 nsew default input
rlabel metal2 s 25580 43312 25636 44112 6 bus_in[10]
port 1 nsew default input
rlabel metal2 s 28064 43312 28120 44112 6 bus_in[11]
port 2 nsew default input
rlabel metal2 s 30548 43312 30604 44112 6 bus_in[12]
port 3 nsew default input
rlabel metal2 s 32940 43312 32996 44112 6 bus_in[13]
port 4 nsew default input
rlabel metal2 s 35424 43312 35480 44112 6 bus_in[14]
port 5 nsew default input
rlabel metal2 s 37816 43312 37872 44112 6 bus_in[15]
port 6 nsew default input
rlabel metal2 s 40300 43312 40356 44112 6 bus_in[16]
port 7 nsew default input
rlabel metal2 s 42692 43312 42748 44112 6 bus_in[17]
port 8 nsew default input
rlabel metal2 s 45176 43312 45232 44112 6 bus_in[18]
port 9 nsew default input
rlabel metal2 s 47660 43312 47716 44112 6 bus_in[19]
port 10 nsew default input
rlabel metal2 s 3592 43312 3648 44112 6 bus_in[1]
port 11 nsew default input
rlabel metal2 s 50052 43312 50108 44112 6 bus_in[20]
port 12 nsew default input
rlabel metal2 s 52536 43312 52592 44112 6 bus_in[21]
port 13 nsew default input
rlabel metal2 s 54928 43312 54984 44112 6 bus_in[22]
port 14 nsew default input
rlabel metal2 s 57412 43312 57468 44112 6 bus_in[23]
port 15 nsew default input
rlabel metal2 s 59804 43312 59860 44112 6 bus_in[24]
port 16 nsew default input
rlabel metal2 s 62288 43312 62344 44112 6 bus_in[25]
port 17 nsew default input
rlabel metal2 s 64680 43312 64736 44112 6 bus_in[26]
port 18 nsew default input
rlabel metal2 s 67164 43312 67220 44112 6 bus_in[27]
port 19 nsew default input
rlabel metal2 s 69648 43312 69704 44112 6 bus_in[28]
port 20 nsew default input
rlabel metal2 s 72040 43312 72096 44112 6 bus_in[29]
port 21 nsew default input
rlabel metal2 s 6076 43312 6132 44112 6 bus_in[2]
port 22 nsew default input
rlabel metal2 s 74524 43312 74580 44112 6 bus_in[30]
port 23 nsew default input
rlabel metal2 s 76916 43312 76972 44112 6 bus_in[31]
port 24 nsew default input
rlabel metal2 s 79400 43312 79456 44112 6 bus_in[32]
port 25 nsew default input
rlabel metal2 s 81792 43312 81848 44112 6 bus_in[33]
port 26 nsew default input
rlabel metal2 s 84276 43312 84332 44112 6 bus_in[34]
port 27 nsew default input
rlabel metal2 s 86760 43312 86816 44112 6 bus_in[35]
port 28 nsew default input
rlabel metal2 s 87956 43312 88012 44112 6 bus_in[36]
port 29 nsew default input
rlabel metal2 s 89152 43312 89208 44112 6 bus_in[37]
port 30 nsew default input
rlabel metal2 s 90348 43312 90404 44112 6 bus_in[38]
port 31 nsew default input
rlabel metal2 s 91636 43312 91692 44112 6 bus_in[39]
port 32 nsew default input
rlabel metal2 s 8468 43312 8524 44112 6 bus_in[3]
port 33 nsew default input
rlabel metal2 s 92832 43312 92888 44112 6 bus_in[40]
port 34 nsew default input
rlabel metal2 s 94028 43312 94084 44112 6 bus_in[41]
port 35 nsew default input
rlabel metal2 s 10952 43312 11008 44112 6 bus_in[4]
port 36 nsew default input
rlabel metal2 s 13436 43312 13492 44112 6 bus_in[5]
port 37 nsew default input
rlabel metal2 s 15828 43312 15884 44112 6 bus_in[6]
port 38 nsew default input
rlabel metal2 s 18312 43312 18368 44112 6 bus_in[7]
port 39 nsew default input
rlabel metal2 s 20704 43312 20760 44112 6 bus_in[8]
port 40 nsew default input
rlabel metal2 s 23188 43312 23244 44112 6 bus_in[9]
port 41 nsew default input
rlabel metal2 s 2396 43312 2452 44112 6 bus_out[0]
port 42 nsew default tristate
rlabel metal2 s 26868 43312 26924 44112 6 bus_out[10]
port 43 nsew default tristate
rlabel metal2 s 29260 43312 29316 44112 6 bus_out[11]
port 44 nsew default tristate
rlabel metal2 s 31744 43312 31800 44112 6 bus_out[12]
port 45 nsew default tristate
rlabel metal2 s 34136 43312 34192 44112 6 bus_out[13]
port 46 nsew default tristate
rlabel metal2 s 36620 43312 36676 44112 6 bus_out[14]
port 47 nsew default tristate
rlabel metal2 s 39104 43312 39160 44112 6 bus_out[15]
port 48 nsew default tristate
rlabel metal2 s 41496 43312 41552 44112 6 bus_out[16]
port 49 nsew default tristate
rlabel metal2 s 43980 43312 44036 44112 6 bus_out[17]
port 50 nsew default tristate
rlabel metal2 s 46372 43312 46428 44112 6 bus_out[18]
port 51 nsew default tristate
rlabel metal2 s 48856 43312 48912 44112 6 bus_out[19]
port 52 nsew default tristate
rlabel metal2 s 4880 43312 4936 44112 6 bus_out[1]
port 53 nsew default tristate
rlabel metal2 s 51248 43312 51304 44112 6 bus_out[20]
port 54 nsew default tristate
rlabel metal2 s 53732 43312 53788 44112 6 bus_out[21]
port 55 nsew default tristate
rlabel metal2 s 56124 43312 56180 44112 6 bus_out[22]
port 56 nsew default tristate
rlabel metal2 s 58608 43312 58664 44112 6 bus_out[23]
port 57 nsew default tristate
rlabel metal2 s 61092 43312 61148 44112 6 bus_out[24]
port 58 nsew default tristate
rlabel metal2 s 63484 43312 63540 44112 6 bus_out[25]
port 59 nsew default tristate
rlabel metal2 s 65968 43312 66024 44112 6 bus_out[26]
port 60 nsew default tristate
rlabel metal2 s 68360 43312 68416 44112 6 bus_out[27]
port 61 nsew default tristate
rlabel metal2 s 70844 43312 70900 44112 6 bus_out[28]
port 62 nsew default tristate
rlabel metal2 s 73236 43312 73292 44112 6 bus_out[29]
port 63 nsew default tristate
rlabel metal2 s 7272 43312 7328 44112 6 bus_out[2]
port 64 nsew default tristate
rlabel metal2 s 75720 43312 75776 44112 6 bus_out[30]
port 65 nsew default tristate
rlabel metal2 s 78204 43312 78260 44112 6 bus_out[31]
port 66 nsew default tristate
rlabel metal2 s 80596 43312 80652 44112 6 bus_out[32]
port 67 nsew default tristate
rlabel metal2 s 83080 43312 83136 44112 6 bus_out[33]
port 68 nsew default tristate
rlabel metal2 s 85472 43312 85528 44112 6 bus_out[34]
port 69 nsew default tristate
rlabel metal2 s 9756 43312 9812 44112 6 bus_out[3]
port 70 nsew default tristate
rlabel metal2 s 12148 43312 12204 44112 6 bus_out[4]
port 71 nsew default tristate
rlabel metal2 s 14632 43312 14688 44112 6 bus_out[5]
port 72 nsew default tristate
rlabel metal2 s 17024 43312 17080 44112 6 bus_out[6]
port 73 nsew default tristate
rlabel metal2 s 19508 43312 19564 44112 6 bus_out[7]
port 74 nsew default tristate
rlabel metal2 s 21992 43312 22048 44112 6 bus_out[8]
port 75 nsew default tristate
rlabel metal2 s 24384 43312 24440 44112 6 bus_out[9]
port 76 nsew default tristate
rlabel metal3 s 93946 9440 94746 9560 6 clk_i
port 77 nsew default input
rlabel metal3 s 93946 32560 94746 32680 6 out_o
port 78 nsew default tristate
rlabel metal2 s 4 43312 60 44112 6 rst_n_i
port 79 nsew default input
rlabel metal5 s 538 3748 93642 4348 6 VPWR
port 80 nsew default input
rlabel metal5 s 538 21748 93642 22348 6 VGND
port 81 nsew default input
<< properties >>
string FIXED_BBOX 0 0 94746 44112
<< end >>
