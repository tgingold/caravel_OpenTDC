magic
tech sky130A
magscale 1 2
timestamp 1607276814
<< locali >>
rect 19165 21471 19199 21641
rect 46489 21471 46523 21641
rect 4445 19703 4479 20009
rect 15025 17051 15059 17289
rect 41245 17119 41279 17289
rect 48973 14399 49007 14569
rect 26341 5559 26375 5729
<< viali >>
rect 38853 24837 38887 24871
rect 8585 24769 8619 24803
rect 22845 24769 22879 24803
rect 42625 24769 42659 24803
rect 49985 24769 50019 24803
rect 6929 24701 6963 24735
rect 7205 24701 7239 24735
rect 21465 24701 21499 24735
rect 21741 24701 21775 24735
rect 38669 24701 38703 24735
rect 39773 24701 39807 24735
rect 41245 24701 41279 24735
rect 41521 24701 41555 24735
rect 44005 24701 44039 24735
rect 44281 24701 44315 24735
rect 49709 24701 49743 24735
rect 8677 24565 8711 24599
rect 21373 24565 21407 24599
rect 38485 24565 38519 24599
rect 39957 24565 39991 24599
rect 42993 24565 43027 24599
rect 43729 24565 43763 24599
rect 45569 24565 45603 24599
rect 49433 24565 49467 24599
rect 51089 24565 51123 24599
rect 2789 24361 2823 24395
rect 7941 24361 7975 24395
rect 13829 24361 13863 24395
rect 16681 24361 16715 24395
rect 19349 24361 19383 24395
rect 22293 24361 22327 24395
rect 24961 24361 24995 24395
rect 27905 24361 27939 24395
rect 30389 24361 30423 24395
rect 33701 24361 33735 24395
rect 36185 24361 36219 24395
rect 39865 24361 39899 24395
rect 52561 24361 52595 24395
rect 5733 24293 5767 24327
rect 11621 24293 11655 24327
rect 50629 24293 50663 24327
rect 1685 24225 1719 24259
rect 5917 24225 5951 24259
rect 6561 24225 6595 24259
rect 8401 24225 8435 24259
rect 9965 24225 9999 24259
rect 11805 24225 11839 24259
rect 12449 24225 12483 24259
rect 14197 24225 14231 24259
rect 15025 24225 15059 24259
rect 15301 24225 15335 24259
rect 15577 24225 15611 24259
rect 20729 24225 20763 24259
rect 20913 24225 20947 24259
rect 23213 24225 23247 24259
rect 23397 24225 23431 24259
rect 26249 24225 26283 24259
rect 26525 24225 26559 24259
rect 26801 24225 26835 24259
rect 34069 24225 34103 24259
rect 34805 24225 34839 24259
rect 36553 24225 36587 24259
rect 38485 24225 38519 24259
rect 40233 24225 40267 24259
rect 50997 24225 51031 24259
rect 51273 24225 51307 24259
rect 1409 24157 1443 24191
rect 4077 24157 4111 24191
rect 4353 24157 4387 24191
rect 6837 24157 6871 24191
rect 10241 24157 10275 24191
rect 12725 24157 12759 24191
rect 17693 24157 17727 24191
rect 17785 24157 17819 24191
rect 18061 24157 18095 24191
rect 21189 24157 21223 24191
rect 23673 24157 23707 24191
rect 29009 24157 29043 24191
rect 29285 24157 29319 24191
rect 32321 24157 32355 24191
rect 32597 24157 32631 24191
rect 35081 24157 35115 24191
rect 38761 24157 38795 24191
rect 45937 24157 45971 24191
rect 46213 24157 46247 24191
rect 50905 24157 50939 24191
rect 3249 24021 3283 24055
rect 30757 24021 30791 24055
rect 45753 24021 45787 24055
rect 47317 24021 47351 24055
rect 10057 23817 10091 23851
rect 15025 23817 15059 23851
rect 15393 23817 15427 23851
rect 19441 23817 19475 23851
rect 22477 23817 22511 23851
rect 25237 23817 25271 23851
rect 26801 23817 26835 23851
rect 31953 23817 31987 23851
rect 33701 23817 33735 23851
rect 35909 23817 35943 23851
rect 37473 23817 37507 23851
rect 39313 23817 39347 23851
rect 41981 23817 42015 23851
rect 44281 23817 44315 23851
rect 46581 23817 46615 23851
rect 49525 23817 49559 23851
rect 47777 23749 47811 23783
rect 7389 23681 7423 23715
rect 8493 23681 8527 23715
rect 10241 23681 10275 23715
rect 13645 23681 13679 23715
rect 13921 23681 13955 23715
rect 25421 23681 25455 23715
rect 30573 23681 30607 23715
rect 30849 23681 30883 23715
rect 36093 23681 36127 23715
rect 38853 23681 38887 23715
rect 41521 23681 41555 23715
rect 43821 23681 43855 23715
rect 48145 23681 48179 23715
rect 5457 23613 5491 23647
rect 5733 23613 5767 23647
rect 6929 23613 6963 23647
rect 7297 23613 7331 23647
rect 8769 23613 8803 23647
rect 12541 23613 12575 23647
rect 12633 23613 12667 23647
rect 17877 23613 17911 23647
rect 18061 23613 18095 23647
rect 18337 23613 18371 23647
rect 21925 23613 21959 23647
rect 22017 23613 22051 23647
rect 22293 23613 22327 23647
rect 25697 23613 25731 23647
rect 32321 23613 32355 23647
rect 33333 23613 33367 23647
rect 33517 23613 33551 23647
rect 34989 23613 35023 23647
rect 36369 23613 36403 23647
rect 39129 23613 39163 23647
rect 40509 23613 40543 23647
rect 41797 23613 41831 23647
rect 44097 23613 44131 23647
rect 46213 23613 46247 23647
rect 46397 23613 46431 23647
rect 48421 23613 48455 23647
rect 52101 23613 52135 23647
rect 52377 23613 52411 23647
rect 22201 23545 22235 23579
rect 33425 23545 33459 23579
rect 39037 23545 39071 23579
rect 41705 23545 41739 23579
rect 44005 23545 44039 23579
rect 46305 23545 46339 23579
rect 5457 23477 5491 23511
rect 12725 23477 12759 23511
rect 22937 23477 22971 23511
rect 35173 23477 35207 23511
rect 40601 23477 40635 23511
rect 47961 23477 47995 23511
rect 51917 23477 51951 23511
rect 53481 23477 53515 23511
rect 13277 23273 13311 23307
rect 21925 23273 21959 23307
rect 37013 23273 37047 23307
rect 5917 23205 5951 23239
rect 8769 23205 8803 23239
rect 11713 23205 11747 23239
rect 18337 23205 18371 23239
rect 21741 23205 21775 23239
rect 23857 23205 23891 23239
rect 30665 23205 30699 23239
rect 36277 23205 36311 23239
rect 44557 23205 44591 23239
rect 46305 23205 46339 23239
rect 48053 23205 48087 23239
rect 52377 23205 52411 23239
rect 8033 23137 8067 23171
rect 8585 23137 8619 23171
rect 11069 23137 11103 23171
rect 11437 23137 11471 23171
rect 13369 23137 13403 23171
rect 15301 23137 15335 23171
rect 15853 23137 15887 23171
rect 18521 23137 18555 23171
rect 18705 23137 18739 23171
rect 18797 23137 18831 23171
rect 21189 23137 21223 23171
rect 21281 23137 21315 23171
rect 23305 23137 23339 23171
rect 23397 23137 23431 23171
rect 24593 23137 24627 23171
rect 24685 23137 24719 23171
rect 26525 23137 26559 23171
rect 27721 23137 27755 23171
rect 27997 23137 28031 23171
rect 30757 23137 30791 23171
rect 32137 23137 32171 23171
rect 33977 23137 34011 23171
rect 34069 23137 34103 23171
rect 36093 23137 36127 23171
rect 36369 23137 36403 23171
rect 41061 23137 41095 23171
rect 41245 23137 41279 23171
rect 41797 23137 41831 23171
rect 41981 23137 42015 23171
rect 47501 23137 47535 23171
rect 47593 23137 47627 23171
rect 51273 23137 51307 23171
rect 51825 23137 51859 23171
rect 51917 23137 51951 23171
rect 4077 23069 4111 23103
rect 4353 23069 4387 23103
rect 5549 23069 5583 23103
rect 16129 23069 16163 23103
rect 29101 23069 29135 23103
rect 30481 23069 30515 23103
rect 38577 23069 38611 23103
rect 38853 23069 38887 23103
rect 44649 23069 44683 23103
rect 44925 23069 44959 23103
rect 47317 23069 47351 23103
rect 13553 23001 13587 23035
rect 15393 23001 15427 23035
rect 22937 23001 22971 23035
rect 23121 23001 23155 23035
rect 33793 23001 33827 23035
rect 34713 23001 34747 23035
rect 15025 22933 15059 22967
rect 18981 22933 19015 22967
rect 21005 22933 21039 22967
rect 22017 22933 22051 22967
rect 24869 22933 24903 22967
rect 26709 22933 26743 22967
rect 29469 22933 29503 22967
rect 30941 22933 30975 22967
rect 32321 22933 32355 22967
rect 34253 22933 34287 22967
rect 36553 22933 36587 22967
rect 38393 22933 38427 22967
rect 40141 22933 40175 22967
rect 42257 22933 42291 22967
rect 47133 22933 47167 22967
rect 48145 22933 48179 22967
rect 51457 22933 51491 22967
rect 51641 22933 51675 22967
rect 18981 22729 19015 22763
rect 19165 22729 19199 22763
rect 20085 22729 20119 22763
rect 31861 22729 31895 22763
rect 33241 22729 33275 22763
rect 33701 22729 33735 22763
rect 34897 22729 34931 22763
rect 35357 22729 35391 22763
rect 36645 22729 36679 22763
rect 38761 22729 38795 22763
rect 6929 22661 6963 22695
rect 15025 22661 15059 22695
rect 16681 22661 16715 22695
rect 20729 22661 20763 22695
rect 21649 22661 21683 22695
rect 25789 22661 25823 22695
rect 31401 22661 31435 22695
rect 40693 22661 40727 22695
rect 3157 22593 3191 22627
rect 3341 22593 3375 22627
rect 4537 22593 4571 22627
rect 4905 22593 4939 22627
rect 10241 22593 10275 22627
rect 15393 22593 15427 22627
rect 19901 22593 19935 22627
rect 21465 22593 21499 22627
rect 26985 22593 27019 22627
rect 37565 22593 37599 22627
rect 48881 22593 48915 22627
rect 53481 22593 53515 22627
rect 1501 22525 1535 22559
rect 1777 22525 1811 22559
rect 4261 22525 4295 22559
rect 4445 22525 4479 22559
rect 7205 22525 7239 22559
rect 9689 22525 9723 22559
rect 9965 22525 9999 22559
rect 11069 22525 11103 22559
rect 12909 22525 12943 22559
rect 15117 22525 15151 22559
rect 19349 22525 19383 22559
rect 19441 22525 19475 22559
rect 21005 22525 21039 22559
rect 24041 22525 24075 22559
rect 24225 22525 24259 22559
rect 24317 22525 24351 22559
rect 25605 22525 25639 22559
rect 27077 22525 27111 22559
rect 27629 22525 27663 22559
rect 27813 22525 27847 22559
rect 29285 22525 29319 22559
rect 31677 22525 31711 22559
rect 33517 22525 33551 22559
rect 35173 22525 35207 22559
rect 36461 22525 36495 22559
rect 37749 22525 37783 22559
rect 38301 22525 38335 22559
rect 38485 22525 38519 22559
rect 40509 22525 40543 22559
rect 42441 22525 42475 22559
rect 42533 22525 42567 22559
rect 42901 22525 42935 22559
rect 42993 22525 43027 22559
rect 46121 22525 46155 22559
rect 48513 22525 48547 22559
rect 48605 22525 48639 22559
rect 52101 22525 52135 22559
rect 52377 22525 52411 22559
rect 7113 22457 7147 22491
rect 7665 22457 7699 22491
rect 20913 22457 20947 22491
rect 24777 22457 24811 22491
rect 28181 22457 28215 22491
rect 31585 22457 31619 22491
rect 33425 22457 33459 22491
rect 35081 22457 35115 22491
rect 35817 22457 35851 22491
rect 42073 22457 42107 22491
rect 43545 22457 43579 22491
rect 51917 22457 51951 22491
rect 11161 22389 11195 22423
rect 13093 22389 13127 22423
rect 23857 22389 23891 22423
rect 28365 22389 28399 22423
rect 29377 22389 29411 22423
rect 46213 22389 46247 22423
rect 49985 22389 50019 22423
rect 2053 22185 2087 22219
rect 4169 22185 4203 22219
rect 4905 22185 4939 22219
rect 21925 22185 21959 22219
rect 42349 22185 42383 22219
rect 51917 22185 51951 22219
rect 2881 22117 2915 22151
rect 21741 22117 21775 22151
rect 23489 22117 23523 22151
rect 44649 22117 44683 22151
rect 51733 22117 51767 22151
rect 2237 22049 2271 22083
rect 2513 22049 2547 22083
rect 4353 22049 4387 22083
rect 4629 22049 4663 22083
rect 5917 22049 5951 22083
rect 6929 22049 6963 22083
rect 7205 22049 7239 22083
rect 7665 22049 7699 22083
rect 8585 22049 8619 22083
rect 9873 22049 9907 22083
rect 10425 22049 10459 22083
rect 10609 22049 10643 22083
rect 10793 22049 10827 22083
rect 10977 22049 11011 22083
rect 11161 22049 11195 22083
rect 12541 22049 12575 22083
rect 13645 22049 13679 22083
rect 18889 22049 18923 22083
rect 21097 22049 21131 22083
rect 21230 22049 21264 22083
rect 22569 22049 22603 22083
rect 23765 22049 23799 22083
rect 24317 22049 24351 22083
rect 26985 22049 27019 22083
rect 28641 22049 28675 22083
rect 33977 22049 34011 22083
rect 34161 22049 34195 22083
rect 34713 22049 34747 22083
rect 34897 22049 34931 22083
rect 42257 22049 42291 22083
rect 43545 22049 43579 22083
rect 44097 22049 44131 22083
rect 44281 22049 44315 22083
rect 44833 22049 44867 22083
rect 46581 22049 46615 22083
rect 49893 22049 49927 22083
rect 50077 22049 50111 22083
rect 50629 22049 50663 22083
rect 50813 22049 50847 22083
rect 52101 22049 52135 22083
rect 52285 22049 52319 22083
rect 52377 22049 52411 22083
rect 17141 21981 17175 22015
rect 17417 21981 17451 22015
rect 18797 21981 18831 22015
rect 24409 21981 24443 22015
rect 24869 21981 24903 22015
rect 28365 21981 28399 22015
rect 30113 21981 30147 22015
rect 39589 21981 39623 22015
rect 39865 21981 39899 22015
rect 43361 21981 43395 22015
rect 46305 21981 46339 22015
rect 47685 21981 47719 22015
rect 6009 21913 6043 21947
rect 7021 21913 7055 21947
rect 12725 21913 12759 21947
rect 20913 21913 20947 21947
rect 23213 21913 23247 21947
rect 23673 21913 23707 21947
rect 52929 21913 52963 21947
rect 8677 21845 8711 21879
rect 11529 21845 11563 21879
rect 13737 21845 13771 21879
rect 21373 21845 21407 21879
rect 22661 21845 22695 21879
rect 26801 21845 26835 21879
rect 27169 21845 27203 21879
rect 29745 21845 29779 21879
rect 35173 21845 35207 21879
rect 39405 21845 39439 21879
rect 41153 21845 41187 21879
rect 42625 21845 42659 21879
rect 45937 21845 45971 21879
rect 46121 21845 46155 21879
rect 51089 21845 51123 21879
rect 52561 21845 52595 21879
rect 5825 21641 5859 21675
rect 9689 21641 9723 21675
rect 12725 21641 12759 21675
rect 14841 21641 14875 21675
rect 17693 21641 17727 21675
rect 19165 21641 19199 21675
rect 19257 21641 19291 21675
rect 21005 21641 21039 21675
rect 22385 21641 22419 21675
rect 46489 21641 46523 21675
rect 46581 21641 46615 21675
rect 51457 21641 51491 21675
rect 7113 21573 7147 21607
rect 11161 21573 11195 21607
rect 13185 21573 13219 21607
rect 15301 21573 15335 21607
rect 2145 21505 2179 21539
rect 3893 21505 3927 21539
rect 7757 21505 7791 21539
rect 9413 21505 9447 21539
rect 27721 21573 27755 21607
rect 32781 21573 32815 21607
rect 33885 21573 33919 21607
rect 23765 21505 23799 21539
rect 24133 21505 24167 21539
rect 26709 21505 26743 21539
rect 38301 21505 38335 21539
rect 39497 21505 39531 21539
rect 43545 21505 43579 21539
rect 51733 21505 51767 21539
rect 52009 21505 52043 21539
rect 53113 21505 53147 21539
rect 2421 21437 2455 21471
rect 5733 21437 5767 21471
rect 7021 21437 7055 21471
rect 7297 21437 7331 21471
rect 9505 21437 9539 21471
rect 10057 21437 10091 21471
rect 11069 21437 11103 21471
rect 12449 21437 12483 21471
rect 12561 21437 12595 21471
rect 13829 21437 13863 21471
rect 15025 21437 15059 21471
rect 15577 21437 15611 21471
rect 16037 21437 16071 21471
rect 17877 21437 17911 21471
rect 19165 21437 19199 21471
rect 19441 21437 19475 21471
rect 19717 21437 19751 21471
rect 22569 21437 22603 21471
rect 23673 21437 23707 21471
rect 23949 21437 23983 21471
rect 25237 21437 25271 21471
rect 26801 21437 26835 21471
rect 27353 21437 27387 21471
rect 27537 21437 27571 21471
rect 29745 21437 29779 21471
rect 31033 21437 31067 21471
rect 31309 21437 31343 21471
rect 33793 21437 33827 21471
rect 35357 21437 35391 21471
rect 35633 21437 35667 21471
rect 37105 21437 37139 21471
rect 38393 21437 38427 21471
rect 38853 21437 38887 21471
rect 38945 21437 38979 21471
rect 40785 21437 40819 21471
rect 40877 21437 40911 21471
rect 43269 21437 43303 21471
rect 46489 21437 46523 21471
rect 46765 21437 46799 21471
rect 47041 21437 47075 21471
rect 13921 21369 13955 21403
rect 22661 21369 22695 21403
rect 37013 21369 37047 21403
rect 3709 21301 3743 21335
rect 23489 21301 23523 21335
rect 25421 21301 25455 21335
rect 29837 21301 29871 21335
rect 32413 21301 32447 21335
rect 41061 21301 41095 21335
rect 43085 21301 43119 21335
rect 44649 21301 44683 21335
rect 48329 21301 48363 21335
rect 5641 21097 5675 21131
rect 8125 21097 8159 21131
rect 13737 21097 13771 21131
rect 14197 21097 14231 21131
rect 14841 21097 14875 21131
rect 16129 21097 16163 21131
rect 17049 21097 17083 21131
rect 19809 21097 19843 21131
rect 20177 21097 20211 21131
rect 21005 21097 21039 21131
rect 36001 21097 36035 21131
rect 40233 21097 40267 21131
rect 41889 21097 41923 21131
rect 51825 21097 51859 21131
rect 7205 21029 7239 21063
rect 10241 21029 10275 21063
rect 22293 21029 22327 21063
rect 24133 21029 24167 21063
rect 24777 21029 24811 21063
rect 28825 21029 28859 21063
rect 31125 21029 31159 21063
rect 47041 21029 47075 21063
rect 4629 20961 4663 20995
rect 5181 20961 5215 20995
rect 5365 20961 5399 20995
rect 7352 20961 7386 20995
rect 9781 20961 9815 20995
rect 11069 20961 11103 20995
rect 12357 20961 12391 20995
rect 15025 20961 15059 20995
rect 15853 20961 15887 20995
rect 16037 20961 16071 20995
rect 17325 20961 17359 20995
rect 17877 20961 17911 20995
rect 18797 20961 18831 20995
rect 18889 20961 18923 20995
rect 19349 20961 19383 20995
rect 19533 20961 19567 20995
rect 20913 20961 20947 20995
rect 22477 20961 22511 20995
rect 22753 20961 22787 20995
rect 24961 20961 24995 20995
rect 29837 20961 29871 20995
rect 30021 20961 30055 20995
rect 30573 20961 30607 20995
rect 30757 20961 30791 20995
rect 33241 20961 33275 20995
rect 33425 20961 33459 20995
rect 33885 20961 33919 20995
rect 33977 20961 34011 20995
rect 36177 20961 36211 20995
rect 36277 20961 36311 20995
rect 41521 20961 41555 20995
rect 41705 20961 41739 20995
rect 44649 20961 44683 20995
rect 45937 20961 45971 20995
rect 46029 20961 46063 20995
rect 46489 20961 46523 20995
rect 46673 20961 46707 20995
rect 49525 20961 49559 20995
rect 49709 20961 49743 20995
rect 50169 20961 50203 20995
rect 50261 20961 50295 20995
rect 52009 20961 52043 20995
rect 4537 20893 4571 20927
rect 7573 20893 7607 20927
rect 9689 20893 9723 20927
rect 12633 20893 12667 20927
rect 17233 20893 17267 20927
rect 27077 20893 27111 20927
rect 27353 20893 27387 20927
rect 34805 20893 34839 20927
rect 36645 20893 36679 20927
rect 38669 20893 38703 20927
rect 38945 20893 38979 20927
rect 52285 20893 52319 20927
rect 7481 20825 7515 20859
rect 16589 20825 16623 20859
rect 25053 20825 25087 20859
rect 44833 20825 44867 20859
rect 50721 20825 50755 20859
rect 7849 20757 7883 20791
rect 11253 20757 11287 20791
rect 17509 20757 17543 20791
rect 28641 20757 28675 20791
rect 34437 20757 34471 20791
rect 36461 20757 36495 20791
rect 40417 20757 40451 20791
rect 44465 20757 44499 20791
rect 47225 20757 47259 20791
rect 53389 20757 53423 20791
rect 5825 20553 5859 20587
rect 11345 20553 11379 20587
rect 15117 20553 15151 20587
rect 16037 20553 16071 20587
rect 17141 20553 17175 20587
rect 24961 20553 24995 20587
rect 49709 20553 49743 20587
rect 11713 20485 11747 20519
rect 24298 20485 24332 20519
rect 26801 20485 26835 20519
rect 30205 20485 30239 20519
rect 39221 20485 39255 20519
rect 41245 20485 41279 20519
rect 42073 20485 42107 20519
rect 50721 20485 50755 20519
rect 7297 20417 7331 20451
rect 10149 20417 10183 20451
rect 19257 20417 19291 20451
rect 24501 20417 24535 20451
rect 25697 20417 25731 20451
rect 31493 20417 31527 20451
rect 35909 20417 35943 20451
rect 38117 20417 38151 20451
rect 43637 20417 43671 20451
rect 46121 20417 46155 20451
rect 51733 20417 51767 20451
rect 3525 20349 3559 20383
rect 3709 20349 3743 20383
rect 4169 20349 4203 20383
rect 4261 20349 4295 20383
rect 5733 20349 5767 20383
rect 7481 20349 7515 20383
rect 7941 20349 7975 20383
rect 8033 20349 8067 20383
rect 10333 20349 10367 20383
rect 10885 20349 10919 20383
rect 11069 20349 11103 20383
rect 13277 20349 13311 20383
rect 13553 20349 13587 20383
rect 15761 20349 15795 20383
rect 15945 20349 15979 20383
rect 17325 20349 17359 20383
rect 18061 20349 18095 20383
rect 19349 20349 19383 20383
rect 19901 20349 19935 20383
rect 20085 20349 20119 20383
rect 20637 20349 20671 20383
rect 21741 20349 21775 20383
rect 24363 20349 24397 20383
rect 25881 20349 25915 20383
rect 26341 20349 26375 20383
rect 26433 20349 26467 20383
rect 30021 20349 30055 20383
rect 31677 20349 31711 20383
rect 32229 20349 32263 20383
rect 32413 20349 32447 20383
rect 35633 20349 35667 20383
rect 38301 20349 38335 20383
rect 38853 20349 38887 20383
rect 39037 20349 39071 20383
rect 41429 20349 41463 20383
rect 42257 20349 42291 20383
rect 42533 20349 42567 20383
rect 46305 20349 46339 20383
rect 46765 20349 46799 20383
rect 46857 20349 46891 20383
rect 48421 20349 48455 20383
rect 49617 20349 49651 20383
rect 50629 20349 50663 20383
rect 51917 20349 51951 20383
rect 52377 20349 52411 20383
rect 52469 20349 52503 20383
rect 4813 20281 4847 20315
rect 16497 20281 16531 20315
rect 21833 20281 21867 20315
rect 24133 20281 24167 20315
rect 24869 20281 24903 20315
rect 32781 20281 32815 20315
rect 37289 20281 37323 20315
rect 49893 20281 49927 20315
rect 8493 20213 8527 20247
rect 11805 20213 11839 20247
rect 11989 20213 12023 20247
rect 14657 20213 14691 20247
rect 18245 20213 18279 20247
rect 20361 20213 20395 20247
rect 29929 20213 29963 20247
rect 37381 20213 37415 20247
rect 47317 20213 47351 20247
rect 48513 20213 48547 20247
rect 52929 20213 52963 20247
rect 3065 20009 3099 20043
rect 4445 20009 4479 20043
rect 7297 20009 7331 20043
rect 8401 20009 8435 20043
rect 9781 20009 9815 20043
rect 16865 20009 16899 20043
rect 22293 20009 22327 20043
rect 23397 20009 23431 20043
rect 31033 20009 31067 20043
rect 34529 20009 34563 20043
rect 38485 20009 38519 20043
rect 45845 20009 45879 20043
rect 53389 20009 53423 20043
rect 1501 19873 1535 19907
rect 3341 19873 3375 19907
rect 1771 19805 1805 19839
rect 4629 19941 4663 19975
rect 13277 19941 13311 19975
rect 26893 19941 26927 19975
rect 29561 19941 29595 19975
rect 50629 19941 50663 19975
rect 51825 19941 51859 19975
rect 4537 19873 4571 19907
rect 6285 19873 6319 19907
rect 6837 19873 6871 19907
rect 7021 19873 7055 19907
rect 8309 19873 8343 19907
rect 10149 19873 10183 19907
rect 10333 19873 10367 19907
rect 10701 19873 10735 19907
rect 10885 19873 10919 19907
rect 12173 19873 12207 19907
rect 12725 19873 12759 19907
rect 12909 19873 12943 19907
rect 14197 19873 14231 19907
rect 15577 19873 15611 19907
rect 16681 19873 16715 19907
rect 18061 19873 18095 19907
rect 18153 19873 18187 19907
rect 18613 19873 18647 19907
rect 18797 19873 18831 19907
rect 19349 19873 19383 19907
rect 21189 19873 21223 19907
rect 23489 19873 23523 19907
rect 25145 19873 25179 19907
rect 26525 19873 26559 19907
rect 28089 19873 28123 19907
rect 30941 19873 30975 19907
rect 32965 19873 32999 19907
rect 33241 19873 33275 19907
rect 38669 19873 38703 19907
rect 39221 19873 39255 19907
rect 39313 19873 39347 19907
rect 39681 19873 39715 19907
rect 39773 19873 39807 19907
rect 41245 19873 41279 19907
rect 46305 19873 46339 19907
rect 48789 19873 48823 19907
rect 48973 19873 49007 19907
rect 49249 19873 49283 19907
rect 52009 19873 52043 19907
rect 6193 19805 6227 19839
rect 11989 19805 12023 19839
rect 13737 19805 13771 19839
rect 13921 19805 13955 19839
rect 19165 19805 19199 19839
rect 20729 19805 20763 19839
rect 20913 19805 20947 19839
rect 25053 19805 25087 19839
rect 26617 19805 26651 19839
rect 27813 19805 27847 19839
rect 29193 19805 29227 19839
rect 34713 19805 34747 19839
rect 46029 19805 46063 19839
rect 52285 19805 52319 19839
rect 11069 19737 11103 19771
rect 13461 19737 13495 19771
rect 14289 19737 14323 19771
rect 25789 19737 25823 19771
rect 40141 19737 40175 19771
rect 40601 19737 40635 19771
rect 4445 19669 4479 19703
rect 15761 19669 15795 19703
rect 23673 19669 23707 19703
rect 25329 19669 25363 19703
rect 41061 19669 41095 19703
rect 41429 19669 41463 19703
rect 47409 19669 47443 19703
rect 3065 19465 3099 19499
rect 10517 19465 10551 19499
rect 16497 19465 16531 19499
rect 18521 19465 18555 19499
rect 30481 19465 30515 19499
rect 42901 19465 42935 19499
rect 17417 19397 17451 19431
rect 8125 19329 8159 19363
rect 3249 19261 3283 19295
rect 4077 19261 4111 19295
rect 5917 19261 5951 19295
rect 6837 19261 6871 19295
rect 8217 19261 8251 19295
rect 8769 19261 8803 19295
rect 8953 19261 8987 19295
rect 10701 19261 10735 19295
rect 10885 19261 10919 19295
rect 11253 19261 11287 19295
rect 11437 19261 11471 19295
rect 15209 19261 15243 19295
rect 16313 19261 16347 19295
rect 17601 19261 17635 19295
rect 18337 19261 18371 19295
rect 19349 19261 19383 19295
rect 19441 19261 19475 19295
rect 19717 19261 19751 19295
rect 21097 19261 21131 19295
rect 23857 19261 23891 19295
rect 23949 19261 23983 19295
rect 24409 19261 24443 19295
rect 24593 19261 24627 19295
rect 26433 19261 26467 19295
rect 26617 19261 26651 19295
rect 27169 19261 27203 19295
rect 27353 19261 27387 19295
rect 30665 19261 30699 19295
rect 30849 19261 30883 19295
rect 31171 19261 31205 19295
rect 31309 19261 31343 19295
rect 32321 19261 32355 19295
rect 36277 19261 36311 19295
rect 36369 19261 36403 19295
rect 36737 19261 36771 19295
rect 36829 19261 36863 19295
rect 38301 19261 38335 19295
rect 38393 19261 38427 19295
rect 39313 19261 39347 19295
rect 41889 19261 41923 19295
rect 41981 19261 42015 19295
rect 42349 19261 42383 19295
rect 42441 19261 42475 19295
rect 45017 19261 45051 19295
rect 46121 19261 46155 19295
rect 46397 19261 46431 19295
rect 47961 19261 47995 19295
rect 48605 19261 48639 19295
rect 48697 19261 48731 19295
rect 48973 19261 49007 19295
rect 49065 19261 49099 19295
rect 49985 19261 50019 19295
rect 52101 19261 52135 19295
rect 53297 19261 53331 19295
rect 27721 19193 27755 19227
rect 37841 19193 37875 19227
rect 45109 19193 45143 19227
rect 51917 19193 51951 19227
rect 52469 19193 52503 19227
rect 4169 19125 4203 19159
rect 5733 19125 5767 19159
rect 7021 19125 7055 19159
rect 9229 19125 9263 19159
rect 15393 19125 15427 19159
rect 17785 19125 17819 19159
rect 18245 19125 18279 19159
rect 24869 19125 24903 19159
rect 32413 19125 32447 19159
rect 37289 19125 37323 19159
rect 37657 19125 37691 19159
rect 39405 19125 39439 19159
rect 39681 19125 39715 19159
rect 43177 19125 43211 19159
rect 46213 19125 46247 19159
rect 50077 19125 50111 19159
rect 53389 19125 53423 19159
rect 2973 18921 3007 18955
rect 9965 18921 9999 18955
rect 17233 18921 17267 18955
rect 17509 18921 17543 18955
rect 25513 18921 25547 18955
rect 29745 18921 29779 18955
rect 33701 18921 33735 18955
rect 36185 18921 36219 18955
rect 41705 18921 41739 18955
rect 4353 18853 4387 18887
rect 29285 18853 29319 18887
rect 39865 18853 39899 18887
rect 41981 18853 42015 18887
rect 49617 18853 49651 18887
rect 3157 18785 3191 18819
rect 4261 18785 4295 18819
rect 6377 18785 6411 18819
rect 6929 18785 6963 18819
rect 7113 18785 7147 18819
rect 10149 18785 10183 18819
rect 10333 18785 10367 18819
rect 10701 18785 10735 18819
rect 10885 18785 10919 18819
rect 12909 18785 12943 18819
rect 13461 18785 13495 18819
rect 13645 18785 13679 18819
rect 15853 18785 15887 18819
rect 17049 18785 17083 18819
rect 21741 18785 21775 18819
rect 24225 18785 24259 18819
rect 26525 18785 26559 18819
rect 28365 18785 28399 18819
rect 29929 18785 29963 18819
rect 30021 18785 30055 18819
rect 32321 18785 32355 18819
rect 32413 18785 32447 18819
rect 32781 18785 32815 18819
rect 32873 18785 32907 18819
rect 36553 18785 36587 18819
rect 38761 18785 38795 18819
rect 39313 18785 39347 18819
rect 39497 18785 39531 18819
rect 41889 18785 41923 18819
rect 44097 18785 44131 18819
rect 44557 18785 44591 18819
rect 44649 18785 44683 18819
rect 47869 18785 47903 18819
rect 48145 18785 48179 18819
rect 49065 18785 49099 18819
rect 49249 18785 49283 18819
rect 50629 18785 50663 18819
rect 50721 18785 50755 18819
rect 50905 18785 50939 18819
rect 51365 18785 51399 18819
rect 51457 18785 51491 18819
rect 52929 18785 52963 18819
rect 53113 18785 53147 18819
rect 6101 18717 6135 18751
rect 6285 18717 6319 18751
rect 12725 18717 12759 18751
rect 23765 18717 23799 18751
rect 23949 18717 23983 18751
rect 28733 18717 28767 18751
rect 31861 18717 31895 18751
rect 33425 18717 33459 18751
rect 38209 18717 38243 18751
rect 38577 18717 38611 18751
rect 44005 18717 44039 18751
rect 15761 18649 15795 18683
rect 26617 18649 26651 18683
rect 28641 18649 28675 18683
rect 38393 18649 38427 18683
rect 45017 18649 45051 18683
rect 51825 18649 51859 18683
rect 7389 18581 7423 18615
rect 13921 18581 13955 18615
rect 16037 18581 16071 18615
rect 21833 18581 21867 18615
rect 28503 18581 28537 18615
rect 29009 18581 29043 18615
rect 33885 18581 33919 18615
rect 36369 18581 36403 18615
rect 47961 18581 47995 18615
rect 53205 18581 53239 18615
rect 10977 18377 11011 18411
rect 32505 18377 32539 18411
rect 33517 18377 33551 18411
rect 36553 18377 36587 18411
rect 39018 18377 39052 18411
rect 39773 18377 39807 18411
rect 44170 18377 44204 18411
rect 48145 18377 48179 18411
rect 52837 18377 52871 18411
rect 4169 18309 4203 18343
rect 12265 18309 12299 18343
rect 19901 18309 19935 18343
rect 21005 18309 21039 18343
rect 28089 18309 28123 18343
rect 29561 18309 29595 18343
rect 32229 18309 32263 18343
rect 32965 18309 32999 18343
rect 33406 18309 33440 18343
rect 39129 18309 39163 18343
rect 43361 18309 43395 18343
rect 48421 18309 48455 18343
rect 49709 18309 49743 18343
rect 1869 18241 1903 18275
rect 8677 18241 8711 18275
rect 12449 18241 12483 18275
rect 13737 18241 13771 18275
rect 15025 18241 15059 18275
rect 18337 18241 18371 18275
rect 21097 18241 21131 18275
rect 21373 18241 21407 18275
rect 25237 18241 25271 18275
rect 25697 18241 25731 18275
rect 29432 18241 29466 18275
rect 29653 18241 29687 18275
rect 29745 18241 29779 18275
rect 33609 18241 33643 18275
rect 33701 18241 33735 18275
rect 39221 18241 39255 18275
rect 41797 18241 41831 18275
rect 43085 18241 43119 18275
rect 44373 18241 44407 18275
rect 44465 18241 44499 18275
rect 46121 18241 46155 18275
rect 49065 18241 49099 18275
rect 1593 18173 1627 18207
rect 3341 18173 3375 18207
rect 4353 18173 4387 18207
rect 4629 18173 4663 18207
rect 5089 18173 5123 18207
rect 5273 18173 5307 18207
rect 6837 18173 6871 18207
rect 8401 18173 8435 18207
rect 10057 18173 10091 18207
rect 10885 18173 10919 18207
rect 12633 18173 12667 18207
rect 13093 18173 13127 18207
rect 13185 18173 13219 18207
rect 14749 18173 14783 18207
rect 18061 18173 18095 18207
rect 25421 18173 25455 18207
rect 25789 18173 25823 18207
rect 31033 18173 31067 18207
rect 31217 18173 31251 18207
rect 31769 18173 31803 18207
rect 31953 18173 31987 18207
rect 34989 18173 35023 18207
rect 35173 18173 35207 18207
rect 35633 18173 35667 18207
rect 35725 18173 35759 18207
rect 36737 18173 36771 18207
rect 40785 18173 40819 18207
rect 41981 18173 42015 18207
rect 42533 18173 42567 18207
rect 42717 18173 42751 18207
rect 44235 18173 44269 18207
rect 46305 18173 46339 18207
rect 46765 18173 46799 18207
rect 46857 18173 46891 18207
rect 48329 18173 48363 18207
rect 48605 18173 48639 18207
rect 50077 18173 50111 18207
rect 52377 18173 52411 18207
rect 52653 18173 52687 18207
rect 3249 18105 3283 18139
rect 10149 18105 10183 18139
rect 16405 18105 16439 18139
rect 19717 18105 19751 18139
rect 22753 18105 22787 18139
rect 26709 18105 26743 18139
rect 26801 18105 26835 18139
rect 29285 18105 29319 18139
rect 33241 18105 33275 18139
rect 36277 18105 36311 18139
rect 38853 18105 38887 18139
rect 44005 18105 44039 18139
rect 45937 18105 45971 18139
rect 49893 18105 49927 18139
rect 50445 18105 50479 18139
rect 52561 18105 52595 18139
rect 7021 18037 7055 18071
rect 14565 18037 14599 18071
rect 25053 18037 25087 18071
rect 32781 18037 32815 18071
rect 39497 18037 39531 18071
rect 40877 18037 40911 18071
rect 47317 18037 47351 18071
rect 2973 17833 3007 17867
rect 4813 17833 4847 17867
rect 11621 17833 11655 17867
rect 14197 17833 14231 17867
rect 19257 17833 19291 17867
rect 21189 17833 21223 17867
rect 23673 17833 23707 17867
rect 38945 17833 38979 17867
rect 53021 17833 53055 17867
rect 16129 17765 16163 17799
rect 24869 17765 24903 17799
rect 25789 17765 25823 17799
rect 29745 17765 29779 17799
rect 29929 17765 29963 17799
rect 36277 17765 36311 17799
rect 40049 17765 40083 17799
rect 45477 17765 45511 17799
rect 49525 17765 49559 17799
rect 3157 17697 3191 17731
rect 4997 17697 5031 17731
rect 6009 17697 6043 17731
rect 6653 17697 6687 17731
rect 7849 17697 7883 17731
rect 10517 17697 10551 17731
rect 11805 17697 11839 17731
rect 11989 17697 12023 17731
rect 12449 17697 12483 17731
rect 12541 17697 12575 17731
rect 14381 17697 14415 17731
rect 16037 17697 16071 17731
rect 17049 17697 17083 17731
rect 18245 17697 18279 17731
rect 19165 17697 19199 17731
rect 21097 17697 21131 17731
rect 22017 17697 22051 17731
rect 22109 17697 22143 17731
rect 22293 17697 22327 17731
rect 22845 17697 22879 17731
rect 23029 17697 23063 17731
rect 28733 17697 28767 17731
rect 29101 17697 29135 17731
rect 29469 17697 29503 17731
rect 32321 17697 32355 17731
rect 32781 17697 32815 17731
rect 32873 17697 32907 17731
rect 34345 17697 34379 17731
rect 36093 17697 36127 17731
rect 36185 17697 36219 17731
rect 37565 17697 37599 17731
rect 37749 17697 37783 17731
rect 37933 17697 37967 17731
rect 38393 17697 38427 17731
rect 38485 17697 38519 17731
rect 39221 17697 39255 17731
rect 40325 17697 40359 17731
rect 40417 17697 40451 17731
rect 40877 17697 40911 17731
rect 41061 17697 41095 17731
rect 41613 17697 41647 17731
rect 47041 17697 47075 17731
rect 47409 17697 47443 17731
rect 47593 17697 47627 17731
rect 48973 17697 49007 17731
rect 49157 17697 49191 17731
rect 50353 17697 50387 17731
rect 51549 17697 51583 17731
rect 51641 17697 51675 17731
rect 52929 17697 52963 17731
rect 25016 17629 25050 17663
rect 25237 17629 25271 17663
rect 31953 17629 31987 17663
rect 32137 17629 32171 17663
rect 34437 17629 34471 17663
rect 43821 17629 43855 17663
rect 44097 17629 44131 17663
rect 47133 17629 47167 17663
rect 51365 17629 51399 17663
rect 52101 17629 52135 17663
rect 5825 17561 5859 17595
rect 25145 17561 25179 17595
rect 25513 17561 25547 17595
rect 35909 17561 35943 17595
rect 37381 17561 37415 17595
rect 41245 17561 41279 17595
rect 50445 17561 50479 17595
rect 6837 17493 6871 17527
rect 8033 17493 8067 17527
rect 10701 17493 10735 17527
rect 13001 17493 13035 17527
rect 14565 17493 14599 17527
rect 17141 17493 17175 17527
rect 18061 17493 18095 17527
rect 23305 17493 23339 17527
rect 33333 17493 33367 17527
rect 43729 17493 43763 17527
rect 46489 17493 46523 17527
rect 2145 17289 2179 17323
rect 4813 17289 4847 17323
rect 15025 17289 15059 17323
rect 24869 17289 24903 17323
rect 28273 17289 28307 17323
rect 28549 17289 28583 17323
rect 30757 17289 30791 17323
rect 31861 17289 31895 17323
rect 41245 17289 41279 17323
rect 41521 17289 41555 17323
rect 44097 17289 44131 17323
rect 45109 17289 45143 17323
rect 46857 17289 46891 17323
rect 14289 17221 14323 17255
rect 7205 17153 7239 17187
rect 9781 17153 9815 17187
rect 13001 17153 13035 17187
rect 2329 17085 2363 17119
rect 3341 17085 3375 17119
rect 3801 17085 3835 17119
rect 3893 17085 3927 17119
rect 4353 17085 4387 17119
rect 4537 17085 4571 17119
rect 7573 17085 7607 17119
rect 7757 17085 7791 17119
rect 8125 17085 8159 17119
rect 8309 17085 8343 17119
rect 10241 17085 10275 17119
rect 10425 17085 10459 17119
rect 10793 17085 10827 17119
rect 10885 17085 10919 17119
rect 12725 17085 12759 17119
rect 21189 17221 21223 17255
rect 24501 17221 24535 17255
rect 27905 17221 27939 17255
rect 36001 17221 36035 17255
rect 39865 17221 39899 17255
rect 18889 17153 18923 17187
rect 20177 17153 20211 17187
rect 24593 17153 24627 17187
rect 27997 17153 28031 17187
rect 29469 17153 29503 17187
rect 30389 17153 30423 17187
rect 34621 17153 34655 17187
rect 34897 17153 34931 17187
rect 37565 17153 37599 17187
rect 37657 17153 37691 17187
rect 41613 17153 41647 17187
rect 46949 17153 46983 17187
rect 50813 17153 50847 17187
rect 50905 17153 50939 17187
rect 52377 17153 52411 17187
rect 53481 17153 53515 17187
rect 15301 17085 15335 17119
rect 15485 17085 15519 17119
rect 16037 17085 16071 17119
rect 16221 17085 16255 17119
rect 19073 17085 19107 17119
rect 19533 17085 19567 17119
rect 19625 17085 19659 17119
rect 21097 17085 21131 17119
rect 24225 17085 24259 17119
rect 24372 17085 24406 17119
rect 27776 17085 27810 17119
rect 29929 17085 29963 17119
rect 30113 17085 30147 17119
rect 30481 17085 30515 17119
rect 31769 17085 31803 17119
rect 35081 17085 35115 17119
rect 35633 17085 35667 17119
rect 35817 17085 35851 17119
rect 36369 17085 36403 17119
rect 37841 17085 37875 17119
rect 38301 17085 38335 17119
rect 38393 17085 38427 17119
rect 39221 17085 39255 17119
rect 40049 17085 40083 17119
rect 41245 17085 41279 17119
rect 41797 17085 41831 17119
rect 42257 17085 42291 17119
rect 42349 17085 42383 17119
rect 44005 17085 44039 17119
rect 45017 17085 45051 17119
rect 47225 17085 47259 17119
rect 50261 17085 50295 17119
rect 50425 17085 50459 17119
rect 52101 17085 52135 17119
rect 15025 17017 15059 17051
rect 27629 17017 27663 17051
rect 38945 17017 38979 17051
rect 42901 17017 42935 17051
rect 3157 16949 3191 16983
rect 14473 16949 14507 16983
rect 15117 16949 15151 16983
rect 16497 16949 16531 16983
rect 29285 16949 29319 16983
rect 48513 16949 48547 16983
rect 51917 16949 51951 16983
rect 2605 16745 2639 16779
rect 4169 16745 4203 16779
rect 10793 16745 10827 16779
rect 13461 16745 13495 16779
rect 17785 16745 17819 16779
rect 25789 16745 25823 16779
rect 28733 16745 28767 16779
rect 30665 16745 30699 16779
rect 33609 16745 33643 16779
rect 42257 16745 42291 16779
rect 47501 16745 47535 16779
rect 21649 16677 21683 16711
rect 21833 16677 21867 16711
rect 39957 16677 39991 16711
rect 40601 16677 40635 16711
rect 53297 16677 53331 16711
rect 2789 16609 2823 16643
rect 3801 16609 3835 16643
rect 4077 16609 4111 16643
rect 5549 16609 5583 16643
rect 5641 16609 5675 16643
rect 5825 16609 5859 16643
rect 6377 16609 6411 16643
rect 6561 16609 6595 16643
rect 8033 16609 8067 16643
rect 11161 16609 11195 16643
rect 11529 16609 11563 16643
rect 11713 16609 11747 16643
rect 13369 16609 13403 16643
rect 14565 16609 14599 16643
rect 16037 16609 16071 16643
rect 16221 16609 16255 16643
rect 16497 16609 16531 16643
rect 18889 16609 18923 16643
rect 19349 16609 19383 16643
rect 22017 16609 22051 16643
rect 22201 16609 22235 16643
rect 22661 16609 22695 16643
rect 22753 16609 22787 16643
rect 24409 16609 24443 16643
rect 24501 16609 24535 16643
rect 24869 16609 24903 16643
rect 24961 16609 24995 16643
rect 26525 16609 26559 16643
rect 26709 16609 26743 16643
rect 27169 16609 27203 16643
rect 27261 16609 27295 16643
rect 29101 16609 29135 16643
rect 29193 16609 29227 16643
rect 29653 16609 29687 16643
rect 29837 16609 29871 16643
rect 30481 16609 30515 16643
rect 32229 16609 32263 16643
rect 34069 16609 34103 16643
rect 35173 16609 35207 16643
rect 40748 16609 40782 16643
rect 41337 16609 41371 16643
rect 42165 16609 42199 16643
rect 43361 16609 43395 16643
rect 47409 16609 47443 16643
rect 48973 16609 49007 16643
rect 50261 16609 50295 16643
rect 50445 16609 50479 16643
rect 51641 16609 51675 16643
rect 51825 16609 51859 16643
rect 51917 16609 51951 16643
rect 53205 16609 53239 16643
rect 11253 16541 11287 16575
rect 32505 16541 32539 16575
rect 35449 16541 35483 16575
rect 38117 16541 38151 16575
rect 38393 16541 38427 16575
rect 39497 16541 39531 16575
rect 40969 16541 41003 16575
rect 50813 16541 50847 16575
rect 52377 16541 52411 16575
rect 18705 16473 18739 16507
rect 25329 16473 25363 16507
rect 27997 16473 28031 16507
rect 30021 16473 30055 16507
rect 36553 16473 36587 16507
rect 53481 16473 53515 16507
rect 3617 16405 3651 16439
rect 6837 16405 6871 16439
rect 7849 16405 7883 16439
rect 14381 16405 14415 16439
rect 19441 16405 19475 16439
rect 23213 16405 23247 16439
rect 25973 16405 26007 16439
rect 27721 16405 27755 16439
rect 36921 16405 36955 16439
rect 40417 16405 40451 16439
rect 40877 16405 40911 16439
rect 43453 16405 43487 16439
rect 49065 16405 49099 16439
rect 4721 16201 4755 16235
rect 8861 16201 8895 16235
rect 14841 16201 14875 16235
rect 25697 16201 25731 16235
rect 26985 16201 27019 16235
rect 27353 16201 27387 16235
rect 29377 16201 29411 16235
rect 32873 16201 32907 16235
rect 35909 16201 35943 16235
rect 39221 16201 39255 16235
rect 47685 16201 47719 16235
rect 53481 16201 53515 16235
rect 32413 16133 32447 16167
rect 2421 16065 2455 16099
rect 21465 16065 21499 16099
rect 24593 16065 24627 16099
rect 27077 16065 27111 16099
rect 31585 16065 31619 16099
rect 43361 16065 43395 16099
rect 48145 16065 48179 16099
rect 52377 16065 52411 16099
rect 2145 15997 2179 16031
rect 3801 15997 3835 16031
rect 4629 15997 4663 16031
rect 5825 15997 5859 16031
rect 7113 15997 7147 16031
rect 9045 15997 9079 16031
rect 9229 15997 9263 16031
rect 9597 15997 9631 16031
rect 9781 15997 9815 16031
rect 10793 15997 10827 16031
rect 13277 15997 13311 16031
rect 13553 15997 13587 16031
rect 15761 15997 15795 16031
rect 15945 15997 15979 16031
rect 16405 15997 16439 16031
rect 16497 15997 16531 16031
rect 18981 15997 19015 16031
rect 19349 15997 19383 16031
rect 19441 15997 19475 16031
rect 19809 15997 19843 16031
rect 19901 15997 19935 16031
rect 21557 15997 21591 16031
rect 22017 15997 22051 16031
rect 22109 15997 22143 16031
rect 24685 15997 24719 16031
rect 25145 15997 25179 16031
rect 25237 15997 25271 16031
rect 26856 15997 26890 16031
rect 29285 15997 29319 16031
rect 31217 15997 31251 16031
rect 32689 15997 32723 16031
rect 35541 15997 35575 16031
rect 35725 15997 35759 16031
rect 39129 15997 39163 16031
rect 42073 15997 42107 16031
rect 43269 15997 43303 16031
rect 43545 15997 43579 16031
rect 48237 15997 48271 16031
rect 48605 15997 48639 16031
rect 48697 15997 48731 16031
rect 49801 15997 49835 16031
rect 52101 15997 52135 16031
rect 3985 15929 4019 15963
rect 17049 15929 17083 15963
rect 20453 15929 20487 15963
rect 26709 15929 26743 15963
rect 31033 15929 31067 15963
rect 32597 15929 32631 15963
rect 35633 15929 35667 15963
rect 41889 15929 41923 15963
rect 44005 15929 44039 15963
rect 49617 15929 49651 15963
rect 50169 15929 50203 15963
rect 5641 15861 5675 15895
rect 7297 15861 7331 15895
rect 9965 15861 9999 15895
rect 10425 15861 10459 15895
rect 10609 15861 10643 15895
rect 15025 15861 15059 15895
rect 15669 15861 15703 15895
rect 18613 15861 18647 15895
rect 18797 15861 18831 15895
rect 22569 15861 22603 15895
rect 42165 15861 42199 15895
rect 51917 15861 51951 15895
rect 2145 15657 2179 15691
rect 3157 15657 3191 15691
rect 7665 15657 7699 15691
rect 11437 15657 11471 15691
rect 18521 15657 18555 15691
rect 21005 15657 21039 15691
rect 29285 15657 29319 15691
rect 33977 15657 34011 15691
rect 44005 15657 44039 15691
rect 45477 15657 45511 15691
rect 13185 15589 13219 15623
rect 19349 15589 19383 15623
rect 32321 15589 32355 15623
rect 38209 15589 38243 15623
rect 41889 15589 41923 15623
rect 51733 15589 51767 15623
rect 2329 15521 2363 15555
rect 3341 15521 3375 15555
rect 4997 15521 5031 15555
rect 5549 15521 5583 15555
rect 6101 15521 6135 15555
rect 6285 15521 6319 15555
rect 8217 15521 8251 15555
rect 8585 15521 8619 15555
rect 8769 15521 8803 15555
rect 10609 15521 10643 15555
rect 11621 15521 11655 15555
rect 12081 15521 12115 15555
rect 12633 15521 12667 15555
rect 12817 15521 12851 15555
rect 14289 15521 14323 15555
rect 15301 15521 15335 15555
rect 16773 15521 16807 15555
rect 17049 15521 17083 15555
rect 19533 15521 19567 15555
rect 20913 15521 20947 15555
rect 24593 15521 24627 15555
rect 30389 15521 30423 15555
rect 32505 15521 32539 15555
rect 33701 15521 33735 15555
rect 33885 15521 33919 15555
rect 35449 15521 35483 15555
rect 35817 15521 35851 15555
rect 36185 15521 36219 15555
rect 39037 15521 39071 15555
rect 39221 15521 39255 15555
rect 40325 15521 40359 15555
rect 40509 15521 40543 15555
rect 40877 15521 40911 15555
rect 41981 15521 42015 15555
rect 42441 15521 42475 15555
rect 44373 15521 44407 15555
rect 46765 15521 46799 15555
rect 46949 15521 46983 15555
rect 48973 15521 49007 15555
rect 49065 15521 49099 15555
rect 49249 15521 49283 15555
rect 51181 15521 51215 15555
rect 51365 15521 51399 15555
rect 51825 15521 51859 15555
rect 5273 15453 5307 15487
rect 5365 15453 5399 15487
rect 8033 15453 8067 15487
rect 11805 15453 11839 15487
rect 11989 15453 12023 15487
rect 18429 15453 18463 15487
rect 21925 15453 21959 15487
rect 22201 15453 22235 15487
rect 27905 15453 27939 15487
rect 28181 15453 28215 15487
rect 32873 15453 32907 15487
rect 38761 15453 38795 15487
rect 44097 15453 44131 15487
rect 49617 15453 49651 15487
rect 4813 15385 4847 15419
rect 6469 15385 6503 15419
rect 14105 15385 14139 15419
rect 10425 15317 10459 15351
rect 13461 15317 13495 15351
rect 15393 15317 15427 15351
rect 19625 15317 19659 15351
rect 21741 15317 21775 15351
rect 23489 15317 23523 15351
rect 24225 15317 24259 15351
rect 24409 15317 24443 15351
rect 29653 15317 29687 15351
rect 30481 15317 30515 15351
rect 41705 15317 41739 15351
rect 47041 15317 47075 15351
rect 11345 15113 11379 15147
rect 14657 15113 14691 15147
rect 22477 15113 22511 15147
rect 33333 15113 33367 15147
rect 36507 15113 36541 15147
rect 36645 15113 36679 15147
rect 47087 15113 47121 15147
rect 47593 15113 47627 15147
rect 50629 15113 50663 15147
rect 51733 15113 51767 15147
rect 2145 15045 2179 15079
rect 24685 15045 24719 15079
rect 38577 15045 38611 15079
rect 47225 15045 47259 15079
rect 3709 14977 3743 15011
rect 8953 14977 8987 15011
rect 9137 14977 9171 15011
rect 12265 14977 12299 15011
rect 12541 14977 12575 15011
rect 13645 14977 13679 15011
rect 24869 14977 24903 15011
rect 27629 14977 27663 15011
rect 32689 14977 32723 15011
rect 35541 14977 35575 15011
rect 36737 14977 36771 15011
rect 39129 14977 39163 15011
rect 42073 14977 42107 15011
rect 43821 14977 43855 15011
rect 45293 14977 45327 15011
rect 47317 14977 47351 15011
rect 2329 14909 2363 14943
rect 3249 14909 3283 14943
rect 3893 14909 3927 14943
rect 4169 14909 4203 14943
rect 4445 14909 4479 14943
rect 5641 14909 5675 14943
rect 6653 14909 6687 14943
rect 6837 14909 6871 14943
rect 7021 14909 7055 14943
rect 7481 14909 7515 14943
rect 7573 14909 7607 14943
rect 9229 14909 9263 14943
rect 9689 14909 9723 14943
rect 9781 14909 9815 14943
rect 11529 14909 11563 14943
rect 12633 14909 12667 14943
rect 13093 14909 13127 14943
rect 13185 14909 13219 14943
rect 14841 14909 14875 14943
rect 15853 14909 15887 14943
rect 16865 14909 16899 14943
rect 18981 14909 19015 14943
rect 19717 14909 19751 14943
rect 20913 14909 20947 14943
rect 22201 14909 22235 14943
rect 22293 14909 22327 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 27537 14909 27571 14943
rect 30757 14909 30791 14943
rect 30849 14909 30883 14943
rect 31125 14909 31159 14943
rect 31309 14909 31343 14943
rect 32137 14909 32171 14943
rect 32321 14909 32355 14943
rect 33517 14909 33551 14943
rect 34989 14909 35023 14943
rect 35173 14909 35207 14943
rect 38485 14909 38519 14943
rect 38945 14909 38979 14943
rect 40509 14909 40543 14943
rect 40601 14909 40635 14943
rect 42165 14909 42199 14943
rect 42533 14909 42567 14943
rect 42717 14909 42751 14943
rect 43729 14909 43763 14943
rect 45017 14909 45051 14943
rect 49249 14909 49283 14943
rect 50537 14909 50571 14943
rect 52009 14909 52043 14943
rect 10333 14841 10367 14875
rect 19533 14841 19567 14875
rect 21005 14841 21039 14875
rect 30113 14841 30147 14875
rect 36369 14841 36403 14875
rect 41521 14841 41555 14875
rect 45109 14841 45143 14875
rect 46949 14841 46983 14875
rect 51917 14841 51951 14875
rect 52469 14841 52503 14875
rect 5457 14773 5491 14807
rect 8033 14773 8067 14807
rect 15669 14773 15703 14807
rect 16681 14773 16715 14807
rect 18797 14773 18831 14807
rect 19809 14773 19843 14807
rect 22937 14773 22971 14807
rect 24409 14773 24443 14807
rect 26433 14773 26467 14807
rect 31493 14773 31527 14807
rect 33609 14773 33643 14807
rect 37013 14773 37047 14807
rect 39589 14773 39623 14807
rect 49341 14773 49375 14807
rect 2237 14569 2271 14603
rect 3249 14569 3283 14603
rect 5825 14569 5859 14603
rect 6561 14569 6595 14603
rect 12817 14569 12851 14603
rect 13829 14569 13863 14603
rect 15393 14569 15427 14603
rect 24133 14569 24167 14603
rect 29193 14569 29227 14603
rect 31125 14569 31159 14603
rect 35725 14569 35759 14603
rect 41429 14569 41463 14603
rect 44097 14569 44131 14603
rect 48973 14569 49007 14603
rect 10517 14501 10551 14535
rect 18429 14501 18463 14535
rect 20085 14501 20119 14535
rect 22017 14501 22051 14535
rect 23397 14501 23431 14535
rect 37749 14501 37783 14535
rect 41153 14501 41187 14535
rect 45661 14501 45695 14535
rect 47593 14501 47627 14535
rect 2421 14433 2455 14467
rect 3433 14433 3467 14467
rect 4077 14433 4111 14467
rect 4353 14433 4387 14467
rect 6745 14433 6779 14467
rect 7757 14433 7791 14467
rect 8769 14433 8803 14467
rect 10793 14433 10827 14467
rect 10885 14433 10919 14467
rect 11345 14433 11379 14467
rect 11529 14433 11563 14467
rect 13001 14433 13035 14467
rect 14013 14433 14047 14467
rect 15301 14433 15335 14467
rect 19349 14433 19383 14467
rect 19441 14433 19475 14467
rect 19574 14433 19608 14467
rect 21833 14433 21867 14467
rect 22109 14433 22143 14467
rect 23581 14433 23615 14467
rect 25145 14433 25179 14467
rect 26525 14433 26559 14467
rect 27813 14433 27847 14467
rect 31033 14433 31067 14467
rect 33701 14433 33735 14467
rect 34069 14433 34103 14467
rect 35265 14433 35299 14467
rect 35541 14433 35575 14467
rect 37933 14433 37967 14467
rect 40141 14433 40175 14467
rect 41337 14433 41371 14467
rect 44005 14433 44039 14467
rect 44281 14433 44315 14467
rect 45845 14433 45879 14467
rect 47041 14433 47075 14467
rect 47225 14433 47259 14467
rect 49709 14433 49743 14467
rect 50077 14433 50111 14467
rect 50169 14433 50203 14467
rect 52285 14433 52319 14467
rect 16589 14365 16623 14399
rect 16865 14365 16899 14399
rect 19993 14365 20027 14399
rect 23857 14365 23891 14399
rect 28089 14365 28123 14399
rect 33793 14365 33827 14399
rect 34161 14365 34195 14399
rect 46213 14365 46247 14399
rect 48973 14365 49007 14399
rect 49617 14365 49651 14399
rect 52009 14365 52043 14399
rect 8585 14297 8619 14331
rect 18153 14297 18187 14331
rect 34437 14297 34471 14331
rect 35357 14297 35391 14331
rect 5457 14229 5491 14263
rect 7573 14229 7607 14263
rect 11805 14229 11839 14263
rect 22293 14229 22327 14263
rect 22753 14229 22787 14263
rect 25237 14229 25271 14263
rect 26617 14229 26651 14263
rect 29653 14229 29687 14263
rect 33149 14229 33183 14263
rect 38025 14229 38059 14263
rect 38485 14229 38519 14263
rect 40233 14229 40267 14263
rect 49157 14229 49191 14263
rect 51825 14229 51859 14263
rect 53389 14229 53423 14263
rect 5457 14025 5491 14059
rect 8125 14025 8159 14059
rect 10793 14025 10827 14059
rect 14841 14025 14875 14059
rect 18797 14025 18831 14059
rect 20821 14025 20855 14059
rect 21281 14025 21315 14059
rect 24317 14025 24351 14059
rect 26433 14025 26467 14059
rect 28273 14025 28307 14059
rect 29377 14025 29411 14059
rect 43729 14025 43763 14059
rect 44741 14025 44775 14059
rect 46305 14025 46339 14059
rect 47225 14025 47259 14059
rect 50721 14025 50755 14059
rect 52009 14025 52043 14059
rect 52469 14025 52503 14059
rect 4261 13957 4295 13991
rect 7573 13957 7607 13991
rect 9781 13957 9815 13991
rect 16957 13957 16991 13991
rect 21649 13957 21683 13991
rect 22569 13957 22603 13991
rect 32597 13957 32631 13991
rect 32965 13957 32999 13991
rect 33885 13957 33919 13991
rect 37381 13957 37415 13991
rect 45017 13957 45051 13991
rect 13553 13889 13587 13923
rect 15761 13889 15795 13923
rect 19625 13889 19659 13923
rect 25237 13889 25271 13923
rect 31217 13889 31251 13923
rect 42625 13889 42659 13923
rect 2329 13821 2363 13855
rect 3433 13821 3467 13855
rect 4445 13821 4479 13855
rect 5365 13821 5399 13855
rect 7757 13821 7791 13855
rect 8033 13821 8067 13855
rect 9965 13821 9999 13855
rect 10977 13821 11011 13855
rect 13277 13821 13311 13855
rect 15945 13821 15979 13855
rect 16405 13821 16439 13855
rect 16497 13821 16531 13855
rect 18981 13821 19015 13855
rect 19441 13821 19475 13855
rect 19809 13821 19843 13855
rect 21097 13821 21131 13855
rect 22753 13821 22787 13855
rect 24225 13821 24259 13855
rect 25053 13821 25087 13855
rect 25421 13821 25455 13855
rect 25881 13821 25915 13855
rect 25973 13821 26007 13855
rect 28181 13821 28215 13855
rect 29285 13821 29319 13855
rect 31493 13821 31527 13855
rect 33793 13821 33827 13855
rect 34069 13821 34103 13855
rect 35265 13821 35299 13855
rect 35449 13821 35483 13855
rect 35817 13821 35851 13855
rect 37565 13821 37599 13855
rect 37657 13821 37691 13855
rect 39405 13821 39439 13855
rect 39497 13821 39531 13855
rect 41245 13821 41279 13855
rect 42257 13821 42291 13855
rect 42349 13821 42383 13855
rect 44833 13821 44867 13855
rect 46121 13821 46155 13855
rect 46489 13821 46523 13855
rect 47501 13821 47535 13855
rect 49617 13821 49651 13855
rect 50629 13821 50663 13855
rect 51733 13821 51767 13855
rect 51917 13821 51951 13855
rect 21005 13753 21039 13787
rect 38117 13753 38151 13787
rect 39313 13753 39347 13787
rect 47409 13753 47443 13787
rect 47961 13753 47995 13787
rect 2145 13685 2179 13719
rect 3249 13685 3283 13719
rect 15025 13685 15059 13719
rect 41429 13685 41463 13719
rect 49709 13685 49743 13719
rect 4445 13481 4479 13515
rect 8677 13481 8711 13515
rect 16037 13481 16071 13515
rect 20729 13481 20763 13515
rect 22385 13481 22419 13515
rect 26801 13481 26835 13515
rect 29561 13481 29595 13515
rect 30021 13481 30055 13515
rect 31125 13481 31159 13515
rect 42165 13481 42199 13515
rect 45569 13481 45603 13515
rect 51457 13481 51491 13515
rect 16773 13413 16807 13447
rect 19257 13413 19291 13447
rect 24409 13413 24443 13447
rect 25697 13413 25731 13447
rect 32873 13413 32907 13447
rect 36553 13413 36587 13447
rect 2329 13345 2363 13379
rect 4997 13345 5031 13379
rect 5365 13345 5399 13379
rect 5457 13345 5491 13379
rect 6929 13345 6963 13379
rect 7205 13345 7239 13379
rect 9689 13345 9723 13379
rect 9965 13345 9999 13379
rect 12449 13345 12483 13379
rect 16221 13345 16255 13379
rect 16681 13345 16715 13379
rect 17877 13345 17911 13379
rect 18061 13345 18095 13379
rect 21281 13345 21315 13379
rect 25053 13345 25087 13379
rect 25421 13345 25455 13379
rect 26525 13345 26559 13379
rect 26709 13345 26743 13379
rect 28181 13345 28215 13379
rect 31033 13345 31067 13379
rect 32137 13345 32171 13379
rect 32413 13345 32447 13379
rect 34437 13345 34471 13379
rect 34529 13345 34563 13379
rect 36001 13345 36035 13379
rect 36185 13345 36219 13379
rect 38209 13345 38243 13379
rect 40877 13345 40911 13379
rect 41981 13345 42015 13379
rect 42349 13345 42383 13379
rect 44465 13345 44499 13379
rect 45477 13345 45511 13379
rect 45753 13345 45787 13379
rect 46949 13345 46983 13379
rect 47317 13345 47351 13379
rect 47501 13345 47535 13379
rect 50353 13345 50387 13379
rect 5089 13277 5123 13311
rect 11437 13277 11471 13311
rect 12173 13277 12207 13311
rect 13921 13277 13955 13311
rect 18429 13277 18463 13311
rect 19625 13277 19659 13311
rect 21005 13277 21039 13311
rect 25145 13277 25179 13311
rect 25513 13277 25547 13311
rect 28457 13277 28491 13311
rect 32229 13277 32263 13311
rect 34989 13277 35023 13311
rect 37933 13277 37967 13311
rect 39313 13277 39347 13311
rect 43637 13277 43671 13311
rect 44189 13277 44223 13311
rect 44649 13277 44683 13311
rect 49985 13277 50019 13311
rect 50077 13277 50111 13311
rect 19533 13209 19567 13243
rect 34253 13209 34287 13243
rect 2145 13141 2179 13175
rect 8309 13141 8343 13175
rect 11069 13141 11103 13175
rect 13553 13141 13587 13175
rect 19422 13141 19456 13175
rect 19901 13141 19935 13175
rect 39773 13141 39807 13175
rect 41061 13141 41095 13175
rect 2237 12937 2271 12971
rect 7113 12937 7147 12971
rect 10425 12937 10459 12971
rect 13093 12937 13127 12971
rect 14933 12937 14967 12971
rect 16681 12937 16715 12971
rect 19809 12937 19843 12971
rect 21373 12937 21407 12971
rect 25697 12937 25731 12971
rect 29653 12937 29687 12971
rect 30941 12937 30975 12971
rect 41705 12937 41739 12971
rect 47869 12937 47903 12971
rect 49341 12937 49375 12971
rect 8861 12869 8895 12903
rect 18797 12869 18831 12903
rect 19349 12869 19383 12903
rect 20269 12869 20303 12903
rect 25237 12869 25271 12903
rect 26065 12869 26099 12903
rect 36829 12869 36863 12903
rect 37657 12869 37691 12903
rect 39957 12869 39991 12903
rect 44097 12869 44131 12903
rect 7389 12801 7423 12835
rect 15117 12801 15151 12835
rect 30113 12801 30147 12835
rect 33977 12801 34011 12835
rect 35357 12801 35391 12835
rect 44833 12801 44867 12835
rect 47133 12801 47167 12835
rect 47961 12801 47995 12835
rect 48237 12801 48271 12835
rect 2413 12733 2447 12767
rect 3433 12733 3467 12767
rect 4445 12733 4479 12767
rect 5457 12733 5491 12767
rect 7481 12733 7515 12767
rect 7849 12733 7883 12767
rect 8033 12733 8067 12767
rect 9045 12733 9079 12767
rect 10333 12733 10367 12767
rect 11529 12733 11563 12767
rect 13001 12733 13035 12767
rect 14197 12733 14231 12767
rect 15393 12733 15427 12767
rect 18981 12733 19015 12767
rect 19625 12733 19659 12767
rect 21565 12733 21599 12767
rect 22569 12733 22603 12767
rect 24041 12733 24075 12767
rect 25513 12733 25547 12767
rect 26801 12733 26835 12767
rect 27997 12733 28031 12767
rect 30205 12733 30239 12767
rect 30573 12733 30607 12767
rect 30757 12733 30791 12767
rect 31769 12733 31803 12767
rect 31953 12733 31987 12767
rect 33425 12733 33459 12767
rect 33609 12733 33643 12767
rect 35081 12733 35115 12767
rect 37565 12733 37599 12767
rect 39129 12733 39163 12767
rect 39405 12733 39439 12767
rect 40693 12733 40727 12767
rect 41061 12733 41095 12767
rect 41797 12733 41831 12767
rect 43729 12733 43763 12767
rect 43821 12733 43855 12767
rect 44373 12733 44407 12767
rect 46581 12733 46615 12767
rect 46765 12733 46799 12767
rect 19533 12665 19567 12699
rect 23857 12665 23891 12699
rect 24409 12665 24443 12699
rect 25421 12665 25455 12699
rect 27813 12665 27847 12699
rect 28365 12665 28399 12699
rect 32321 12665 32355 12699
rect 39589 12665 39623 12699
rect 39773 12665 39807 12699
rect 3249 12597 3283 12631
rect 4261 12597 4295 12631
rect 5273 12597 5307 12631
rect 11345 12597 11379 12631
rect 14013 12597 14047 12631
rect 22385 12597 22419 12631
rect 26893 12597 26927 12631
rect 36461 12597 36495 12631
rect 40877 12597 40911 12631
rect 41981 12597 42015 12631
rect 2881 12393 2915 12427
rect 4813 12393 4847 12427
rect 7849 12393 7883 12427
rect 9965 12393 9999 12427
rect 21189 12393 21223 12427
rect 26801 12393 26835 12427
rect 29101 12393 29135 12427
rect 34253 12393 34287 12427
rect 40785 12393 40819 12427
rect 41245 12393 41279 12427
rect 43085 12393 43119 12427
rect 44741 12393 44775 12427
rect 13829 12325 13863 12359
rect 20913 12325 20947 12359
rect 26525 12325 26559 12359
rect 28365 12325 28399 12359
rect 31217 12325 31251 12359
rect 3065 12257 3099 12291
rect 4997 12257 5031 12291
rect 6009 12257 6043 12291
rect 7021 12257 7055 12291
rect 8033 12257 8067 12291
rect 9045 12257 9079 12291
rect 10333 12257 10367 12291
rect 10701 12257 10735 12291
rect 13093 12257 13127 12291
rect 13461 12257 13495 12291
rect 16221 12257 16255 12291
rect 16681 12257 16715 12291
rect 17141 12257 17175 12291
rect 17509 12257 17543 12291
rect 19441 12257 19475 12291
rect 19625 12257 19659 12291
rect 19809 12257 19843 12291
rect 21097 12257 21131 12291
rect 22569 12257 22603 12291
rect 25145 12257 25179 12291
rect 25605 12257 25639 12291
rect 26709 12257 26743 12291
rect 28457 12257 28491 12291
rect 30481 12257 30515 12291
rect 32965 12257 32999 12291
rect 34161 12257 34195 12291
rect 34437 12257 34471 12291
rect 35357 12257 35391 12291
rect 35449 12257 35483 12291
rect 39405 12257 39439 12291
rect 43361 12257 43395 12291
rect 43637 12257 43671 12291
rect 10425 12189 10459 12223
rect 10609 12189 10643 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 22201 12189 22235 12223
rect 22293 12189 22327 12223
rect 23857 12189 23891 12223
rect 30628 12189 30662 12223
rect 30849 12189 30883 12223
rect 32137 12189 32171 12223
rect 32689 12189 32723 12223
rect 32827 12189 32861 12223
rect 39681 12189 39715 12223
rect 12725 12121 12759 12155
rect 16589 12121 16623 12155
rect 28181 12121 28215 12155
rect 30757 12121 30791 12155
rect 35173 12121 35207 12155
rect 5825 12053 5859 12087
rect 6837 12053 6871 12087
rect 8861 12053 8895 12087
rect 16037 12053 16071 12087
rect 17785 12053 17819 12087
rect 24961 12053 24995 12087
rect 28641 12053 28675 12087
rect 35633 12053 35667 12087
rect 36093 12053 36127 12087
rect 2145 11849 2179 11883
rect 7573 11849 7607 11883
rect 8585 11849 8619 11883
rect 14197 11849 14231 11883
rect 15209 11849 15243 11883
rect 18797 11849 18831 11883
rect 30021 11849 30055 11883
rect 33609 11849 33643 11883
rect 36829 11849 36863 11883
rect 11621 11781 11655 11815
rect 24317 11781 24351 11815
rect 31033 11781 31067 11815
rect 31861 11781 31895 11815
rect 32873 11781 32907 11815
rect 16037 11713 16071 11747
rect 16589 11713 16623 11747
rect 17049 11713 17083 11747
rect 19165 11713 19199 11747
rect 19257 11713 19291 11747
rect 19533 11713 19567 11747
rect 24501 11713 24535 11747
rect 35265 11713 35299 11747
rect 37013 11713 37047 11747
rect 2329 11645 2363 11679
rect 3525 11645 3559 11679
rect 4537 11645 4571 11679
rect 5549 11645 5583 11679
rect 7757 11645 7791 11679
rect 8769 11645 8803 11679
rect 9781 11645 9815 11679
rect 10793 11645 10827 11679
rect 11805 11645 11839 11679
rect 13369 11645 13403 11679
rect 14381 11645 14415 11679
rect 15393 11645 15427 11679
rect 16865 11645 16899 11679
rect 18981 11645 19015 11679
rect 21925 11645 21959 11679
rect 24777 11645 24811 11679
rect 27169 11645 27203 11679
rect 30205 11645 30239 11679
rect 31217 11645 31251 11679
rect 31585 11645 31619 11679
rect 32321 11645 32355 11679
rect 32597 11645 32631 11679
rect 33517 11645 33551 11679
rect 34897 11645 34931 11679
rect 35449 11645 35483 11679
rect 37289 11645 37323 11679
rect 20913 11577 20947 11611
rect 26985 11577 27019 11611
rect 3341 11509 3375 11543
rect 4353 11509 4387 11543
rect 5365 11509 5399 11543
rect 9597 11509 9631 11543
rect 10609 11509 10643 11543
rect 13185 11509 13219 11543
rect 21741 11509 21775 11543
rect 25881 11509 25915 11543
rect 27261 11509 27295 11543
rect 38393 11509 38427 11543
rect 2145 11305 2179 11339
rect 6837 11305 6871 11339
rect 7849 11305 7883 11339
rect 8861 11305 8895 11339
rect 11437 11305 11471 11339
rect 13461 11305 13495 11339
rect 21005 11305 21039 11339
rect 27261 11305 27295 11339
rect 32229 11305 32263 11339
rect 25421 11237 25455 11271
rect 25605 11237 25639 11271
rect 29561 11237 29595 11271
rect 30113 11237 30147 11271
rect 33149 11237 33183 11271
rect 33701 11237 33735 11271
rect 35081 11237 35115 11271
rect 2329 11169 2363 11203
rect 4997 11169 5031 11203
rect 6009 11169 6043 11203
rect 7021 11169 7055 11203
rect 8033 11169 8067 11203
rect 9045 11169 9079 11203
rect 10609 11169 10643 11203
rect 11621 11169 11655 11203
rect 12633 11169 12667 11203
rect 13645 11169 13679 11203
rect 16221 11169 16255 11203
rect 17233 11169 17267 11203
rect 18245 11169 18279 11203
rect 19257 11169 19291 11203
rect 20269 11169 20303 11203
rect 20913 11169 20947 11203
rect 22109 11169 22143 11203
rect 23121 11169 23155 11203
rect 24133 11169 24167 11203
rect 24685 11169 24719 11203
rect 24869 11169 24903 11203
rect 24961 11169 24995 11203
rect 27445 11169 27479 11203
rect 27997 11169 28031 11203
rect 28365 11169 28399 11203
rect 28549 11169 28583 11203
rect 29745 11169 29779 11203
rect 32137 11169 32171 11203
rect 33333 11169 33367 11203
rect 34529 11169 34563 11203
rect 34713 11169 34747 11203
rect 4813 11033 4847 11067
rect 10425 11033 10459 11067
rect 16037 11033 16071 11067
rect 19073 11033 19107 11067
rect 21925 11033 21959 11067
rect 22937 11033 22971 11067
rect 5825 10965 5859 10999
rect 12449 10965 12483 10999
rect 17049 10965 17083 10999
rect 18061 10965 18095 10999
rect 20085 10965 20119 10999
rect 23949 10965 23983 10999
rect 2145 10761 2179 10795
rect 6193 10761 6227 10795
rect 8585 10761 8619 10795
rect 11437 10761 11471 10795
rect 13185 10761 13219 10795
rect 14197 10761 14231 10795
rect 17233 10761 17267 10795
rect 25697 10761 25731 10795
rect 32137 10761 32171 10795
rect 32597 10761 32631 10795
rect 18797 10693 18831 10727
rect 21833 10693 21867 10727
rect 30757 10625 30791 10659
rect 2329 10557 2363 10591
rect 3341 10557 3375 10591
rect 4353 10557 4387 10591
rect 5365 10557 5399 10591
rect 6377 10557 6411 10591
rect 7757 10557 7791 10591
rect 8769 10557 8803 10591
rect 10609 10557 10643 10591
rect 11621 10557 11655 10591
rect 13369 10557 13403 10591
rect 14381 10557 14415 10591
rect 15393 10557 15427 10591
rect 16405 10557 16439 10591
rect 17417 10557 17451 10591
rect 18981 10557 19015 10591
rect 19993 10557 20027 10591
rect 21005 10557 21039 10591
rect 22017 10557 22051 10591
rect 23029 10557 23063 10591
rect 24777 10557 24811 10591
rect 25605 10557 25639 10591
rect 27445 10557 27479 10591
rect 30205 10557 30239 10591
rect 31033 10557 31067 10591
rect 35817 10557 35851 10591
rect 3157 10421 3191 10455
rect 4169 10421 4203 10455
rect 5181 10421 5215 10455
rect 7573 10421 7607 10455
rect 10425 10421 10459 10455
rect 15209 10421 15243 10455
rect 16221 10421 16255 10455
rect 19809 10421 19843 10455
rect 20821 10421 20855 10455
rect 22845 10421 22879 10455
rect 24593 10421 24627 10455
rect 27261 10421 27295 10455
rect 30021 10421 30055 10455
rect 35633 10421 35667 10455
rect 2237 10217 2271 10251
rect 7021 10217 7055 10251
rect 8033 10217 8067 10251
rect 11529 10217 11563 10251
rect 12541 10217 12575 10251
rect 13553 10217 13587 10251
rect 16037 10217 16071 10251
rect 17049 10217 17083 10251
rect 18061 10217 18095 10251
rect 20085 10217 20119 10251
rect 21649 10217 21683 10251
rect 22661 10217 22695 10251
rect 25421 10217 25455 10251
rect 29285 10217 29319 10251
rect 2421 10081 2455 10115
rect 3433 10081 3467 10115
rect 4997 10081 5031 10115
rect 6009 10081 6043 10115
rect 7205 10081 7239 10115
rect 8217 10081 8251 10115
rect 9505 10081 9539 10115
rect 10701 10081 10735 10115
rect 11713 10081 11747 10115
rect 12725 10081 12759 10115
rect 13737 10081 13771 10115
rect 16221 10081 16255 10115
rect 17233 10081 17267 10115
rect 18245 10081 18279 10115
rect 19257 10081 19291 10115
rect 20269 10081 20303 10115
rect 21833 10081 21867 10115
rect 22845 10081 22879 10115
rect 24593 10081 24627 10115
rect 25605 10081 25639 10115
rect 27445 10081 27479 10115
rect 28457 10081 28491 10115
rect 29469 10081 29503 10115
rect 30481 10081 30515 10115
rect 33241 10081 33275 10115
rect 34253 10081 34287 10115
rect 35265 10081 35299 10115
rect 36277 10081 36311 10115
rect 5825 9945 5859 9979
rect 9321 9945 9355 9979
rect 3249 9877 3283 9911
rect 4813 9877 4847 9911
rect 10517 9877 10551 9911
rect 19073 9877 19107 9911
rect 24409 9877 24443 9911
rect 27261 9877 27295 9911
rect 28273 9877 28307 9911
rect 30297 9877 30331 9911
rect 33057 9877 33091 9911
rect 34069 9877 34103 9911
rect 35081 9877 35115 9911
rect 36093 9877 36127 9911
rect 7573 9673 7607 9707
rect 13185 9673 13219 9707
rect 27445 9673 27479 9707
rect 3433 9605 3467 9639
rect 4445 9605 4479 9639
rect 14197 9605 14231 9639
rect 17233 9605 17267 9639
rect 21833 9605 21867 9639
rect 24409 9605 24443 9639
rect 28917 9605 28951 9639
rect 32781 9605 32815 9639
rect 36645 9605 36679 9639
rect 37657 9605 37691 9639
rect 2605 9469 2639 9503
rect 3617 9469 3651 9503
rect 4629 9469 4663 9503
rect 5917 9469 5951 9503
rect 7757 9469 7791 9503
rect 8769 9469 8803 9503
rect 10701 9469 10735 9503
rect 13369 9469 13403 9503
rect 14381 9469 14415 9503
rect 15393 9469 15427 9503
rect 16405 9469 16439 9503
rect 17417 9469 17451 9503
rect 18981 9469 19015 9503
rect 19993 9469 20027 9503
rect 21005 9469 21039 9503
rect 22017 9469 22051 9503
rect 23029 9469 23063 9503
rect 24593 9469 24627 9503
rect 25605 9469 25639 9503
rect 26617 9469 26651 9503
rect 27629 9469 27663 9503
rect 29101 9469 29135 9503
rect 30941 9469 30975 9503
rect 31953 9469 31987 9503
rect 32965 9469 32999 9503
rect 33977 9469 34011 9503
rect 35817 9469 35851 9503
rect 36829 9469 36863 9503
rect 37841 9469 37875 9503
rect 2421 9333 2455 9367
rect 5733 9333 5767 9367
rect 8585 9333 8619 9367
rect 10517 9333 10551 9367
rect 15209 9333 15243 9367
rect 16221 9333 16255 9367
rect 18797 9333 18831 9367
rect 19809 9333 19843 9367
rect 20821 9333 20855 9367
rect 22845 9333 22879 9367
rect 25421 9333 25455 9367
rect 26433 9333 26467 9367
rect 30757 9333 30791 9367
rect 31769 9333 31803 9367
rect 33793 9333 33827 9367
rect 35633 9333 35667 9367
rect 4813 9129 4847 9163
rect 7481 9129 7515 9163
rect 12449 9129 12483 9163
rect 13461 9129 13495 9163
rect 16037 9129 16071 9163
rect 20085 9129 20119 9163
rect 21649 9129 21683 9163
rect 24133 9129 24167 9163
rect 25145 9129 25179 9163
rect 28733 9129 28767 9163
rect 29745 9129 29779 9163
rect 31769 9129 31803 9163
rect 33149 9129 33183 9163
rect 38485 9129 38519 9163
rect 16865 9061 16899 9095
rect 3157 8993 3191 9027
rect 4997 8993 5031 9027
rect 6653 8993 6687 9027
rect 7665 8993 7699 9027
rect 8677 8993 8711 9027
rect 10609 8993 10643 9027
rect 11621 8993 11655 9027
rect 12633 8993 12667 9027
rect 13645 8993 13679 9027
rect 16221 8993 16255 9027
rect 17233 8993 17267 9027
rect 18245 8993 18279 9027
rect 19257 8993 19291 9027
rect 20269 8993 20303 9027
rect 21833 8993 21867 9027
rect 23305 8993 23339 9027
rect 24317 8993 24351 9027
rect 25329 8993 25363 9027
rect 26341 8993 26375 9027
rect 27905 8993 27939 9027
rect 28917 8993 28951 9027
rect 29929 8993 29963 9027
rect 30941 8993 30975 9027
rect 31953 8993 31987 9027
rect 33333 8993 33367 9027
rect 34345 8993 34379 9027
rect 35357 8993 35391 9027
rect 36369 8993 36403 9027
rect 38669 8993 38703 9027
rect 2973 8857 3007 8891
rect 11437 8857 11471 8891
rect 17049 8857 17083 8891
rect 19073 8857 19107 8891
rect 36185 8857 36219 8891
rect 6469 8789 6503 8823
rect 8493 8789 8527 8823
rect 10425 8789 10459 8823
rect 18061 8789 18095 8823
rect 23121 8789 23155 8823
rect 26157 8789 26191 8823
rect 27721 8789 27755 8823
rect 30757 8789 30791 8823
rect 34161 8789 34195 8823
rect 35173 8789 35207 8823
rect 2881 8585 2915 8619
rect 5457 8585 5491 8619
rect 8585 8585 8619 8619
rect 13185 8585 13219 8619
rect 16957 8585 16991 8619
rect 21833 8585 21867 8619
rect 25145 8585 25179 8619
rect 27169 8585 27203 8619
rect 30573 8585 30607 8619
rect 31769 8585 31803 8619
rect 32781 8585 32815 8619
rect 33793 8585 33827 8619
rect 37657 8585 37691 8619
rect 4445 8517 4479 8551
rect 6469 8517 6503 8551
rect 7573 8517 7607 8551
rect 10609 8517 10643 8551
rect 14197 8517 14231 8551
rect 15209 8517 15243 8551
rect 19809 8517 19843 8551
rect 20821 8517 20855 8551
rect 26157 8517 26191 8551
rect 28181 8517 28215 8551
rect 36645 8517 36679 8551
rect 3065 8381 3099 8415
rect 4629 8381 4663 8415
rect 5641 8381 5675 8415
rect 6653 8381 6687 8415
rect 7757 8381 7791 8415
rect 8769 8381 8803 8415
rect 9781 8381 9815 8415
rect 10793 8381 10827 8415
rect 13369 8381 13403 8415
rect 14381 8381 14415 8415
rect 15393 8381 15427 8415
rect 17141 8381 17175 8415
rect 18981 8381 19015 8415
rect 19993 8381 20027 8415
rect 21005 8381 21039 8415
rect 22017 8381 22051 8415
rect 23029 8381 23063 8415
rect 25329 8381 25363 8415
rect 26341 8381 26375 8415
rect 27353 8381 27387 8415
rect 28365 8381 28399 8415
rect 30757 8381 30791 8415
rect 31953 8381 31987 8415
rect 32965 8381 32999 8415
rect 33977 8381 34011 8415
rect 35817 8381 35851 8415
rect 36829 8381 36863 8415
rect 37841 8381 37875 8415
rect 9597 8245 9631 8279
rect 18797 8245 18831 8279
rect 22845 8245 22879 8279
rect 35633 8245 35667 8279
rect 2145 8041 2179 8075
rect 5549 8041 5583 8075
rect 7573 8041 7607 8075
rect 11437 8041 11471 8075
rect 12449 8041 12483 8075
rect 13461 8041 13495 8075
rect 14933 8041 14967 8075
rect 19625 8041 19659 8075
rect 21649 8041 21683 8075
rect 23121 8041 23155 8075
rect 24133 8041 24167 8075
rect 25145 8041 25179 8075
rect 27537 8041 27571 8075
rect 28549 8041 28583 8075
rect 29561 8041 29595 8075
rect 33793 8041 33827 8075
rect 2329 7905 2363 7939
rect 3341 7905 3375 7939
rect 5733 7905 5767 7939
rect 6745 7905 6779 7939
rect 7757 7905 7791 7939
rect 8769 7905 8803 7939
rect 10609 7905 10643 7939
rect 11621 7905 11655 7939
rect 12633 7905 12667 7939
rect 13645 7905 13679 7939
rect 15117 7905 15151 7939
rect 16221 7905 16255 7939
rect 17233 7905 17267 7939
rect 18797 7905 18831 7939
rect 19809 7905 19843 7939
rect 21833 7905 21867 7939
rect 23305 7905 23339 7939
rect 24317 7905 24351 7939
rect 25329 7905 25363 7939
rect 26341 7905 26375 7939
rect 27721 7905 27755 7939
rect 28733 7905 28767 7939
rect 29745 7905 29779 7939
rect 33977 7905 34011 7939
rect 34989 7905 35023 7939
rect 36001 7905 36035 7939
rect 37013 7905 37047 7939
rect 8585 7769 8619 7803
rect 3157 7701 3191 7735
rect 6561 7701 6595 7735
rect 10425 7701 10459 7735
rect 16037 7701 16071 7735
rect 17049 7701 17083 7735
rect 18613 7701 18647 7735
rect 26157 7701 26191 7735
rect 34805 7701 34839 7735
rect 35817 7701 35851 7735
rect 36829 7701 36863 7735
rect 3525 7497 3559 7531
rect 5733 7497 5767 7531
rect 7573 7497 7607 7531
rect 13185 7497 13219 7531
rect 20821 7497 20855 7531
rect 22569 7497 22603 7531
rect 27353 7497 27387 7531
rect 30021 7497 30055 7531
rect 32781 7497 32815 7531
rect 33793 7497 33827 7531
rect 2145 7429 2179 7463
rect 25421 7429 25455 7463
rect 2329 7293 2363 7327
rect 3717 7293 3751 7327
rect 4721 7293 4755 7327
rect 5917 7293 5951 7327
rect 7757 7293 7791 7327
rect 8769 7293 8803 7327
rect 9781 7293 9815 7327
rect 10793 7293 10827 7327
rect 13369 7293 13403 7327
rect 14381 7293 14415 7327
rect 15393 7293 15427 7327
rect 16405 7293 16439 7327
rect 17785 7293 17819 7327
rect 18981 7293 19015 7327
rect 19993 7293 20027 7327
rect 21005 7293 21039 7327
rect 22753 7293 22787 7327
rect 24593 7293 24627 7327
rect 25605 7293 25639 7327
rect 27537 7293 27571 7327
rect 30205 7293 30239 7327
rect 32965 7293 32999 7327
rect 33977 7293 34011 7327
rect 35817 7293 35851 7327
rect 36829 7293 36863 7327
rect 38025 7293 38059 7327
rect 4537 7157 4571 7191
rect 8585 7157 8619 7191
rect 9597 7157 9631 7191
rect 10609 7157 10643 7191
rect 14197 7157 14231 7191
rect 15209 7157 15243 7191
rect 16221 7157 16255 7191
rect 17601 7157 17635 7191
rect 18797 7157 18831 7191
rect 19809 7157 19843 7191
rect 24409 7157 24443 7191
rect 35633 7157 35667 7191
rect 36645 7157 36679 7191
rect 37841 7157 37875 7191
rect 5641 6953 5675 6987
rect 16037 6953 16071 6987
rect 21649 6953 21683 6987
rect 22753 6953 22787 6987
rect 24777 6953 24811 6987
rect 29561 6953 29595 6987
rect 33609 6953 33643 6987
rect 2881 6817 2915 6851
rect 3893 6817 3927 6851
rect 5825 6817 5859 6851
rect 7665 6817 7699 6851
rect 8677 6817 8711 6851
rect 10609 6817 10643 6851
rect 11621 6817 11655 6851
rect 12725 6817 12759 6851
rect 13737 6817 13771 6851
rect 16221 6817 16255 6851
rect 17233 6817 17267 6851
rect 18245 6817 18279 6851
rect 19257 6817 19291 6851
rect 20269 6817 20303 6851
rect 21833 6817 21867 6851
rect 22937 6817 22971 6851
rect 23949 6817 23983 6851
rect 24961 6817 24995 6851
rect 25973 6817 26007 6851
rect 27445 6817 27479 6851
rect 29745 6817 29779 6851
rect 33793 6817 33827 6851
rect 34805 6817 34839 6851
rect 35817 6817 35851 6851
rect 36921 6817 36955 6851
rect 38669 6817 38703 6851
rect 39681 6817 39715 6851
rect 7481 6681 7515 6715
rect 8493 6681 8527 6715
rect 12541 6681 12575 6715
rect 35633 6681 35667 6715
rect 36737 6681 36771 6715
rect 2697 6613 2731 6647
rect 3709 6613 3743 6647
rect 10425 6613 10459 6647
rect 11437 6613 11471 6647
rect 13553 6613 13587 6647
rect 17049 6613 17083 6647
rect 18061 6613 18095 6647
rect 19073 6613 19107 6647
rect 20085 6613 20119 6647
rect 23765 6613 23799 6647
rect 25789 6613 25823 6647
rect 27261 6613 27295 6647
rect 34621 6613 34655 6647
rect 38485 6613 38519 6647
rect 39497 6613 39531 6647
rect 4721 6409 4755 6443
rect 5733 6409 5767 6443
rect 8217 6409 8251 6443
rect 9229 6409 9263 6443
rect 15209 6409 15243 6443
rect 16221 6409 16255 6443
rect 22569 6409 22603 6443
rect 33793 6409 33827 6443
rect 35633 6409 35667 6443
rect 36645 6409 36679 6443
rect 2697 6341 2731 6375
rect 25421 6341 25455 6375
rect 2881 6205 2915 6239
rect 3893 6205 3927 6239
rect 4905 6205 4939 6239
rect 5917 6205 5951 6239
rect 8401 6205 8435 6239
rect 9413 6205 9447 6239
rect 10425 6205 10459 6239
rect 11437 6205 11471 6239
rect 13369 6205 13403 6239
rect 14381 6205 14415 6239
rect 15393 6205 15427 6239
rect 16405 6205 16439 6239
rect 17417 6205 17451 6239
rect 18981 6205 19015 6239
rect 19993 6205 20027 6239
rect 21005 6205 21039 6239
rect 22753 6205 22787 6239
rect 24593 6205 24627 6239
rect 25605 6205 25639 6239
rect 26617 6205 26651 6239
rect 27629 6205 27663 6239
rect 28641 6205 28675 6239
rect 30205 6205 30239 6239
rect 33977 6205 34011 6239
rect 35817 6205 35851 6239
rect 36829 6205 36863 6239
rect 37933 6205 37967 6239
rect 38945 6205 38979 6239
rect 3709 6069 3743 6103
rect 10241 6069 10275 6103
rect 11253 6069 11287 6103
rect 13185 6069 13219 6103
rect 14197 6069 14231 6103
rect 17233 6069 17267 6103
rect 18797 6069 18831 6103
rect 19809 6069 19843 6103
rect 20821 6069 20855 6103
rect 24409 6069 24443 6103
rect 26433 6069 26467 6103
rect 27445 6069 27479 6103
rect 28457 6069 28491 6103
rect 30021 6069 30055 6103
rect 37749 6069 37783 6103
rect 38761 6069 38795 6103
rect 2145 5865 2179 5899
rect 7849 5865 7883 5899
rect 10425 5865 10459 5899
rect 13461 5865 13495 5899
rect 14473 5865 14507 5899
rect 16037 5865 16071 5899
rect 17049 5865 17083 5899
rect 18061 5865 18095 5899
rect 20085 5865 20119 5899
rect 21649 5865 21683 5899
rect 22661 5865 22695 5899
rect 24685 5865 24719 5899
rect 35357 5865 35391 5899
rect 36369 5865 36403 5899
rect 37381 5865 37415 5899
rect 40509 5865 40543 5899
rect 2329 5729 2363 5763
rect 4997 5729 5031 5763
rect 6009 5729 6043 5763
rect 7021 5729 7055 5763
rect 8033 5729 8067 5763
rect 9045 5729 9079 5763
rect 10609 5729 10643 5763
rect 11621 5729 11655 5763
rect 12633 5729 12667 5763
rect 13645 5729 13679 5763
rect 14657 5729 14691 5763
rect 16221 5729 16255 5763
rect 17233 5729 17267 5763
rect 18245 5729 18279 5763
rect 19257 5729 19291 5763
rect 20269 5729 20303 5763
rect 21833 5729 21867 5763
rect 22845 5729 22879 5763
rect 23865 5729 23899 5763
rect 24869 5729 24903 5763
rect 25881 5729 25915 5763
rect 26341 5729 26375 5763
rect 27445 5729 27479 5763
rect 28457 5729 28491 5763
rect 29469 5729 29503 5763
rect 30481 5729 30515 5763
rect 35541 5729 35575 5763
rect 36553 5729 36587 5763
rect 37565 5729 37599 5763
rect 38669 5729 38703 5763
rect 39681 5729 39715 5763
rect 40693 5729 40727 5763
rect 4813 5593 4847 5627
rect 5825 5593 5859 5627
rect 6837 5593 6871 5627
rect 8861 5593 8895 5627
rect 19073 5593 19107 5627
rect 25697 5593 25731 5627
rect 39497 5593 39531 5627
rect 11437 5525 11471 5559
rect 12449 5525 12483 5559
rect 23673 5525 23707 5559
rect 26341 5525 26375 5559
rect 27261 5525 27295 5559
rect 28273 5525 28307 5559
rect 29285 5525 29319 5559
rect 30297 5525 30331 5559
rect 38485 5525 38519 5559
rect 2145 5321 2179 5355
rect 5181 5321 5215 5355
rect 8585 5321 8619 5355
rect 10609 5321 10643 5355
rect 11621 5321 11655 5355
rect 16129 5321 16163 5355
rect 18797 5321 18831 5355
rect 21097 5321 21131 5355
rect 24409 5321 24443 5355
rect 36369 5321 36403 5355
rect 41245 5321 41279 5355
rect 13185 5253 13219 5287
rect 15117 5253 15151 5287
rect 22109 5253 22143 5287
rect 30021 5253 30055 5287
rect 2329 5117 2363 5151
rect 5365 5117 5399 5151
rect 7757 5117 7791 5151
rect 8769 5117 8803 5151
rect 9781 5117 9815 5151
rect 10793 5117 10827 5151
rect 11805 5117 11839 5151
rect 13369 5117 13403 5151
rect 15301 5117 15335 5151
rect 16313 5117 16347 5151
rect 18981 5117 19015 5151
rect 19993 5117 20027 5151
rect 21281 5117 21315 5151
rect 22293 5117 22327 5151
rect 23305 5117 23339 5151
rect 24593 5117 24627 5151
rect 25605 5117 25639 5151
rect 26617 5117 26651 5151
rect 27629 5117 27663 5151
rect 28641 5117 28675 5151
rect 30205 5117 30239 5151
rect 31217 5117 31251 5151
rect 36553 5117 36587 5151
rect 37565 5117 37599 5151
rect 38577 5117 38611 5151
rect 39589 5117 39623 5151
rect 41429 5117 41463 5151
rect 7573 4981 7607 5015
rect 9597 4981 9631 5015
rect 19809 4981 19843 5015
rect 23121 4981 23155 5015
rect 25421 4981 25455 5015
rect 26433 4981 26467 5015
rect 27445 4981 27479 5015
rect 28457 4981 28491 5015
rect 31033 4981 31067 5015
rect 37381 4981 37415 5015
rect 38393 4981 38427 5015
rect 39405 4981 39439 5015
rect 6377 4777 6411 4811
rect 8401 4777 8435 4811
rect 14105 4777 14139 4811
rect 15945 4777 15979 4811
rect 17877 4777 17911 4811
rect 18889 4777 18923 4811
rect 22661 4777 22695 4811
rect 24961 4777 24995 4811
rect 31309 4777 31343 4811
rect 38761 4777 38795 4811
rect 40785 4777 40819 4811
rect 5549 4641 5583 4675
rect 6561 4641 6595 4675
rect 7573 4641 7607 4675
rect 8585 4641 8619 4675
rect 13277 4641 13311 4675
rect 14289 4641 14323 4675
rect 16221 4641 16255 4675
rect 18061 4641 18095 4675
rect 19073 4641 19107 4675
rect 20637 4641 20671 4675
rect 21833 4641 21867 4675
rect 22845 4641 22879 4675
rect 23857 4641 23891 4675
rect 25145 4641 25179 4675
rect 26157 4641 26191 4675
rect 27445 4641 27479 4675
rect 28457 4641 28491 4675
rect 29469 4641 29503 4675
rect 30481 4641 30515 4675
rect 31493 4641 31527 4675
rect 33057 4641 33091 4675
rect 35817 4641 35851 4675
rect 37565 4641 37599 4675
rect 38945 4641 38979 4675
rect 39957 4641 39991 4675
rect 40969 4641 41003 4675
rect 5365 4505 5399 4539
rect 7389 4505 7423 4539
rect 16037 4505 16071 4539
rect 20453 4505 20487 4539
rect 37381 4505 37415 4539
rect 13093 4437 13127 4471
rect 21649 4437 21683 4471
rect 23673 4437 23707 4471
rect 25973 4437 26007 4471
rect 27261 4437 27295 4471
rect 28273 4437 28307 4471
rect 29285 4437 29319 4471
rect 30297 4437 30331 4471
rect 32873 4437 32907 4471
rect 35633 4437 35667 4471
rect 39773 4437 39807 4471
rect 6469 4233 6503 4267
rect 13185 4233 13219 4267
rect 14197 4233 14231 4267
rect 18797 4233 18831 4267
rect 22477 4233 22511 4267
rect 32689 4233 32723 4267
rect 7849 4165 7883 4199
rect 6653 4029 6687 4063
rect 8033 4029 8067 4063
rect 13369 4029 13403 4063
rect 14381 4029 14415 4063
rect 15577 4029 15611 4063
rect 16589 4029 16623 4063
rect 18981 4029 19015 4063
rect 19993 4029 20027 4063
rect 21005 4029 21039 4063
rect 22661 4029 22695 4063
rect 24593 4029 24627 4063
rect 25605 4029 25639 4063
rect 26617 4029 26651 4063
rect 27629 4029 27663 4063
rect 28641 4029 28675 4063
rect 30849 4029 30883 4063
rect 31861 4029 31895 4063
rect 32873 4029 32907 4063
rect 33885 4029 33919 4063
rect 35817 4029 35851 4063
rect 36829 4029 36863 4063
rect 38577 4029 38611 4063
rect 39589 4029 39623 4063
rect 41429 4029 41463 4063
rect 15393 3893 15427 3927
rect 16405 3893 16439 3927
rect 19809 3893 19843 3927
rect 20821 3893 20855 3927
rect 24409 3893 24443 3927
rect 25421 3893 25455 3927
rect 26433 3893 26467 3927
rect 27445 3893 27479 3927
rect 28457 3893 28491 3927
rect 30665 3893 30699 3927
rect 31677 3893 31711 3927
rect 33701 3893 33735 3927
rect 35633 3893 35667 3927
rect 36645 3893 36679 3927
rect 38393 3893 38427 3927
rect 39405 3893 39439 3927
rect 41245 3893 41279 3927
rect 14013 3689 14047 3723
rect 16405 3689 16439 3723
rect 21649 3689 21683 3723
rect 24777 3689 24811 3723
rect 28273 3689 28307 3723
rect 35909 3689 35943 3723
rect 42533 3689 42567 3723
rect 14197 3553 14231 3587
rect 16589 3553 16623 3587
rect 18889 3553 18923 3587
rect 21833 3553 21867 3587
rect 22937 3553 22971 3587
rect 23949 3553 23983 3587
rect 24961 3553 24995 3587
rect 25973 3553 26007 3587
rect 27445 3553 27479 3587
rect 28457 3553 28491 3587
rect 29469 3553 29503 3587
rect 30573 3553 30607 3587
rect 33057 3553 33091 3587
rect 34069 3553 34103 3587
rect 35081 3553 35115 3587
rect 36093 3553 36127 3587
rect 37105 3553 37139 3587
rect 38669 3553 38703 3587
rect 39681 3553 39715 3587
rect 40693 3553 40727 3587
rect 41705 3553 41739 3587
rect 42717 3553 42751 3587
rect 22753 3417 22787 3451
rect 23765 3417 23799 3451
rect 34897 3417 34931 3451
rect 41521 3417 41555 3451
rect 18705 3349 18739 3383
rect 25789 3349 25823 3383
rect 27261 3349 27295 3383
rect 29285 3349 29319 3383
rect 30389 3349 30423 3383
rect 32873 3349 32907 3383
rect 33885 3349 33919 3383
rect 36921 3349 36955 3383
rect 38485 3349 38519 3383
rect 39497 3349 39531 3383
rect 40509 3349 40543 3383
rect 21741 3145 21775 3179
rect 25789 3145 25823 3179
rect 26801 3145 26835 3179
rect 32045 3145 32079 3179
rect 33057 3145 33091 3179
rect 34069 3145 34103 3179
rect 35633 3145 35667 3179
rect 36645 3145 36679 3179
rect 39681 3145 39715 3179
rect 41245 3145 41279 3179
rect 42257 3145 42291 3179
rect 20729 3077 20763 3111
rect 24777 3077 24811 3111
rect 20913 2941 20947 2975
rect 21925 2941 21959 2975
rect 22937 2941 22971 2975
rect 24961 2941 24995 2975
rect 25973 2941 26007 2975
rect 26985 2941 27019 2975
rect 27997 2941 28031 2975
rect 30205 2941 30239 2975
rect 31217 2941 31251 2975
rect 32229 2941 32263 2975
rect 33241 2941 33275 2975
rect 34253 2941 34287 2975
rect 35817 2941 35851 2975
rect 36829 2941 36863 2975
rect 37841 2941 37875 2975
rect 38853 2941 38887 2975
rect 39865 2941 39899 2975
rect 41429 2941 41463 2975
rect 42441 2941 42475 2975
rect 22753 2805 22787 2839
rect 27813 2805 27847 2839
rect 30021 2805 30055 2839
rect 31033 2805 31067 2839
rect 37657 2805 37691 2839
rect 38669 2805 38703 2839
rect 20821 2601 20855 2635
rect 22661 2601 22695 2635
rect 27629 2601 27663 2635
rect 28641 2601 28675 2635
rect 30481 2601 30515 2635
rect 31493 2601 31527 2635
rect 34345 2601 34379 2635
rect 36185 2601 36219 2635
rect 37197 2601 37231 2635
rect 39037 2601 39071 2635
rect 40049 2601 40083 2635
rect 41889 2601 41923 2635
rect 19993 2465 20027 2499
rect 21005 2465 21039 2499
rect 22845 2465 22879 2499
rect 23857 2465 23891 2499
rect 24961 2465 24995 2499
rect 25973 2465 26007 2499
rect 27813 2465 27847 2499
rect 28825 2465 28859 2499
rect 30665 2465 30699 2499
rect 31677 2465 31711 2499
rect 33517 2465 33551 2499
rect 34529 2465 34563 2499
rect 36369 2465 36403 2499
rect 37381 2465 37415 2499
rect 39221 2465 39255 2499
rect 40233 2465 40267 2499
rect 42073 2465 42107 2499
rect 43085 2465 43119 2499
rect 23673 2329 23707 2363
rect 24777 2329 24811 2363
rect 25789 2329 25823 2363
rect 42901 2329 42935 2363
rect 19809 2261 19843 2295
rect 33333 2261 33367 2295
<< metal1 >>
rect 1104 25050 54832 25072
rect 1104 24998 9947 25050
rect 9999 24998 10011 25050
rect 10063 24998 10075 25050
rect 10127 24998 10139 25050
rect 10191 24998 27878 25050
rect 27930 24998 27942 25050
rect 27994 24998 28006 25050
rect 28058 24998 28070 25050
rect 28122 24998 45808 25050
rect 45860 24998 45872 25050
rect 45924 24998 45936 25050
rect 45988 24998 46000 25050
rect 46052 24998 54832 25050
rect 1104 24976 54832 24998
rect 38841 24871 38899 24877
rect 38841 24837 38853 24871
rect 38887 24837 38899 24871
rect 38841 24831 38899 24837
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24800 8631 24803
rect 8846 24800 8852 24812
rect 8619 24772 8852 24800
rect 8619 24769 8631 24772
rect 8573 24763 8631 24769
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 21818 24760 21824 24812
rect 21876 24800 21882 24812
rect 22833 24803 22891 24809
rect 22833 24800 22845 24803
rect 21876 24772 22845 24800
rect 21876 24760 21882 24772
rect 22833 24769 22845 24772
rect 22879 24769 22891 24803
rect 22833 24763 22891 24769
rect 34974 24760 34980 24812
rect 35032 24800 35038 24812
rect 38856 24800 38884 24831
rect 35032 24772 38884 24800
rect 35032 24760 35038 24772
rect 6917 24735 6975 24741
rect 6917 24701 6929 24735
rect 6963 24701 6975 24735
rect 7190 24732 7196 24744
rect 7151 24704 7196 24732
rect 6917 24695 6975 24701
rect 6546 24556 6552 24608
rect 6604 24596 6610 24608
rect 6932 24596 6960 24695
rect 7190 24692 7196 24704
rect 7248 24692 7254 24744
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24701 21511 24735
rect 21453 24695 21511 24701
rect 21729 24735 21787 24741
rect 21729 24701 21741 24735
rect 21775 24732 21787 24735
rect 22462 24732 22468 24744
rect 21775 24704 22468 24732
rect 21775 24701 21787 24704
rect 21729 24695 21787 24701
rect 8662 24596 8668 24608
rect 6604 24568 8668 24596
rect 6604 24556 6610 24568
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 21361 24599 21419 24605
rect 21361 24565 21373 24599
rect 21407 24596 21419 24599
rect 21468 24596 21496 24695
rect 22462 24692 22468 24704
rect 22520 24692 22526 24744
rect 38657 24735 38715 24741
rect 38657 24732 38669 24735
rect 38488 24704 38669 24732
rect 38488 24664 38516 24704
rect 38657 24701 38669 24704
rect 38703 24701 38715 24735
rect 38856 24732 38884 24772
rect 40494 24760 40500 24812
rect 40552 24800 40558 24812
rect 42613 24803 42671 24809
rect 42613 24800 42625 24803
rect 40552 24772 42625 24800
rect 40552 24760 40558 24772
rect 42613 24769 42625 24772
rect 42659 24769 42671 24803
rect 42613 24763 42671 24769
rect 43346 24760 43352 24812
rect 43404 24800 43410 24812
rect 47486 24800 47492 24812
rect 43404 24772 47492 24800
rect 43404 24760 43410 24772
rect 47486 24760 47492 24772
rect 47544 24760 47550 24812
rect 48498 24760 48504 24812
rect 48556 24800 48562 24812
rect 49973 24803 50031 24809
rect 49973 24800 49985 24803
rect 48556 24772 49985 24800
rect 48556 24760 48562 24772
rect 49973 24769 49985 24772
rect 50019 24769 50031 24803
rect 49973 24763 50031 24769
rect 39761 24735 39819 24741
rect 39761 24732 39773 24735
rect 38856 24704 39773 24732
rect 38657 24695 38715 24701
rect 39761 24701 39773 24704
rect 39807 24732 39819 24735
rect 40402 24732 40408 24744
rect 39807 24704 40408 24732
rect 39807 24701 39819 24704
rect 39761 24695 39819 24701
rect 40402 24692 40408 24704
rect 40460 24692 40466 24744
rect 41230 24732 41236 24744
rect 41191 24704 41236 24732
rect 41230 24692 41236 24704
rect 41288 24692 41294 24744
rect 41509 24735 41567 24741
rect 41509 24701 41521 24735
rect 41555 24732 41567 24735
rect 41966 24732 41972 24744
rect 41555 24704 41972 24732
rect 41555 24701 41567 24704
rect 41509 24695 41567 24701
rect 41966 24692 41972 24704
rect 42024 24692 42030 24744
rect 43993 24735 44051 24741
rect 43993 24732 44005 24735
rect 43732 24704 44005 24732
rect 38488 24636 40080 24664
rect 21542 24596 21548 24608
rect 21407 24568 21548 24596
rect 21407 24565 21419 24568
rect 21361 24559 21419 24565
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 24394 24556 24400 24608
rect 24452 24596 24458 24608
rect 38488 24605 38516 24636
rect 38473 24599 38531 24605
rect 38473 24596 38485 24599
rect 24452 24568 38485 24596
rect 24452 24556 24458 24568
rect 38473 24565 38485 24568
rect 38519 24565 38531 24599
rect 39942 24596 39948 24608
rect 39903 24568 39948 24596
rect 38473 24559 38531 24565
rect 39942 24556 39948 24568
rect 40000 24556 40006 24608
rect 40052 24596 40080 24636
rect 42886 24596 42892 24608
rect 40052 24568 42892 24596
rect 42886 24556 42892 24568
rect 42944 24556 42950 24608
rect 42978 24556 42984 24608
rect 43036 24596 43042 24608
rect 43732 24605 43760 24704
rect 43993 24701 44005 24704
rect 44039 24701 44051 24735
rect 44266 24732 44272 24744
rect 44227 24704 44272 24732
rect 43993 24695 44051 24701
rect 44266 24692 44272 24704
rect 44324 24692 44330 24744
rect 49697 24735 49755 24741
rect 49697 24732 49709 24735
rect 49436 24704 49709 24732
rect 43717 24599 43775 24605
rect 43717 24596 43729 24599
rect 43036 24568 43729 24596
rect 43036 24556 43042 24568
rect 43717 24565 43729 24568
rect 43763 24596 43775 24599
rect 44542 24596 44548 24608
rect 43763 24568 44548 24596
rect 43763 24565 43775 24568
rect 43717 24559 43775 24565
rect 44542 24556 44548 24568
rect 44600 24556 44606 24608
rect 45554 24596 45560 24608
rect 45515 24568 45560 24596
rect 45554 24556 45560 24568
rect 45612 24556 45618 24608
rect 48590 24556 48596 24608
rect 48648 24596 48654 24608
rect 49436 24605 49464 24704
rect 49697 24701 49709 24704
rect 49743 24732 49755 24735
rect 50614 24732 50620 24744
rect 49743 24704 50620 24732
rect 49743 24701 49755 24704
rect 49697 24695 49755 24701
rect 50614 24692 50620 24704
rect 50672 24692 50678 24744
rect 49421 24599 49479 24605
rect 49421 24596 49433 24599
rect 48648 24568 49433 24596
rect 48648 24556 48654 24568
rect 49421 24565 49433 24568
rect 49467 24565 49479 24599
rect 51074 24596 51080 24608
rect 51035 24568 51080 24596
rect 49421 24559 49479 24565
rect 51074 24556 51080 24568
rect 51132 24556 51138 24608
rect 1104 24506 54832 24528
rect 1104 24454 18912 24506
rect 18964 24454 18976 24506
rect 19028 24454 19040 24506
rect 19092 24454 19104 24506
rect 19156 24454 36843 24506
rect 36895 24454 36907 24506
rect 36959 24454 36971 24506
rect 37023 24454 37035 24506
rect 37087 24454 54832 24506
rect 1104 24432 54832 24454
rect 1670 24352 1676 24404
rect 1728 24392 1734 24404
rect 2777 24395 2835 24401
rect 2777 24392 2789 24395
rect 1728 24364 2789 24392
rect 1728 24352 1734 24364
rect 2777 24361 2789 24364
rect 2823 24361 2835 24395
rect 2777 24355 2835 24361
rect 7466 24352 7472 24404
rect 7524 24392 7530 24404
rect 7929 24395 7987 24401
rect 7929 24392 7941 24395
rect 7524 24364 7941 24392
rect 7524 24352 7530 24364
rect 7929 24361 7941 24364
rect 7975 24361 7987 24395
rect 7929 24355 7987 24361
rect 13170 24352 13176 24404
rect 13228 24392 13234 24404
rect 13817 24395 13875 24401
rect 13817 24392 13829 24395
rect 13228 24364 13829 24392
rect 13228 24352 13234 24364
rect 13817 24361 13829 24364
rect 13863 24361 13875 24395
rect 13817 24355 13875 24361
rect 16022 24352 16028 24404
rect 16080 24392 16086 24404
rect 16669 24395 16727 24401
rect 16669 24392 16681 24395
rect 16080 24364 16681 24392
rect 16080 24352 16086 24364
rect 16669 24361 16681 24364
rect 16715 24361 16727 24395
rect 16669 24355 16727 24361
rect 17494 24352 17500 24404
rect 17552 24392 17558 24404
rect 19337 24395 19395 24401
rect 19337 24392 19349 24395
rect 17552 24364 19349 24392
rect 17552 24352 17558 24364
rect 19337 24361 19349 24364
rect 19383 24361 19395 24395
rect 19337 24355 19395 24361
rect 20346 24352 20352 24404
rect 20404 24392 20410 24404
rect 22281 24395 22339 24401
rect 22281 24392 22293 24395
rect 20404 24364 22293 24392
rect 20404 24352 20410 24364
rect 22281 24361 22293 24364
rect 22327 24361 22339 24395
rect 22281 24355 22339 24361
rect 23474 24352 23480 24404
rect 23532 24392 23538 24404
rect 24949 24395 25007 24401
rect 24949 24392 24961 24395
rect 23532 24364 24961 24392
rect 23532 24352 23538 24364
rect 24949 24361 24961 24364
rect 24995 24361 25007 24395
rect 24949 24355 25007 24361
rect 27614 24352 27620 24404
rect 27672 24392 27678 24404
rect 27893 24395 27951 24401
rect 27893 24392 27905 24395
rect 27672 24364 27905 24392
rect 27672 24352 27678 24364
rect 27893 24361 27905 24364
rect 27939 24361 27951 24395
rect 30374 24392 30380 24404
rect 30335 24364 30380 24392
rect 27893 24355 27951 24361
rect 30374 24352 30380 24364
rect 30432 24352 30438 24404
rect 33318 24352 33324 24404
rect 33376 24392 33382 24404
rect 33689 24395 33747 24401
rect 33689 24392 33701 24395
rect 33376 24364 33701 24392
rect 33376 24352 33382 24364
rect 33689 24361 33701 24364
rect 33735 24361 33747 24395
rect 33689 24355 33747 24361
rect 34698 24352 34704 24404
rect 34756 24392 34762 24404
rect 36173 24395 36231 24401
rect 36173 24392 36185 24395
rect 34756 24364 36185 24392
rect 34756 24352 34762 24364
rect 36173 24361 36185 24364
rect 36219 24361 36231 24395
rect 36173 24355 36231 24361
rect 39022 24352 39028 24404
rect 39080 24392 39086 24404
rect 39853 24395 39911 24401
rect 39853 24392 39865 24395
rect 39080 24364 39865 24392
rect 39080 24352 39086 24364
rect 39853 24361 39865 24364
rect 39899 24361 39911 24395
rect 39853 24355 39911 24361
rect 50522 24352 50528 24404
rect 50580 24392 50586 24404
rect 52549 24395 52607 24401
rect 52549 24392 52561 24395
rect 50580 24364 52561 24392
rect 50580 24352 50586 24364
rect 52549 24361 52561 24364
rect 52595 24361 52607 24395
rect 52549 24355 52607 24361
rect 5721 24327 5779 24333
rect 5721 24293 5733 24327
rect 5767 24324 5779 24327
rect 5994 24324 6000 24336
rect 5767 24296 6000 24324
rect 5767 24293 5779 24296
rect 5721 24287 5779 24293
rect 5994 24284 6000 24296
rect 6052 24284 6058 24336
rect 11609 24327 11667 24333
rect 11609 24293 11621 24327
rect 11655 24324 11667 24327
rect 11698 24324 11704 24336
rect 11655 24296 11704 24324
rect 11655 24293 11667 24296
rect 11609 24287 11667 24293
rect 11698 24284 11704 24296
rect 11756 24284 11762 24336
rect 42886 24284 42892 24336
rect 42944 24324 42950 24336
rect 50614 24324 50620 24336
rect 42944 24296 46060 24324
rect 50575 24296 50620 24324
rect 42944 24284 42950 24296
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24256 1731 24259
rect 1719 24228 5856 24256
rect 1719 24225 1731 24228
rect 1673 24219 1731 24225
rect 1397 24191 1455 24197
rect 1397 24157 1409 24191
rect 1443 24188 1455 24191
rect 4065 24191 4123 24197
rect 1443 24160 3280 24188
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 3252 24061 3280 24160
rect 4065 24157 4077 24191
rect 4111 24157 4123 24191
rect 4065 24151 4123 24157
rect 4080 24064 4108 24151
rect 4246 24148 4252 24200
rect 4304 24188 4310 24200
rect 4341 24191 4399 24197
rect 4341 24188 4353 24191
rect 4304 24160 4353 24188
rect 4304 24148 4310 24160
rect 4341 24157 4353 24160
rect 4387 24157 4399 24191
rect 5828 24188 5856 24228
rect 5902 24216 5908 24268
rect 5960 24256 5966 24268
rect 6546 24256 6552 24268
rect 5960 24228 6552 24256
rect 5960 24216 5966 24228
rect 6546 24216 6552 24228
rect 6604 24216 6610 24268
rect 8389 24259 8447 24265
rect 8389 24225 8401 24259
rect 8435 24256 8447 24259
rect 8662 24256 8668 24268
rect 8435 24228 8668 24256
rect 8435 24225 8447 24228
rect 8389 24219 8447 24225
rect 8662 24216 8668 24228
rect 8720 24256 8726 24268
rect 9766 24256 9772 24268
rect 8720 24228 9772 24256
rect 8720 24216 8726 24228
rect 9766 24216 9772 24228
rect 9824 24256 9830 24268
rect 9953 24259 10011 24265
rect 9953 24256 9965 24259
rect 9824 24228 9965 24256
rect 9824 24216 9830 24228
rect 9953 24225 9965 24228
rect 9999 24256 10011 24259
rect 11793 24259 11851 24265
rect 11793 24256 11805 24259
rect 9999 24228 11805 24256
rect 9999 24225 10011 24228
rect 9953 24219 10011 24225
rect 11793 24225 11805 24228
rect 11839 24256 11851 24259
rect 12437 24259 12495 24265
rect 12437 24256 12449 24259
rect 11839 24228 12449 24256
rect 11839 24225 11851 24228
rect 11793 24219 11851 24225
rect 12437 24225 12449 24228
rect 12483 24256 12495 24259
rect 13630 24256 13636 24268
rect 12483 24228 13636 24256
rect 12483 24225 12495 24228
rect 12437 24219 12495 24225
rect 13630 24216 13636 24228
rect 13688 24256 13694 24268
rect 14185 24259 14243 24265
rect 14185 24256 14197 24259
rect 13688 24228 14197 24256
rect 13688 24216 13694 24228
rect 14185 24225 14197 24228
rect 14231 24256 14243 24259
rect 15013 24259 15071 24265
rect 15013 24256 15025 24259
rect 14231 24228 15025 24256
rect 14231 24225 14243 24228
rect 14185 24219 14243 24225
rect 15013 24225 15025 24228
rect 15059 24256 15071 24259
rect 15289 24259 15347 24265
rect 15289 24256 15301 24259
rect 15059 24228 15301 24256
rect 15059 24225 15071 24228
rect 15013 24219 15071 24225
rect 15289 24225 15301 24228
rect 15335 24256 15347 24259
rect 15378 24256 15384 24268
rect 15335 24228 15384 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15378 24216 15384 24228
rect 15436 24216 15442 24268
rect 15565 24259 15623 24265
rect 15565 24225 15577 24259
rect 15611 24256 15623 24259
rect 19426 24256 19432 24268
rect 15611 24228 19432 24256
rect 15611 24225 15623 24228
rect 15565 24219 15623 24225
rect 19426 24216 19432 24228
rect 19484 24216 19490 24268
rect 20717 24259 20775 24265
rect 20717 24225 20729 24259
rect 20763 24256 20775 24259
rect 20901 24259 20959 24265
rect 20901 24256 20913 24259
rect 20763 24228 20913 24256
rect 20763 24225 20775 24228
rect 20717 24219 20775 24225
rect 20901 24225 20913 24228
rect 20947 24256 20959 24259
rect 21542 24256 21548 24268
rect 20947 24228 21548 24256
rect 20947 24225 20959 24228
rect 20901 24219 20959 24225
rect 21542 24216 21548 24228
rect 21600 24256 21606 24268
rect 23201 24259 23259 24265
rect 23201 24256 23213 24259
rect 21600 24228 23213 24256
rect 21600 24216 21606 24228
rect 23201 24225 23213 24228
rect 23247 24256 23259 24259
rect 23385 24259 23443 24265
rect 23385 24256 23397 24259
rect 23247 24228 23397 24256
rect 23247 24225 23259 24228
rect 23201 24219 23259 24225
rect 23385 24225 23397 24228
rect 23431 24256 23443 24259
rect 25222 24256 25228 24268
rect 23431 24228 25228 24256
rect 23431 24225 23443 24228
rect 23385 24219 23443 24225
rect 25222 24216 25228 24228
rect 25280 24256 25286 24268
rect 26237 24259 26295 24265
rect 26237 24256 26249 24259
rect 25280 24228 26249 24256
rect 25280 24216 25286 24228
rect 26237 24225 26249 24228
rect 26283 24256 26295 24259
rect 26513 24259 26571 24265
rect 26513 24256 26525 24259
rect 26283 24228 26525 24256
rect 26283 24225 26295 24228
rect 26237 24219 26295 24225
rect 26513 24225 26525 24228
rect 26559 24225 26571 24259
rect 26513 24219 26571 24225
rect 26789 24259 26847 24265
rect 26789 24225 26801 24259
rect 26835 24256 26847 24259
rect 31478 24256 31484 24268
rect 26835 24228 31484 24256
rect 26835 24225 26847 24228
rect 26789 24219 26847 24225
rect 31478 24216 31484 24228
rect 31536 24216 31542 24268
rect 34057 24259 34115 24265
rect 34057 24256 34069 24259
rect 32324 24228 34069 24256
rect 32324 24200 32352 24228
rect 34057 24225 34069 24228
rect 34103 24256 34115 24259
rect 34793 24259 34851 24265
rect 34793 24256 34805 24259
rect 34103 24228 34805 24256
rect 34103 24225 34115 24228
rect 34057 24219 34115 24225
rect 34793 24225 34805 24228
rect 34839 24256 34851 24259
rect 35894 24256 35900 24268
rect 34839 24228 35900 24256
rect 34839 24225 34851 24228
rect 34793 24219 34851 24225
rect 35894 24216 35900 24228
rect 35952 24256 35958 24268
rect 36541 24259 36599 24265
rect 36541 24256 36553 24259
rect 35952 24228 36553 24256
rect 35952 24216 35958 24228
rect 36541 24225 36553 24228
rect 36587 24225 36599 24259
rect 36541 24219 36599 24225
rect 38473 24259 38531 24265
rect 38473 24225 38485 24259
rect 38519 24256 38531 24259
rect 40221 24259 40279 24265
rect 40221 24256 40233 24259
rect 38519 24228 40233 24256
rect 38519 24225 38531 24228
rect 38473 24219 38531 24225
rect 40221 24225 40233 24228
rect 40267 24256 40279 24259
rect 41230 24256 41236 24268
rect 40267 24228 41236 24256
rect 40267 24225 40279 24228
rect 40221 24219 40279 24225
rect 41230 24216 41236 24228
rect 41288 24256 41294 24268
rect 42978 24256 42984 24268
rect 41288 24228 42984 24256
rect 41288 24216 41294 24228
rect 42978 24216 42984 24228
rect 43036 24216 43042 24268
rect 46032 24256 46060 24296
rect 50614 24284 50620 24296
rect 50672 24324 50678 24336
rect 50672 24296 51028 24324
rect 50672 24284 50678 24296
rect 51000 24265 51028 24296
rect 50985 24259 51043 24265
rect 46032 24228 47808 24256
rect 6822 24188 6828 24200
rect 5828 24160 5948 24188
rect 6783 24160 6828 24188
rect 4341 24151 4399 24157
rect 3237 24055 3295 24061
rect 3237 24021 3249 24055
rect 3283 24052 3295 24055
rect 4062 24052 4068 24064
rect 3283 24024 4068 24052
rect 3283 24021 3295 24024
rect 3237 24015 3295 24021
rect 4062 24012 4068 24024
rect 4120 24052 4126 24064
rect 5810 24052 5816 24064
rect 4120 24024 5816 24052
rect 4120 24012 4126 24024
rect 5810 24012 5816 24024
rect 5868 24012 5874 24064
rect 5920 24052 5948 24160
rect 6822 24148 6828 24160
rect 6880 24148 6886 24200
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10410 24188 10416 24200
rect 10275 24160 10416 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 10410 24148 10416 24160
rect 10468 24148 10474 24200
rect 12618 24148 12624 24200
rect 12676 24188 12682 24200
rect 12713 24191 12771 24197
rect 12713 24188 12725 24191
rect 12676 24160 12725 24188
rect 12676 24148 12682 24160
rect 12713 24157 12725 24160
rect 12759 24157 12771 24191
rect 12713 24151 12771 24157
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24188 17739 24191
rect 17770 24188 17776 24200
rect 17727 24160 17776 24188
rect 17727 24157 17739 24160
rect 17681 24151 17739 24157
rect 17770 24148 17776 24160
rect 17828 24148 17834 24200
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 20806 24188 20812 24200
rect 18095 24160 20812 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 20806 24148 20812 24160
rect 20864 24148 20870 24200
rect 21174 24188 21180 24200
rect 21135 24160 21180 24188
rect 21174 24148 21180 24160
rect 21232 24148 21238 24200
rect 23658 24188 23664 24200
rect 23619 24160 23664 24188
rect 23658 24148 23664 24160
rect 23716 24148 23722 24200
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24157 29055 24191
rect 28997 24151 29055 24157
rect 29273 24191 29331 24197
rect 29273 24157 29285 24191
rect 29319 24188 29331 24191
rect 32214 24188 32220 24200
rect 29319 24160 32220 24188
rect 29319 24157 29331 24160
rect 29273 24151 29331 24157
rect 9674 24120 9680 24132
rect 7484 24092 9680 24120
rect 7484 24052 7512 24092
rect 9674 24080 9680 24092
rect 9732 24080 9738 24132
rect 5920 24024 7512 24052
rect 29012 24052 29040 24151
rect 32214 24148 32220 24160
rect 32272 24148 32278 24200
rect 32306 24148 32312 24200
rect 32364 24188 32370 24200
rect 32585 24191 32643 24197
rect 32364 24160 32409 24188
rect 32364 24148 32370 24160
rect 32585 24157 32597 24191
rect 32631 24188 32643 24191
rect 33686 24188 33692 24200
rect 32631 24160 33692 24188
rect 32631 24157 32643 24160
rect 32585 24151 32643 24157
rect 33686 24148 33692 24160
rect 33744 24148 33750 24200
rect 35066 24188 35072 24200
rect 35027 24160 35072 24188
rect 35066 24148 35072 24160
rect 35124 24148 35130 24200
rect 38746 24188 38752 24200
rect 38707 24160 38752 24188
rect 38746 24148 38752 24160
rect 38804 24148 38810 24200
rect 45925 24191 45983 24197
rect 45925 24188 45937 24191
rect 45756 24160 45937 24188
rect 29362 24052 29368 24064
rect 29012 24024 29368 24052
rect 29362 24012 29368 24024
rect 29420 24012 29426 24064
rect 30742 24052 30748 24064
rect 30703 24024 30748 24052
rect 30742 24012 30748 24024
rect 30800 24012 30806 24064
rect 44542 24012 44548 24064
rect 44600 24052 44606 24064
rect 45370 24052 45376 24064
rect 44600 24024 45376 24052
rect 44600 24012 44606 24024
rect 45370 24012 45376 24024
rect 45428 24052 45434 24064
rect 45756 24061 45784 24160
rect 45925 24157 45937 24160
rect 45971 24157 45983 24191
rect 45925 24151 45983 24157
rect 46201 24191 46259 24197
rect 46201 24157 46213 24191
rect 46247 24188 46259 24191
rect 46566 24188 46572 24200
rect 46247 24160 46572 24188
rect 46247 24157 46259 24160
rect 46201 24151 46259 24157
rect 46566 24148 46572 24160
rect 46624 24148 46630 24200
rect 47780 24120 47808 24228
rect 50985 24225 50997 24259
rect 51031 24225 51043 24259
rect 50985 24219 51043 24225
rect 51261 24259 51319 24265
rect 51261 24225 51273 24259
rect 51307 24256 51319 24259
rect 54846 24256 54852 24268
rect 51307 24228 54852 24256
rect 51307 24225 51319 24228
rect 51261 24219 51319 24225
rect 50893 24191 50951 24197
rect 50893 24157 50905 24191
rect 50939 24188 50951 24191
rect 51276 24188 51304 24219
rect 54846 24216 54852 24228
rect 54904 24216 54910 24268
rect 50939 24160 51304 24188
rect 50939 24157 50951 24160
rect 50893 24151 50951 24157
rect 50908 24120 50936 24151
rect 47780 24092 50936 24120
rect 45741 24055 45799 24061
rect 45741 24052 45753 24055
rect 45428 24024 45753 24052
rect 45428 24012 45434 24024
rect 45741 24021 45753 24024
rect 45787 24021 45799 24055
rect 45741 24015 45799 24021
rect 46658 24012 46664 24064
rect 46716 24052 46722 24064
rect 47305 24055 47363 24061
rect 47305 24052 47317 24055
rect 46716 24024 47317 24052
rect 46716 24012 46722 24024
rect 47305 24021 47317 24024
rect 47351 24021 47363 24055
rect 47305 24015 47363 24021
rect 1104 23962 54832 23984
rect 1104 23910 9947 23962
rect 9999 23910 10011 23962
rect 10063 23910 10075 23962
rect 10127 23910 10139 23962
rect 10191 23910 27878 23962
rect 27930 23910 27942 23962
rect 27994 23910 28006 23962
rect 28058 23910 28070 23962
rect 28122 23910 45808 23962
rect 45860 23910 45872 23962
rect 45924 23910 45936 23962
rect 45988 23910 46000 23962
rect 46052 23910 54832 23962
rect 1104 23888 54832 23910
rect 10045 23851 10103 23857
rect 10045 23817 10057 23851
rect 10091 23848 10103 23851
rect 10318 23848 10324 23860
rect 10091 23820 10324 23848
rect 10091 23817 10103 23820
rect 10045 23811 10103 23817
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 14642 23808 14648 23860
rect 14700 23848 14706 23860
rect 15013 23851 15071 23857
rect 15013 23848 15025 23851
rect 14700 23820 15025 23848
rect 14700 23808 14706 23820
rect 15013 23817 15025 23820
rect 15059 23817 15071 23851
rect 15013 23811 15071 23817
rect 15102 23808 15108 23860
rect 15160 23848 15166 23860
rect 15378 23848 15384 23860
rect 15160 23820 15384 23848
rect 15160 23808 15166 23820
rect 15378 23808 15384 23820
rect 15436 23808 15442 23860
rect 18064 23820 19288 23848
rect 18064 23780 18092 23820
rect 14660 23752 18092 23780
rect 19260 23780 19288 23820
rect 19334 23808 19340 23860
rect 19392 23848 19398 23860
rect 19429 23851 19487 23857
rect 19429 23848 19441 23851
rect 19392 23820 19441 23848
rect 19392 23808 19398 23820
rect 19429 23817 19441 23820
rect 19475 23817 19487 23851
rect 22462 23848 22468 23860
rect 22423 23820 22468 23848
rect 19429 23811 19487 23817
rect 22462 23808 22468 23820
rect 22520 23808 22526 23860
rect 25222 23848 25228 23860
rect 25183 23820 25228 23848
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 26142 23808 26148 23860
rect 26200 23848 26206 23860
rect 26789 23851 26847 23857
rect 26789 23848 26801 23851
rect 26200 23820 26801 23848
rect 26200 23808 26206 23820
rect 26789 23817 26801 23820
rect 26835 23817 26847 23851
rect 26789 23811 26847 23817
rect 31846 23808 31852 23860
rect 31904 23848 31910 23860
rect 31941 23851 31999 23857
rect 31941 23848 31953 23851
rect 31904 23820 31953 23848
rect 31904 23808 31910 23820
rect 31941 23817 31953 23820
rect 31987 23817 31999 23851
rect 31941 23811 31999 23817
rect 32214 23808 32220 23860
rect 32272 23848 32278 23860
rect 33689 23851 33747 23857
rect 33689 23848 33701 23851
rect 32272 23820 33701 23848
rect 32272 23808 32278 23820
rect 33689 23817 33701 23820
rect 33735 23817 33747 23851
rect 35894 23848 35900 23860
rect 35855 23820 35900 23848
rect 33689 23811 33747 23817
rect 35894 23808 35900 23820
rect 35952 23808 35958 23860
rect 36262 23808 36268 23860
rect 36320 23848 36326 23860
rect 37461 23851 37519 23857
rect 37461 23848 37473 23851
rect 36320 23820 37473 23848
rect 36320 23808 36326 23820
rect 37461 23817 37473 23820
rect 37507 23817 37519 23851
rect 37461 23811 37519 23817
rect 38746 23808 38752 23860
rect 38804 23848 38810 23860
rect 39301 23851 39359 23857
rect 39301 23848 39313 23851
rect 38804 23820 39313 23848
rect 38804 23808 38810 23820
rect 39301 23817 39313 23820
rect 39347 23817 39359 23851
rect 41966 23848 41972 23860
rect 41927 23820 41972 23848
rect 39301 23811 39359 23817
rect 41966 23808 41972 23820
rect 42024 23808 42030 23860
rect 44266 23848 44272 23860
rect 44227 23820 44272 23848
rect 44266 23808 44272 23820
rect 44324 23808 44330 23860
rect 46566 23848 46572 23860
rect 46527 23820 46572 23848
rect 46566 23808 46572 23820
rect 46624 23808 46630 23860
rect 49050 23808 49056 23860
rect 49108 23848 49114 23860
rect 49513 23851 49571 23857
rect 49513 23848 49525 23851
rect 49108 23820 49525 23848
rect 49108 23808 49114 23820
rect 49513 23817 49525 23820
rect 49559 23817 49571 23851
rect 49513 23811 49571 23817
rect 21358 23780 21364 23792
rect 19260 23752 21364 23780
rect 5460 23684 5856 23712
rect 5460 23653 5488 23684
rect 5445 23647 5503 23653
rect 5445 23613 5457 23647
rect 5491 23613 5503 23647
rect 5445 23607 5503 23613
rect 5721 23647 5779 23653
rect 5721 23613 5733 23647
rect 5767 23613 5779 23647
rect 5828 23644 5856 23684
rect 7190 23672 7196 23724
rect 7248 23712 7254 23724
rect 7377 23715 7435 23721
rect 7377 23712 7389 23715
rect 7248 23684 7389 23712
rect 7248 23672 7254 23684
rect 7377 23681 7389 23684
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23712 8539 23715
rect 9766 23712 9772 23724
rect 8527 23684 9772 23712
rect 8527 23681 8539 23684
rect 8481 23675 8539 23681
rect 9766 23672 9772 23684
rect 9824 23712 9830 23724
rect 10229 23715 10287 23721
rect 10229 23712 10241 23715
rect 9824 23684 10241 23712
rect 9824 23672 9830 23684
rect 10229 23681 10241 23684
rect 10275 23681 10287 23715
rect 13630 23712 13636 23724
rect 13591 23684 13636 23712
rect 10229 23675 10287 23681
rect 13630 23672 13636 23684
rect 13688 23672 13694 23724
rect 13909 23715 13967 23721
rect 13909 23681 13921 23715
rect 13955 23712 13967 23715
rect 14660 23712 14688 23752
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 24394 23712 24400 23724
rect 13955 23684 14688 23712
rect 14752 23684 24400 23712
rect 13955 23681 13967 23684
rect 13909 23675 13967 23681
rect 6917 23647 6975 23653
rect 6917 23644 6929 23647
rect 5828 23616 6929 23644
rect 5721 23607 5779 23613
rect 6917 23613 6929 23616
rect 6963 23644 6975 23647
rect 7098 23644 7104 23656
rect 6963 23616 7104 23644
rect 6963 23613 6975 23616
rect 6917 23607 6975 23613
rect 5736 23576 5764 23607
rect 7098 23604 7104 23616
rect 7156 23604 7162 23656
rect 7285 23647 7343 23653
rect 7285 23613 7297 23647
rect 7331 23644 7343 23647
rect 7650 23644 7656 23656
rect 7331 23616 7656 23644
rect 7331 23613 7343 23616
rect 7285 23607 7343 23613
rect 7650 23604 7656 23616
rect 7708 23604 7714 23656
rect 8754 23644 8760 23656
rect 8715 23616 8760 23644
rect 8754 23604 8760 23616
rect 8812 23604 8818 23656
rect 12529 23647 12587 23653
rect 12529 23613 12541 23647
rect 12575 23644 12587 23647
rect 12621 23647 12679 23653
rect 12621 23644 12633 23647
rect 12575 23616 12633 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 12621 23613 12633 23616
rect 12667 23644 12679 23647
rect 12667 23616 13308 23644
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 7190 23576 7196 23588
rect 5736 23548 7196 23576
rect 7190 23536 7196 23548
rect 7248 23536 7254 23588
rect 13280 23520 13308 23616
rect 5445 23511 5503 23517
rect 5445 23477 5457 23511
rect 5491 23508 5503 23511
rect 6822 23508 6828 23520
rect 5491 23480 6828 23508
rect 5491 23477 5503 23480
rect 5445 23471 5503 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 12710 23508 12716 23520
rect 12671 23480 12716 23508
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 13262 23468 13268 23520
rect 13320 23508 13326 23520
rect 14752 23508 14780 23684
rect 24394 23672 24400 23684
rect 24452 23672 24458 23724
rect 25240 23712 25268 23808
rect 25409 23715 25467 23721
rect 25409 23712 25421 23715
rect 25240 23684 25421 23712
rect 25409 23681 25421 23684
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 29362 23672 29368 23724
rect 29420 23712 29426 23724
rect 30561 23715 30619 23721
rect 30561 23712 30573 23715
rect 29420 23684 30573 23712
rect 29420 23672 29426 23684
rect 30561 23681 30573 23684
rect 30607 23712 30619 23715
rect 30742 23712 30748 23724
rect 30607 23684 30748 23712
rect 30607 23681 30619 23684
rect 30561 23675 30619 23681
rect 30742 23672 30748 23684
rect 30800 23672 30806 23724
rect 30837 23715 30895 23721
rect 30837 23681 30849 23715
rect 30883 23712 30895 23715
rect 34238 23712 34244 23724
rect 30883 23684 34244 23712
rect 30883 23681 30895 23684
rect 30837 23675 30895 23681
rect 34238 23672 34244 23684
rect 34296 23672 34302 23724
rect 35912 23712 35940 23808
rect 45370 23740 45376 23792
rect 45428 23780 45434 23792
rect 47765 23783 47823 23789
rect 47765 23780 47777 23783
rect 45428 23752 47777 23780
rect 45428 23740 45434 23752
rect 47765 23749 47777 23752
rect 47811 23780 47823 23783
rect 47811 23752 48176 23780
rect 47811 23749 47823 23752
rect 47765 23743 47823 23749
rect 36081 23715 36139 23721
rect 36081 23712 36093 23715
rect 35912 23684 36093 23712
rect 36081 23681 36093 23684
rect 36127 23681 36139 23715
rect 36081 23675 36139 23681
rect 38841 23715 38899 23721
rect 38841 23681 38853 23715
rect 38887 23712 38899 23715
rect 39942 23712 39948 23724
rect 38887 23684 39948 23712
rect 38887 23681 38899 23684
rect 38841 23675 38899 23681
rect 39942 23672 39948 23684
rect 40000 23712 40006 23724
rect 48148 23721 48176 23752
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 40000 23684 41521 23712
rect 40000 23672 40006 23684
rect 41509 23681 41521 23684
rect 41555 23712 41567 23715
rect 43809 23715 43867 23721
rect 43809 23712 43821 23715
rect 41555 23684 43821 23712
rect 41555 23681 41567 23684
rect 41509 23675 41567 23681
rect 43809 23681 43821 23684
rect 43855 23712 43867 23715
rect 48133 23715 48191 23721
rect 43855 23684 46244 23712
rect 43855 23681 43867 23684
rect 43809 23675 43867 23681
rect 17770 23604 17776 23656
rect 17828 23644 17834 23656
rect 17865 23647 17923 23653
rect 17865 23644 17877 23647
rect 17828 23616 17877 23644
rect 17828 23604 17834 23616
rect 17865 23613 17877 23616
rect 17911 23644 17923 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17911 23616 18061 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 18325 23647 18383 23653
rect 18095 23616 18184 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 13320 23480 14780 23508
rect 18156 23508 18184 23616
rect 18325 23613 18337 23647
rect 18371 23644 18383 23647
rect 18598 23644 18604 23656
rect 18371 23616 18604 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 21913 23647 21971 23653
rect 21913 23613 21925 23647
rect 21959 23644 21971 23647
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21959 23616 22017 23644
rect 21959 23613 21971 23616
rect 21913 23607 21971 23613
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22281 23647 22339 23653
rect 22281 23613 22293 23647
rect 22327 23613 22339 23647
rect 22281 23607 22339 23613
rect 25685 23647 25743 23653
rect 25685 23613 25697 23647
rect 25731 23644 25743 23647
rect 29546 23644 29552 23656
rect 25731 23616 29552 23644
rect 25731 23613 25743 23616
rect 25685 23607 25743 23613
rect 21542 23576 21548 23588
rect 18984 23548 21548 23576
rect 18984 23508 19012 23548
rect 21542 23536 21548 23548
rect 21600 23536 21606 23588
rect 18156 23480 19012 23508
rect 13320 23468 13326 23480
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 21726 23508 21732 23520
rect 19576 23480 21732 23508
rect 19576 23468 19582 23480
rect 21726 23468 21732 23480
rect 21784 23468 21790 23520
rect 22020 23508 22048 23607
rect 22186 23576 22192 23588
rect 22147 23548 22192 23576
rect 22186 23536 22192 23548
rect 22244 23536 22250 23588
rect 22094 23508 22100 23520
rect 22020 23480 22100 23508
rect 22094 23468 22100 23480
rect 22152 23468 22158 23520
rect 22296 23508 22324 23607
rect 29546 23604 29552 23616
rect 29604 23604 29610 23656
rect 30760 23644 30788 23672
rect 46216 23656 46244 23684
rect 48133 23681 48145 23715
rect 48179 23712 48191 23715
rect 48590 23712 48596 23724
rect 48179 23684 48596 23712
rect 48179 23681 48191 23684
rect 48133 23675 48191 23681
rect 48590 23672 48596 23684
rect 48648 23672 48654 23724
rect 32306 23644 32312 23656
rect 30760 23616 32312 23644
rect 32306 23604 32312 23616
rect 32364 23604 32370 23656
rect 33318 23644 33324 23656
rect 33279 23616 33324 23644
rect 33318 23604 33324 23616
rect 33376 23604 33382 23656
rect 33505 23647 33563 23653
rect 33505 23613 33517 23647
rect 33551 23644 33563 23647
rect 33778 23644 33784 23656
rect 33551 23616 33784 23644
rect 33551 23613 33563 23616
rect 33505 23607 33563 23613
rect 33778 23604 33784 23616
rect 33836 23604 33842 23656
rect 34974 23644 34980 23656
rect 34935 23616 34980 23644
rect 34974 23604 34980 23616
rect 35032 23604 35038 23656
rect 36354 23644 36360 23656
rect 36315 23616 36360 23644
rect 36354 23604 36360 23616
rect 36412 23604 36418 23656
rect 39117 23647 39175 23653
rect 39117 23613 39129 23647
rect 39163 23644 39175 23647
rect 40034 23644 40040 23656
rect 39163 23616 40040 23644
rect 39163 23613 39175 23616
rect 39117 23607 39175 23613
rect 40034 23604 40040 23616
rect 40092 23604 40098 23656
rect 40126 23604 40132 23656
rect 40184 23644 40190 23656
rect 40497 23647 40555 23653
rect 40497 23644 40509 23647
rect 40184 23616 40509 23644
rect 40184 23604 40190 23616
rect 40497 23613 40509 23616
rect 40543 23613 40555 23647
rect 41782 23644 41788 23656
rect 41743 23616 41788 23644
rect 40497 23607 40555 23613
rect 41782 23604 41788 23616
rect 41840 23604 41846 23656
rect 44085 23647 44143 23653
rect 44085 23613 44097 23647
rect 44131 23644 44143 23647
rect 44174 23644 44180 23656
rect 44131 23616 44180 23644
rect 44131 23613 44143 23616
rect 44085 23607 44143 23613
rect 44174 23604 44180 23616
rect 44232 23604 44238 23656
rect 46198 23644 46204 23656
rect 46159 23616 46204 23644
rect 46198 23604 46204 23616
rect 46256 23604 46262 23656
rect 46382 23644 46388 23656
rect 46343 23616 46388 23644
rect 46382 23604 46388 23616
rect 46440 23604 46446 23656
rect 48409 23647 48467 23653
rect 48409 23644 48421 23647
rect 47964 23616 48421 23644
rect 33410 23576 33416 23588
rect 33371 23548 33416 23576
rect 33410 23536 33416 23548
rect 33468 23536 33474 23588
rect 34992 23576 35020 23604
rect 33520 23548 35020 23576
rect 22925 23511 22983 23517
rect 22925 23508 22937 23511
rect 22296 23480 22937 23508
rect 22925 23477 22937 23480
rect 22971 23508 22983 23511
rect 28626 23508 28632 23520
rect 22971 23480 28632 23508
rect 22971 23477 22983 23480
rect 22925 23471 22983 23477
rect 28626 23468 28632 23480
rect 28684 23468 28690 23520
rect 31570 23468 31576 23520
rect 31628 23508 31634 23520
rect 33520 23508 33548 23548
rect 37366 23536 37372 23588
rect 37424 23576 37430 23588
rect 39025 23579 39083 23585
rect 39025 23576 39037 23579
rect 37424 23548 39037 23576
rect 37424 23536 37430 23548
rect 39025 23545 39037 23548
rect 39071 23576 39083 23579
rect 41693 23579 41751 23585
rect 41693 23576 41705 23579
rect 39071 23548 41705 23576
rect 39071 23545 39083 23548
rect 39025 23539 39083 23545
rect 41693 23545 41705 23548
rect 41739 23576 41751 23579
rect 43993 23579 44051 23585
rect 43993 23576 44005 23579
rect 41739 23548 44005 23576
rect 41739 23545 41751 23548
rect 41693 23539 41751 23545
rect 43993 23545 44005 23548
rect 44039 23576 44051 23579
rect 46293 23579 46351 23585
rect 46293 23576 46305 23579
rect 44039 23548 46305 23576
rect 44039 23545 44051 23548
rect 43993 23539 44051 23545
rect 46293 23545 46305 23548
rect 46339 23545 46351 23579
rect 46293 23539 46351 23545
rect 31628 23480 33548 23508
rect 31628 23468 31634 23480
rect 34514 23468 34520 23520
rect 34572 23508 34578 23520
rect 35158 23508 35164 23520
rect 34572 23480 35164 23508
rect 34572 23468 34578 23480
rect 35158 23468 35164 23480
rect 35216 23468 35222 23520
rect 38838 23468 38844 23520
rect 38896 23508 38902 23520
rect 40589 23511 40647 23517
rect 40589 23508 40601 23511
rect 38896 23480 40601 23508
rect 38896 23468 38902 23480
rect 40589 23477 40601 23480
rect 40635 23477 40647 23511
rect 40589 23471 40647 23477
rect 41046 23468 41052 23520
rect 41104 23508 41110 23520
rect 47964 23517 47992 23616
rect 48409 23613 48421 23616
rect 48455 23613 48467 23647
rect 52089 23647 52147 23653
rect 52089 23644 52101 23647
rect 48409 23607 48467 23613
rect 51920 23616 52101 23644
rect 47949 23511 48007 23517
rect 47949 23508 47961 23511
rect 41104 23480 47961 23508
rect 41104 23468 41110 23480
rect 47949 23477 47961 23480
rect 47995 23477 48007 23511
rect 47949 23471 48007 23477
rect 51810 23468 51816 23520
rect 51868 23508 51874 23520
rect 51920 23517 51948 23616
rect 52089 23613 52101 23616
rect 52135 23613 52147 23647
rect 52362 23644 52368 23656
rect 52323 23616 52368 23644
rect 52089 23607 52147 23613
rect 52362 23604 52368 23616
rect 52420 23604 52426 23656
rect 51905 23511 51963 23517
rect 51905 23508 51917 23511
rect 51868 23480 51917 23508
rect 51868 23468 51874 23480
rect 51905 23477 51917 23480
rect 51951 23477 51963 23511
rect 53466 23508 53472 23520
rect 53427 23480 53472 23508
rect 51905 23471 51963 23477
rect 53466 23468 53472 23480
rect 53524 23468 53530 23520
rect 1104 23418 54832 23440
rect 1104 23366 18912 23418
rect 18964 23366 18976 23418
rect 19028 23366 19040 23418
rect 19092 23366 19104 23418
rect 19156 23366 36843 23418
rect 36895 23366 36907 23418
rect 36959 23366 36971 23418
rect 37023 23366 37035 23418
rect 37087 23366 54832 23418
rect 1104 23344 54832 23366
rect 3878 23264 3884 23316
rect 3936 23304 3942 23316
rect 7006 23304 7012 23316
rect 3936 23276 7012 23304
rect 3936 23264 3942 23276
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 13262 23304 13268 23316
rect 13223 23276 13268 23304
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 19518 23304 19524 23316
rect 18524 23276 19524 23304
rect 5902 23236 5908 23248
rect 5863 23208 5908 23236
rect 5902 23196 5908 23208
rect 5960 23196 5966 23248
rect 8754 23236 8760 23248
rect 8715 23208 8760 23236
rect 8754 23196 8760 23208
rect 8812 23196 8818 23248
rect 11701 23239 11759 23245
rect 11701 23205 11713 23239
rect 11747 23236 11759 23239
rect 12618 23236 12624 23248
rect 11747 23208 12624 23236
rect 11747 23205 11759 23208
rect 11701 23199 11759 23205
rect 12618 23196 12624 23208
rect 12676 23196 12682 23248
rect 934 23128 940 23180
rect 992 23168 998 23180
rect 6914 23168 6920 23180
rect 992 23140 6920 23168
rect 992 23128 998 23140
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 7098 23128 7104 23180
rect 7156 23168 7162 23180
rect 8018 23168 8024 23180
rect 7156 23140 8024 23168
rect 7156 23128 7162 23140
rect 8018 23128 8024 23140
rect 8076 23128 8082 23180
rect 8573 23171 8631 23177
rect 8573 23137 8585 23171
rect 8619 23168 8631 23171
rect 11054 23168 11060 23180
rect 8619 23140 8800 23168
rect 11015 23140 11060 23168
rect 8619 23137 8631 23140
rect 8573 23131 8631 23137
rect 8772 23112 8800 23140
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 11422 23168 11428 23180
rect 11383 23140 11428 23168
rect 11422 23128 11428 23140
rect 11480 23128 11486 23180
rect 13280 23168 13308 23264
rect 18325 23239 18383 23245
rect 18325 23236 18337 23239
rect 13556 23208 18337 23236
rect 13357 23171 13415 23177
rect 13357 23168 13369 23171
rect 13280 23140 13369 23168
rect 13357 23137 13369 23140
rect 13403 23137 13415 23171
rect 13357 23131 13415 23137
rect 4062 23100 4068 23112
rect 4023 23072 4068 23100
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 4338 23100 4344 23112
rect 4299 23072 4344 23100
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 4522 23060 4528 23112
rect 4580 23100 4586 23112
rect 5537 23103 5595 23109
rect 5537 23100 5549 23103
rect 4580 23072 5549 23100
rect 4580 23060 4586 23072
rect 5537 23069 5549 23072
rect 5583 23069 5595 23103
rect 5537 23063 5595 23069
rect 8754 23060 8760 23112
rect 8812 23060 8818 23112
rect 11514 22992 11520 23044
rect 11572 23032 11578 23044
rect 13556 23041 13584 23208
rect 18325 23205 18337 23208
rect 18371 23236 18383 23239
rect 18524 23236 18552 23276
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 19702 23264 19708 23316
rect 19760 23304 19766 23316
rect 21082 23304 21088 23316
rect 19760 23276 21088 23304
rect 19760 23264 19766 23276
rect 21082 23264 21088 23276
rect 21140 23264 21146 23316
rect 21634 23264 21640 23316
rect 21692 23304 21698 23316
rect 21913 23307 21971 23313
rect 21913 23304 21925 23307
rect 21692 23276 21925 23304
rect 21692 23264 21698 23276
rect 21913 23273 21925 23276
rect 21959 23304 21971 23307
rect 32490 23304 32496 23316
rect 21959 23276 32496 23304
rect 21959 23273 21971 23276
rect 21913 23267 21971 23273
rect 32490 23264 32496 23276
rect 32548 23264 32554 23316
rect 32582 23264 32588 23316
rect 32640 23304 32646 23316
rect 33226 23304 33232 23316
rect 32640 23276 33232 23304
rect 32640 23264 32646 23276
rect 33226 23264 33232 23276
rect 33284 23264 33290 23316
rect 37001 23307 37059 23313
rect 37001 23273 37013 23307
rect 37047 23304 37059 23307
rect 41598 23304 41604 23316
rect 37047 23276 41604 23304
rect 37047 23273 37059 23276
rect 37001 23267 37059 23273
rect 18371 23208 18552 23236
rect 18371 23205 18383 23208
rect 18325 23199 18383 23205
rect 18524 23180 18552 23208
rect 19426 23196 19432 23248
rect 19484 23236 19490 23248
rect 21729 23239 21787 23245
rect 21729 23236 21741 23239
rect 19484 23208 21741 23236
rect 19484 23196 19490 23208
rect 21729 23205 21741 23208
rect 21775 23205 21787 23239
rect 23474 23236 23480 23248
rect 21729 23199 21787 23205
rect 21836 23208 23480 23236
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 15028 23140 15301 23168
rect 13541 23035 13599 23041
rect 13541 23032 13553 23035
rect 11572 23004 13553 23032
rect 11572 22992 11578 23004
rect 13541 23001 13553 23004
rect 13587 23001 13599 23035
rect 13541 22995 13599 23001
rect 2406 22924 2412 22976
rect 2464 22964 2470 22976
rect 5718 22964 5724 22976
rect 2464 22936 5724 22964
rect 2464 22924 2470 22936
rect 5718 22924 5724 22936
rect 5776 22924 5782 22976
rect 14826 22924 14832 22976
rect 14884 22964 14890 22976
rect 15028 22973 15056 23140
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15838 23168 15844 23180
rect 15799 23140 15844 23168
rect 15289 23131 15347 23137
rect 15838 23128 15844 23140
rect 15896 23128 15902 23180
rect 18506 23168 18512 23180
rect 18419 23140 18512 23168
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 18693 23171 18751 23177
rect 18693 23137 18705 23171
rect 18739 23137 18751 23171
rect 18693 23131 18751 23137
rect 18785 23171 18843 23177
rect 18785 23137 18797 23171
rect 18831 23168 18843 23171
rect 21082 23168 21088 23180
rect 18831 23140 21088 23168
rect 18831 23137 18843 23140
rect 18785 23131 18843 23137
rect 16114 23100 16120 23112
rect 16075 23072 16120 23100
rect 16114 23060 16120 23072
rect 16172 23060 16178 23112
rect 18708 23100 18736 23131
rect 21082 23128 21088 23140
rect 21140 23128 21146 23180
rect 21177 23171 21235 23177
rect 21177 23137 21189 23171
rect 21223 23137 21235 23171
rect 21177 23131 21235 23137
rect 19334 23100 19340 23112
rect 18708 23072 19340 23100
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 20898 23060 20904 23112
rect 20956 23100 20962 23112
rect 21192 23100 21220 23131
rect 21266 23128 21272 23180
rect 21324 23168 21330 23180
rect 21324 23140 21369 23168
rect 21324 23128 21330 23140
rect 21836 23100 21864 23208
rect 23474 23196 23480 23208
rect 23532 23196 23538 23248
rect 23658 23196 23664 23248
rect 23716 23236 23722 23248
rect 23845 23239 23903 23245
rect 23845 23236 23857 23239
rect 23716 23208 23857 23236
rect 23716 23196 23722 23208
rect 23845 23205 23857 23208
rect 23891 23205 23903 23239
rect 23845 23199 23903 23205
rect 23934 23196 23940 23248
rect 23992 23236 23998 23248
rect 25314 23236 25320 23248
rect 23992 23208 25320 23236
rect 23992 23196 23998 23208
rect 25314 23196 25320 23208
rect 25372 23196 25378 23248
rect 27614 23236 27620 23248
rect 26528 23208 27620 23236
rect 23290 23168 23296 23180
rect 23251 23140 23296 23168
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 23385 23171 23443 23177
rect 23385 23137 23397 23171
rect 23431 23137 23443 23171
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 23385 23131 23443 23137
rect 23860 23140 24593 23168
rect 20956 23072 21220 23100
rect 21560 23072 21864 23100
rect 20956 23060 20962 23072
rect 15378 23032 15384 23044
rect 15339 23004 15384 23032
rect 15378 22992 15384 23004
rect 15436 22992 15442 23044
rect 16666 22992 16672 23044
rect 16724 23032 16730 23044
rect 21560 23032 21588 23072
rect 16724 23004 21588 23032
rect 16724 22992 16730 23004
rect 21726 22992 21732 23044
rect 21784 23032 21790 23044
rect 22094 23032 22100 23044
rect 21784 23004 22100 23032
rect 21784 22992 21790 23004
rect 22094 22992 22100 23004
rect 22152 23032 22158 23044
rect 22925 23035 22983 23041
rect 22925 23032 22937 23035
rect 22152 23004 22937 23032
rect 22152 22992 22158 23004
rect 22925 23001 22937 23004
rect 22971 23032 22983 23035
rect 23109 23035 23167 23041
rect 23109 23032 23121 23035
rect 22971 23004 23121 23032
rect 22971 23001 22983 23004
rect 22925 22995 22983 23001
rect 23109 23001 23121 23004
rect 23155 23001 23167 23035
rect 23400 23032 23428 23131
rect 23860 23112 23888 23140
rect 24581 23137 24593 23140
rect 24627 23168 24639 23171
rect 24673 23171 24731 23177
rect 24673 23168 24685 23171
rect 24627 23140 24685 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24673 23137 24685 23140
rect 24719 23137 24731 23171
rect 24673 23131 24731 23137
rect 25590 23128 25596 23180
rect 25648 23168 25654 23180
rect 26528 23177 26556 23208
rect 27614 23196 27620 23208
rect 27672 23196 27678 23248
rect 30653 23239 30711 23245
rect 30653 23236 30665 23239
rect 28644 23208 30665 23236
rect 26513 23171 26571 23177
rect 26513 23168 26525 23171
rect 25648 23140 26525 23168
rect 25648 23128 25654 23140
rect 26513 23137 26525 23140
rect 26559 23137 26571 23171
rect 27709 23171 27767 23177
rect 27709 23168 27721 23171
rect 26513 23131 26571 23137
rect 27632 23140 27721 23168
rect 27632 23112 27660 23140
rect 27709 23137 27721 23140
rect 27755 23137 27767 23171
rect 27709 23131 27767 23137
rect 27798 23128 27804 23180
rect 27856 23168 27862 23180
rect 27985 23171 28043 23177
rect 27985 23168 27997 23171
rect 27856 23140 27997 23168
rect 27856 23128 27862 23140
rect 27985 23137 27997 23140
rect 28031 23137 28043 23171
rect 27985 23131 28043 23137
rect 28074 23128 28080 23180
rect 28132 23168 28138 23180
rect 28644 23168 28672 23208
rect 30653 23205 30665 23208
rect 30699 23236 30711 23239
rect 36265 23239 36323 23245
rect 30699 23208 30880 23236
rect 30699 23205 30711 23208
rect 30653 23199 30711 23205
rect 30742 23168 30748 23180
rect 28132 23140 28672 23168
rect 30703 23140 30748 23168
rect 28132 23128 28138 23140
rect 30742 23128 30748 23140
rect 30800 23128 30806 23180
rect 30852 23168 30880 23208
rect 36265 23205 36277 23239
rect 36311 23236 36323 23239
rect 37366 23236 37372 23248
rect 36311 23208 37372 23236
rect 36311 23205 36323 23208
rect 36265 23199 36323 23205
rect 37366 23196 37372 23208
rect 37424 23196 37430 23248
rect 32122 23168 32128 23180
rect 30852 23140 32128 23168
rect 32122 23128 32128 23140
rect 32180 23128 32186 23180
rect 33410 23128 33416 23180
rect 33468 23168 33474 23180
rect 33965 23171 34023 23177
rect 33965 23168 33977 23171
rect 33468 23140 33977 23168
rect 33468 23128 33474 23140
rect 33965 23137 33977 23140
rect 34011 23137 34023 23171
rect 33965 23131 34023 23137
rect 34057 23171 34115 23177
rect 34057 23137 34069 23171
rect 34103 23168 34115 23171
rect 34103 23140 34744 23168
rect 34103 23137 34115 23140
rect 34057 23131 34115 23137
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 27614 23060 27620 23112
rect 27672 23060 27678 23112
rect 29089 23103 29147 23109
rect 29089 23100 29101 23103
rect 27724 23072 29101 23100
rect 27724 23032 27752 23072
rect 29089 23069 29101 23072
rect 29135 23100 29147 23103
rect 29270 23100 29276 23112
rect 29135 23072 29276 23100
rect 29135 23069 29147 23072
rect 29089 23063 29147 23069
rect 29270 23060 29276 23072
rect 29328 23060 29334 23112
rect 30469 23103 30527 23109
rect 30469 23069 30481 23103
rect 30515 23100 30527 23103
rect 31570 23100 31576 23112
rect 30515 23072 31576 23100
rect 30515 23069 30527 23072
rect 30469 23063 30527 23069
rect 31570 23060 31576 23072
rect 31628 23060 31634 23112
rect 23400 23004 27752 23032
rect 23109 22995 23167 23001
rect 33318 22992 33324 23044
rect 33376 23032 33382 23044
rect 33781 23035 33839 23041
rect 33781 23032 33793 23035
rect 33376 23004 33793 23032
rect 33376 22992 33382 23004
rect 33781 23001 33793 23004
rect 33827 23032 33839 23035
rect 34514 23032 34520 23044
rect 33827 23004 34520 23032
rect 33827 23001 33839 23004
rect 33781 22995 33839 23001
rect 34514 22992 34520 23004
rect 34572 22992 34578 23044
rect 34716 23041 34744 23140
rect 35158 23128 35164 23180
rect 35216 23168 35222 23180
rect 36081 23171 36139 23177
rect 36081 23168 36093 23171
rect 35216 23140 36093 23168
rect 35216 23128 35222 23140
rect 36081 23137 36093 23140
rect 36127 23137 36139 23171
rect 36081 23131 36139 23137
rect 36357 23171 36415 23177
rect 36357 23137 36369 23171
rect 36403 23168 36415 23171
rect 37476 23168 37504 23276
rect 41598 23264 41604 23276
rect 41656 23264 41662 23316
rect 41874 23264 41880 23316
rect 41932 23304 41938 23316
rect 45554 23304 45560 23316
rect 41932 23276 45560 23304
rect 41932 23264 41938 23276
rect 45554 23264 45560 23276
rect 45612 23264 45618 23316
rect 46106 23264 46112 23316
rect 46164 23304 46170 23316
rect 53466 23304 53472 23316
rect 46164 23276 53472 23304
rect 46164 23264 46170 23276
rect 53466 23264 53472 23276
rect 53524 23264 53530 23316
rect 37642 23196 37648 23248
rect 37700 23236 37706 23248
rect 44542 23236 44548 23248
rect 37700 23208 38700 23236
rect 37700 23196 37706 23208
rect 36403 23140 37504 23168
rect 38672 23168 38700 23208
rect 39500 23208 43024 23236
rect 44503 23208 44548 23236
rect 39500 23168 39528 23208
rect 38672 23140 39528 23168
rect 36403 23137 36415 23140
rect 36357 23131 36415 23137
rect 39758 23128 39764 23180
rect 39816 23168 39822 23180
rect 41049 23171 41107 23177
rect 41049 23168 41061 23171
rect 39816 23140 41061 23168
rect 39816 23128 39822 23140
rect 41049 23137 41061 23140
rect 41095 23137 41107 23171
rect 41049 23131 41107 23137
rect 41138 23128 41144 23180
rect 41196 23168 41202 23180
rect 41233 23171 41291 23177
rect 41233 23168 41245 23171
rect 41196 23140 41245 23168
rect 41196 23128 41202 23140
rect 41233 23137 41245 23140
rect 41279 23137 41291 23171
rect 41233 23131 41291 23137
rect 41785 23171 41843 23177
rect 41785 23137 41797 23171
rect 41831 23168 41843 23171
rect 41874 23168 41880 23180
rect 41831 23140 41880 23168
rect 41831 23137 41843 23140
rect 41785 23131 41843 23137
rect 41874 23128 41880 23140
rect 41932 23128 41938 23180
rect 41969 23171 42027 23177
rect 41969 23137 41981 23171
rect 42015 23168 42027 23171
rect 42334 23168 42340 23180
rect 42015 23140 42340 23168
rect 42015 23137 42027 23140
rect 41969 23131 42027 23137
rect 42334 23128 42340 23140
rect 42392 23128 42398 23180
rect 42996 23168 43024 23208
rect 44542 23196 44548 23208
rect 44600 23196 44606 23248
rect 46293 23239 46351 23245
rect 46293 23205 46305 23239
rect 46339 23236 46351 23239
rect 46382 23236 46388 23248
rect 46339 23208 46388 23236
rect 46339 23205 46351 23208
rect 46293 23199 46351 23205
rect 46382 23196 46388 23208
rect 46440 23196 46446 23248
rect 48041 23239 48099 23245
rect 48041 23205 48053 23239
rect 48087 23236 48099 23239
rect 48498 23236 48504 23248
rect 48087 23208 48504 23236
rect 48087 23205 48099 23208
rect 48041 23199 48099 23205
rect 48498 23196 48504 23208
rect 48556 23196 48562 23248
rect 52362 23236 52368 23248
rect 52323 23208 52368 23236
rect 52362 23196 52368 23208
rect 52420 23196 52426 23248
rect 46658 23168 46664 23180
rect 42996 23140 46664 23168
rect 46658 23128 46664 23140
rect 46716 23128 46722 23180
rect 47394 23128 47400 23180
rect 47452 23168 47458 23180
rect 47489 23171 47547 23177
rect 47489 23168 47501 23171
rect 47452 23140 47501 23168
rect 47452 23128 47458 23140
rect 47489 23137 47501 23140
rect 47535 23137 47547 23171
rect 47489 23131 47547 23137
rect 47581 23171 47639 23177
rect 47581 23137 47593 23171
rect 47627 23168 47639 23171
rect 47854 23168 47860 23180
rect 47627 23140 47860 23168
rect 47627 23137 47639 23140
rect 47581 23131 47639 23137
rect 35434 23060 35440 23112
rect 35492 23100 35498 23112
rect 38102 23100 38108 23112
rect 35492 23072 38108 23100
rect 35492 23060 35498 23072
rect 38102 23060 38108 23072
rect 38160 23060 38166 23112
rect 38565 23103 38623 23109
rect 38565 23100 38577 23103
rect 38396 23072 38577 23100
rect 34701 23035 34759 23041
rect 34701 23001 34713 23035
rect 34747 23032 34759 23035
rect 37274 23032 37280 23044
rect 34747 23004 37280 23032
rect 34747 23001 34759 23004
rect 34701 22995 34759 23001
rect 37274 22992 37280 23004
rect 37332 22992 37338 23044
rect 15013 22967 15071 22973
rect 15013 22964 15025 22967
rect 14884 22936 15025 22964
rect 14884 22924 14890 22936
rect 15013 22933 15025 22936
rect 15059 22933 15071 22967
rect 15013 22927 15071 22933
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 18969 22967 19027 22973
rect 18969 22964 18981 22967
rect 18656 22936 18981 22964
rect 18656 22924 18662 22936
rect 18969 22933 18981 22936
rect 19015 22933 19027 22967
rect 18969 22927 19027 22933
rect 20714 22924 20720 22976
rect 20772 22964 20778 22976
rect 20993 22967 21051 22973
rect 20993 22964 21005 22967
rect 20772 22936 21005 22964
rect 20772 22924 20778 22936
rect 20993 22933 21005 22936
rect 21039 22964 21051 22967
rect 21634 22964 21640 22976
rect 21039 22936 21640 22964
rect 21039 22933 21051 22936
rect 20993 22927 21051 22933
rect 21634 22924 21640 22936
rect 21692 22924 21698 22976
rect 21910 22924 21916 22976
rect 21968 22964 21974 22976
rect 22005 22967 22063 22973
rect 22005 22964 22017 22967
rect 21968 22936 22017 22964
rect 21968 22924 21974 22936
rect 22005 22933 22017 22936
rect 22051 22933 22063 22967
rect 22005 22927 22063 22933
rect 22554 22924 22560 22976
rect 22612 22964 22618 22976
rect 23934 22964 23940 22976
rect 22612 22936 23940 22964
rect 22612 22924 22618 22936
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 24857 22967 24915 22973
rect 24857 22933 24869 22967
rect 24903 22964 24915 22967
rect 25590 22964 25596 22976
rect 24903 22936 25596 22964
rect 24903 22933 24915 22936
rect 24857 22927 24915 22933
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 26694 22964 26700 22976
rect 26607 22936 26700 22964
rect 26694 22924 26700 22936
rect 26752 22964 26758 22976
rect 28166 22964 28172 22976
rect 26752 22936 28172 22964
rect 26752 22924 26758 22936
rect 28166 22924 28172 22936
rect 28224 22924 28230 22976
rect 29362 22924 29368 22976
rect 29420 22964 29426 22976
rect 29457 22967 29515 22973
rect 29457 22964 29469 22967
rect 29420 22936 29469 22964
rect 29420 22924 29426 22936
rect 29457 22933 29469 22936
rect 29503 22933 29515 22967
rect 29457 22927 29515 22933
rect 29546 22924 29552 22976
rect 29604 22964 29610 22976
rect 30929 22967 30987 22973
rect 30929 22964 30941 22967
rect 29604 22936 30941 22964
rect 29604 22924 29610 22936
rect 30929 22933 30941 22936
rect 30975 22933 30987 22967
rect 30929 22927 30987 22933
rect 32214 22924 32220 22976
rect 32272 22964 32278 22976
rect 32309 22967 32367 22973
rect 32309 22964 32321 22967
rect 32272 22936 32321 22964
rect 32272 22924 32278 22936
rect 32309 22933 32321 22936
rect 32355 22933 32367 22967
rect 34238 22964 34244 22976
rect 34199 22936 34244 22964
rect 32309 22927 32367 22933
rect 34238 22924 34244 22936
rect 34296 22924 34302 22976
rect 36354 22924 36360 22976
rect 36412 22964 36418 22976
rect 36541 22967 36599 22973
rect 36541 22964 36553 22967
rect 36412 22936 36553 22964
rect 36412 22924 36418 22936
rect 36541 22933 36553 22936
rect 36587 22933 36599 22967
rect 36541 22927 36599 22933
rect 38194 22924 38200 22976
rect 38252 22964 38258 22976
rect 38396 22973 38424 23072
rect 38565 23069 38577 23072
rect 38611 23069 38623 23103
rect 38565 23063 38623 23069
rect 38746 23060 38752 23112
rect 38804 23100 38810 23112
rect 38841 23103 38899 23109
rect 38841 23100 38853 23103
rect 38804 23072 38853 23100
rect 38804 23060 38810 23072
rect 38841 23069 38853 23072
rect 38887 23069 38899 23103
rect 38841 23063 38899 23069
rect 44542 23060 44548 23112
rect 44600 23100 44606 23112
rect 44637 23103 44695 23109
rect 44637 23100 44649 23103
rect 44600 23072 44649 23100
rect 44600 23060 44606 23072
rect 44637 23069 44649 23072
rect 44683 23069 44695 23103
rect 44910 23100 44916 23112
rect 44871 23072 44916 23100
rect 44637 23063 44695 23069
rect 44910 23060 44916 23072
rect 44968 23060 44974 23112
rect 46198 23060 46204 23112
rect 46256 23100 46262 23112
rect 47305 23103 47363 23109
rect 47305 23100 47317 23103
rect 46256 23072 47317 23100
rect 46256 23060 46262 23072
rect 47305 23069 47317 23072
rect 47351 23069 47363 23103
rect 47504 23100 47532 23131
rect 47854 23128 47860 23140
rect 47912 23128 47918 23180
rect 51261 23171 51319 23177
rect 51261 23168 51273 23171
rect 47964 23140 51273 23168
rect 47964 23100 47992 23140
rect 51261 23137 51273 23140
rect 51307 23168 51319 23171
rect 51718 23168 51724 23180
rect 51307 23140 51724 23168
rect 51307 23137 51319 23140
rect 51261 23131 51319 23137
rect 51718 23128 51724 23140
rect 51776 23168 51782 23180
rect 51813 23171 51871 23177
rect 51813 23168 51825 23171
rect 51776 23140 51825 23168
rect 51776 23128 51782 23140
rect 51813 23137 51825 23140
rect 51859 23137 51871 23171
rect 51813 23131 51871 23137
rect 51905 23171 51963 23177
rect 51905 23137 51917 23171
rect 51951 23168 51963 23171
rect 51994 23168 52000 23180
rect 51951 23140 52000 23168
rect 51951 23137 51963 23140
rect 51905 23131 51963 23137
rect 51994 23128 52000 23140
rect 52052 23128 52058 23180
rect 47504 23072 47992 23100
rect 47305 23063 47363 23069
rect 40586 22992 40592 23044
rect 40644 23032 40650 23044
rect 40644 23004 44680 23032
rect 40644 22992 40650 23004
rect 38381 22967 38439 22973
rect 38381 22964 38393 22967
rect 38252 22936 38393 22964
rect 38252 22924 38258 22936
rect 38381 22933 38393 22936
rect 38427 22933 38439 22967
rect 40126 22964 40132 22976
rect 40087 22936 40132 22964
rect 38381 22927 38439 22933
rect 40126 22924 40132 22936
rect 40184 22924 40190 22976
rect 42245 22967 42303 22973
rect 42245 22933 42257 22967
rect 42291 22964 42303 22967
rect 44358 22964 44364 22976
rect 42291 22936 44364 22964
rect 42291 22933 42303 22936
rect 42245 22927 42303 22933
rect 44358 22924 44364 22936
rect 44416 22924 44422 22976
rect 44652 22964 44680 23004
rect 47486 22992 47492 23044
rect 47544 23032 47550 23044
rect 51074 23032 51080 23044
rect 47544 23004 51080 23032
rect 47544 22992 47550 23004
rect 51074 22992 51080 23004
rect 51132 22992 51138 23044
rect 47121 22967 47179 22973
rect 47121 22964 47133 22967
rect 44652 22936 47133 22964
rect 47121 22933 47133 22936
rect 47167 22964 47179 22967
rect 47394 22964 47400 22976
rect 47167 22936 47400 22964
rect 47167 22933 47179 22936
rect 47121 22927 47179 22933
rect 47394 22924 47400 22936
rect 47452 22924 47458 22976
rect 47854 22924 47860 22976
rect 47912 22964 47918 22976
rect 48133 22967 48191 22973
rect 48133 22964 48145 22967
rect 47912 22936 48145 22964
rect 47912 22924 47918 22936
rect 48133 22933 48145 22936
rect 48179 22933 48191 22967
rect 51442 22964 51448 22976
rect 51403 22936 51448 22964
rect 48133 22927 48191 22933
rect 51442 22924 51448 22936
rect 51500 22964 51506 22976
rect 51629 22967 51687 22973
rect 51629 22964 51641 22967
rect 51500 22936 51641 22964
rect 51500 22924 51506 22936
rect 51629 22933 51641 22936
rect 51675 22933 51687 22967
rect 51629 22927 51687 22933
rect 1104 22874 54832 22896
rect 1104 22822 9947 22874
rect 9999 22822 10011 22874
rect 10063 22822 10075 22874
rect 10127 22822 10139 22874
rect 10191 22822 27878 22874
rect 27930 22822 27942 22874
rect 27994 22822 28006 22874
rect 28058 22822 28070 22874
rect 28122 22822 45808 22874
rect 45860 22822 45872 22874
rect 45924 22822 45936 22874
rect 45988 22822 46000 22874
rect 46052 22822 54832 22874
rect 1104 22800 54832 22822
rect 290 22720 296 22772
rect 348 22760 354 22772
rect 348 22732 17264 22760
rect 348 22720 354 22732
rect 6914 22692 6920 22704
rect 6875 22664 6920 22692
rect 6914 22652 6920 22664
rect 6972 22652 6978 22704
rect 11054 22692 11060 22704
rect 9692 22664 11060 22692
rect 3142 22624 3148 22636
rect 3103 22596 3148 22624
rect 3142 22584 3148 22596
rect 3200 22584 3206 22636
rect 3329 22627 3387 22633
rect 3329 22593 3341 22627
rect 3375 22624 3387 22627
rect 4062 22624 4068 22636
rect 3375 22596 4068 22624
rect 3375 22593 3387 22596
rect 3329 22587 3387 22593
rect 1489 22559 1547 22565
rect 1489 22525 1501 22559
rect 1535 22525 1547 22559
rect 1489 22519 1547 22525
rect 1765 22559 1823 22565
rect 1765 22525 1777 22559
rect 1811 22556 1823 22559
rect 2038 22556 2044 22568
rect 1811 22528 2044 22556
rect 1811 22525 1823 22528
rect 1765 22519 1823 22525
rect 1504 22420 1532 22519
rect 2038 22516 2044 22528
rect 2096 22516 2102 22568
rect 3344 22432 3372 22587
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4338 22584 4344 22636
rect 4396 22624 4402 22636
rect 4525 22627 4583 22633
rect 4525 22624 4537 22627
rect 4396 22596 4537 22624
rect 4396 22584 4402 22596
rect 4525 22593 4537 22596
rect 4571 22593 4583 22627
rect 4890 22624 4896 22636
rect 4803 22596 4896 22624
rect 4525 22587 4583 22593
rect 4890 22584 4896 22596
rect 4948 22624 4954 22636
rect 7098 22624 7104 22636
rect 4948 22596 7104 22624
rect 4948 22584 4954 22596
rect 7098 22584 7104 22596
rect 7156 22584 7162 22636
rect 4249 22559 4307 22565
rect 4249 22525 4261 22559
rect 4295 22525 4307 22559
rect 4249 22519 4307 22525
rect 4433 22559 4491 22565
rect 4433 22525 4445 22559
rect 4479 22556 4491 22559
rect 4479 22528 5672 22556
rect 4479 22525 4491 22528
rect 4433 22519 4491 22525
rect 4264 22488 4292 22519
rect 4890 22488 4896 22500
rect 4264 22460 4896 22488
rect 4890 22448 4896 22460
rect 4948 22448 4954 22500
rect 3326 22420 3332 22432
rect 1504 22392 3332 22420
rect 3326 22380 3332 22392
rect 3384 22380 3390 22432
rect 5644 22420 5672 22528
rect 7006 22516 7012 22568
rect 7064 22556 7070 22568
rect 7193 22559 7251 22565
rect 7193 22556 7205 22559
rect 7064 22528 7205 22556
rect 7064 22516 7070 22528
rect 7193 22525 7205 22528
rect 7239 22525 7251 22559
rect 7193 22519 7251 22525
rect 8018 22516 8024 22568
rect 8076 22556 8082 22568
rect 9692 22565 9720 22664
rect 11054 22652 11060 22664
rect 11112 22692 11118 22704
rect 11238 22692 11244 22704
rect 11112 22664 11244 22692
rect 11112 22652 11118 22664
rect 11238 22652 11244 22664
rect 11296 22652 11302 22704
rect 15013 22695 15071 22701
rect 15013 22661 15025 22695
rect 15059 22692 15071 22695
rect 15102 22692 15108 22704
rect 15059 22664 15108 22692
rect 15059 22661 15071 22664
rect 15013 22655 15071 22661
rect 10229 22627 10287 22633
rect 10229 22593 10241 22627
rect 10275 22624 10287 22627
rect 10410 22624 10416 22636
rect 10275 22596 10416 22624
rect 10275 22593 10287 22596
rect 10229 22587 10287 22593
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 9677 22559 9735 22565
rect 9677 22556 9689 22559
rect 8076 22528 9689 22556
rect 8076 22516 8082 22528
rect 9677 22525 9689 22528
rect 9723 22525 9735 22559
rect 9677 22519 9735 22525
rect 9766 22516 9772 22568
rect 9824 22556 9830 22568
rect 9953 22559 10011 22565
rect 9953 22556 9965 22559
rect 9824 22528 9965 22556
rect 9824 22516 9830 22528
rect 9953 22525 9965 22528
rect 9999 22525 10011 22559
rect 9953 22519 10011 22525
rect 11057 22559 11115 22565
rect 11057 22525 11069 22559
rect 11103 22556 11115 22559
rect 11146 22556 11152 22568
rect 11103 22528 11152 22556
rect 11103 22525 11115 22528
rect 11057 22519 11115 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12768 22528 12909 22556
rect 12768 22516 12774 22528
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 15028 22556 15056 22655
rect 15102 22652 15108 22664
rect 15160 22652 15166 22704
rect 16666 22692 16672 22704
rect 16627 22664 16672 22692
rect 16666 22652 16672 22664
rect 16724 22652 16730 22704
rect 15378 22624 15384 22636
rect 15339 22596 15384 22624
rect 15378 22584 15384 22596
rect 15436 22584 15442 22636
rect 15105 22559 15163 22565
rect 15105 22556 15117 22559
rect 15028 22528 15117 22556
rect 12897 22519 12955 22525
rect 15105 22525 15117 22528
rect 15151 22525 15163 22559
rect 15105 22519 15163 22525
rect 5718 22448 5724 22500
rect 5776 22488 5782 22500
rect 7101 22491 7159 22497
rect 7101 22488 7113 22491
rect 5776 22460 7113 22488
rect 5776 22448 5782 22460
rect 7101 22457 7113 22460
rect 7147 22488 7159 22491
rect 7374 22488 7380 22500
rect 7147 22460 7380 22488
rect 7147 22457 7159 22460
rect 7101 22451 7159 22457
rect 7374 22448 7380 22460
rect 7432 22448 7438 22500
rect 7653 22491 7711 22497
rect 7653 22457 7665 22491
rect 7699 22488 7711 22491
rect 9582 22488 9588 22500
rect 7699 22460 9588 22488
rect 7699 22457 7711 22460
rect 7653 22451 7711 22457
rect 9582 22448 9588 22460
rect 9640 22448 9646 22500
rect 10502 22420 10508 22432
rect 5644 22392 10508 22420
rect 10502 22380 10508 22392
rect 10560 22380 10566 22432
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 11149 22423 11207 22429
rect 11149 22420 11161 22423
rect 11112 22392 11161 22420
rect 11112 22380 11118 22392
rect 11149 22389 11161 22392
rect 11195 22389 11207 22423
rect 13078 22420 13084 22432
rect 13039 22392 13084 22420
rect 11149 22383 11207 22389
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 17236 22420 17264 22732
rect 18506 22720 18512 22772
rect 18564 22760 18570 22772
rect 18969 22763 19027 22769
rect 18969 22760 18981 22763
rect 18564 22732 18981 22760
rect 18564 22720 18570 22732
rect 18969 22729 18981 22732
rect 19015 22760 19027 22763
rect 19153 22763 19211 22769
rect 19153 22760 19165 22763
rect 19015 22732 19165 22760
rect 19015 22729 19027 22732
rect 18969 22723 19027 22729
rect 19153 22729 19165 22732
rect 19199 22729 19211 22763
rect 20073 22763 20131 22769
rect 20073 22760 20085 22763
rect 19153 22723 19211 22729
rect 19444 22732 20085 22760
rect 19334 22556 19340 22568
rect 19295 22528 19340 22556
rect 19334 22516 19340 22528
rect 19392 22516 19398 22568
rect 19444 22565 19472 22732
rect 20073 22729 20085 22732
rect 20119 22760 20131 22763
rect 23198 22760 23204 22772
rect 20119 22732 23204 22760
rect 20119 22729 20131 22732
rect 20073 22723 20131 22729
rect 23198 22720 23204 22732
rect 23256 22720 23262 22772
rect 23474 22720 23480 22772
rect 23532 22760 23538 22772
rect 24670 22760 24676 22772
rect 23532 22732 24676 22760
rect 23532 22720 23538 22732
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 31478 22720 31484 22772
rect 31536 22760 31542 22772
rect 31849 22763 31907 22769
rect 31849 22760 31861 22763
rect 31536 22732 31861 22760
rect 31536 22720 31542 22732
rect 31849 22729 31861 22732
rect 31895 22729 31907 22763
rect 31849 22723 31907 22729
rect 33229 22763 33287 22769
rect 33229 22729 33241 22763
rect 33275 22760 33287 22763
rect 33318 22760 33324 22772
rect 33275 22732 33324 22760
rect 33275 22729 33287 22732
rect 33229 22723 33287 22729
rect 33318 22720 33324 22732
rect 33376 22720 33382 22772
rect 33686 22760 33692 22772
rect 33647 22732 33692 22760
rect 33686 22720 33692 22732
rect 33744 22720 33750 22772
rect 34514 22720 34520 22772
rect 34572 22760 34578 22772
rect 34885 22763 34943 22769
rect 34885 22760 34897 22763
rect 34572 22732 34897 22760
rect 34572 22720 34578 22732
rect 34885 22729 34897 22732
rect 34931 22729 34943 22763
rect 34885 22723 34943 22729
rect 35066 22720 35072 22772
rect 35124 22760 35130 22772
rect 35345 22763 35403 22769
rect 35345 22760 35357 22763
rect 35124 22732 35357 22760
rect 35124 22720 35130 22732
rect 35345 22729 35357 22732
rect 35391 22729 35403 22763
rect 35345 22723 35403 22729
rect 36633 22763 36691 22769
rect 36633 22729 36645 22763
rect 36679 22760 36691 22763
rect 37366 22760 37372 22772
rect 36679 22732 37372 22760
rect 36679 22729 36691 22732
rect 36633 22723 36691 22729
rect 37366 22720 37372 22732
rect 37424 22720 37430 22772
rect 37734 22720 37740 22772
rect 37792 22760 37798 22772
rect 38378 22760 38384 22772
rect 37792 22732 38384 22760
rect 37792 22720 37798 22732
rect 38378 22720 38384 22732
rect 38436 22720 38442 22772
rect 38746 22760 38752 22772
rect 38707 22732 38752 22760
rect 38746 22720 38752 22732
rect 38804 22720 38810 22772
rect 41874 22720 41880 22772
rect 41932 22760 41938 22772
rect 42794 22760 42800 22772
rect 41932 22732 42800 22760
rect 41932 22720 41938 22732
rect 42794 22720 42800 22732
rect 42852 22760 42858 22772
rect 43070 22760 43076 22772
rect 42852 22732 43076 22760
rect 42852 22720 42858 22732
rect 43070 22720 43076 22732
rect 43128 22720 43134 22772
rect 51442 22760 51448 22772
rect 46492 22732 51448 22760
rect 20714 22692 20720 22704
rect 20675 22664 20720 22692
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 20806 22652 20812 22704
rect 20864 22692 20870 22704
rect 21634 22692 21640 22704
rect 20864 22664 21496 22692
rect 21595 22664 21640 22692
rect 20864 22652 20870 22664
rect 19889 22627 19947 22633
rect 19889 22593 19901 22627
rect 19935 22624 19947 22627
rect 21174 22624 21180 22636
rect 19935 22596 21180 22624
rect 19935 22593 19947 22596
rect 19889 22587 19947 22593
rect 21174 22584 21180 22596
rect 21232 22584 21238 22636
rect 21468 22633 21496 22664
rect 21634 22652 21640 22664
rect 21692 22652 21698 22704
rect 23290 22652 23296 22704
rect 23348 22692 23354 22704
rect 25777 22695 25835 22701
rect 25777 22692 25789 22695
rect 23348 22664 25789 22692
rect 23348 22652 23354 22664
rect 25777 22661 25789 22664
rect 25823 22661 25835 22695
rect 28258 22692 28264 22704
rect 25777 22655 25835 22661
rect 26988 22664 28264 22692
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 26694 22624 26700 22636
rect 21968 22596 26700 22624
rect 21968 22584 21974 22596
rect 26694 22584 26700 22596
rect 26752 22584 26758 22636
rect 26988 22633 27016 22664
rect 28258 22652 28264 22664
rect 28316 22652 28322 22704
rect 31389 22695 31447 22701
rect 31389 22661 31401 22695
rect 31435 22692 31447 22695
rect 31570 22692 31576 22704
rect 31435 22664 31576 22692
rect 31435 22661 31447 22664
rect 31389 22655 31447 22661
rect 31570 22652 31576 22664
rect 31628 22652 31634 22704
rect 40586 22692 40592 22704
rect 32048 22664 40592 22692
rect 26973 22627 27031 22633
rect 26973 22593 26985 22627
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 28166 22584 28172 22636
rect 28224 22624 28230 22636
rect 32048 22624 32076 22664
rect 40586 22652 40592 22664
rect 40644 22652 40650 22704
rect 40681 22695 40739 22701
rect 40681 22661 40693 22695
rect 40727 22692 40739 22695
rect 46492 22692 46520 22732
rect 51442 22720 51448 22732
rect 51500 22720 51506 22772
rect 40727 22664 46520 22692
rect 40727 22661 40739 22664
rect 40681 22655 40739 22661
rect 28224 22596 32076 22624
rect 28224 22584 28230 22596
rect 32122 22584 32128 22636
rect 32180 22624 32186 22636
rect 32180 22596 36492 22624
rect 32180 22584 32186 22596
rect 19429 22559 19487 22565
rect 19429 22525 19441 22559
rect 19475 22525 19487 22559
rect 20990 22556 20996 22568
rect 20951 22528 20996 22556
rect 19429 22519 19487 22525
rect 20990 22516 20996 22528
rect 21048 22516 21054 22568
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 24026 22556 24032 22568
rect 21140 22528 23428 22556
rect 23987 22528 24032 22556
rect 21140 22516 21146 22528
rect 19352 22488 19380 22516
rect 20901 22491 20959 22497
rect 20901 22488 20913 22491
rect 19352 22460 20913 22488
rect 20901 22457 20913 22460
rect 20947 22488 20959 22491
rect 22186 22488 22192 22500
rect 20947 22460 22192 22488
rect 20947 22457 20959 22460
rect 20901 22451 20959 22457
rect 22186 22448 22192 22460
rect 22244 22488 22250 22500
rect 23290 22488 23296 22500
rect 22244 22460 23296 22488
rect 22244 22448 22250 22460
rect 23290 22448 23296 22460
rect 23348 22448 23354 22500
rect 23400 22488 23428 22528
rect 24026 22516 24032 22528
rect 24084 22516 24090 22568
rect 24210 22556 24216 22568
rect 24171 22528 24216 22556
rect 24210 22516 24216 22528
rect 24268 22516 24274 22568
rect 24302 22516 24308 22568
rect 24360 22556 24366 22568
rect 25590 22556 25596 22568
rect 24360 22528 24405 22556
rect 25551 22528 25596 22556
rect 24360 22516 24366 22528
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 27065 22559 27123 22565
rect 27065 22525 27077 22559
rect 27111 22556 27123 22559
rect 27154 22556 27160 22568
rect 27111 22528 27160 22556
rect 27111 22525 27123 22528
rect 27065 22519 27123 22525
rect 27154 22516 27160 22528
rect 27212 22556 27218 22568
rect 27617 22559 27675 22565
rect 27617 22556 27629 22559
rect 27212 22528 27629 22556
rect 27212 22516 27218 22528
rect 27617 22525 27629 22528
rect 27663 22525 27675 22559
rect 27617 22519 27675 22525
rect 27801 22559 27859 22565
rect 27801 22525 27813 22559
rect 27847 22525 27859 22559
rect 29270 22556 29276 22568
rect 29231 22528 29276 22556
rect 27801 22519 27859 22525
rect 24765 22491 24823 22497
rect 23400 22460 24348 22488
rect 22370 22420 22376 22432
rect 17236 22392 22376 22420
rect 22370 22380 22376 22392
rect 22428 22420 22434 22432
rect 23845 22423 23903 22429
rect 23845 22420 23857 22423
rect 22428 22392 23857 22420
rect 22428 22380 22434 22392
rect 23845 22389 23857 22392
rect 23891 22420 23903 22423
rect 24210 22420 24216 22432
rect 23891 22392 24216 22420
rect 23891 22389 23903 22392
rect 23845 22383 23903 22389
rect 24210 22380 24216 22392
rect 24268 22380 24274 22432
rect 24320 22420 24348 22460
rect 24765 22457 24777 22491
rect 24811 22488 24823 22491
rect 25222 22488 25228 22500
rect 24811 22460 25228 22488
rect 24811 22457 24823 22460
rect 24765 22451 24823 22457
rect 25222 22448 25228 22460
rect 25280 22448 25286 22500
rect 25498 22420 25504 22432
rect 24320 22392 25504 22420
rect 25498 22380 25504 22392
rect 25556 22380 25562 22432
rect 26510 22380 26516 22432
rect 26568 22420 26574 22432
rect 27816 22420 27844 22519
rect 29270 22516 29276 22528
rect 29328 22516 29334 22568
rect 31665 22559 31723 22565
rect 31665 22525 31677 22559
rect 31711 22525 31723 22559
rect 33502 22556 33508 22568
rect 33463 22528 33508 22556
rect 31665 22519 31723 22525
rect 28166 22488 28172 22500
rect 28127 22460 28172 22488
rect 28166 22448 28172 22460
rect 28224 22448 28230 22500
rect 28258 22448 28264 22500
rect 28316 22488 28322 22500
rect 29454 22488 29460 22500
rect 28316 22460 29460 22488
rect 28316 22448 28322 22460
rect 29454 22448 29460 22460
rect 29512 22448 29518 22500
rect 31573 22491 31631 22497
rect 31573 22457 31585 22491
rect 31619 22457 31631 22491
rect 31680 22488 31708 22519
rect 33502 22516 33508 22528
rect 33560 22516 33566 22568
rect 36464 22565 36492 22596
rect 37182 22584 37188 22636
rect 37240 22624 37246 22636
rect 37553 22627 37611 22633
rect 37553 22624 37565 22627
rect 37240 22596 37565 22624
rect 37240 22584 37246 22596
rect 37553 22593 37565 22596
rect 37599 22593 37611 22627
rect 37553 22587 37611 22593
rect 38746 22584 38752 22636
rect 38804 22624 38810 22636
rect 40696 22624 40724 22655
rect 38804 22596 40724 22624
rect 38804 22584 38810 22596
rect 41598 22584 41604 22636
rect 41656 22624 41662 22636
rect 42242 22624 42248 22636
rect 41656 22596 42248 22624
rect 41656 22584 41662 22596
rect 42242 22584 42248 22596
rect 42300 22584 42306 22636
rect 44358 22584 44364 22636
rect 44416 22624 44422 22636
rect 48869 22627 48927 22633
rect 48869 22624 48881 22627
rect 44416 22596 48881 22624
rect 44416 22584 44422 22596
rect 48869 22593 48881 22596
rect 48915 22593 48927 22627
rect 48869 22587 48927 22593
rect 48958 22584 48964 22636
rect 49016 22624 49022 22636
rect 53469 22627 53527 22633
rect 53469 22624 53481 22627
rect 49016 22596 53481 22624
rect 49016 22584 49022 22596
rect 53469 22593 53481 22596
rect 53515 22593 53527 22627
rect 53469 22587 53527 22593
rect 35161 22559 35219 22565
rect 35161 22525 35173 22559
rect 35207 22525 35219 22559
rect 35161 22519 35219 22525
rect 36449 22559 36507 22565
rect 36449 22525 36461 22559
rect 36495 22525 36507 22559
rect 37734 22556 37740 22568
rect 37695 22528 37740 22556
rect 36449 22519 36507 22525
rect 32306 22488 32312 22500
rect 31680 22460 32312 22488
rect 31573 22451 31631 22457
rect 28350 22420 28356 22432
rect 26568 22392 28356 22420
rect 26568 22380 26574 22392
rect 28350 22380 28356 22392
rect 28408 22380 28414 22432
rect 28810 22380 28816 22432
rect 28868 22420 28874 22432
rect 29365 22423 29423 22429
rect 29365 22420 29377 22423
rect 28868 22392 29377 22420
rect 28868 22380 28874 22392
rect 29365 22389 29377 22392
rect 29411 22389 29423 22423
rect 31588 22420 31616 22451
rect 32306 22448 32312 22460
rect 32364 22448 32370 22500
rect 33410 22488 33416 22500
rect 33323 22460 33416 22488
rect 33410 22448 33416 22460
rect 33468 22488 33474 22500
rect 35069 22491 35127 22497
rect 35069 22488 35081 22491
rect 33468 22460 35081 22488
rect 33468 22448 33474 22460
rect 35069 22457 35081 22460
rect 35115 22457 35127 22491
rect 35176 22488 35204 22519
rect 37734 22516 37740 22528
rect 37792 22556 37798 22568
rect 38289 22559 38347 22565
rect 38289 22556 38301 22559
rect 37792 22528 38301 22556
rect 37792 22516 37798 22528
rect 38289 22525 38301 22528
rect 38335 22525 38347 22559
rect 38289 22519 38347 22525
rect 38473 22559 38531 22565
rect 38473 22525 38485 22559
rect 38519 22556 38531 22559
rect 38838 22556 38844 22568
rect 38519 22528 38844 22556
rect 38519 22525 38531 22528
rect 38473 22519 38531 22525
rect 38838 22516 38844 22528
rect 38896 22556 38902 22568
rect 39482 22556 39488 22568
rect 38896 22528 39488 22556
rect 38896 22516 38902 22528
rect 39482 22516 39488 22528
rect 39540 22516 39546 22568
rect 40402 22516 40408 22568
rect 40460 22556 40466 22568
rect 40497 22559 40555 22565
rect 40497 22556 40509 22559
rect 40460 22528 40509 22556
rect 40460 22516 40466 22528
rect 40497 22525 40509 22528
rect 40543 22525 40555 22559
rect 40497 22519 40555 22525
rect 41874 22516 41880 22568
rect 41932 22556 41938 22568
rect 42429 22559 42487 22565
rect 42429 22556 42441 22559
rect 41932 22528 42441 22556
rect 41932 22516 41938 22528
rect 42429 22525 42441 22528
rect 42475 22525 42487 22559
rect 42429 22519 42487 22525
rect 42521 22559 42579 22565
rect 42521 22525 42533 22559
rect 42567 22556 42579 22559
rect 42610 22556 42616 22568
rect 42567 22528 42616 22556
rect 42567 22525 42579 22528
rect 42521 22519 42579 22525
rect 42610 22516 42616 22528
rect 42668 22516 42674 22568
rect 42889 22559 42947 22565
rect 42889 22525 42901 22559
rect 42935 22525 42947 22559
rect 42889 22519 42947 22525
rect 42981 22559 43039 22565
rect 42981 22525 42993 22559
rect 43027 22556 43039 22559
rect 43070 22556 43076 22568
rect 43027 22528 43076 22556
rect 43027 22525 43039 22528
rect 42981 22519 43039 22525
rect 35805 22491 35863 22497
rect 35805 22488 35817 22491
rect 35176 22460 35817 22488
rect 35069 22451 35127 22457
rect 35805 22457 35817 22460
rect 35851 22488 35863 22491
rect 35851 22460 37136 22488
rect 35851 22457 35863 22460
rect 35805 22451 35863 22457
rect 32214 22420 32220 22432
rect 31588 22392 32220 22420
rect 29365 22383 29423 22389
rect 32214 22380 32220 22392
rect 32272 22420 32278 22432
rect 33428 22420 33456 22448
rect 32272 22392 33456 22420
rect 37108 22420 37136 22460
rect 37274 22448 37280 22500
rect 37332 22488 37338 22500
rect 40218 22488 40224 22500
rect 37332 22460 40224 22488
rect 37332 22448 37338 22460
rect 40218 22448 40224 22460
rect 40276 22448 40282 22500
rect 41966 22448 41972 22500
rect 42024 22488 42030 22500
rect 42061 22491 42119 22497
rect 42061 22488 42073 22491
rect 42024 22460 42073 22488
rect 42024 22448 42030 22460
rect 42061 22457 42073 22460
rect 42107 22488 42119 22491
rect 42904 22488 42932 22519
rect 43070 22516 43076 22528
rect 43128 22516 43134 22568
rect 46109 22559 46167 22565
rect 46109 22525 46121 22559
rect 46155 22556 46167 22559
rect 46382 22556 46388 22568
rect 46155 22528 46388 22556
rect 46155 22525 46167 22528
rect 46109 22519 46167 22525
rect 46382 22516 46388 22528
rect 46440 22516 46446 22568
rect 48501 22559 48559 22565
rect 48501 22525 48513 22559
rect 48547 22556 48559 22559
rect 48590 22556 48596 22568
rect 48547 22528 48596 22556
rect 48547 22525 48559 22528
rect 48501 22519 48559 22525
rect 48590 22516 48596 22528
rect 48648 22516 48654 22568
rect 52089 22559 52147 22565
rect 52089 22525 52101 22559
rect 52135 22525 52147 22559
rect 52089 22519 52147 22525
rect 52365 22559 52423 22565
rect 52365 22525 52377 22559
rect 52411 22556 52423 22559
rect 52454 22556 52460 22568
rect 52411 22528 52460 22556
rect 52411 22525 52423 22528
rect 52365 22519 52423 22525
rect 43530 22488 43536 22500
rect 42107 22460 42932 22488
rect 43491 22460 43536 22488
rect 42107 22457 42119 22460
rect 42061 22451 42119 22457
rect 43530 22448 43536 22460
rect 43588 22448 43594 22500
rect 49528 22460 50108 22488
rect 41230 22420 41236 22432
rect 37108 22392 41236 22420
rect 32272 22380 32278 22392
rect 41230 22380 41236 22392
rect 41288 22380 41294 22432
rect 44818 22380 44824 22432
rect 44876 22420 44882 22432
rect 46201 22423 46259 22429
rect 46201 22420 46213 22423
rect 44876 22392 46213 22420
rect 44876 22380 44882 22392
rect 46201 22389 46213 22392
rect 46247 22389 46259 22423
rect 46201 22383 46259 22389
rect 46290 22380 46296 22432
rect 46348 22420 46354 22432
rect 49528 22420 49556 22460
rect 49970 22420 49976 22432
rect 46348 22392 49556 22420
rect 49931 22392 49976 22420
rect 46348 22380 46354 22392
rect 49970 22380 49976 22392
rect 50028 22380 50034 22432
rect 50080 22420 50108 22460
rect 51810 22448 51816 22500
rect 51868 22488 51874 22500
rect 51905 22491 51963 22497
rect 51905 22488 51917 22491
rect 51868 22460 51917 22488
rect 51868 22448 51874 22460
rect 51905 22457 51917 22460
rect 51951 22488 51963 22491
rect 52104 22488 52132 22519
rect 52454 22516 52460 22528
rect 52512 22516 52518 22568
rect 51951 22460 52132 22488
rect 51951 22457 51963 22460
rect 51905 22451 51963 22457
rect 54110 22420 54116 22432
rect 50080 22392 54116 22420
rect 54110 22380 54116 22392
rect 54168 22380 54174 22432
rect 1104 22330 54832 22352
rect 1104 22278 18912 22330
rect 18964 22278 18976 22330
rect 19028 22278 19040 22330
rect 19092 22278 19104 22330
rect 19156 22278 36843 22330
rect 36895 22278 36907 22330
rect 36959 22278 36971 22330
rect 37023 22278 37035 22330
rect 37087 22278 54832 22330
rect 1104 22256 54832 22278
rect 2038 22216 2044 22228
rect 1999 22188 2044 22216
rect 2038 22176 2044 22188
rect 2096 22176 2102 22228
rect 4157 22219 4215 22225
rect 4157 22185 4169 22219
rect 4203 22216 4215 22219
rect 4246 22216 4252 22228
rect 4203 22188 4252 22216
rect 4203 22185 4215 22188
rect 4157 22179 4215 22185
rect 4246 22176 4252 22188
rect 4304 22176 4310 22228
rect 4890 22216 4896 22228
rect 4851 22188 4896 22216
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 6914 22216 6920 22228
rect 6696 22188 6920 22216
rect 6696 22176 6702 22188
rect 6914 22176 6920 22188
rect 6972 22176 6978 22228
rect 7098 22176 7104 22228
rect 7156 22216 7162 22228
rect 13078 22216 13084 22228
rect 7156 22188 13084 22216
rect 7156 22176 7162 22188
rect 13078 22176 13084 22188
rect 13136 22216 13142 22228
rect 14826 22216 14832 22228
rect 13136 22188 14832 22216
rect 13136 22176 13142 22188
rect 14826 22176 14832 22188
rect 14884 22176 14890 22228
rect 20898 22176 20904 22228
rect 20956 22216 20962 22228
rect 21910 22216 21916 22228
rect 20956 22188 21916 22216
rect 20956 22176 20962 22188
rect 2869 22151 2927 22157
rect 2869 22148 2881 22151
rect 2240 22120 2881 22148
rect 2240 22089 2268 22120
rect 2869 22117 2881 22120
rect 2915 22148 2927 22151
rect 4908 22148 4936 22176
rect 2915 22120 4936 22148
rect 2915 22117 2927 22120
rect 2869 22111 2927 22117
rect 2225 22083 2283 22089
rect 2225 22049 2237 22083
rect 2271 22049 2283 22083
rect 2498 22080 2504 22092
rect 2459 22052 2504 22080
rect 2225 22043 2283 22049
rect 2498 22040 2504 22052
rect 2556 22040 2562 22092
rect 4356 22089 4384 22120
rect 5718 22108 5724 22160
rect 5776 22148 5782 22160
rect 5776 22120 5948 22148
rect 5776 22108 5782 22120
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22049 4399 22083
rect 4614 22080 4620 22092
rect 4575 22052 4620 22080
rect 4341 22043 4399 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 5920 22089 5948 22120
rect 10428 22120 11560 22148
rect 5905 22083 5963 22089
rect 5905 22049 5917 22083
rect 5951 22049 5963 22083
rect 5905 22043 5963 22049
rect 6178 22040 6184 22092
rect 6236 22080 6242 22092
rect 6730 22080 6736 22092
rect 6236 22052 6736 22080
rect 6236 22040 6242 22052
rect 6730 22040 6736 22052
rect 6788 22040 6794 22092
rect 6917 22083 6975 22089
rect 6917 22049 6929 22083
rect 6963 22080 6975 22083
rect 7006 22080 7012 22092
rect 6963 22052 7012 22080
rect 6963 22049 6975 22052
rect 6917 22043 6975 22049
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 7193 22083 7251 22089
rect 7193 22049 7205 22083
rect 7239 22049 7251 22083
rect 7193 22043 7251 22049
rect 7653 22083 7711 22089
rect 7653 22049 7665 22083
rect 7699 22080 7711 22083
rect 8570 22080 8576 22092
rect 7699 22052 8576 22080
rect 7699 22049 7711 22052
rect 7653 22043 7711 22049
rect 5810 21972 5816 22024
rect 5868 22012 5874 22024
rect 7208 22012 7236 22043
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 9674 22040 9680 22092
rect 9732 22080 9738 22092
rect 10428 22089 10456 22120
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 9732 22052 9873 22080
rect 9732 22040 9738 22052
rect 9861 22049 9873 22052
rect 9907 22049 9919 22083
rect 9861 22043 9919 22049
rect 10413 22083 10471 22089
rect 10413 22049 10425 22083
rect 10459 22080 10471 22083
rect 10594 22080 10600 22092
rect 10459 22052 10493 22080
rect 10555 22052 10600 22080
rect 10459 22049 10471 22052
rect 10413 22043 10471 22049
rect 10594 22040 10600 22052
rect 10652 22040 10658 22092
rect 10781 22083 10839 22089
rect 10781 22049 10793 22083
rect 10827 22080 10839 22083
rect 10870 22080 10876 22092
rect 10827 22052 10876 22080
rect 10827 22049 10839 22052
rect 10781 22043 10839 22049
rect 10870 22040 10876 22052
rect 10928 22040 10934 22092
rect 10965 22083 11023 22089
rect 10965 22049 10977 22083
rect 11011 22080 11023 22083
rect 11054 22080 11060 22092
rect 11011 22052 11060 22080
rect 11011 22049 11023 22052
rect 10965 22043 11023 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11149 22083 11207 22089
rect 11149 22049 11161 22083
rect 11195 22049 11207 22083
rect 11532 22080 11560 22120
rect 11606 22080 11612 22092
rect 11532 22052 11612 22080
rect 11149 22043 11207 22049
rect 11164 22012 11192 22043
rect 11606 22040 11612 22052
rect 11664 22040 11670 22092
rect 12529 22083 12587 22089
rect 12529 22049 12541 22083
rect 12575 22080 12587 22083
rect 12710 22080 12716 22092
rect 12575 22052 12716 22080
rect 12575 22049 12587 22052
rect 12529 22043 12587 22049
rect 12710 22040 12716 22052
rect 12768 22040 12774 22092
rect 21100 22089 21128 22188
rect 21910 22176 21916 22188
rect 21968 22176 21974 22228
rect 23198 22176 23204 22228
rect 23256 22216 23262 22228
rect 29086 22216 29092 22228
rect 23256 22188 29092 22216
rect 23256 22176 23262 22188
rect 29086 22176 29092 22188
rect 29144 22176 29150 22228
rect 29454 22176 29460 22228
rect 29512 22216 29518 22228
rect 42150 22216 42156 22228
rect 29512 22188 42156 22216
rect 29512 22176 29518 22188
rect 42150 22176 42156 22188
rect 42208 22176 42214 22228
rect 42334 22216 42340 22228
rect 42295 22188 42340 22216
rect 42334 22176 42340 22188
rect 42392 22176 42398 22228
rect 45002 22176 45008 22228
rect 45060 22216 45066 22228
rect 48958 22216 48964 22228
rect 45060 22188 48964 22216
rect 45060 22176 45066 22188
rect 48958 22176 48964 22188
rect 49016 22176 49022 22228
rect 51442 22176 51448 22228
rect 51500 22216 51506 22228
rect 51905 22219 51963 22225
rect 51905 22216 51917 22219
rect 51500 22188 51917 22216
rect 51500 22176 51506 22188
rect 51905 22185 51917 22188
rect 51951 22185 51963 22219
rect 51905 22179 51963 22185
rect 21634 22108 21640 22160
rect 21692 22148 21698 22160
rect 21729 22151 21787 22157
rect 21729 22148 21741 22151
rect 21692 22120 21741 22148
rect 21692 22108 21698 22120
rect 21729 22117 21741 22120
rect 21775 22117 21787 22151
rect 21729 22111 21787 22117
rect 23477 22151 23535 22157
rect 23477 22117 23489 22151
rect 23523 22148 23535 22151
rect 23523 22120 24311 22148
rect 23523 22117 23535 22120
rect 23477 22111 23535 22117
rect 24283 22092 24311 22120
rect 33502 22108 33508 22160
rect 33560 22148 33566 22160
rect 33560 22120 39712 22148
rect 33560 22108 33566 22120
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22049 13691 22083
rect 18877 22083 18935 22089
rect 18877 22080 18889 22083
rect 13633 22043 13691 22049
rect 17144 22052 18889 22080
rect 13648 22012 13676 22043
rect 17144 22024 17172 22052
rect 18877 22049 18889 22052
rect 18923 22049 18935 22083
rect 18877 22043 18935 22049
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22049 21143 22083
rect 21085 22043 21143 22049
rect 21218 22083 21276 22089
rect 21218 22049 21230 22083
rect 21264 22080 21276 22083
rect 21450 22080 21456 22092
rect 21264 22052 21456 22080
rect 21264 22049 21276 22052
rect 21218 22043 21276 22049
rect 21450 22040 21456 22052
rect 21508 22040 21514 22092
rect 22554 22080 22560 22092
rect 22515 22052 22560 22080
rect 22554 22040 22560 22052
rect 22612 22040 22618 22092
rect 23750 22080 23756 22092
rect 23711 22052 23756 22080
rect 23750 22040 23756 22052
rect 23808 22040 23814 22092
rect 24283 22080 24308 22092
rect 24263 22052 24308 22080
rect 24302 22040 24308 22052
rect 24360 22040 24366 22092
rect 26694 22040 26700 22092
rect 26752 22080 26758 22092
rect 26973 22083 27031 22089
rect 26973 22080 26985 22083
rect 26752 22052 26985 22080
rect 26752 22040 26758 22052
rect 26973 22049 26985 22052
rect 27019 22049 27031 22083
rect 26973 22043 27031 22049
rect 28166 22040 28172 22092
rect 28224 22080 28230 22092
rect 28629 22083 28687 22089
rect 28629 22080 28641 22083
rect 28224 22052 28641 22080
rect 28224 22040 28230 22052
rect 28629 22049 28641 22052
rect 28675 22049 28687 22083
rect 33962 22080 33968 22092
rect 33923 22052 33968 22080
rect 28629 22043 28687 22049
rect 33962 22040 33968 22052
rect 34020 22040 34026 22092
rect 34146 22080 34152 22092
rect 34107 22052 34152 22080
rect 34146 22040 34152 22052
rect 34204 22080 34210 22092
rect 34701 22083 34759 22089
rect 34701 22080 34713 22083
rect 34204 22052 34713 22080
rect 34204 22040 34210 22052
rect 34701 22049 34713 22052
rect 34747 22049 34759 22083
rect 34882 22080 34888 22092
rect 34843 22052 34888 22080
rect 34701 22043 34759 22049
rect 34882 22040 34888 22052
rect 34940 22040 34946 22092
rect 39684 22080 39712 22120
rect 41322 22108 41328 22160
rect 41380 22148 41386 22160
rect 44637 22151 44695 22157
rect 41380 22120 42196 22148
rect 41380 22108 41386 22120
rect 40126 22080 40132 22092
rect 39684 22052 40132 22080
rect 40126 22040 40132 22052
rect 40184 22040 40190 22092
rect 17126 22012 17132 22024
rect 5868 21984 7236 22012
rect 11072 21984 13676 22012
rect 17087 21984 17132 22012
rect 5868 21972 5874 21984
rect 5997 21947 6055 21953
rect 5997 21913 6009 21947
rect 6043 21944 6055 21947
rect 7009 21947 7067 21953
rect 7009 21944 7021 21947
rect 6043 21916 7021 21944
rect 6043 21913 6055 21916
rect 5997 21907 6055 21913
rect 7009 21913 7021 21916
rect 7055 21944 7067 21947
rect 7098 21944 7104 21956
rect 7055 21916 7104 21944
rect 7055 21913 7067 21916
rect 7009 21907 7067 21913
rect 7098 21904 7104 21916
rect 7156 21904 7162 21956
rect 7282 21904 7288 21956
rect 7340 21944 7346 21956
rect 7340 21916 9536 21944
rect 7340 21904 7346 21916
rect 8665 21879 8723 21885
rect 8665 21845 8677 21879
rect 8711 21876 8723 21879
rect 9398 21876 9404 21888
rect 8711 21848 9404 21876
rect 8711 21845 8723 21848
rect 8665 21839 8723 21845
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9508 21876 9536 21916
rect 9582 21904 9588 21956
rect 9640 21944 9646 21956
rect 11072 21944 11100 21984
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 17402 22012 17408 22024
rect 17363 21984 17408 22012
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 18785 22015 18843 22021
rect 18785 21981 18797 22015
rect 18831 22012 18843 22015
rect 18831 21984 23796 22012
rect 18831 21981 18843 21984
rect 18785 21975 18843 21981
rect 9640 21916 11100 21944
rect 9640 21904 9646 21916
rect 11238 21904 11244 21956
rect 11296 21944 11302 21956
rect 12713 21947 12771 21953
rect 12713 21944 12725 21947
rect 11296 21916 12725 21944
rect 11296 21904 11302 21916
rect 12713 21913 12725 21916
rect 12759 21913 12771 21947
rect 12713 21907 12771 21913
rect 20901 21947 20959 21953
rect 20901 21913 20913 21947
rect 20947 21944 20959 21947
rect 21634 21944 21640 21956
rect 20947 21916 21640 21944
rect 20947 21913 20959 21916
rect 20901 21907 20959 21913
rect 21634 21904 21640 21916
rect 21692 21904 21698 21956
rect 22278 21904 22284 21956
rect 22336 21944 22342 21956
rect 23201 21947 23259 21953
rect 23201 21944 23213 21947
rect 22336 21916 23213 21944
rect 22336 21904 22342 21916
rect 23201 21913 23213 21916
rect 23247 21944 23259 21947
rect 23474 21944 23480 21956
rect 23247 21916 23480 21944
rect 23247 21913 23259 21916
rect 23201 21907 23259 21913
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 23658 21944 23664 21956
rect 23619 21916 23664 21944
rect 23658 21904 23664 21916
rect 23716 21904 23722 21956
rect 23768 21944 23796 21984
rect 23842 21972 23848 22024
rect 23900 22012 23906 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 23900 21984 24409 22012
rect 23900 21972 23906 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 24857 22015 24915 22021
rect 24857 22012 24869 22015
rect 24820 21984 24869 22012
rect 24820 21972 24826 21984
rect 24857 21981 24869 21984
rect 24903 22012 24915 22015
rect 28258 22012 28264 22024
rect 24903 21984 28264 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 28258 21972 28264 21984
rect 28316 21972 28322 22024
rect 28353 22015 28411 22021
rect 28353 21981 28365 22015
rect 28399 22012 28411 22015
rect 28994 22012 29000 22024
rect 28399 21984 29000 22012
rect 28399 21981 28411 21984
rect 28353 21975 28411 21981
rect 23768 21916 27292 21944
rect 9674 21876 9680 21888
rect 9508 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 11514 21876 11520 21888
rect 11475 21848 11520 21876
rect 11514 21836 11520 21848
rect 11572 21836 11578 21888
rect 13725 21879 13783 21885
rect 13725 21845 13737 21879
rect 13771 21876 13783 21879
rect 15562 21876 15568 21888
rect 13771 21848 15568 21876
rect 13771 21845 13783 21848
rect 13725 21839 13783 21845
rect 15562 21836 15568 21848
rect 15620 21876 15626 21888
rect 15838 21876 15844 21888
rect 15620 21848 15844 21876
rect 15620 21836 15626 21848
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 21358 21876 21364 21888
rect 21319 21848 21364 21876
rect 21358 21836 21364 21848
rect 21416 21836 21422 21888
rect 22649 21879 22707 21885
rect 22649 21845 22661 21879
rect 22695 21876 22707 21879
rect 22738 21876 22744 21888
rect 22695 21848 22744 21876
rect 22695 21845 22707 21848
rect 22649 21839 22707 21845
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 26694 21836 26700 21888
rect 26752 21876 26758 21888
rect 26789 21879 26847 21885
rect 26789 21876 26801 21879
rect 26752 21848 26801 21876
rect 26752 21836 26758 21848
rect 26789 21845 26801 21848
rect 26835 21845 26847 21879
rect 27154 21876 27160 21888
rect 27115 21848 27160 21876
rect 26789 21839 26847 21845
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 27264 21876 27292 21916
rect 27614 21904 27620 21956
rect 27672 21944 27678 21956
rect 28368 21944 28396 21975
rect 28994 21972 29000 21984
rect 29052 22012 29058 22024
rect 29362 22012 29368 22024
rect 29052 21984 29368 22012
rect 29052 21972 29058 21984
rect 29362 21972 29368 21984
rect 29420 22012 29426 22024
rect 30101 22015 30159 22021
rect 30101 22012 30113 22015
rect 29420 21984 30113 22012
rect 29420 21972 29426 21984
rect 30101 21981 30113 21984
rect 30147 22012 30159 22015
rect 31018 22012 31024 22024
rect 30147 21984 31024 22012
rect 30147 21981 30159 21984
rect 30101 21975 30159 21981
rect 31018 21972 31024 21984
rect 31076 22012 31082 22024
rect 32766 22012 32772 22024
rect 31076 21984 32772 22012
rect 31076 21972 31082 21984
rect 32766 21972 32772 21984
rect 32824 21972 32830 22024
rect 39577 22015 39635 22021
rect 39577 22012 39589 22015
rect 39408 21984 39589 22012
rect 27672 21916 28396 21944
rect 27672 21904 27678 21916
rect 29086 21876 29092 21888
rect 27264 21848 29092 21876
rect 29086 21836 29092 21848
rect 29144 21836 29150 21888
rect 29730 21876 29736 21888
rect 29691 21848 29736 21876
rect 29730 21836 29736 21848
rect 29788 21836 29794 21888
rect 35161 21879 35219 21885
rect 35161 21845 35173 21879
rect 35207 21876 35219 21879
rect 35618 21876 35624 21888
rect 35207 21848 35624 21876
rect 35207 21845 35219 21848
rect 35161 21839 35219 21845
rect 35618 21836 35624 21848
rect 35676 21836 35682 21888
rect 38194 21836 38200 21888
rect 38252 21876 38258 21888
rect 39408 21885 39436 21984
rect 39577 21981 39589 21984
rect 39623 21981 39635 22015
rect 39850 22012 39856 22024
rect 39811 21984 39856 22012
rect 39577 21975 39635 21981
rect 39850 21972 39856 21984
rect 39908 21972 39914 22024
rect 42168 22012 42196 22120
rect 44637 22117 44649 22151
rect 44683 22148 44695 22151
rect 44910 22148 44916 22160
rect 44683 22120 44916 22148
rect 44683 22117 44695 22120
rect 44637 22111 44695 22117
rect 44910 22108 44916 22120
rect 44968 22108 44974 22160
rect 51718 22148 51724 22160
rect 51679 22120 51724 22148
rect 51718 22108 51724 22120
rect 51776 22108 51782 22160
rect 42242 22040 42248 22092
rect 42300 22080 42306 22092
rect 42610 22080 42616 22092
rect 42300 22052 42616 22080
rect 42300 22040 42306 22052
rect 42610 22040 42616 22052
rect 42668 22040 42674 22092
rect 42794 22040 42800 22092
rect 42852 22080 42858 22092
rect 43533 22083 43591 22089
rect 43533 22080 43545 22083
rect 42852 22052 43545 22080
rect 42852 22040 42858 22052
rect 43533 22049 43545 22052
rect 43579 22080 43591 22083
rect 44085 22083 44143 22089
rect 44085 22080 44097 22083
rect 43579 22052 44097 22080
rect 43579 22049 43591 22052
rect 43533 22043 43591 22049
rect 44085 22049 44097 22052
rect 44131 22049 44143 22083
rect 44266 22080 44272 22092
rect 44227 22052 44272 22080
rect 44085 22043 44143 22049
rect 44266 22040 44272 22052
rect 44324 22080 44330 22092
rect 44818 22080 44824 22092
rect 44324 22052 44824 22080
rect 44324 22040 44330 22052
rect 44818 22040 44824 22052
rect 44876 22040 44882 22092
rect 46106 22040 46112 22092
rect 46164 22080 46170 22092
rect 46569 22083 46627 22089
rect 46569 22080 46581 22083
rect 46164 22052 46581 22080
rect 46164 22040 46170 22052
rect 46569 22049 46581 22052
rect 46615 22049 46627 22083
rect 46569 22043 46627 22049
rect 49786 22040 49792 22092
rect 49844 22080 49850 22092
rect 49881 22083 49939 22089
rect 49881 22080 49893 22083
rect 49844 22052 49893 22080
rect 49844 22040 49850 22052
rect 49881 22049 49893 22052
rect 49927 22049 49939 22083
rect 50062 22080 50068 22092
rect 50023 22052 50068 22080
rect 49881 22043 49939 22049
rect 50062 22040 50068 22052
rect 50120 22080 50126 22092
rect 50617 22083 50675 22089
rect 50617 22080 50629 22083
rect 50120 22052 50629 22080
rect 50120 22040 50126 22052
rect 50617 22049 50629 22052
rect 50663 22049 50675 22083
rect 50617 22043 50675 22049
rect 50706 22040 50712 22092
rect 50764 22080 50770 22092
rect 50801 22083 50859 22089
rect 50801 22080 50813 22083
rect 50764 22052 50813 22080
rect 50764 22040 50770 22052
rect 50801 22049 50813 22052
rect 50847 22049 50859 22083
rect 50801 22043 50859 22049
rect 43349 22015 43407 22021
rect 43349 22012 43361 22015
rect 42168 21984 43361 22012
rect 43349 21981 43361 21984
rect 43395 21981 43407 22015
rect 46290 22012 46296 22024
rect 43349 21975 43407 21981
rect 45940 21984 46296 22012
rect 39393 21879 39451 21885
rect 39393 21876 39405 21879
rect 38252 21848 39405 21876
rect 38252 21836 38258 21848
rect 39393 21845 39405 21848
rect 39439 21845 39451 21879
rect 39393 21839 39451 21845
rect 41141 21879 41199 21885
rect 41141 21845 41153 21879
rect 41187 21876 41199 21879
rect 41322 21876 41328 21888
rect 41187 21848 41328 21876
rect 41187 21845 41199 21848
rect 41141 21839 41199 21845
rect 41322 21836 41328 21848
rect 41380 21836 41386 21888
rect 42610 21876 42616 21888
rect 42571 21848 42616 21876
rect 42610 21836 42616 21848
rect 42668 21836 42674 21888
rect 45370 21836 45376 21888
rect 45428 21876 45434 21888
rect 45940 21885 45968 21984
rect 46290 21972 46296 21984
rect 46348 21972 46354 22024
rect 47670 22012 47676 22024
rect 47631 21984 47676 22012
rect 47670 21972 47676 21984
rect 47728 21972 47734 22024
rect 51736 22012 51764 22108
rect 51920 22080 51948 22179
rect 52089 22083 52147 22089
rect 52089 22080 52101 22083
rect 51920 22052 52101 22080
rect 52089 22049 52101 22052
rect 52135 22049 52147 22083
rect 52089 22043 52147 22049
rect 52273 22083 52331 22089
rect 52273 22049 52285 22083
rect 52319 22049 52331 22083
rect 52273 22043 52331 22049
rect 52365 22083 52423 22089
rect 52365 22049 52377 22083
rect 52411 22049 52423 22083
rect 52365 22043 52423 22049
rect 52288 22012 52316 22043
rect 51736 21984 52316 22012
rect 52270 21904 52276 21956
rect 52328 21944 52334 21956
rect 52380 21944 52408 22043
rect 52917 21947 52975 21953
rect 52917 21944 52929 21947
rect 52328 21916 52929 21944
rect 52328 21904 52334 21916
rect 52917 21913 52929 21916
rect 52963 21913 52975 21947
rect 52917 21907 52975 21913
rect 45925 21879 45983 21885
rect 45925 21876 45937 21879
rect 45428 21848 45937 21876
rect 45428 21836 45434 21848
rect 45925 21845 45937 21848
rect 45971 21845 45983 21879
rect 46106 21876 46112 21888
rect 46067 21848 46112 21876
rect 45925 21839 45983 21845
rect 46106 21836 46112 21848
rect 46164 21836 46170 21888
rect 51077 21879 51135 21885
rect 51077 21845 51089 21879
rect 51123 21876 51135 21879
rect 51994 21876 52000 21888
rect 51123 21848 52000 21876
rect 51123 21845 51135 21848
rect 51077 21839 51135 21845
rect 51994 21836 52000 21848
rect 52052 21836 52058 21888
rect 52454 21836 52460 21888
rect 52512 21876 52518 21888
rect 52549 21879 52607 21885
rect 52549 21876 52561 21879
rect 52512 21848 52561 21876
rect 52512 21836 52518 21848
rect 52549 21845 52561 21848
rect 52595 21845 52607 21879
rect 52549 21839 52607 21845
rect 1104 21786 54832 21808
rect 1104 21734 9947 21786
rect 9999 21734 10011 21786
rect 10063 21734 10075 21786
rect 10127 21734 10139 21786
rect 10191 21734 27878 21786
rect 27930 21734 27942 21786
rect 27994 21734 28006 21786
rect 28058 21734 28070 21786
rect 28122 21734 45808 21786
rect 45860 21734 45872 21786
rect 45924 21734 45936 21786
rect 45988 21734 46000 21786
rect 46052 21734 54832 21786
rect 1104 21712 54832 21734
rect 5810 21672 5816 21684
rect 5771 21644 5816 21672
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 6822 21632 6828 21684
rect 6880 21672 6886 21684
rect 9677 21675 9735 21681
rect 9677 21672 9689 21675
rect 6880 21644 9689 21672
rect 6880 21632 6886 21644
rect 9677 21641 9689 21644
rect 9723 21641 9735 21675
rect 9677 21635 9735 21641
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 12713 21675 12771 21681
rect 12713 21672 12725 21675
rect 10652 21644 12725 21672
rect 10652 21632 10658 21644
rect 12713 21641 12725 21644
rect 12759 21641 12771 21675
rect 14826 21672 14832 21684
rect 14787 21644 14832 21672
rect 12713 21635 12771 21641
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 17034 21672 17040 21684
rect 15028 21644 17040 21672
rect 7098 21604 7104 21616
rect 7059 21576 7104 21604
rect 7098 21564 7104 21576
rect 7156 21564 7162 21616
rect 10962 21604 10968 21616
rect 7760 21576 10968 21604
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 3326 21536 3332 21548
rect 2179 21508 3332 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 3326 21496 3332 21508
rect 3384 21536 3390 21548
rect 3881 21539 3939 21545
rect 3881 21536 3893 21539
rect 3384 21508 3893 21536
rect 3384 21496 3390 21508
rect 3881 21505 3893 21508
rect 3927 21505 3939 21539
rect 6914 21536 6920 21548
rect 3881 21499 3939 21505
rect 5736 21508 6920 21536
rect 2409 21471 2467 21477
rect 2409 21437 2421 21471
rect 2455 21468 2467 21471
rect 5626 21468 5632 21480
rect 2455 21440 5632 21468
rect 2455 21437 2467 21440
rect 2409 21431 2467 21437
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 5736 21477 5764 21508
rect 6914 21496 6920 21508
rect 6972 21536 6978 21548
rect 7760 21545 7788 21576
rect 10962 21564 10968 21576
rect 11020 21564 11026 21616
rect 11149 21607 11207 21613
rect 11149 21573 11161 21607
rect 11195 21604 11207 21607
rect 13173 21607 13231 21613
rect 13173 21604 13185 21607
rect 11195 21576 13185 21604
rect 11195 21573 11207 21576
rect 11149 21567 11207 21573
rect 7745 21539 7803 21545
rect 6972 21508 7328 21536
rect 6972 21496 6978 21508
rect 5721 21471 5779 21477
rect 5721 21437 5733 21471
rect 5767 21437 5779 21471
rect 7006 21468 7012 21480
rect 6967 21440 7012 21468
rect 5721 21431 5779 21437
rect 7006 21428 7012 21440
rect 7064 21428 7070 21480
rect 7300 21477 7328 21508
rect 7745 21505 7757 21539
rect 7791 21505 7803 21539
rect 9398 21536 9404 21548
rect 9359 21508 9404 21536
rect 7745 21499 7803 21505
rect 9398 21496 9404 21508
rect 9456 21496 9462 21548
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 12250 21536 12256 21548
rect 9640 21508 12256 21536
rect 9640 21496 9646 21508
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 7285 21471 7343 21477
rect 7285 21437 7297 21471
rect 7331 21468 7343 21471
rect 7466 21468 7472 21480
rect 7331 21440 7472 21468
rect 7331 21437 7343 21440
rect 7285 21431 7343 21437
rect 7466 21428 7472 21440
rect 7524 21428 7530 21480
rect 9493 21471 9551 21477
rect 9493 21437 9505 21471
rect 9539 21468 9551 21471
rect 10045 21471 10103 21477
rect 10045 21468 10057 21471
rect 9539 21440 10057 21468
rect 9539 21437 9551 21440
rect 9493 21431 9551 21437
rect 10045 21437 10057 21440
rect 10091 21468 10103 21471
rect 10091 21440 10916 21468
rect 10091 21437 10103 21440
rect 10045 21431 10103 21437
rect 4614 21360 4620 21412
rect 4672 21400 4678 21412
rect 10318 21400 10324 21412
rect 4672 21372 10324 21400
rect 4672 21360 4678 21372
rect 10318 21360 10324 21372
rect 10376 21360 10382 21412
rect 3697 21335 3755 21341
rect 3697 21301 3709 21335
rect 3743 21332 3755 21335
rect 5718 21332 5724 21344
rect 3743 21304 5724 21332
rect 3743 21301 3755 21304
rect 3697 21295 3755 21301
rect 5718 21292 5724 21304
rect 5776 21292 5782 21344
rect 10888 21332 10916 21440
rect 10962 21428 10968 21480
rect 11020 21468 11026 21480
rect 11057 21471 11115 21477
rect 11057 21468 11069 21471
rect 11020 21440 11069 21468
rect 11020 21428 11026 21440
rect 11057 21437 11069 21440
rect 11103 21437 11115 21471
rect 11057 21431 11115 21437
rect 12342 21428 12348 21480
rect 12400 21468 12406 21480
rect 12544 21477 12572 21576
rect 13173 21573 13185 21576
rect 13219 21604 13231 21607
rect 15028 21604 15056 21644
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 17126 21632 17132 21684
rect 17184 21672 17190 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 17184 21644 17693 21672
rect 17184 21632 17190 21644
rect 17681 21641 17693 21644
rect 17727 21672 17739 21675
rect 19153 21675 19211 21681
rect 19153 21672 19165 21675
rect 17727 21644 19165 21672
rect 17727 21641 17739 21644
rect 17681 21635 17739 21641
rect 19153 21641 19165 21644
rect 19199 21672 19211 21675
rect 19245 21675 19303 21681
rect 19245 21672 19257 21675
rect 19199 21644 19257 21672
rect 19199 21641 19211 21644
rect 19153 21635 19211 21641
rect 19245 21641 19257 21644
rect 19291 21641 19303 21675
rect 20990 21672 20996 21684
rect 20951 21644 20996 21672
rect 19245 21635 19303 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 22370 21672 22376 21684
rect 22331 21644 22376 21672
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 28258 21632 28264 21684
rect 28316 21672 28322 21684
rect 46106 21672 46112 21684
rect 28316 21644 46112 21672
rect 28316 21632 28322 21644
rect 46106 21632 46112 21644
rect 46164 21632 46170 21684
rect 46290 21632 46296 21684
rect 46348 21672 46354 21684
rect 46477 21675 46535 21681
rect 46477 21672 46489 21675
rect 46348 21644 46489 21672
rect 46348 21632 46354 21644
rect 46477 21641 46489 21644
rect 46523 21672 46535 21675
rect 46569 21675 46627 21681
rect 46569 21672 46581 21675
rect 46523 21644 46581 21672
rect 46523 21641 46535 21644
rect 46477 21635 46535 21641
rect 46569 21641 46581 21644
rect 46615 21641 46627 21675
rect 46569 21635 46627 21641
rect 48590 21632 48596 21684
rect 48648 21672 48654 21684
rect 51445 21675 51503 21681
rect 51445 21672 51457 21675
rect 48648 21644 51457 21672
rect 48648 21632 48654 21644
rect 51445 21641 51457 21644
rect 51491 21641 51503 21675
rect 51445 21635 51503 21641
rect 13219 21576 15056 21604
rect 15289 21607 15347 21613
rect 13219 21573 13231 21576
rect 13173 21567 13231 21573
rect 15289 21573 15301 21607
rect 15335 21604 15347 21607
rect 17402 21604 17408 21616
rect 15335 21576 17408 21604
rect 15335 21573 15347 21576
rect 15289 21567 15347 21573
rect 17402 21564 17408 21576
rect 17460 21564 17466 21616
rect 22554 21564 22560 21616
rect 22612 21604 22618 21616
rect 22612 21576 24164 21604
rect 22612 21564 22618 21576
rect 12710 21496 12716 21548
rect 12768 21536 12774 21548
rect 23753 21539 23811 21545
rect 12768 21508 23520 21536
rect 12768 21496 12774 21508
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 12400 21440 12449 21468
rect 12400 21428 12406 21440
rect 12437 21437 12449 21440
rect 12483 21437 12495 21471
rect 12544 21471 12607 21477
rect 12544 21440 12561 21471
rect 12437 21431 12495 21437
rect 12549 21437 12561 21440
rect 12595 21437 12607 21471
rect 13814 21468 13820 21480
rect 13775 21440 13820 21468
rect 12549 21431 12607 21437
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 14826 21428 14832 21480
rect 14884 21468 14890 21480
rect 15013 21471 15071 21477
rect 15013 21468 15025 21471
rect 14884 21440 15025 21468
rect 14884 21428 14890 21440
rect 15013 21437 15025 21440
rect 15059 21437 15071 21471
rect 15562 21468 15568 21480
rect 15523 21440 15568 21468
rect 15013 21431 15071 21437
rect 15562 21428 15568 21440
rect 15620 21428 15626 21480
rect 16022 21468 16028 21480
rect 15983 21440 16028 21468
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 17126 21428 17132 21480
rect 17184 21468 17190 21480
rect 17865 21471 17923 21477
rect 17865 21468 17877 21471
rect 17184 21440 17877 21468
rect 17184 21428 17190 21440
rect 17865 21437 17877 21440
rect 17911 21437 17923 21471
rect 17865 21431 17923 21437
rect 19153 21471 19211 21477
rect 19153 21437 19165 21471
rect 19199 21468 19211 21471
rect 19426 21468 19432 21480
rect 19199 21440 19432 21468
rect 19199 21437 19211 21440
rect 19153 21431 19211 21437
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21468 19763 21471
rect 19794 21468 19800 21480
rect 19751 21440 19800 21468
rect 19751 21437 19763 21440
rect 19705 21431 19763 21437
rect 19794 21428 19800 21440
rect 19852 21428 19858 21480
rect 22370 21428 22376 21480
rect 22428 21468 22434 21480
rect 22557 21471 22615 21477
rect 22557 21468 22569 21471
rect 22428 21440 22569 21468
rect 22428 21428 22434 21440
rect 22557 21437 22569 21440
rect 22603 21437 22615 21471
rect 23492 21468 23520 21508
rect 23753 21505 23765 21539
rect 23799 21536 23811 21539
rect 23842 21536 23848 21548
rect 23799 21508 23848 21536
rect 23799 21505 23811 21508
rect 23753 21499 23811 21505
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 24136 21545 24164 21576
rect 26786 21564 26792 21616
rect 26844 21564 26850 21616
rect 27706 21604 27712 21616
rect 27667 21576 27712 21604
rect 27706 21564 27712 21576
rect 27764 21564 27770 21616
rect 32766 21604 32772 21616
rect 32727 21576 32772 21604
rect 32766 21564 32772 21576
rect 32824 21564 32830 21616
rect 33873 21607 33931 21613
rect 33873 21573 33885 21607
rect 33919 21604 33931 21607
rect 34882 21604 34888 21616
rect 33919 21576 34888 21604
rect 33919 21573 33931 21576
rect 33873 21567 33931 21573
rect 34882 21564 34888 21576
rect 34940 21564 34946 21616
rect 41046 21604 41052 21616
rect 36556 21576 41052 21604
rect 24121 21539 24179 21545
rect 24121 21505 24133 21539
rect 24167 21505 24179 21539
rect 24121 21499 24179 21505
rect 26697 21539 26755 21545
rect 26697 21505 26709 21539
rect 26743 21536 26755 21539
rect 26804 21536 26832 21564
rect 26743 21508 26832 21536
rect 26743 21505 26755 21508
rect 26697 21499 26755 21505
rect 27798 21496 27804 21548
rect 27856 21536 27862 21548
rect 36556 21536 36584 21576
rect 41046 21564 41052 21576
rect 41104 21564 41110 21616
rect 38286 21536 38292 21548
rect 27856 21508 36584 21536
rect 38247 21508 38292 21536
rect 27856 21496 27862 21508
rect 38286 21496 38292 21508
rect 38344 21496 38350 21548
rect 39485 21539 39543 21545
rect 39485 21505 39497 21539
rect 39531 21536 39543 21539
rect 39850 21536 39856 21548
rect 39531 21508 39856 21536
rect 39531 21505 39543 21508
rect 39485 21499 39543 21505
rect 39850 21496 39856 21508
rect 39908 21496 39914 21548
rect 43530 21536 43536 21548
rect 43491 21508 43536 21536
rect 43530 21496 43536 21508
rect 43588 21496 43594 21548
rect 51460 21536 51488 21635
rect 51718 21536 51724 21548
rect 51460 21508 51724 21536
rect 51718 21496 51724 21508
rect 51776 21496 51782 21548
rect 51994 21536 52000 21548
rect 51955 21508 52000 21536
rect 51994 21496 52000 21508
rect 52052 21496 52058 21548
rect 52086 21496 52092 21548
rect 52144 21536 52150 21548
rect 53101 21539 53159 21545
rect 53101 21536 53113 21539
rect 52144 21508 53113 21536
rect 52144 21496 52150 21508
rect 53101 21505 53113 21508
rect 53147 21505 53159 21539
rect 53101 21499 53159 21505
rect 23566 21468 23572 21480
rect 23492 21440 23572 21468
rect 22557 21431 22615 21437
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 23658 21428 23664 21480
rect 23716 21468 23722 21480
rect 23937 21471 23995 21477
rect 23716 21440 23761 21468
rect 23716 21428 23722 21440
rect 23937 21437 23949 21471
rect 23983 21437 23995 21471
rect 25222 21468 25228 21480
rect 25183 21440 25228 21468
rect 23937 21431 23995 21437
rect 12710 21360 12716 21412
rect 12768 21400 12774 21412
rect 13909 21403 13967 21409
rect 13909 21400 13921 21403
rect 12768 21372 13921 21400
rect 12768 21360 12774 21372
rect 13909 21369 13921 21372
rect 13955 21400 13967 21403
rect 18598 21400 18604 21412
rect 13955 21372 18604 21400
rect 13955 21369 13967 21372
rect 13909 21363 13967 21369
rect 18598 21360 18604 21372
rect 18656 21360 18662 21412
rect 22649 21403 22707 21409
rect 22649 21369 22661 21403
rect 22695 21400 22707 21403
rect 23952 21400 23980 21431
rect 25222 21428 25228 21440
rect 25280 21428 25286 21480
rect 26418 21428 26424 21480
rect 26476 21468 26482 21480
rect 26789 21471 26847 21477
rect 26789 21468 26801 21471
rect 26476 21440 26801 21468
rect 26476 21428 26482 21440
rect 26789 21437 26801 21440
rect 26835 21468 26847 21471
rect 27154 21468 27160 21480
rect 26835 21440 27160 21468
rect 26835 21437 26847 21440
rect 26789 21431 26847 21437
rect 27154 21428 27160 21440
rect 27212 21468 27218 21480
rect 27341 21471 27399 21477
rect 27341 21468 27353 21471
rect 27212 21440 27353 21468
rect 27212 21428 27218 21440
rect 27341 21437 27353 21440
rect 27387 21437 27399 21471
rect 27341 21431 27399 21437
rect 27525 21471 27583 21477
rect 27525 21437 27537 21471
rect 27571 21468 27583 21471
rect 28810 21468 28816 21480
rect 27571 21440 28816 21468
rect 27571 21437 27583 21440
rect 27525 21431 27583 21437
rect 28810 21428 28816 21440
rect 28868 21428 28874 21480
rect 29730 21468 29736 21480
rect 29691 21440 29736 21468
rect 29730 21428 29736 21440
rect 29788 21428 29794 21480
rect 31018 21468 31024 21480
rect 30979 21440 31024 21468
rect 31018 21428 31024 21440
rect 31076 21428 31082 21480
rect 31110 21428 31116 21480
rect 31168 21468 31174 21480
rect 31297 21471 31355 21477
rect 31297 21468 31309 21471
rect 31168 21440 31309 21468
rect 31168 21428 31174 21440
rect 31297 21437 31309 21440
rect 31343 21437 31355 21471
rect 33778 21468 33784 21480
rect 33691 21440 33784 21468
rect 31297 21431 31355 21437
rect 33778 21428 33784 21440
rect 33836 21428 33842 21480
rect 35342 21468 35348 21480
rect 35303 21440 35348 21468
rect 35342 21428 35348 21440
rect 35400 21428 35406 21480
rect 35618 21468 35624 21480
rect 35579 21440 35624 21468
rect 35618 21428 35624 21440
rect 35676 21428 35682 21480
rect 35986 21428 35992 21480
rect 36044 21468 36050 21480
rect 37093 21471 37151 21477
rect 37093 21468 37105 21471
rect 36044 21440 37105 21468
rect 36044 21428 36050 21440
rect 37093 21437 37105 21440
rect 37139 21468 37151 21471
rect 38194 21468 38200 21480
rect 37139 21440 38200 21468
rect 37139 21437 37151 21440
rect 37093 21431 37151 21437
rect 38194 21428 38200 21440
rect 38252 21428 38258 21480
rect 38378 21468 38384 21480
rect 38291 21440 38384 21468
rect 38378 21428 38384 21440
rect 38436 21428 38442 21480
rect 38746 21428 38752 21480
rect 38804 21468 38810 21480
rect 38841 21471 38899 21477
rect 38841 21468 38853 21471
rect 38804 21440 38853 21468
rect 38804 21428 38810 21440
rect 38841 21437 38853 21440
rect 38887 21437 38899 21471
rect 38841 21431 38899 21437
rect 38933 21471 38991 21477
rect 38933 21437 38945 21471
rect 38979 21437 38991 21471
rect 38933 21431 38991 21437
rect 40773 21471 40831 21477
rect 40773 21437 40785 21471
rect 40819 21468 40831 21471
rect 40865 21471 40923 21477
rect 40865 21468 40877 21471
rect 40819 21440 40877 21468
rect 40819 21437 40831 21440
rect 40773 21431 40831 21437
rect 40865 21437 40877 21440
rect 40911 21468 40923 21471
rect 41046 21468 41052 21480
rect 40911 21440 41052 21468
rect 40911 21437 40923 21440
rect 40865 21431 40923 21437
rect 24118 21400 24124 21412
rect 22695 21372 24124 21400
rect 22695 21369 22707 21372
rect 22649 21363 22707 21369
rect 24118 21360 24124 21372
rect 24176 21360 24182 21412
rect 28902 21360 28908 21412
rect 28960 21360 28966 21412
rect 16942 21332 16948 21344
rect 10888 21304 16948 21332
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 22278 21332 22284 21344
rect 17092 21304 22284 21332
rect 17092 21292 17098 21304
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 23474 21332 23480 21344
rect 23435 21304 23480 21332
rect 23474 21292 23480 21304
rect 23532 21332 23538 21344
rect 23842 21332 23848 21344
rect 23532 21304 23848 21332
rect 23532 21292 23538 21304
rect 23842 21292 23848 21304
rect 23900 21292 23906 21344
rect 25222 21292 25228 21344
rect 25280 21332 25286 21344
rect 25409 21335 25467 21341
rect 25409 21332 25421 21335
rect 25280 21304 25421 21332
rect 25280 21292 25286 21304
rect 25409 21301 25421 21304
rect 25455 21332 25467 21335
rect 27798 21332 27804 21344
rect 25455 21304 27804 21332
rect 25455 21301 25467 21304
rect 25409 21295 25467 21301
rect 27798 21292 27804 21304
rect 27856 21292 27862 21344
rect 28920 21332 28948 21360
rect 29825 21335 29883 21341
rect 29825 21332 29837 21335
rect 28920 21304 29837 21332
rect 29825 21301 29837 21304
rect 29871 21301 29883 21335
rect 29825 21295 29883 21301
rect 30742 21292 30748 21344
rect 30800 21332 30806 21344
rect 30926 21332 30932 21344
rect 30800 21304 30932 21332
rect 30800 21292 30806 21304
rect 30926 21292 30932 21304
rect 30984 21332 30990 21344
rect 32401 21335 32459 21341
rect 32401 21332 32413 21335
rect 30984 21304 32413 21332
rect 30984 21292 30990 21304
rect 32401 21301 32413 21304
rect 32447 21301 32459 21335
rect 33796 21332 33824 21428
rect 37001 21403 37059 21409
rect 37001 21369 37013 21403
rect 37047 21400 37059 21403
rect 37182 21400 37188 21412
rect 37047 21372 37188 21400
rect 37047 21369 37059 21372
rect 37001 21363 37059 21369
rect 37016 21332 37044 21363
rect 37182 21360 37188 21372
rect 37240 21360 37246 21412
rect 38396 21400 38424 21428
rect 38948 21400 38976 21431
rect 41046 21428 41052 21440
rect 41104 21428 41110 21480
rect 43257 21471 43315 21477
rect 43257 21468 43269 21471
rect 43088 21440 43269 21468
rect 38396 21372 41092 21400
rect 41064 21341 41092 21372
rect 33796 21304 37044 21332
rect 41049 21335 41107 21341
rect 32401 21295 32459 21301
rect 41049 21301 41061 21335
rect 41095 21332 41107 21335
rect 41138 21332 41144 21344
rect 41095 21304 41144 21332
rect 41095 21301 41107 21304
rect 41049 21295 41107 21301
rect 41138 21292 41144 21304
rect 41196 21292 41202 21344
rect 42978 21292 42984 21344
rect 43036 21332 43042 21344
rect 43088 21341 43116 21440
rect 43257 21437 43269 21440
rect 43303 21437 43315 21471
rect 43257 21431 43315 21437
rect 46477 21471 46535 21477
rect 46477 21437 46489 21471
rect 46523 21468 46535 21471
rect 46753 21471 46811 21477
rect 46753 21468 46765 21471
rect 46523 21440 46765 21468
rect 46523 21437 46535 21440
rect 46477 21431 46535 21437
rect 46753 21437 46765 21440
rect 46799 21437 46811 21471
rect 47026 21468 47032 21480
rect 46987 21440 47032 21468
rect 46753 21431 46811 21437
rect 47026 21428 47032 21440
rect 47084 21428 47090 21480
rect 43073 21335 43131 21341
rect 43073 21332 43085 21335
rect 43036 21304 43085 21332
rect 43036 21292 43042 21304
rect 43073 21301 43085 21304
rect 43119 21301 43131 21335
rect 43073 21295 43131 21301
rect 43162 21292 43168 21344
rect 43220 21332 43226 21344
rect 44637 21335 44695 21341
rect 44637 21332 44649 21335
rect 43220 21304 44649 21332
rect 43220 21292 43226 21304
rect 44637 21301 44649 21304
rect 44683 21301 44695 21335
rect 44637 21295 44695 21301
rect 47854 21292 47860 21344
rect 47912 21332 47918 21344
rect 48317 21335 48375 21341
rect 48317 21332 48329 21335
rect 47912 21304 48329 21332
rect 47912 21292 47918 21304
rect 48317 21301 48329 21304
rect 48363 21301 48375 21335
rect 48317 21295 48375 21301
rect 1104 21242 54832 21264
rect 1104 21190 18912 21242
rect 18964 21190 18976 21242
rect 19028 21190 19040 21242
rect 19092 21190 19104 21242
rect 19156 21190 36843 21242
rect 36895 21190 36907 21242
rect 36959 21190 36971 21242
rect 37023 21190 37035 21242
rect 37087 21190 54832 21242
rect 1104 21168 54832 21190
rect 5626 21128 5632 21140
rect 5587 21100 5632 21128
rect 5626 21088 5632 21100
rect 5684 21088 5690 21140
rect 8113 21131 8171 21137
rect 8113 21097 8125 21131
rect 8159 21128 8171 21131
rect 9582 21128 9588 21140
rect 8159 21100 9588 21128
rect 8159 21097 8171 21100
rect 8113 21091 8171 21097
rect 6638 21060 6644 21072
rect 5184 21032 6644 21060
rect 5184 21001 5212 21032
rect 6638 21020 6644 21032
rect 6696 21020 6702 21072
rect 7006 21020 7012 21072
rect 7064 21060 7070 21072
rect 7193 21063 7251 21069
rect 7193 21060 7205 21063
rect 7064 21032 7205 21060
rect 7064 21020 7070 21032
rect 7193 21029 7205 21032
rect 7239 21029 7251 21063
rect 7193 21023 7251 21029
rect 4617 20995 4675 21001
rect 4617 20961 4629 20995
rect 4663 20992 4675 20995
rect 5169 20995 5227 21001
rect 5169 20992 5181 20995
rect 4663 20964 5181 20992
rect 4663 20961 4675 20964
rect 4617 20955 4675 20961
rect 5169 20961 5181 20964
rect 5215 20961 5227 20995
rect 5169 20955 5227 20961
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5810 20992 5816 21004
rect 5399 20964 5816 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 5810 20952 5816 20964
rect 5868 20952 5874 21004
rect 7374 21001 7380 21004
rect 7340 20995 7380 21001
rect 7340 20961 7352 20995
rect 7340 20955 7380 20961
rect 7374 20952 7380 20955
rect 7432 20952 7438 21004
rect 4525 20927 4583 20933
rect 4525 20893 4537 20927
rect 4571 20924 4583 20927
rect 4798 20924 4804 20936
rect 4571 20896 4804 20924
rect 4571 20893 4583 20896
rect 4525 20887 4583 20893
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 7561 20927 7619 20933
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 8128 20924 8156 21091
rect 9582 21088 9588 21100
rect 9640 21088 9646 21140
rect 12342 21088 12348 21140
rect 12400 21128 12406 21140
rect 13725 21131 13783 21137
rect 13725 21128 13737 21131
rect 12400 21100 13737 21128
rect 12400 21088 12406 21100
rect 13725 21097 13737 21100
rect 13771 21128 13783 21131
rect 13814 21128 13820 21140
rect 13771 21100 13820 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 14185 21131 14243 21137
rect 14185 21097 14197 21131
rect 14231 21128 14243 21131
rect 14829 21131 14887 21137
rect 14829 21128 14841 21131
rect 14231 21100 14841 21128
rect 14231 21097 14243 21100
rect 14185 21091 14243 21097
rect 14829 21097 14841 21100
rect 14875 21128 14887 21131
rect 15102 21128 15108 21140
rect 14875 21100 15108 21128
rect 14875 21097 14887 21100
rect 14829 21091 14887 21097
rect 10229 21063 10287 21069
rect 10229 21029 10241 21063
rect 10275 21060 10287 21063
rect 10870 21060 10876 21072
rect 10275 21032 10876 21060
rect 10275 21029 10287 21032
rect 10229 21023 10287 21029
rect 10870 21020 10876 21032
rect 10928 21020 10934 21072
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 9769 20995 9827 21001
rect 9769 20992 9781 20995
rect 9456 20964 9781 20992
rect 9456 20952 9462 20964
rect 9769 20961 9781 20964
rect 9815 20961 9827 20995
rect 9769 20955 9827 20961
rect 10962 20952 10968 21004
rect 11020 20992 11026 21004
rect 11057 20995 11115 21001
rect 11057 20992 11069 20995
rect 11020 20964 11069 20992
rect 11020 20952 11026 20964
rect 11057 20961 11069 20964
rect 11103 20961 11115 20995
rect 11057 20955 11115 20961
rect 12345 20995 12403 21001
rect 12345 20961 12357 20995
rect 12391 20992 12403 20995
rect 13262 20992 13268 21004
rect 12391 20964 13268 20992
rect 12391 20961 12403 20964
rect 12345 20955 12403 20961
rect 13262 20952 13268 20964
rect 13320 20992 13326 21004
rect 14200 20992 14228 21091
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 16117 21131 16175 21137
rect 16117 21128 16129 21131
rect 16080 21100 16129 21128
rect 16080 21088 16086 21100
rect 16117 21097 16129 21100
rect 16163 21097 16175 21131
rect 17034 21128 17040 21140
rect 16995 21100 17040 21128
rect 16117 21091 16175 21097
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 19794 21128 19800 21140
rect 19755 21100 19800 21128
rect 19794 21088 19800 21100
rect 19852 21088 19858 21140
rect 20165 21131 20223 21137
rect 20165 21097 20177 21131
rect 20211 21128 20223 21131
rect 20993 21131 21051 21137
rect 20993 21128 21005 21131
rect 20211 21100 21005 21128
rect 20211 21097 20223 21100
rect 20165 21091 20223 21097
rect 20993 21097 21005 21100
rect 21039 21128 21051 21131
rect 25682 21128 25688 21140
rect 21039 21100 25688 21128
rect 21039 21097 21051 21100
rect 20993 21091 21051 21097
rect 17126 21060 17132 21072
rect 15028 21032 17132 21060
rect 15028 21001 15056 21032
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 19702 21060 19708 21072
rect 18892 21032 19708 21060
rect 13320 20964 14228 20992
rect 15013 20995 15071 21001
rect 13320 20952 13326 20964
rect 15013 20961 15025 20995
rect 15059 20961 15071 20995
rect 15838 20992 15844 21004
rect 15799 20964 15844 20992
rect 15013 20955 15071 20961
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 16025 20995 16083 21001
rect 16025 20961 16037 20995
rect 16071 20992 16083 20995
rect 16071 20964 16620 20992
rect 16071 20961 16083 20964
rect 16025 20955 16083 20961
rect 7607 20896 8156 20924
rect 9677 20927 9735 20933
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 12618 20924 12624 20936
rect 12579 20896 12624 20924
rect 9677 20887 9735 20893
rect 7466 20856 7472 20868
rect 7427 20828 7472 20856
rect 7466 20816 7472 20828
rect 7524 20816 7530 20868
rect 7926 20816 7932 20868
rect 7984 20856 7990 20868
rect 9692 20856 9720 20887
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 16592 20865 16620 20964
rect 16942 20952 16948 21004
rect 17000 20992 17006 21004
rect 17313 20995 17371 21001
rect 17313 20992 17325 20995
rect 17000 20964 17325 20992
rect 17000 20952 17006 20964
rect 17313 20961 17325 20964
rect 17359 20992 17371 20995
rect 17865 20995 17923 21001
rect 17865 20992 17877 20995
rect 17359 20964 17877 20992
rect 17359 20961 17371 20964
rect 17313 20955 17371 20961
rect 17865 20961 17877 20964
rect 17911 20992 17923 20995
rect 18046 20992 18052 21004
rect 17911 20964 18052 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 18506 20952 18512 21004
rect 18564 20992 18570 21004
rect 18892 21001 18920 21032
rect 19702 21020 19708 21032
rect 19760 21020 19766 21072
rect 18785 20995 18843 21001
rect 18785 20992 18797 20995
rect 18564 20964 18797 20992
rect 18564 20952 18570 20964
rect 18785 20961 18797 20964
rect 18831 20961 18843 20995
rect 18785 20955 18843 20961
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20961 18935 20995
rect 19337 20995 19395 21001
rect 19337 20992 19349 20995
rect 18877 20955 18935 20961
rect 18984 20964 19349 20992
rect 17034 20884 17040 20936
rect 17092 20924 17098 20936
rect 17221 20927 17279 20933
rect 17221 20924 17233 20927
rect 17092 20896 17233 20924
rect 17092 20884 17098 20896
rect 17221 20893 17233 20896
rect 17267 20893 17279 20927
rect 18800 20924 18828 20955
rect 18984 20924 19012 20964
rect 19337 20961 19349 20964
rect 19383 20961 19395 20995
rect 19337 20955 19395 20961
rect 19521 20995 19579 21001
rect 19521 20961 19533 20995
rect 19567 20992 19579 20995
rect 20180 20992 20208 21091
rect 25682 21088 25688 21100
rect 25740 21088 25746 21140
rect 25792 21100 31708 21128
rect 21542 21020 21548 21072
rect 21600 21060 21606 21072
rect 22281 21063 22339 21069
rect 22281 21060 22293 21063
rect 21600 21032 22293 21060
rect 21600 21020 21606 21032
rect 22281 21029 22293 21032
rect 22327 21060 22339 21063
rect 22327 21032 22508 21060
rect 22327 21029 22339 21032
rect 22281 21023 22339 21029
rect 19567 20964 20208 20992
rect 20901 20995 20959 21001
rect 19567 20961 19579 20964
rect 19521 20955 19579 20961
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 20990 20992 20996 21004
rect 20947 20964 20996 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 20990 20952 20996 20964
rect 21048 20952 21054 21004
rect 22480 21001 22508 21032
rect 23750 21020 23756 21072
rect 23808 21060 23814 21072
rect 24121 21063 24179 21069
rect 24121 21060 24133 21063
rect 23808 21032 24133 21060
rect 23808 21020 23814 21032
rect 24121 21029 24133 21032
rect 24167 21060 24179 21063
rect 24762 21060 24768 21072
rect 24167 21032 24768 21060
rect 24167 21029 24179 21032
rect 24121 21023 24179 21029
rect 24762 21020 24768 21032
rect 24820 21020 24826 21072
rect 22465 20995 22523 21001
rect 22465 20961 22477 20995
rect 22511 20961 22523 20995
rect 22738 20992 22744 21004
rect 22699 20964 22744 20992
rect 22465 20955 22523 20961
rect 22738 20952 22744 20964
rect 22796 20952 22802 21004
rect 24780 20992 24808 21020
rect 24949 20995 25007 21001
rect 24949 20992 24961 20995
rect 24780 20964 24961 20992
rect 24949 20961 24961 20964
rect 24995 20961 25007 20995
rect 24949 20955 25007 20961
rect 25792 20924 25820 21100
rect 26786 21020 26792 21072
rect 26844 21060 26850 21072
rect 26844 21032 27200 21060
rect 26844 21020 26850 21032
rect 26878 20952 26884 21004
rect 26936 20992 26942 21004
rect 26936 20964 27016 20992
rect 26936 20952 26942 20964
rect 18800 20896 19012 20924
rect 22480 20896 25820 20924
rect 26988 20924 27016 20964
rect 27065 20927 27123 20933
rect 27065 20924 27077 20927
rect 26988 20896 27077 20924
rect 17221 20887 17279 20893
rect 7984 20828 9720 20856
rect 16577 20859 16635 20865
rect 7984 20816 7990 20828
rect 16577 20825 16589 20859
rect 16623 20856 16635 20859
rect 17770 20856 17776 20868
rect 16623 20828 17776 20856
rect 16623 20825 16635 20828
rect 16577 20819 16635 20825
rect 17770 20816 17776 20828
rect 17828 20816 17834 20868
rect 17954 20816 17960 20868
rect 18012 20856 18018 20868
rect 22480 20856 22508 20896
rect 27065 20893 27077 20896
rect 27111 20893 27123 20927
rect 27172 20924 27200 21032
rect 28718 21020 28724 21072
rect 28776 21060 28782 21072
rect 28813 21063 28871 21069
rect 28813 21060 28825 21063
rect 28776 21032 28825 21060
rect 28776 21020 28782 21032
rect 28813 21029 28825 21032
rect 28859 21060 28871 21063
rect 28994 21060 29000 21072
rect 28859 21032 29000 21060
rect 28859 21029 28871 21032
rect 28813 21023 28871 21029
rect 28994 21020 29000 21032
rect 29052 21020 29058 21072
rect 31110 21060 31116 21072
rect 30576 21032 30972 21060
rect 31071 21032 31116 21060
rect 29822 20992 29828 21004
rect 29783 20964 29828 20992
rect 29822 20952 29828 20964
rect 29880 20952 29886 21004
rect 30009 20995 30067 21001
rect 30009 20961 30021 20995
rect 30055 20992 30067 20995
rect 30190 20992 30196 21004
rect 30055 20964 30196 20992
rect 30055 20961 30067 20964
rect 30009 20955 30067 20961
rect 30190 20952 30196 20964
rect 30248 20992 30254 21004
rect 30576 21001 30604 21032
rect 30561 20995 30619 21001
rect 30561 20992 30573 20995
rect 30248 20964 30573 20992
rect 30248 20952 30254 20964
rect 30561 20961 30573 20964
rect 30607 20961 30619 20995
rect 30742 20992 30748 21004
rect 30703 20964 30748 20992
rect 30561 20955 30619 20961
rect 30742 20952 30748 20964
rect 30800 20952 30806 21004
rect 27341 20927 27399 20933
rect 27341 20924 27353 20927
rect 27172 20896 27353 20924
rect 27065 20887 27123 20893
rect 27341 20893 27353 20896
rect 27387 20893 27399 20927
rect 30944 20924 30972 21032
rect 31110 21020 31116 21032
rect 31168 21020 31174 21072
rect 31680 20992 31708 21100
rect 35342 21088 35348 21140
rect 35400 21128 35406 21140
rect 35986 21128 35992 21140
rect 35400 21100 35992 21128
rect 35400 21088 35406 21100
rect 35986 21088 35992 21100
rect 36044 21088 36050 21140
rect 36446 21128 36452 21140
rect 36096 21100 36452 21128
rect 34790 21060 34796 21072
rect 31864 21032 34796 21060
rect 31864 20992 31892 21032
rect 33226 20992 33232 21004
rect 31680 20964 31892 20992
rect 33187 20964 33232 20992
rect 33226 20952 33232 20964
rect 33284 20952 33290 21004
rect 33888 21001 33916 21032
rect 34790 21020 34796 21032
rect 34848 21020 34854 21072
rect 33413 20995 33471 21001
rect 33413 20961 33425 20995
rect 33459 20961 33471 20995
rect 33413 20955 33471 20961
rect 33873 20995 33931 21001
rect 33873 20961 33885 20995
rect 33919 20961 33931 20995
rect 33873 20955 33931 20961
rect 33965 20995 34023 21001
rect 33965 20961 33977 20995
rect 34011 20992 34023 20995
rect 34146 20992 34152 21004
rect 34011 20964 34152 20992
rect 34011 20961 34023 20964
rect 33965 20955 34023 20961
rect 32030 20924 32036 20936
rect 30944 20896 32036 20924
rect 27341 20887 27399 20893
rect 32030 20884 32036 20896
rect 32088 20924 32094 20936
rect 33428 20924 33456 20955
rect 34146 20952 34152 20964
rect 34204 20992 34210 21004
rect 36096 20992 36124 21100
rect 36446 21088 36452 21100
rect 36504 21088 36510 21140
rect 40218 21128 40224 21140
rect 40179 21100 40224 21128
rect 40218 21088 40224 21100
rect 40276 21128 40282 21140
rect 41690 21128 41696 21140
rect 40276 21100 41696 21128
rect 40276 21088 40282 21100
rect 41690 21088 41696 21100
rect 41748 21088 41754 21140
rect 41877 21131 41935 21137
rect 41877 21097 41889 21131
rect 41923 21128 41935 21131
rect 42794 21128 42800 21140
rect 41923 21100 42800 21128
rect 41923 21097 41935 21100
rect 41877 21091 41935 21097
rect 42794 21088 42800 21100
rect 42852 21088 42858 21140
rect 42978 21088 42984 21140
rect 43036 21128 43042 21140
rect 45370 21128 45376 21140
rect 43036 21100 45376 21128
rect 43036 21088 43042 21100
rect 45370 21088 45376 21100
rect 45428 21128 45434 21140
rect 45646 21128 45652 21140
rect 45428 21100 45652 21128
rect 45428 21088 45434 21100
rect 45646 21088 45652 21100
rect 45704 21088 45710 21140
rect 46934 21128 46940 21140
rect 46032 21100 46940 21128
rect 40034 21020 40040 21072
rect 40092 21060 40098 21072
rect 40770 21060 40776 21072
rect 40092 21032 40776 21060
rect 40092 21020 40098 21032
rect 40770 21020 40776 21032
rect 40828 21060 40834 21072
rect 43162 21060 43168 21072
rect 40828 21032 43168 21060
rect 40828 21020 40834 21032
rect 43162 21020 43168 21032
rect 43220 21020 43226 21072
rect 34204 20964 36124 20992
rect 36165 20995 36223 21001
rect 34204 20952 34210 20964
rect 36165 20961 36177 20995
rect 36211 20961 36223 20995
rect 36165 20955 36223 20961
rect 36265 20995 36323 21001
rect 36265 20961 36277 20995
rect 36311 20961 36323 20995
rect 41509 20995 41567 21001
rect 41509 20992 41521 20995
rect 36265 20955 36323 20961
rect 36648 20964 41521 20992
rect 34790 20924 34796 20936
rect 32088 20896 33456 20924
rect 34751 20896 34796 20924
rect 32088 20884 32094 20896
rect 34790 20884 34796 20896
rect 34848 20884 34854 20936
rect 36188 20868 36216 20955
rect 36280 20924 36308 20955
rect 36648 20933 36676 20964
rect 41509 20961 41521 20964
rect 41555 20992 41567 20995
rect 41693 20995 41751 21001
rect 41693 20992 41705 20995
rect 41555 20964 41705 20992
rect 41555 20961 41567 20964
rect 41509 20955 41567 20961
rect 41693 20961 41705 20964
rect 41739 20961 41751 20995
rect 41693 20955 41751 20961
rect 44450 20952 44456 21004
rect 44508 20992 44514 21004
rect 44637 20995 44695 21001
rect 44637 20992 44649 20995
rect 44508 20964 44649 20992
rect 44508 20952 44514 20964
rect 44637 20961 44649 20964
rect 44683 20961 44695 20995
rect 45922 20992 45928 21004
rect 45883 20964 45928 20992
rect 44637 20955 44695 20961
rect 45922 20952 45928 20964
rect 45980 20952 45986 21004
rect 46032 21001 46060 21100
rect 46934 21088 46940 21100
rect 46992 21088 46998 21140
rect 51718 21088 51724 21140
rect 51776 21128 51782 21140
rect 51813 21131 51871 21137
rect 51813 21128 51825 21131
rect 51776 21100 51825 21128
rect 51776 21088 51782 21100
rect 51813 21097 51825 21100
rect 51859 21097 51871 21131
rect 51813 21091 51871 21097
rect 47026 21060 47032 21072
rect 46492 21032 46888 21060
rect 46987 21032 47032 21060
rect 46492 21001 46520 21032
rect 46017 20995 46075 21001
rect 46017 20961 46029 20995
rect 46063 20961 46075 20995
rect 46477 20995 46535 21001
rect 46477 20992 46489 20995
rect 46017 20955 46075 20961
rect 46124 20964 46489 20992
rect 36633 20927 36691 20933
rect 36633 20924 36645 20927
rect 36280 20896 36645 20924
rect 18012 20828 22508 20856
rect 18012 20816 18018 20828
rect 23566 20816 23572 20868
rect 23624 20856 23630 20868
rect 24946 20856 24952 20868
rect 23624 20828 24952 20856
rect 23624 20816 23630 20828
rect 24946 20816 24952 20828
rect 25004 20856 25010 20868
rect 25041 20859 25099 20865
rect 25041 20856 25053 20859
rect 25004 20828 25053 20856
rect 25004 20816 25010 20828
rect 25041 20825 25053 20828
rect 25087 20825 25099 20859
rect 25041 20819 25099 20825
rect 28000 20828 36124 20856
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 11146 20788 11152 20800
rect 7883 20760 11152 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 11146 20748 11152 20760
rect 11204 20748 11210 20800
rect 11241 20791 11299 20797
rect 11241 20757 11253 20791
rect 11287 20788 11299 20791
rect 11330 20788 11336 20800
rect 11287 20760 11336 20788
rect 11287 20757 11299 20760
rect 11241 20751 11299 20757
rect 11330 20748 11336 20760
rect 11388 20748 11394 20800
rect 17494 20788 17500 20800
rect 17455 20760 17500 20788
rect 17494 20748 17500 20760
rect 17552 20748 17558 20800
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 25222 20788 25228 20800
rect 18104 20760 25228 20788
rect 18104 20748 18110 20760
rect 25222 20748 25228 20760
rect 25280 20748 25286 20800
rect 26694 20748 26700 20800
rect 26752 20788 26758 20800
rect 28000 20788 28028 20828
rect 28626 20788 28632 20800
rect 26752 20760 28028 20788
rect 28587 20760 28632 20788
rect 26752 20748 26758 20760
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 34425 20791 34483 20797
rect 34425 20757 34437 20791
rect 34471 20788 34483 20791
rect 35802 20788 35808 20800
rect 34471 20760 35808 20788
rect 34471 20757 34483 20760
rect 34425 20751 34483 20757
rect 35802 20748 35808 20760
rect 35860 20748 35866 20800
rect 36096 20788 36124 20828
rect 36170 20816 36176 20868
rect 36228 20816 36234 20868
rect 36280 20788 36308 20896
rect 36633 20893 36645 20896
rect 36679 20893 36691 20927
rect 36633 20887 36691 20893
rect 38657 20927 38715 20933
rect 38657 20893 38669 20927
rect 38703 20893 38715 20927
rect 38930 20924 38936 20936
rect 38891 20896 38936 20924
rect 38657 20887 38715 20893
rect 36446 20788 36452 20800
rect 36096 20760 36308 20788
rect 36359 20760 36452 20788
rect 36446 20748 36452 20760
rect 36504 20788 36510 20800
rect 38286 20788 38292 20800
rect 36504 20760 38292 20788
rect 36504 20748 36510 20760
rect 38286 20748 38292 20760
rect 38344 20748 38350 20800
rect 38672 20788 38700 20887
rect 38930 20884 38936 20896
rect 38988 20884 38994 20936
rect 40218 20884 40224 20936
rect 40276 20924 40282 20936
rect 44266 20924 44272 20936
rect 40276 20896 44272 20924
rect 40276 20884 40282 20896
rect 44266 20884 44272 20896
rect 44324 20884 44330 20936
rect 46124 20924 46152 20964
rect 46477 20961 46489 20964
rect 46523 20961 46535 20995
rect 46658 20992 46664 21004
rect 46619 20964 46664 20992
rect 46477 20955 46535 20961
rect 46658 20952 46664 20964
rect 46716 20952 46722 21004
rect 44836 20896 46152 20924
rect 46860 20924 46888 21032
rect 47026 21020 47032 21032
rect 47084 21020 47090 21072
rect 50062 21060 50068 21072
rect 49712 21032 50068 21060
rect 48406 20952 48412 21004
rect 48464 20992 48470 21004
rect 49712 21001 49740 21032
rect 50062 21020 50068 21032
rect 50120 21060 50126 21072
rect 51828 21060 51856 21091
rect 50120 21032 50292 21060
rect 51828 21032 52040 21060
rect 50120 21020 50126 21032
rect 49513 20995 49571 21001
rect 49513 20992 49525 20995
rect 48464 20964 49525 20992
rect 48464 20952 48470 20964
rect 49513 20961 49525 20964
rect 49559 20961 49571 20995
rect 49513 20955 49571 20961
rect 49697 20995 49755 21001
rect 49697 20961 49709 20995
rect 49743 20961 49755 20995
rect 50154 20992 50160 21004
rect 50115 20964 50160 20992
rect 49697 20955 49755 20961
rect 49712 20924 49740 20955
rect 50154 20952 50160 20964
rect 50212 20952 50218 21004
rect 50264 21001 50292 21032
rect 52012 21001 52040 21032
rect 50249 20995 50307 21001
rect 50249 20961 50261 20995
rect 50295 20961 50307 20995
rect 50249 20955 50307 20961
rect 51997 20995 52055 21001
rect 51997 20961 52009 20995
rect 52043 20961 52055 20995
rect 51997 20955 52055 20961
rect 52273 20927 52331 20933
rect 52273 20924 52285 20927
rect 46860 20896 49740 20924
rect 52012 20896 52285 20924
rect 44836 20865 44864 20896
rect 44821 20859 44879 20865
rect 44821 20825 44833 20859
rect 44867 20825 44879 20859
rect 44821 20819 44879 20825
rect 50709 20859 50767 20865
rect 50709 20825 50721 20859
rect 50755 20856 50767 20859
rect 52012 20856 52040 20896
rect 52273 20893 52285 20896
rect 52319 20893 52331 20927
rect 52273 20887 52331 20893
rect 50755 20828 52040 20856
rect 50755 20825 50767 20828
rect 50709 20819 50767 20825
rect 39114 20788 39120 20800
rect 38672 20760 39120 20788
rect 39114 20748 39120 20760
rect 39172 20788 39178 20800
rect 40405 20791 40463 20797
rect 40405 20788 40417 20791
rect 39172 20760 40417 20788
rect 39172 20748 39178 20760
rect 40405 20757 40417 20760
rect 40451 20757 40463 20791
rect 44450 20788 44456 20800
rect 44411 20760 44456 20788
rect 40405 20751 40463 20757
rect 44450 20748 44456 20760
rect 44508 20748 44514 20800
rect 46658 20748 46664 20800
rect 46716 20788 46722 20800
rect 47213 20791 47271 20797
rect 47213 20788 47225 20791
rect 46716 20760 47225 20788
rect 46716 20748 46722 20760
rect 47213 20757 47225 20760
rect 47259 20757 47271 20791
rect 47213 20751 47271 20757
rect 52270 20748 52276 20800
rect 52328 20788 52334 20800
rect 53377 20791 53435 20797
rect 53377 20788 53389 20791
rect 52328 20760 53389 20788
rect 52328 20748 52334 20760
rect 53377 20757 53389 20760
rect 53423 20757 53435 20791
rect 53377 20751 53435 20757
rect 1104 20698 54832 20720
rect 1104 20646 9947 20698
rect 9999 20646 10011 20698
rect 10063 20646 10075 20698
rect 10127 20646 10139 20698
rect 10191 20646 27878 20698
rect 27930 20646 27942 20698
rect 27994 20646 28006 20698
rect 28058 20646 28070 20698
rect 28122 20646 45808 20698
rect 45860 20646 45872 20698
rect 45924 20646 45936 20698
rect 45988 20646 46000 20698
rect 46052 20646 54832 20698
rect 1104 20624 54832 20646
rect 5810 20584 5816 20596
rect 5771 20556 5816 20584
rect 5810 20544 5816 20556
rect 5868 20544 5874 20596
rect 11333 20587 11391 20593
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 12618 20584 12624 20596
rect 11379 20556 12624 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 15102 20584 15108 20596
rect 15063 20556 15108 20584
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 16025 20587 16083 20593
rect 16025 20553 16037 20587
rect 16071 20584 16083 20587
rect 16114 20584 16120 20596
rect 16071 20556 16120 20584
rect 16071 20553 16083 20556
rect 16025 20547 16083 20553
rect 16114 20544 16120 20556
rect 16172 20544 16178 20596
rect 17126 20584 17132 20596
rect 17087 20556 17132 20584
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 24946 20584 24952 20596
rect 24907 20556 24952 20584
rect 24946 20544 24952 20556
rect 25004 20544 25010 20596
rect 26970 20544 26976 20596
rect 27028 20584 27034 20596
rect 44450 20584 44456 20596
rect 27028 20556 44456 20584
rect 27028 20544 27034 20556
rect 44450 20544 44456 20556
rect 44508 20544 44514 20596
rect 49697 20587 49755 20593
rect 49697 20553 49709 20587
rect 49743 20584 49755 20587
rect 50154 20584 50160 20596
rect 49743 20556 50160 20584
rect 49743 20553 49755 20556
rect 49697 20547 49755 20553
rect 50154 20544 50160 20556
rect 50212 20544 50218 20596
rect 4798 20476 4804 20528
rect 4856 20516 4862 20528
rect 5258 20516 5264 20528
rect 4856 20488 5264 20516
rect 4856 20476 4862 20488
rect 5258 20476 5264 20488
rect 5316 20516 5322 20528
rect 11701 20519 11759 20525
rect 11701 20516 11713 20519
rect 5316 20488 10180 20516
rect 5316 20476 5322 20488
rect 10152 20457 10180 20488
rect 11256 20488 11713 20516
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 5736 20420 7297 20448
rect 5736 20392 5764 20420
rect 7285 20417 7297 20420
rect 7331 20448 7343 20451
rect 10137 20451 10195 20457
rect 7331 20420 7604 20448
rect 7331 20417 7343 20420
rect 7285 20411 7343 20417
rect 3510 20380 3516 20392
rect 3471 20352 3516 20380
rect 3510 20340 3516 20352
rect 3568 20340 3574 20392
rect 3694 20380 3700 20392
rect 3655 20352 3700 20380
rect 3694 20340 3700 20352
rect 3752 20340 3758 20392
rect 4157 20383 4215 20389
rect 4157 20349 4169 20383
rect 4203 20349 4215 20383
rect 4157 20343 4215 20349
rect 3528 20312 3556 20340
rect 4172 20312 4200 20343
rect 4246 20340 4252 20392
rect 4304 20380 4310 20392
rect 5718 20380 5724 20392
rect 4304 20352 4349 20380
rect 5679 20352 5724 20380
rect 4304 20340 4310 20352
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7469 20383 7527 20389
rect 7469 20380 7481 20383
rect 6972 20352 7481 20380
rect 6972 20340 6978 20352
rect 7469 20349 7481 20352
rect 7515 20349 7527 20383
rect 7576 20380 7604 20420
rect 10137 20417 10149 20451
rect 10183 20417 10195 20451
rect 10137 20411 10195 20417
rect 7926 20380 7932 20392
rect 7576 20352 7932 20380
rect 7469 20343 7527 20349
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 8386 20380 8392 20392
rect 8067 20352 8392 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10873 20383 10931 20389
rect 10873 20349 10885 20383
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 11057 20383 11115 20389
rect 11057 20349 11069 20383
rect 11103 20380 11115 20383
rect 11256 20380 11284 20488
rect 11701 20485 11713 20488
rect 11747 20516 11759 20519
rect 12710 20516 12716 20528
rect 11747 20488 12716 20516
rect 11747 20485 11759 20488
rect 11701 20479 11759 20485
rect 12710 20476 12716 20488
rect 12768 20476 12774 20528
rect 16482 20476 16488 20528
rect 16540 20516 16546 20528
rect 24026 20516 24032 20528
rect 16540 20488 24032 20516
rect 16540 20476 16546 20488
rect 24026 20476 24032 20488
rect 24084 20476 24090 20528
rect 24302 20525 24308 20528
rect 24286 20519 24308 20525
rect 24286 20485 24298 20519
rect 24286 20479 24308 20485
rect 24302 20476 24308 20479
rect 24360 20476 24366 20528
rect 26786 20516 26792 20528
rect 26747 20488 26792 20516
rect 26786 20476 26792 20488
rect 26844 20476 26850 20528
rect 30190 20516 30196 20528
rect 30151 20488 30196 20516
rect 30190 20476 30196 20488
rect 30248 20476 30254 20528
rect 30300 20488 35664 20516
rect 11330 20408 11336 20460
rect 11388 20448 11394 20460
rect 15838 20448 15844 20460
rect 11388 20420 15844 20448
rect 11388 20408 11394 20420
rect 13262 20380 13268 20392
rect 11103 20352 11284 20380
rect 13223 20352 13268 20380
rect 11103 20349 11115 20352
rect 11057 20343 11115 20349
rect 3528 20284 4200 20312
rect 4801 20315 4859 20321
rect 4801 20281 4813 20315
rect 4847 20312 4859 20315
rect 5902 20312 5908 20324
rect 4847 20284 5908 20312
rect 4847 20281 4859 20284
rect 4801 20275 4859 20281
rect 5902 20272 5908 20284
rect 5960 20272 5966 20324
rect 10336 20312 10364 20343
rect 10888 20312 10916 20343
rect 13262 20340 13268 20352
rect 13320 20340 13326 20392
rect 13538 20380 13544 20392
rect 13499 20352 13544 20380
rect 13538 20340 13544 20352
rect 13596 20340 13602 20392
rect 15764 20389 15792 20420
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 19242 20448 19248 20460
rect 19203 20420 19248 20448
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 23014 20448 23020 20460
rect 21836 20420 23020 20448
rect 15749 20383 15807 20389
rect 15749 20349 15761 20383
rect 15795 20349 15807 20383
rect 15749 20343 15807 20349
rect 15933 20383 15991 20389
rect 15933 20349 15945 20383
rect 15979 20349 15991 20383
rect 15933 20343 15991 20349
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17954 20380 17960 20392
rect 17359 20352 17960 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 10336 20284 10916 20312
rect 15948 20312 15976 20343
rect 17954 20340 17960 20352
rect 18012 20340 18018 20392
rect 18046 20340 18052 20392
rect 18104 20380 18110 20392
rect 18104 20352 18149 20380
rect 18104 20340 18110 20352
rect 18506 20340 18512 20392
rect 18564 20380 18570 20392
rect 19337 20383 19395 20389
rect 19337 20380 19349 20383
rect 18564 20352 19349 20380
rect 18564 20340 18570 20352
rect 19337 20349 19349 20352
rect 19383 20380 19395 20383
rect 19889 20383 19947 20389
rect 19889 20380 19901 20383
rect 19383 20352 19901 20380
rect 19383 20349 19395 20352
rect 19337 20343 19395 20349
rect 19889 20349 19901 20352
rect 19935 20349 19947 20383
rect 19889 20343 19947 20349
rect 20073 20383 20131 20389
rect 20073 20349 20085 20383
rect 20119 20380 20131 20383
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 20119 20352 20637 20380
rect 20119 20349 20131 20352
rect 20073 20343 20131 20349
rect 20625 20349 20637 20352
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 16485 20315 16543 20321
rect 16485 20312 16497 20315
rect 15948 20284 16497 20312
rect 8481 20247 8539 20253
rect 8481 20213 8493 20247
rect 8527 20244 8539 20247
rect 10410 20244 10416 20256
rect 8527 20216 10416 20244
rect 8527 20213 8539 20216
rect 8481 20207 8539 20213
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 10888 20244 10916 20284
rect 16485 20281 16497 20284
rect 16531 20312 16543 20315
rect 20530 20312 20536 20324
rect 16531 20284 20536 20312
rect 16531 20281 16543 20284
rect 16485 20275 16543 20281
rect 20530 20272 20536 20284
rect 20588 20272 20594 20324
rect 20640 20312 20668 20343
rect 21266 20340 21272 20392
rect 21324 20380 21330 20392
rect 21729 20383 21787 20389
rect 21729 20380 21741 20383
rect 21324 20352 21741 20380
rect 21324 20340 21330 20352
rect 21729 20349 21741 20352
rect 21775 20349 21787 20383
rect 21729 20343 21787 20349
rect 21836 20321 21864 20420
rect 23014 20408 23020 20420
rect 23072 20408 23078 20460
rect 24118 20408 24124 20460
rect 24176 20448 24182 20460
rect 24489 20451 24547 20457
rect 24176 20420 24389 20448
rect 24176 20408 24182 20420
rect 24361 20389 24389 20420
rect 24489 20417 24501 20451
rect 24535 20448 24547 20451
rect 24946 20448 24952 20460
rect 24535 20420 24952 20448
rect 24535 20417 24547 20420
rect 24489 20411 24547 20417
rect 24946 20408 24952 20420
rect 25004 20408 25010 20460
rect 25406 20408 25412 20460
rect 25464 20448 25470 20460
rect 25685 20451 25743 20457
rect 25685 20448 25697 20451
rect 25464 20420 25697 20448
rect 25464 20408 25470 20420
rect 25685 20417 25697 20420
rect 25731 20417 25743 20451
rect 25685 20411 25743 20417
rect 27706 20408 27712 20460
rect 27764 20448 27770 20460
rect 28626 20448 28632 20460
rect 27764 20420 28632 20448
rect 27764 20408 27770 20420
rect 28626 20408 28632 20420
rect 28684 20448 28690 20460
rect 30300 20448 30328 20488
rect 28684 20420 30328 20448
rect 28684 20408 28690 20420
rect 31202 20408 31208 20460
rect 31260 20448 31266 20460
rect 31481 20451 31539 20457
rect 31481 20448 31493 20451
rect 31260 20420 31493 20448
rect 31260 20408 31266 20420
rect 31481 20417 31493 20420
rect 31527 20417 31539 20451
rect 35636 20448 35664 20488
rect 38930 20476 38936 20528
rect 38988 20516 38994 20528
rect 39209 20519 39267 20525
rect 39209 20516 39221 20519
rect 38988 20488 39221 20516
rect 38988 20476 38994 20488
rect 39209 20485 39221 20488
rect 39255 20485 39267 20519
rect 39209 20479 39267 20485
rect 41233 20519 41291 20525
rect 41233 20485 41245 20519
rect 41279 20516 41291 20519
rect 42061 20519 42119 20525
rect 42061 20516 42073 20519
rect 41279 20488 42073 20516
rect 41279 20485 41291 20488
rect 41233 20479 41291 20485
rect 35636 20420 35756 20448
rect 31481 20411 31539 20417
rect 24351 20383 24409 20389
rect 24351 20349 24363 20383
rect 24397 20349 24409 20383
rect 25866 20380 25872 20392
rect 25827 20352 25872 20380
rect 24351 20343 24409 20349
rect 25866 20340 25872 20352
rect 25924 20340 25930 20392
rect 26326 20380 26332 20392
rect 26287 20352 26332 20380
rect 26326 20340 26332 20352
rect 26384 20340 26390 20392
rect 26418 20340 26424 20392
rect 26476 20380 26482 20392
rect 30009 20383 30067 20389
rect 26476 20352 26521 20380
rect 26476 20340 26482 20352
rect 30009 20349 30021 20383
rect 30055 20349 30067 20383
rect 30009 20343 30067 20349
rect 31665 20383 31723 20389
rect 31665 20349 31677 20383
rect 31711 20349 31723 20383
rect 31665 20343 31723 20349
rect 21821 20315 21879 20321
rect 21821 20312 21833 20315
rect 20640 20284 21833 20312
rect 21821 20281 21833 20284
rect 21867 20281 21879 20315
rect 24118 20312 24124 20324
rect 24079 20284 24124 20312
rect 21821 20275 21879 20281
rect 24118 20272 24124 20284
rect 24176 20272 24182 20324
rect 24857 20315 24915 20321
rect 24857 20281 24869 20315
rect 24903 20312 24915 20315
rect 25406 20312 25412 20324
rect 24903 20284 25412 20312
rect 24903 20281 24915 20284
rect 24857 20275 24915 20281
rect 25406 20272 25412 20284
rect 25464 20272 25470 20324
rect 25682 20272 25688 20324
rect 25740 20312 25746 20324
rect 28902 20312 28908 20324
rect 25740 20284 28908 20312
rect 25740 20272 25746 20284
rect 28902 20272 28908 20284
rect 28960 20272 28966 20324
rect 11793 20247 11851 20253
rect 11793 20244 11805 20247
rect 10888 20216 11805 20244
rect 11793 20213 11805 20216
rect 11839 20244 11851 20247
rect 11977 20247 12035 20253
rect 11977 20244 11989 20247
rect 11839 20216 11989 20244
rect 11839 20213 11851 20216
rect 11793 20207 11851 20213
rect 11977 20213 11989 20216
rect 12023 20244 12035 20247
rect 12158 20244 12164 20256
rect 12023 20216 12164 20244
rect 12023 20213 12035 20216
rect 11977 20207 12035 20213
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 14182 20204 14188 20256
rect 14240 20244 14246 20256
rect 14645 20247 14703 20253
rect 14645 20244 14657 20247
rect 14240 20216 14657 20244
rect 14240 20204 14246 20216
rect 14645 20213 14657 20216
rect 14691 20213 14703 20247
rect 14645 20207 14703 20213
rect 18233 20247 18291 20253
rect 18233 20213 18245 20247
rect 18279 20244 18291 20247
rect 18322 20244 18328 20256
rect 18279 20216 18328 20244
rect 18279 20213 18291 20216
rect 18233 20207 18291 20213
rect 18322 20204 18328 20216
rect 18380 20204 18386 20256
rect 20346 20244 20352 20256
rect 20307 20216 20352 20244
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 23382 20204 23388 20256
rect 23440 20244 23446 20256
rect 29917 20247 29975 20253
rect 29917 20244 29929 20247
rect 23440 20216 29929 20244
rect 23440 20204 23446 20216
rect 29917 20213 29929 20216
rect 29963 20244 29975 20247
rect 30024 20244 30052 20343
rect 31680 20312 31708 20343
rect 32030 20340 32036 20392
rect 32088 20380 32094 20392
rect 32217 20383 32275 20389
rect 32217 20380 32229 20383
rect 32088 20352 32229 20380
rect 32088 20340 32094 20352
rect 32217 20349 32229 20352
rect 32263 20349 32275 20383
rect 32398 20380 32404 20392
rect 32359 20352 32404 20380
rect 32217 20343 32275 20349
rect 32398 20340 32404 20352
rect 32456 20340 32462 20392
rect 35621 20383 35679 20389
rect 35621 20349 35633 20383
rect 35667 20349 35679 20383
rect 35728 20380 35756 20420
rect 35802 20408 35808 20460
rect 35860 20448 35866 20460
rect 35897 20451 35955 20457
rect 35897 20448 35909 20451
rect 35860 20420 35909 20448
rect 35860 20408 35866 20420
rect 35897 20417 35909 20420
rect 35943 20417 35955 20451
rect 38102 20448 38108 20460
rect 38063 20420 38108 20448
rect 35897 20411 35955 20417
rect 38102 20408 38108 20420
rect 38160 20408 38166 20460
rect 38010 20380 38016 20392
rect 35728 20352 38016 20380
rect 35621 20343 35679 20349
rect 32048 20312 32076 20340
rect 31680 20284 32076 20312
rect 32769 20315 32827 20321
rect 32769 20281 32781 20315
rect 32815 20312 32827 20315
rect 33226 20312 33232 20324
rect 32815 20284 33232 20312
rect 32815 20281 32827 20284
rect 32769 20275 32827 20281
rect 33226 20272 33232 20284
rect 33284 20272 33290 20324
rect 35636 20312 35664 20343
rect 38010 20340 38016 20352
rect 38068 20340 38074 20392
rect 38286 20380 38292 20392
rect 38199 20352 38292 20380
rect 38286 20340 38292 20352
rect 38344 20380 38350 20392
rect 38841 20383 38899 20389
rect 38841 20380 38853 20383
rect 38344 20352 38853 20380
rect 38344 20340 38350 20352
rect 38841 20349 38853 20352
rect 38887 20349 38899 20383
rect 38841 20343 38899 20349
rect 39025 20383 39083 20389
rect 39025 20349 39037 20383
rect 39071 20380 39083 20383
rect 40034 20380 40040 20392
rect 39071 20352 40040 20380
rect 39071 20349 39083 20352
rect 39025 20343 39083 20349
rect 40034 20340 40040 20352
rect 40092 20340 40098 20392
rect 41417 20383 41475 20389
rect 41417 20349 41429 20383
rect 41463 20349 41475 20383
rect 41708 20380 41736 20488
rect 42061 20485 42073 20488
rect 42107 20485 42119 20519
rect 42061 20479 42119 20485
rect 41782 20408 41788 20460
rect 41840 20448 41846 20460
rect 43625 20451 43683 20457
rect 43625 20448 43637 20451
rect 41840 20420 43637 20448
rect 41840 20408 41846 20420
rect 43625 20417 43637 20420
rect 43671 20417 43683 20451
rect 43625 20411 43683 20417
rect 45554 20408 45560 20460
rect 45612 20448 45618 20460
rect 46109 20451 46167 20457
rect 46109 20448 46121 20451
rect 45612 20420 46121 20448
rect 45612 20408 45618 20420
rect 46109 20417 46121 20420
rect 46155 20417 46167 20451
rect 50172 20448 50200 20544
rect 50706 20516 50712 20528
rect 50667 20488 50712 20516
rect 50706 20476 50712 20488
rect 50764 20476 50770 20528
rect 51721 20451 51779 20457
rect 51721 20448 51733 20451
rect 50172 20420 51733 20448
rect 46109 20411 46167 20417
rect 51721 20417 51733 20420
rect 51767 20417 51779 20451
rect 51721 20411 51779 20417
rect 42245 20383 42303 20389
rect 42245 20380 42257 20383
rect 41708 20352 42257 20380
rect 41417 20343 41475 20349
rect 42245 20349 42257 20352
rect 42291 20349 42303 20383
rect 42245 20343 42303 20349
rect 42521 20383 42579 20389
rect 42521 20349 42533 20383
rect 42567 20380 42579 20383
rect 42886 20380 42892 20392
rect 42567 20352 42892 20380
rect 42567 20349 42579 20352
rect 42521 20343 42579 20349
rect 37274 20312 37280 20324
rect 35636 20284 35756 20312
rect 37235 20284 37280 20312
rect 31110 20244 31116 20256
rect 29963 20216 31116 20244
rect 29963 20213 29975 20216
rect 29917 20207 29975 20213
rect 31110 20204 31116 20216
rect 31168 20204 31174 20256
rect 35728 20244 35756 20284
rect 37274 20272 37280 20284
rect 37332 20272 37338 20324
rect 38470 20272 38476 20324
rect 38528 20312 38534 20324
rect 41432 20312 41460 20343
rect 38528 20284 41460 20312
rect 38528 20272 38534 20284
rect 35894 20244 35900 20256
rect 35728 20216 35900 20244
rect 35894 20204 35900 20216
rect 35952 20244 35958 20256
rect 37369 20247 37427 20253
rect 37369 20244 37381 20247
rect 35952 20216 37381 20244
rect 35952 20204 35958 20216
rect 37369 20213 37381 20216
rect 37415 20213 37427 20247
rect 42260 20244 42288 20343
rect 42886 20340 42892 20352
rect 42944 20340 42950 20392
rect 46293 20383 46351 20389
rect 46293 20349 46305 20383
rect 46339 20349 46351 20383
rect 46750 20380 46756 20392
rect 46711 20352 46756 20380
rect 46293 20343 46351 20349
rect 46106 20272 46112 20324
rect 46164 20312 46170 20324
rect 46308 20312 46336 20343
rect 46750 20340 46756 20352
rect 46808 20340 46814 20392
rect 46845 20383 46903 20389
rect 46845 20349 46857 20383
rect 46891 20349 46903 20383
rect 48406 20380 48412 20392
rect 48367 20352 48412 20380
rect 46845 20343 46903 20349
rect 46860 20312 46888 20343
rect 48406 20340 48412 20352
rect 48464 20340 48470 20392
rect 49605 20383 49663 20389
rect 49605 20349 49617 20383
rect 49651 20349 49663 20383
rect 49605 20343 49663 20349
rect 50617 20383 50675 20389
rect 50617 20349 50629 20383
rect 50663 20349 50675 20383
rect 50617 20343 50675 20349
rect 46164 20284 46888 20312
rect 46164 20272 46170 20284
rect 46934 20272 46940 20324
rect 46992 20312 46998 20324
rect 49620 20312 49648 20343
rect 49881 20315 49939 20321
rect 49881 20312 49893 20315
rect 46992 20284 49893 20312
rect 46992 20272 46998 20284
rect 49881 20281 49893 20284
rect 49927 20281 49939 20315
rect 50632 20312 50660 20343
rect 50706 20340 50712 20392
rect 50764 20380 50770 20392
rect 51905 20383 51963 20389
rect 51905 20380 51917 20383
rect 50764 20352 51917 20380
rect 50764 20340 50770 20352
rect 51905 20349 51917 20352
rect 51951 20349 51963 20383
rect 51905 20343 51963 20349
rect 52086 20340 52092 20392
rect 52144 20380 52150 20392
rect 52365 20383 52423 20389
rect 52365 20380 52377 20383
rect 52144 20352 52377 20380
rect 52144 20340 52150 20352
rect 52365 20349 52377 20352
rect 52411 20349 52423 20383
rect 52365 20343 52423 20349
rect 52457 20383 52515 20389
rect 52457 20349 52469 20383
rect 52503 20380 52515 20383
rect 53374 20380 53380 20392
rect 52503 20352 53380 20380
rect 52503 20349 52515 20352
rect 52457 20343 52515 20349
rect 53374 20340 53380 20352
rect 53432 20340 53438 20392
rect 51350 20312 51356 20324
rect 50632 20284 51356 20312
rect 49881 20275 49939 20281
rect 42978 20244 42984 20256
rect 42260 20216 42984 20244
rect 37369 20207 37427 20213
rect 42978 20204 42984 20216
rect 43036 20204 43042 20256
rect 46290 20204 46296 20256
rect 46348 20244 46354 20256
rect 47305 20247 47363 20253
rect 47305 20244 47317 20247
rect 46348 20216 47317 20244
rect 46348 20204 46354 20216
rect 47305 20213 47317 20216
rect 47351 20213 47363 20247
rect 47305 20207 47363 20213
rect 48501 20247 48559 20253
rect 48501 20213 48513 20247
rect 48547 20244 48559 20247
rect 49234 20244 49240 20256
rect 48547 20216 49240 20244
rect 48547 20213 48559 20216
rect 48501 20207 48559 20213
rect 49234 20204 49240 20216
rect 49292 20204 49298 20256
rect 49896 20244 49924 20275
rect 51350 20272 51356 20284
rect 51408 20312 51414 20324
rect 51994 20312 52000 20324
rect 51408 20284 52000 20312
rect 51408 20272 51414 20284
rect 51994 20272 52000 20284
rect 52052 20272 52058 20324
rect 52270 20244 52276 20256
rect 49896 20216 52276 20244
rect 52270 20204 52276 20216
rect 52328 20204 52334 20256
rect 52914 20244 52920 20256
rect 52875 20216 52920 20244
rect 52914 20204 52920 20216
rect 52972 20204 52978 20256
rect 1104 20154 54832 20176
rect 1104 20102 18912 20154
rect 18964 20102 18976 20154
rect 19028 20102 19040 20154
rect 19092 20102 19104 20154
rect 19156 20102 36843 20154
rect 36895 20102 36907 20154
rect 36959 20102 36971 20154
rect 37023 20102 37035 20154
rect 37087 20102 54832 20154
rect 1104 20080 54832 20102
rect 3053 20043 3111 20049
rect 3053 20009 3065 20043
rect 3099 20040 3111 20043
rect 3510 20040 3516 20052
rect 3099 20012 3516 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 4433 20043 4491 20049
rect 4433 20009 4445 20043
rect 4479 20040 4491 20043
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 4479 20012 7297 20040
rect 4479 20009 4491 20012
rect 4433 20003 4491 20009
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 8386 20040 8392 20052
rect 8347 20012 8392 20040
rect 7285 20003 7343 20009
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 9769 20043 9827 20049
rect 9769 20040 9781 20043
rect 9732 20012 9781 20040
rect 9732 20000 9738 20012
rect 9769 20009 9781 20012
rect 9815 20009 9827 20043
rect 9769 20003 9827 20009
rect 16298 20000 16304 20052
rect 16356 20040 16362 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16356 20012 16865 20040
rect 16356 20000 16362 20012
rect 16853 20009 16865 20012
rect 16899 20040 16911 20043
rect 18046 20040 18052 20052
rect 16899 20012 18052 20040
rect 16899 20009 16911 20012
rect 16853 20003 16911 20009
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 21266 20000 21272 20052
rect 21324 20040 21330 20052
rect 22281 20043 22339 20049
rect 22281 20040 22293 20043
rect 21324 20012 22293 20040
rect 21324 20000 21330 20012
rect 22281 20009 22293 20012
rect 22327 20009 22339 20043
rect 23382 20040 23388 20052
rect 23343 20012 23388 20040
rect 22281 20003 22339 20009
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 30466 20040 30472 20052
rect 24176 20012 30472 20040
rect 24176 20000 24182 20012
rect 30466 20000 30472 20012
rect 30524 20000 30530 20052
rect 30742 20000 30748 20052
rect 30800 20040 30806 20052
rect 31021 20043 31079 20049
rect 31021 20040 31033 20043
rect 30800 20012 31033 20040
rect 30800 20000 30806 20012
rect 31021 20009 31033 20012
rect 31067 20009 31079 20043
rect 31021 20003 31079 20009
rect 31110 20000 31116 20052
rect 31168 20040 31174 20052
rect 32214 20040 32220 20052
rect 31168 20012 32220 20040
rect 31168 20000 31174 20012
rect 32214 20000 32220 20012
rect 32272 20000 32278 20052
rect 32306 20000 32312 20052
rect 32364 20040 32370 20052
rect 34517 20043 34575 20049
rect 34517 20040 34529 20043
rect 32364 20012 34529 20040
rect 32364 20000 32370 20012
rect 34517 20009 34529 20012
rect 34563 20009 34575 20043
rect 34517 20003 34575 20009
rect 36170 20000 36176 20052
rect 36228 20040 36234 20052
rect 38470 20040 38476 20052
rect 36228 20012 38476 20040
rect 36228 20000 36234 20012
rect 38470 20000 38476 20012
rect 38528 20000 38534 20052
rect 45554 20040 45560 20052
rect 39224 20012 45560 20040
rect 1489 19907 1547 19913
rect 1489 19873 1501 19907
rect 1535 19904 1547 19907
rect 3326 19904 3332 19916
rect 1535 19876 3332 19904
rect 1535 19873 1547 19876
rect 1489 19867 1547 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 3528 19904 3556 20000
rect 4617 19975 4675 19981
rect 4617 19941 4629 19975
rect 4663 19972 4675 19975
rect 11330 19972 11336 19984
rect 4663 19944 10180 19972
rect 4663 19941 4675 19944
rect 4617 19935 4675 19941
rect 4525 19907 4583 19913
rect 4525 19904 4537 19907
rect 3528 19876 4537 19904
rect 4525 19873 4537 19876
rect 4571 19873 4583 19907
rect 4525 19867 4583 19873
rect 6273 19907 6331 19913
rect 6273 19873 6285 19907
rect 6319 19904 6331 19907
rect 6638 19904 6644 19916
rect 6319 19876 6644 19904
rect 6319 19873 6331 19876
rect 6273 19867 6331 19873
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 6730 19864 6736 19916
rect 6788 19904 6794 19916
rect 7024 19913 7052 19944
rect 10152 19913 10180 19944
rect 10704 19944 11336 19972
rect 10704 19913 10732 19944
rect 11330 19932 11336 19944
rect 11388 19932 11394 19984
rect 13265 19975 13323 19981
rect 12728 19944 13032 19972
rect 6825 19907 6883 19913
rect 6825 19904 6837 19907
rect 6788 19876 6837 19904
rect 6788 19864 6794 19876
rect 6825 19873 6837 19876
rect 6871 19873 6883 19907
rect 6825 19867 6883 19873
rect 7009 19907 7067 19913
rect 7009 19873 7021 19907
rect 7055 19873 7067 19907
rect 7009 19867 7067 19873
rect 8297 19907 8355 19913
rect 8297 19873 8309 19907
rect 8343 19873 8355 19907
rect 8297 19867 8355 19873
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 10321 19907 10379 19913
rect 10321 19873 10333 19907
rect 10367 19873 10379 19907
rect 10321 19867 10379 19873
rect 10689 19907 10747 19913
rect 10689 19873 10701 19907
rect 10735 19873 10747 19907
rect 10689 19867 10747 19873
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19904 10931 19907
rect 12158 19904 12164 19916
rect 10919 19876 11100 19904
rect 12119 19876 12164 19904
rect 10919 19873 10931 19876
rect 10873 19867 10931 19873
rect 1762 19845 1768 19848
rect 1759 19836 1768 19845
rect 1723 19808 1768 19836
rect 1759 19799 1768 19808
rect 1762 19796 1768 19799
rect 1820 19796 1826 19848
rect 6178 19836 6184 19848
rect 6139 19808 6184 19836
rect 6178 19796 6184 19808
rect 6236 19796 6242 19848
rect 1762 19660 1768 19712
rect 1820 19700 1826 19712
rect 4433 19703 4491 19709
rect 4433 19700 4445 19703
rect 1820 19672 4445 19700
rect 1820 19660 1826 19672
rect 4433 19669 4445 19672
rect 4479 19669 4491 19703
rect 4433 19663 4491 19669
rect 5902 19660 5908 19712
rect 5960 19700 5966 19712
rect 8312 19700 8340 19867
rect 8570 19796 8576 19848
rect 8628 19836 8634 19848
rect 9582 19836 9588 19848
rect 8628 19808 9588 19836
rect 8628 19796 8634 19808
rect 9582 19796 9588 19808
rect 9640 19836 9646 19848
rect 10336 19836 10364 19867
rect 9640 19808 10364 19836
rect 9640 19796 9646 19808
rect 11072 19777 11100 19876
rect 12158 19864 12164 19876
rect 12216 19904 12222 19916
rect 12728 19913 12756 19944
rect 12713 19907 12771 19913
rect 12713 19904 12725 19907
rect 12216 19876 12725 19904
rect 12216 19864 12222 19876
rect 12713 19873 12725 19876
rect 12759 19873 12771 19907
rect 12894 19904 12900 19916
rect 12855 19876 12900 19904
rect 12713 19867 12771 19873
rect 12894 19864 12900 19876
rect 12952 19864 12958 19916
rect 13004 19904 13032 19944
rect 13265 19941 13277 19975
rect 13311 19972 13323 19975
rect 13538 19972 13544 19984
rect 13311 19944 13544 19972
rect 13311 19941 13323 19944
rect 13265 19935 13323 19941
rect 13538 19932 13544 19944
rect 13596 19932 13602 19984
rect 14182 19904 14188 19916
rect 13004 19876 13768 19904
rect 14143 19876 14188 19904
rect 11974 19836 11980 19848
rect 11935 19808 11980 19836
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 13740 19845 13768 19876
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 16298 19904 16304 19916
rect 15611 19876 16304 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19904 16727 19907
rect 17494 19904 17500 19916
rect 16715 19876 17500 19904
rect 16715 19873 16727 19876
rect 16669 19867 16727 19873
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 18141 19907 18199 19913
rect 18141 19873 18153 19907
rect 18187 19904 18199 19907
rect 18230 19904 18236 19916
rect 18187 19876 18236 19904
rect 18187 19873 18199 19876
rect 18141 19867 18199 19873
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19836 13783 19839
rect 13909 19839 13967 19845
rect 13909 19836 13921 19839
rect 13771 19808 13921 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 13909 19805 13921 19808
rect 13955 19836 13967 19839
rect 16482 19836 16488 19848
rect 13955 19808 16488 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 17218 19796 17224 19848
rect 17276 19836 17282 19848
rect 18064 19836 18092 19867
rect 18230 19864 18236 19876
rect 18288 19864 18294 19916
rect 18506 19864 18512 19916
rect 18564 19904 18570 19916
rect 18601 19907 18659 19913
rect 18601 19904 18613 19907
rect 18564 19876 18613 19904
rect 18564 19864 18570 19876
rect 18601 19873 18613 19876
rect 18647 19873 18659 19907
rect 18601 19867 18659 19873
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 19334 19904 19340 19916
rect 18831 19876 19340 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 20346 19864 20352 19916
rect 20404 19904 20410 19916
rect 21177 19907 21235 19913
rect 21177 19904 21189 19907
rect 20404 19876 21189 19904
rect 20404 19864 20410 19876
rect 21177 19873 21189 19876
rect 21223 19873 21235 19907
rect 21177 19867 21235 19873
rect 23400 19904 23428 20000
rect 26881 19975 26939 19981
rect 26881 19972 26893 19975
rect 26528 19944 26893 19972
rect 26528 19913 26556 19944
rect 26881 19941 26893 19944
rect 26927 19972 26939 19975
rect 27706 19972 27712 19984
rect 26927 19944 27712 19972
rect 26927 19941 26939 19944
rect 26881 19935 26939 19941
rect 27706 19932 27712 19944
rect 27764 19932 27770 19984
rect 28994 19932 29000 19984
rect 29052 19972 29058 19984
rect 29549 19975 29607 19981
rect 29549 19972 29561 19975
rect 29052 19944 29561 19972
rect 29052 19932 29058 19944
rect 29549 19941 29561 19944
rect 29595 19941 29607 19975
rect 29549 19935 29607 19941
rect 34790 19932 34796 19984
rect 34848 19972 34854 19984
rect 38378 19972 38384 19984
rect 34848 19944 38384 19972
rect 34848 19932 34854 19944
rect 38378 19932 38384 19944
rect 38436 19932 38442 19984
rect 23477 19907 23535 19913
rect 23477 19904 23489 19907
rect 23400 19876 23489 19904
rect 17276 19808 18092 19836
rect 19153 19839 19211 19845
rect 17276 19796 17282 19808
rect 19153 19805 19165 19839
rect 19199 19836 19211 19839
rect 19702 19836 19708 19848
rect 19199 19808 19708 19836
rect 19199 19805 19211 19808
rect 19153 19799 19211 19805
rect 19702 19796 19708 19808
rect 19760 19796 19766 19848
rect 20714 19836 20720 19848
rect 20675 19808 20720 19836
rect 20714 19796 20720 19808
rect 20772 19836 20778 19848
rect 20901 19839 20959 19845
rect 20901 19836 20913 19839
rect 20772 19808 20913 19836
rect 20772 19796 20778 19808
rect 20901 19805 20913 19808
rect 20947 19836 20959 19839
rect 21542 19836 21548 19848
rect 20947 19808 21548 19836
rect 20947 19805 20959 19808
rect 20901 19799 20959 19805
rect 21542 19796 21548 19808
rect 21600 19796 21606 19848
rect 11057 19771 11115 19777
rect 11057 19737 11069 19771
rect 11103 19768 11115 19771
rect 12894 19768 12900 19780
rect 11103 19740 12900 19768
rect 11103 19737 11115 19740
rect 11057 19731 11115 19737
rect 12894 19728 12900 19740
rect 12952 19768 12958 19780
rect 13449 19771 13507 19777
rect 13449 19768 13461 19771
rect 12952 19740 13461 19768
rect 12952 19728 12958 19740
rect 13449 19737 13461 19740
rect 13495 19768 13507 19771
rect 14277 19771 14335 19777
rect 14277 19768 14289 19771
rect 13495 19740 14289 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 14277 19737 14289 19740
rect 14323 19768 14335 19771
rect 17862 19768 17868 19780
rect 14323 19740 17868 19768
rect 14323 19737 14335 19740
rect 14277 19731 14335 19737
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 15746 19700 15752 19712
rect 5960 19672 8340 19700
rect 15707 19672 15752 19700
rect 5960 19660 5966 19672
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 18046 19660 18052 19712
rect 18104 19700 18110 19712
rect 18322 19700 18328 19712
rect 18104 19672 18328 19700
rect 18104 19660 18110 19672
rect 18322 19660 18328 19672
rect 18380 19700 18386 19712
rect 23400 19700 23428 19876
rect 23477 19873 23489 19876
rect 23523 19873 23535 19907
rect 25133 19907 25191 19913
rect 25133 19904 25145 19907
rect 23477 19867 23535 19873
rect 24964 19876 25145 19904
rect 24964 19768 24992 19876
rect 25133 19873 25145 19876
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 26513 19907 26571 19913
rect 26513 19873 26525 19907
rect 26559 19873 26571 19907
rect 28077 19907 28135 19913
rect 28077 19904 28089 19907
rect 26513 19867 26571 19873
rect 27724 19876 28089 19904
rect 27724 19848 27752 19876
rect 28077 19873 28089 19876
rect 28123 19873 28135 19907
rect 30926 19904 30932 19916
rect 30887 19876 30932 19904
rect 28077 19867 28135 19873
rect 30926 19864 30932 19876
rect 30984 19904 30990 19916
rect 31294 19904 31300 19916
rect 30984 19876 31300 19904
rect 30984 19864 30990 19876
rect 31294 19864 31300 19876
rect 31352 19864 31358 19916
rect 32766 19864 32772 19916
rect 32824 19904 32830 19916
rect 32953 19907 33011 19913
rect 32953 19904 32965 19907
rect 32824 19876 32965 19904
rect 32824 19864 32830 19876
rect 32953 19873 32965 19876
rect 32999 19873 33011 19907
rect 33226 19904 33232 19916
rect 33187 19876 33232 19904
rect 32953 19867 33011 19873
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19836 25099 19839
rect 26326 19836 26332 19848
rect 25087 19808 26332 19836
rect 25087 19805 25099 19808
rect 25041 19799 25099 19805
rect 26326 19796 26332 19808
rect 26384 19836 26390 19848
rect 26605 19839 26663 19845
rect 26605 19836 26617 19839
rect 26384 19808 26617 19836
rect 26384 19796 26390 19808
rect 26605 19805 26617 19808
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 27706 19796 27712 19848
rect 27764 19796 27770 19848
rect 27801 19839 27859 19845
rect 27801 19805 27813 19839
rect 27847 19836 27859 19839
rect 28994 19836 29000 19848
rect 27847 19808 29000 19836
rect 27847 19805 27859 19808
rect 27801 19799 27859 19805
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29178 19836 29184 19848
rect 29139 19808 29184 19836
rect 29178 19796 29184 19808
rect 29236 19796 29242 19848
rect 32968 19836 32996 19867
rect 33226 19864 33232 19876
rect 33284 19864 33290 19916
rect 37366 19864 37372 19916
rect 37424 19904 37430 19916
rect 39224 19913 39252 20012
rect 45554 20000 45560 20012
rect 45612 20000 45618 20052
rect 45646 20000 45652 20052
rect 45704 20040 45710 20052
rect 45833 20043 45891 20049
rect 45833 20040 45845 20043
rect 45704 20012 45845 20040
rect 45704 20000 45710 20012
rect 45833 20009 45845 20012
rect 45879 20040 45891 20043
rect 46014 20040 46020 20052
rect 45879 20012 46020 20040
rect 45879 20009 45891 20012
rect 45833 20003 45891 20009
rect 46014 20000 46020 20012
rect 46072 20000 46078 20052
rect 46382 20000 46388 20052
rect 46440 20040 46446 20052
rect 52914 20040 52920 20052
rect 46440 20012 52920 20040
rect 46440 20000 46446 20012
rect 52914 20000 52920 20012
rect 52972 20000 52978 20052
rect 53374 20040 53380 20052
rect 53335 20012 53380 20040
rect 53374 20000 53380 20012
rect 53432 20000 53438 20052
rect 50617 19975 50675 19981
rect 39316 19944 40540 19972
rect 39316 19913 39344 19944
rect 38657 19907 38715 19913
rect 38657 19904 38669 19907
rect 37424 19876 38669 19904
rect 37424 19864 37430 19876
rect 38657 19873 38669 19876
rect 38703 19873 38715 19907
rect 38657 19867 38715 19873
rect 39209 19907 39267 19913
rect 39209 19873 39221 19907
rect 39255 19873 39267 19907
rect 39209 19867 39267 19873
rect 39301 19907 39359 19913
rect 39301 19873 39313 19907
rect 39347 19873 39359 19907
rect 39669 19907 39727 19913
rect 39669 19904 39681 19907
rect 39301 19867 39359 19873
rect 39408 19876 39681 19904
rect 34701 19839 34759 19845
rect 34701 19836 34713 19839
rect 32968 19808 34713 19836
rect 34701 19805 34713 19808
rect 34747 19836 34759 19839
rect 35342 19836 35348 19848
rect 34747 19808 35348 19836
rect 34747 19805 34759 19808
rect 34701 19799 34759 19805
rect 35342 19796 35348 19808
rect 35400 19796 35406 19848
rect 38286 19796 38292 19848
rect 38344 19836 38350 19848
rect 39408 19836 39436 19876
rect 39669 19873 39681 19876
rect 39715 19873 39727 19907
rect 39669 19867 39727 19873
rect 39758 19864 39764 19916
rect 39816 19904 39822 19916
rect 39816 19876 39861 19904
rect 39816 19864 39822 19876
rect 38344 19808 39436 19836
rect 40512 19836 40540 19944
rect 50617 19941 50629 19975
rect 50663 19972 50675 19975
rect 50706 19972 50712 19984
rect 50663 19944 50712 19972
rect 50663 19941 50675 19944
rect 50617 19935 50675 19941
rect 50706 19932 50712 19944
rect 50764 19932 50770 19984
rect 51718 19932 51724 19984
rect 51776 19972 51782 19984
rect 51813 19975 51871 19981
rect 51813 19972 51825 19975
rect 51776 19944 51825 19972
rect 51776 19932 51782 19944
rect 51813 19941 51825 19944
rect 51859 19972 51871 19975
rect 51859 19944 52040 19972
rect 51859 19941 51871 19944
rect 51813 19935 51871 19941
rect 41046 19864 41052 19916
rect 41104 19904 41110 19916
rect 41233 19907 41291 19913
rect 41233 19904 41245 19907
rect 41104 19876 41245 19904
rect 41104 19864 41110 19876
rect 41233 19873 41245 19876
rect 41279 19873 41291 19907
rect 41233 19867 41291 19873
rect 45738 19864 45744 19916
rect 45796 19904 45802 19916
rect 46290 19904 46296 19916
rect 45796 19876 46152 19904
rect 46251 19876 46296 19904
rect 45796 19864 45802 19876
rect 46014 19836 46020 19848
rect 40512 19808 40632 19836
rect 45975 19808 46020 19836
rect 38344 19796 38350 19808
rect 25777 19771 25835 19777
rect 25777 19768 25789 19771
rect 24964 19740 25789 19768
rect 25777 19737 25789 19740
rect 25823 19768 25835 19771
rect 32582 19768 32588 19780
rect 25823 19740 27568 19768
rect 25823 19737 25835 19740
rect 25777 19731 25835 19737
rect 23658 19700 23664 19712
rect 18380 19672 23428 19700
rect 23619 19672 23664 19700
rect 18380 19660 18386 19672
rect 23658 19660 23664 19672
rect 23716 19660 23722 19712
rect 24302 19660 24308 19712
rect 24360 19700 24366 19712
rect 25317 19703 25375 19709
rect 25317 19700 25329 19703
rect 24360 19672 25329 19700
rect 24360 19660 24366 19672
rect 25317 19669 25329 19672
rect 25363 19669 25375 19703
rect 27540 19700 27568 19740
rect 28736 19740 32588 19768
rect 28736 19700 28764 19740
rect 32582 19728 32588 19740
rect 32640 19728 32646 19780
rect 40126 19768 40132 19780
rect 40087 19740 40132 19768
rect 40126 19728 40132 19740
rect 40184 19728 40190 19780
rect 40604 19777 40632 19808
rect 46014 19796 46020 19808
rect 46072 19796 46078 19848
rect 46124 19836 46152 19876
rect 46290 19864 46296 19876
rect 46348 19864 46354 19916
rect 48590 19864 48596 19916
rect 48648 19904 48654 19916
rect 48777 19907 48835 19913
rect 48777 19904 48789 19907
rect 48648 19876 48789 19904
rect 48648 19864 48654 19876
rect 48777 19873 48789 19876
rect 48823 19904 48835 19907
rect 48961 19907 49019 19913
rect 48961 19904 48973 19907
rect 48823 19876 48973 19904
rect 48823 19873 48835 19876
rect 48777 19867 48835 19873
rect 48961 19873 48973 19876
rect 49007 19873 49019 19907
rect 49234 19904 49240 19916
rect 49195 19876 49240 19904
rect 48961 19867 49019 19873
rect 49234 19864 49240 19876
rect 49292 19864 49298 19916
rect 52012 19913 52040 19944
rect 51997 19907 52055 19913
rect 51997 19873 52009 19907
rect 52043 19873 52055 19907
rect 51997 19867 52055 19873
rect 48498 19836 48504 19848
rect 46124 19808 48504 19836
rect 48498 19796 48504 19808
rect 48556 19796 48562 19848
rect 52273 19839 52331 19845
rect 52273 19805 52285 19839
rect 52319 19836 52331 19839
rect 52730 19836 52736 19848
rect 52319 19808 52736 19836
rect 52319 19805 52331 19808
rect 52273 19799 52331 19805
rect 52730 19796 52736 19808
rect 52788 19796 52794 19848
rect 40589 19771 40647 19777
rect 40589 19737 40601 19771
rect 40635 19768 40647 19771
rect 40635 19740 42656 19768
rect 40635 19737 40647 19740
rect 40589 19731 40647 19737
rect 41046 19700 41052 19712
rect 27540 19672 28764 19700
rect 41007 19672 41052 19700
rect 25317 19663 25375 19669
rect 41046 19660 41052 19672
rect 41104 19660 41110 19712
rect 41414 19660 41420 19712
rect 41472 19700 41478 19712
rect 42628 19700 42656 19740
rect 46934 19700 46940 19712
rect 41472 19672 41517 19700
rect 42628 19672 46940 19700
rect 41472 19660 41478 19672
rect 46934 19660 46940 19672
rect 46992 19660 46998 19712
rect 47394 19700 47400 19712
rect 47355 19672 47400 19700
rect 47394 19660 47400 19672
rect 47452 19660 47458 19712
rect 1104 19610 54832 19632
rect 1104 19558 9947 19610
rect 9999 19558 10011 19610
rect 10063 19558 10075 19610
rect 10127 19558 10139 19610
rect 10191 19558 27878 19610
rect 27930 19558 27942 19610
rect 27994 19558 28006 19610
rect 28058 19558 28070 19610
rect 28122 19558 45808 19610
rect 45860 19558 45872 19610
rect 45924 19558 45936 19610
rect 45988 19558 46000 19610
rect 46052 19558 54832 19610
rect 1104 19536 54832 19558
rect 3053 19499 3111 19505
rect 3053 19465 3065 19499
rect 3099 19496 3111 19499
rect 3694 19496 3700 19508
rect 3099 19468 3700 19496
rect 3099 19465 3111 19468
rect 3053 19459 3111 19465
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 10502 19496 10508 19508
rect 10463 19468 10508 19496
rect 10502 19456 10508 19468
rect 10560 19456 10566 19508
rect 16482 19496 16488 19508
rect 16443 19468 16488 19496
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 18506 19496 18512 19508
rect 18467 19468 18512 19496
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 18598 19456 18604 19508
rect 18656 19496 18662 19508
rect 27338 19496 27344 19508
rect 18656 19468 27344 19496
rect 18656 19456 18662 19468
rect 27338 19456 27344 19468
rect 27396 19456 27402 19508
rect 30466 19496 30472 19508
rect 30427 19468 30472 19496
rect 30466 19456 30472 19468
rect 30524 19456 30530 19508
rect 32214 19456 32220 19508
rect 32272 19496 32278 19508
rect 41046 19496 41052 19508
rect 32272 19468 41052 19496
rect 32272 19456 32278 19468
rect 41046 19456 41052 19468
rect 41104 19456 41110 19508
rect 42886 19496 42892 19508
rect 42847 19468 42892 19496
rect 42886 19456 42892 19468
rect 42944 19456 42950 19508
rect 44818 19456 44824 19508
rect 44876 19496 44882 19508
rect 47394 19496 47400 19508
rect 44876 19468 47400 19496
rect 44876 19456 44882 19468
rect 47394 19456 47400 19468
rect 47452 19456 47458 19508
rect 6178 19388 6184 19440
rect 6236 19428 6242 19440
rect 11974 19428 11980 19440
rect 6236 19400 11980 19428
rect 6236 19388 6242 19400
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 17405 19431 17463 19437
rect 17405 19397 17417 19431
rect 17451 19428 17463 19431
rect 17954 19428 17960 19440
rect 17451 19400 17960 19428
rect 17451 19397 17463 19400
rect 17405 19391 17463 19397
rect 17954 19388 17960 19400
rect 18012 19428 18018 19440
rect 18230 19428 18236 19440
rect 18012 19400 18236 19428
rect 18012 19388 18018 19400
rect 18230 19388 18236 19400
rect 18288 19388 18294 19440
rect 20530 19388 20536 19440
rect 20588 19428 20594 19440
rect 26510 19428 26516 19440
rect 20588 19400 26516 19428
rect 20588 19388 20594 19400
rect 26510 19388 26516 19400
rect 26568 19388 26574 19440
rect 27798 19388 27804 19440
rect 27856 19428 27862 19440
rect 52362 19428 52368 19440
rect 27856 19400 52368 19428
rect 27856 19388 27862 19400
rect 52362 19388 52368 19400
rect 52420 19388 52426 19440
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8159 19332 8340 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 8312 19304 8340 19332
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 22002 19360 22008 19372
rect 10468 19332 22008 19360
rect 10468 19320 10474 19332
rect 22002 19320 22008 19332
rect 22060 19320 22066 19372
rect 27614 19320 27620 19372
rect 27672 19360 27678 19372
rect 34514 19360 34520 19372
rect 27672 19332 34520 19360
rect 27672 19320 27678 19332
rect 34514 19320 34520 19332
rect 34572 19320 34578 19372
rect 36096 19332 36492 19360
rect 2958 19252 2964 19304
rect 3016 19292 3022 19304
rect 3237 19295 3295 19301
rect 3237 19292 3249 19295
rect 3016 19264 3249 19292
rect 3016 19252 3022 19264
rect 3237 19261 3249 19264
rect 3283 19261 3295 19295
rect 3237 19255 3295 19261
rect 4065 19295 4123 19301
rect 4065 19261 4077 19295
rect 4111 19292 4123 19295
rect 4154 19292 4160 19304
rect 4111 19264 4160 19292
rect 4111 19261 4123 19264
rect 4065 19255 4123 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 5902 19292 5908 19304
rect 5863 19264 5908 19292
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6696 19264 6837 19292
rect 6696 19252 6702 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19261 8263 19295
rect 8205 19255 8263 19261
rect 6730 19184 6736 19236
rect 6788 19224 6794 19236
rect 8220 19224 8248 19255
rect 8294 19252 8300 19304
rect 8352 19252 8358 19304
rect 8757 19295 8815 19301
rect 8757 19261 8769 19295
rect 8803 19261 8815 19295
rect 8757 19255 8815 19261
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19292 8999 19295
rect 10134 19292 10140 19304
rect 8987 19264 10140 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 8772 19224 8800 19255
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 10873 19295 10931 19301
rect 10873 19261 10885 19295
rect 10919 19261 10931 19295
rect 10873 19255 10931 19261
rect 11241 19295 11299 19301
rect 11241 19261 11253 19295
rect 11287 19292 11299 19295
rect 11330 19292 11336 19304
rect 11287 19264 11336 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 6788 19196 8800 19224
rect 6788 19184 6794 19196
rect 3142 19116 3148 19168
rect 3200 19156 3206 19168
rect 4157 19159 4215 19165
rect 4157 19156 4169 19159
rect 3200 19128 4169 19156
rect 3200 19116 3206 19128
rect 4157 19125 4169 19128
rect 4203 19125 4215 19159
rect 4157 19119 4215 19125
rect 5721 19159 5779 19165
rect 5721 19125 5733 19159
rect 5767 19156 5779 19159
rect 6914 19156 6920 19168
rect 5767 19128 6920 19156
rect 5767 19125 5779 19128
rect 5721 19119 5779 19125
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7024 19165 7052 19196
rect 8846 19184 8852 19236
rect 8904 19224 8910 19236
rect 10704 19224 10732 19255
rect 8904 19196 10732 19224
rect 8904 19184 8910 19196
rect 7009 19159 7067 19165
rect 7009 19125 7021 19159
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 8662 19116 8668 19168
rect 8720 19156 8726 19168
rect 9217 19159 9275 19165
rect 9217 19156 9229 19159
rect 8720 19128 9229 19156
rect 8720 19116 8726 19128
rect 9217 19125 9229 19128
rect 9263 19125 9275 19159
rect 9217 19119 9275 19125
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 10888 19156 10916 19255
rect 11330 19252 11336 19264
rect 11388 19252 11394 19304
rect 11425 19295 11483 19301
rect 11425 19261 11437 19295
rect 11471 19292 11483 19295
rect 13078 19292 13084 19304
rect 11471 19264 13084 19292
rect 11471 19261 11483 19264
rect 11425 19255 11483 19261
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 15197 19295 15255 19301
rect 15197 19261 15209 19295
rect 15243 19292 15255 19295
rect 16298 19292 16304 19304
rect 15243 19264 16304 19292
rect 15243 19261 15255 19264
rect 15197 19255 15255 19261
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19292 17647 19295
rect 18325 19295 18383 19301
rect 17635 19264 17816 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 17788 19168 17816 19264
rect 18325 19261 18337 19295
rect 18371 19261 18383 19295
rect 18325 19255 18383 19261
rect 19337 19295 19395 19301
rect 19337 19261 19349 19295
rect 19383 19292 19395 19295
rect 19426 19292 19432 19304
rect 19383 19264 19432 19292
rect 19383 19261 19395 19264
rect 19337 19255 19395 19261
rect 18340 19168 18368 19255
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 19702 19292 19708 19304
rect 19663 19264 19708 19292
rect 19702 19252 19708 19264
rect 19760 19252 19766 19304
rect 21082 19292 21088 19304
rect 20995 19264 21088 19292
rect 21082 19252 21088 19264
rect 21140 19292 21146 19304
rect 21450 19292 21456 19304
rect 21140 19264 21456 19292
rect 21140 19252 21146 19264
rect 21450 19252 21456 19264
rect 21508 19252 21514 19304
rect 23658 19252 23664 19304
rect 23716 19292 23722 19304
rect 23845 19295 23903 19301
rect 23845 19292 23857 19295
rect 23716 19264 23857 19292
rect 23716 19252 23722 19264
rect 23845 19261 23857 19264
rect 23891 19261 23903 19295
rect 23845 19255 23903 19261
rect 9640 19128 10916 19156
rect 9640 19116 9646 19128
rect 13446 19116 13452 19168
rect 13504 19156 13510 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 13504 19128 15393 19156
rect 13504 19116 13510 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 15381 19119 15439 19125
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18322 19156 18328 19168
rect 18279 19128 18328 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 19444 19156 19472 19252
rect 23860 19224 23888 19255
rect 23934 19252 23940 19304
rect 23992 19292 23998 19304
rect 24397 19295 24455 19301
rect 23992 19264 24037 19292
rect 23992 19252 23998 19264
rect 24397 19261 24409 19295
rect 24443 19261 24455 19295
rect 24397 19255 24455 19261
rect 24581 19295 24639 19301
rect 24581 19261 24593 19295
rect 24627 19292 24639 19295
rect 25222 19292 25228 19304
rect 24627 19264 25228 19292
rect 24627 19261 24639 19264
rect 24581 19255 24639 19261
rect 24412 19224 24440 19255
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 25314 19252 25320 19304
rect 25372 19292 25378 19304
rect 26421 19295 26479 19301
rect 26421 19292 26433 19295
rect 25372 19264 26433 19292
rect 25372 19252 25378 19264
rect 26421 19261 26433 19264
rect 26467 19261 26479 19295
rect 26421 19255 26479 19261
rect 26605 19295 26663 19301
rect 26605 19261 26617 19295
rect 26651 19292 26663 19295
rect 27157 19295 27215 19301
rect 27157 19292 27169 19295
rect 26651 19264 27169 19292
rect 26651 19261 26663 19264
rect 26605 19255 26663 19261
rect 27157 19261 27169 19264
rect 27203 19261 27215 19295
rect 27157 19255 27215 19261
rect 27341 19295 27399 19301
rect 27341 19261 27353 19295
rect 27387 19292 27399 19295
rect 30006 19292 30012 19304
rect 27387 19264 30012 19292
rect 27387 19261 27399 19264
rect 27341 19255 27399 19261
rect 25866 19224 25872 19236
rect 23860 19196 25872 19224
rect 25866 19184 25872 19196
rect 25924 19224 25930 19236
rect 26620 19224 26648 19255
rect 30006 19252 30012 19264
rect 30064 19252 30070 19304
rect 30653 19295 30711 19301
rect 30653 19261 30665 19295
rect 30699 19292 30711 19295
rect 30742 19292 30748 19304
rect 30699 19264 30748 19292
rect 30699 19261 30711 19264
rect 30653 19255 30711 19261
rect 30742 19252 30748 19264
rect 30800 19252 30806 19304
rect 30837 19295 30895 19301
rect 30837 19261 30849 19295
rect 30883 19261 30895 19295
rect 30837 19255 30895 19261
rect 27706 19224 27712 19236
rect 25924 19196 26648 19224
rect 27667 19196 27712 19224
rect 25924 19184 25930 19196
rect 27706 19184 27712 19196
rect 27764 19184 27770 19236
rect 30852 19224 30880 19255
rect 31110 19252 31116 19304
rect 31168 19301 31174 19304
rect 31168 19295 31217 19301
rect 31168 19261 31171 19295
rect 31205 19261 31217 19295
rect 31294 19292 31300 19304
rect 31255 19264 31300 19292
rect 31168 19255 31217 19261
rect 31168 19252 31174 19255
rect 31294 19252 31300 19264
rect 31352 19252 31358 19304
rect 31386 19252 31392 19304
rect 31444 19292 31450 19304
rect 31444 19264 32260 19292
rect 31444 19252 31450 19264
rect 31938 19224 31944 19236
rect 30852 19196 31944 19224
rect 31938 19184 31944 19196
rect 31996 19184 32002 19236
rect 32232 19224 32260 19264
rect 32306 19252 32312 19304
rect 32364 19292 32370 19304
rect 36096 19292 36124 19332
rect 36262 19292 36268 19304
rect 32364 19264 36124 19292
rect 36223 19264 36268 19292
rect 32364 19252 32370 19264
rect 36262 19252 36268 19264
rect 36320 19252 36326 19304
rect 36357 19295 36415 19301
rect 36357 19261 36369 19295
rect 36403 19261 36415 19295
rect 36464 19292 36492 19332
rect 39390 19320 39396 19372
rect 39448 19360 39454 19372
rect 39666 19360 39672 19372
rect 39448 19332 39672 19360
rect 39448 19320 39454 19332
rect 39666 19320 39672 19332
rect 39724 19320 39730 19372
rect 46014 19360 46020 19372
rect 42812 19332 46020 19360
rect 36725 19295 36783 19301
rect 36725 19292 36737 19295
rect 36464 19264 36737 19292
rect 36357 19255 36415 19261
rect 36725 19261 36737 19264
rect 36771 19261 36783 19295
rect 36725 19255 36783 19261
rect 36170 19224 36176 19236
rect 32232 19196 36176 19224
rect 36170 19184 36176 19196
rect 36228 19184 36234 19236
rect 36372 19224 36400 19255
rect 36814 19252 36820 19304
rect 36872 19292 36878 19304
rect 36872 19264 36917 19292
rect 36872 19252 36878 19264
rect 37274 19252 37280 19304
rect 37332 19292 37338 19304
rect 38286 19292 38292 19304
rect 37332 19264 38292 19292
rect 37332 19252 37338 19264
rect 38286 19252 38292 19264
rect 38344 19252 38350 19304
rect 38378 19252 38384 19304
rect 38436 19292 38442 19304
rect 39301 19295 39359 19301
rect 38436 19264 38481 19292
rect 38436 19252 38442 19264
rect 39301 19261 39313 19295
rect 39347 19292 39359 19295
rect 39758 19292 39764 19304
rect 39347 19264 39764 19292
rect 39347 19261 39359 19264
rect 39301 19255 39359 19261
rect 39758 19252 39764 19264
rect 39816 19252 39822 19304
rect 41414 19252 41420 19304
rect 41472 19292 41478 19304
rect 41877 19295 41935 19301
rect 41877 19292 41889 19295
rect 41472 19264 41889 19292
rect 41472 19252 41478 19264
rect 41877 19261 41889 19264
rect 41923 19261 41935 19295
rect 41877 19255 41935 19261
rect 41969 19295 42027 19301
rect 41969 19261 41981 19295
rect 42015 19261 42027 19295
rect 42334 19292 42340 19304
rect 42295 19264 42340 19292
rect 41969 19255 42027 19261
rect 37829 19227 37887 19233
rect 37829 19224 37841 19227
rect 36372 19196 37841 19224
rect 37829 19193 37841 19196
rect 37875 19224 37887 19227
rect 41598 19224 41604 19236
rect 37875 19196 41604 19224
rect 37875 19193 37887 19196
rect 37829 19187 37887 19193
rect 41598 19184 41604 19196
rect 41656 19184 41662 19236
rect 20714 19156 20720 19168
rect 19444 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 24210 19116 24216 19168
rect 24268 19156 24274 19168
rect 24857 19159 24915 19165
rect 24857 19156 24869 19159
rect 24268 19128 24869 19156
rect 24268 19116 24274 19128
rect 24857 19125 24869 19128
rect 24903 19125 24915 19159
rect 32398 19156 32404 19168
rect 32311 19128 32404 19156
rect 24857 19119 24915 19125
rect 32398 19116 32404 19128
rect 32456 19156 32462 19168
rect 32766 19156 32772 19168
rect 32456 19128 32772 19156
rect 32456 19116 32462 19128
rect 32766 19116 32772 19128
rect 32824 19116 32830 19168
rect 37274 19156 37280 19168
rect 37235 19128 37280 19156
rect 37274 19116 37280 19128
rect 37332 19116 37338 19168
rect 37642 19156 37648 19168
rect 37603 19128 37648 19156
rect 37642 19116 37648 19128
rect 37700 19116 37706 19168
rect 38746 19116 38752 19168
rect 38804 19156 38810 19168
rect 39393 19159 39451 19165
rect 39393 19156 39405 19159
rect 38804 19128 39405 19156
rect 38804 19116 38810 19128
rect 39393 19125 39405 19128
rect 39439 19125 39451 19159
rect 39393 19119 39451 19125
rect 39669 19159 39727 19165
rect 39669 19125 39681 19159
rect 39715 19156 39727 19159
rect 39758 19156 39764 19168
rect 39715 19128 39764 19156
rect 39715 19125 39727 19128
rect 39669 19119 39727 19125
rect 39758 19116 39764 19128
rect 39816 19156 39822 19168
rect 41322 19156 41328 19168
rect 39816 19128 41328 19156
rect 39816 19116 39822 19128
rect 41322 19116 41328 19128
rect 41380 19116 41386 19168
rect 41892 19156 41920 19255
rect 41984 19224 42012 19255
rect 42334 19252 42340 19264
rect 42392 19252 42398 19304
rect 42426 19252 42432 19304
rect 42484 19292 42490 19304
rect 42812 19292 42840 19332
rect 46014 19320 46020 19332
rect 46072 19320 46078 19372
rect 48498 19320 48504 19372
rect 48556 19360 48562 19372
rect 49234 19360 49240 19372
rect 48556 19332 49240 19360
rect 48556 19320 48562 19332
rect 42484 19264 42840 19292
rect 42484 19252 42490 19264
rect 44174 19252 44180 19304
rect 44232 19292 44238 19304
rect 44818 19292 44824 19304
rect 44232 19264 44824 19292
rect 44232 19252 44238 19264
rect 44818 19252 44824 19264
rect 44876 19292 44882 19304
rect 45005 19295 45063 19301
rect 45005 19292 45017 19295
rect 44876 19264 45017 19292
rect 44876 19252 44882 19264
rect 45005 19261 45017 19264
rect 45051 19261 45063 19295
rect 46106 19292 46112 19304
rect 46067 19264 46112 19292
rect 45005 19255 45063 19261
rect 46106 19252 46112 19264
rect 46164 19292 46170 19304
rect 46385 19295 46443 19301
rect 46385 19292 46397 19295
rect 46164 19264 46397 19292
rect 46164 19252 46170 19264
rect 46385 19261 46397 19264
rect 46431 19292 46443 19295
rect 47854 19292 47860 19304
rect 46431 19264 47860 19292
rect 46431 19261 46443 19264
rect 46385 19255 46443 19261
rect 47854 19252 47860 19264
rect 47912 19252 47918 19304
rect 47949 19295 48007 19301
rect 47949 19261 47961 19295
rect 47995 19292 48007 19295
rect 48406 19292 48412 19304
rect 47995 19264 48412 19292
rect 47995 19261 48007 19264
rect 47949 19255 48007 19261
rect 48406 19252 48412 19264
rect 48464 19252 48470 19304
rect 48590 19292 48596 19304
rect 48551 19264 48596 19292
rect 48590 19252 48596 19264
rect 48648 19252 48654 19304
rect 48976 19301 49004 19332
rect 49234 19320 49240 19332
rect 49292 19320 49298 19372
rect 52454 19360 52460 19372
rect 52104 19332 52460 19360
rect 48685 19295 48743 19301
rect 48685 19261 48697 19295
rect 48731 19261 48743 19295
rect 48685 19255 48743 19261
rect 48961 19295 49019 19301
rect 48961 19261 48973 19295
rect 49007 19261 49019 19295
rect 48961 19255 49019 19261
rect 44082 19224 44088 19236
rect 41984 19196 44088 19224
rect 44082 19184 44088 19196
rect 44140 19184 44146 19236
rect 45097 19227 45155 19233
rect 45097 19193 45109 19227
rect 45143 19224 45155 19227
rect 46750 19224 46756 19236
rect 45143 19196 46756 19224
rect 45143 19193 45155 19196
rect 45097 19187 45155 19193
rect 46124 19168 46152 19196
rect 46750 19184 46756 19196
rect 46808 19184 46814 19236
rect 47118 19184 47124 19236
rect 47176 19224 47182 19236
rect 48700 19224 48728 19255
rect 49050 19252 49056 19304
rect 49108 19292 49114 19304
rect 49973 19295 50031 19301
rect 49108 19264 49153 19292
rect 49108 19252 49114 19264
rect 49973 19261 49985 19295
rect 50019 19292 50031 19295
rect 50706 19292 50712 19304
rect 50019 19264 50712 19292
rect 50019 19261 50031 19264
rect 49973 19255 50031 19261
rect 50706 19252 50712 19264
rect 50764 19252 50770 19304
rect 52104 19301 52132 19332
rect 52454 19320 52460 19332
rect 52512 19320 52518 19372
rect 52089 19295 52147 19301
rect 52089 19261 52101 19295
rect 52135 19261 52147 19295
rect 53285 19295 53343 19301
rect 53285 19292 53297 19295
rect 52089 19255 52147 19261
rect 52196 19264 53297 19292
rect 47176 19196 48728 19224
rect 47176 19184 47182 19196
rect 49602 19184 49608 19236
rect 49660 19224 49666 19236
rect 51905 19227 51963 19233
rect 51905 19224 51917 19227
rect 49660 19196 51917 19224
rect 49660 19184 49666 19196
rect 51905 19193 51917 19196
rect 51951 19224 51963 19227
rect 52196 19224 52224 19264
rect 53285 19261 53297 19264
rect 53331 19261 53343 19295
rect 53285 19255 53343 19261
rect 51951 19196 52224 19224
rect 52457 19227 52515 19233
rect 51951 19193 51963 19196
rect 51905 19187 51963 19193
rect 52457 19193 52469 19227
rect 52503 19224 52515 19227
rect 52638 19224 52644 19236
rect 52503 19196 52644 19224
rect 52503 19193 52515 19196
rect 52457 19187 52515 19193
rect 52638 19184 52644 19196
rect 52696 19184 52702 19236
rect 42426 19156 42432 19168
rect 41892 19128 42432 19156
rect 42426 19116 42432 19128
rect 42484 19116 42490 19168
rect 42518 19116 42524 19168
rect 42576 19156 42582 19168
rect 43165 19159 43223 19165
rect 43165 19156 43177 19159
rect 42576 19128 43177 19156
rect 42576 19116 42582 19128
rect 43165 19125 43177 19128
rect 43211 19125 43223 19159
rect 43165 19119 43223 19125
rect 46106 19116 46112 19168
rect 46164 19116 46170 19168
rect 46198 19116 46204 19168
rect 46256 19156 46262 19168
rect 46658 19156 46664 19168
rect 46256 19128 46664 19156
rect 46256 19116 46262 19128
rect 46658 19116 46664 19128
rect 46716 19116 46722 19168
rect 49234 19116 49240 19168
rect 49292 19156 49298 19168
rect 50065 19159 50123 19165
rect 50065 19156 50077 19159
rect 49292 19128 50077 19156
rect 49292 19116 49298 19128
rect 50065 19125 50077 19128
rect 50111 19125 50123 19159
rect 53374 19156 53380 19168
rect 53335 19128 53380 19156
rect 50065 19119 50123 19125
rect 53374 19116 53380 19128
rect 53432 19116 53438 19168
rect 1104 19066 54832 19088
rect 1104 19014 18912 19066
rect 18964 19014 18976 19066
rect 19028 19014 19040 19066
rect 19092 19014 19104 19066
rect 19156 19014 36843 19066
rect 36895 19014 36907 19066
rect 36959 19014 36971 19066
rect 37023 19014 37035 19066
rect 37087 19014 54832 19066
rect 1104 18992 54832 19014
rect 2958 18952 2964 18964
rect 2919 18924 2964 18952
rect 2958 18912 2964 18924
rect 3016 18912 3022 18964
rect 9953 18955 10011 18961
rect 9953 18921 9965 18955
rect 9999 18952 10011 18955
rect 10318 18952 10324 18964
rect 9999 18924 10324 18952
rect 9999 18921 10011 18924
rect 9953 18915 10011 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 17218 18952 17224 18964
rect 16632 18924 17224 18952
rect 16632 18912 16638 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 17497 18955 17555 18961
rect 17497 18921 17509 18955
rect 17543 18952 17555 18955
rect 18046 18952 18052 18964
rect 17543 18924 18052 18952
rect 17543 18921 17555 18924
rect 17497 18915 17555 18921
rect 4341 18887 4399 18893
rect 4341 18853 4353 18887
rect 4387 18884 4399 18887
rect 5074 18884 5080 18896
rect 4387 18856 5080 18884
rect 4387 18853 4399 18856
rect 4341 18847 4399 18853
rect 5074 18844 5080 18856
rect 5132 18884 5138 18896
rect 5132 18856 7144 18884
rect 5132 18844 5138 18856
rect 3142 18816 3148 18828
rect 3103 18788 3148 18816
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 4246 18816 4252 18828
rect 4207 18788 4252 18816
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 6365 18819 6423 18825
rect 6365 18785 6377 18819
rect 6411 18816 6423 18819
rect 6730 18816 6736 18828
rect 6411 18788 6736 18816
rect 6411 18785 6423 18788
rect 6365 18779 6423 18785
rect 6730 18776 6736 18788
rect 6788 18816 6794 18828
rect 7116 18825 7144 18856
rect 9582 18844 9588 18896
rect 9640 18884 9646 18896
rect 9640 18856 10364 18884
rect 9640 18844 9646 18856
rect 6917 18819 6975 18825
rect 6917 18816 6929 18819
rect 6788 18788 6929 18816
rect 6788 18776 6794 18788
rect 6917 18785 6929 18788
rect 6963 18785 6975 18819
rect 6917 18779 6975 18785
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 8846 18816 8852 18828
rect 7147 18788 8852 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 10134 18816 10140 18828
rect 10095 18788 10140 18816
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 10336 18825 10364 18856
rect 10888 18856 13676 18884
rect 10888 18825 10916 18856
rect 10321 18819 10379 18825
rect 10321 18785 10333 18819
rect 10367 18785 10379 18819
rect 10321 18779 10379 18785
rect 10689 18819 10747 18825
rect 10689 18785 10701 18819
rect 10735 18785 10747 18819
rect 10689 18779 10747 18785
rect 10873 18819 10931 18825
rect 10873 18785 10885 18819
rect 10919 18785 10931 18819
rect 10873 18779 10931 18785
rect 12897 18819 12955 18825
rect 12897 18785 12909 18819
rect 12943 18816 12955 18819
rect 13262 18816 13268 18828
rect 12943 18788 13268 18816
rect 12943 18785 12955 18788
rect 12897 18779 12955 18785
rect 6089 18751 6147 18757
rect 6089 18717 6101 18751
rect 6135 18748 6147 18751
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 6135 18720 6285 18748
rect 6135 18717 6147 18720
rect 6089 18711 6147 18717
rect 6273 18717 6285 18720
rect 6319 18717 6331 18751
rect 10704 18748 10732 18779
rect 13262 18776 13268 18788
rect 13320 18816 13326 18828
rect 13446 18816 13452 18828
rect 13320 18788 13452 18816
rect 13320 18776 13326 18788
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 13648 18825 13676 18856
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 13814 18816 13820 18828
rect 13679 18788 13820 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 15841 18819 15899 18825
rect 15841 18816 15853 18819
rect 15804 18788 15853 18816
rect 15804 18776 15810 18788
rect 15841 18785 15853 18788
rect 15887 18785 15899 18819
rect 15841 18779 15899 18785
rect 17037 18819 17095 18825
rect 17037 18785 17049 18819
rect 17083 18816 17095 18819
rect 17512 18816 17540 18915
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 25498 18952 25504 18964
rect 25459 18924 25504 18952
rect 25498 18912 25504 18924
rect 25556 18912 25562 18964
rect 29178 18912 29184 18964
rect 29236 18952 29242 18964
rect 29733 18955 29791 18961
rect 29733 18952 29745 18955
rect 29236 18924 29745 18952
rect 29236 18912 29242 18924
rect 29733 18921 29745 18924
rect 29779 18952 29791 18955
rect 29914 18952 29920 18964
rect 29779 18924 29920 18952
rect 29779 18921 29791 18924
rect 29733 18915 29791 18921
rect 29914 18912 29920 18924
rect 29972 18912 29978 18964
rect 31864 18924 33640 18952
rect 29273 18887 29331 18893
rect 29273 18853 29285 18887
rect 29319 18884 29331 18887
rect 31864 18884 31892 18924
rect 33502 18884 33508 18896
rect 29319 18856 31892 18884
rect 32140 18856 32812 18884
rect 29319 18853 29331 18856
rect 29273 18847 29331 18853
rect 17083 18788 17540 18816
rect 21729 18819 21787 18825
rect 17083 18785 17095 18788
rect 17037 18779 17095 18785
rect 21729 18785 21741 18819
rect 21775 18816 21787 18819
rect 24210 18816 24216 18828
rect 21775 18788 24072 18816
rect 24171 18788 24216 18816
rect 21775 18785 21787 18788
rect 21729 18779 21787 18785
rect 11330 18748 11336 18760
rect 10704 18720 11336 18748
rect 6273 18711 6331 18717
rect 6288 18680 6316 18711
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 12713 18751 12771 18757
rect 12713 18748 12725 18751
rect 12452 18720 12725 18748
rect 6914 18680 6920 18692
rect 6288 18652 6920 18680
rect 6914 18640 6920 18652
rect 6972 18640 6978 18692
rect 7374 18612 7380 18624
rect 7335 18584 7380 18612
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 12452 18612 12480 18720
rect 12713 18717 12725 18720
rect 12759 18717 12771 18751
rect 12713 18711 12771 18717
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 15749 18683 15807 18689
rect 12676 18652 15148 18680
rect 12676 18640 12682 18652
rect 9732 18584 12480 18612
rect 13909 18615 13967 18621
rect 9732 18572 9738 18584
rect 13909 18581 13921 18615
rect 13955 18612 13967 18615
rect 15010 18612 15016 18624
rect 13955 18584 15016 18612
rect 13955 18581 13967 18584
rect 13909 18575 13967 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15120 18612 15148 18652
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 15856 18680 15884 18779
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 21048 18720 23765 18748
rect 21048 18708 21054 18720
rect 23753 18717 23765 18720
rect 23799 18748 23811 18751
rect 23937 18751 23995 18757
rect 23937 18748 23949 18751
rect 23799 18720 23949 18748
rect 23799 18717 23811 18720
rect 23753 18711 23811 18717
rect 23937 18717 23949 18720
rect 23983 18717 23995 18751
rect 24044 18748 24072 18788
rect 24210 18776 24216 18788
rect 24268 18776 24274 18828
rect 25498 18776 25504 18828
rect 25556 18816 25562 18828
rect 26513 18819 26571 18825
rect 26513 18816 26525 18819
rect 25556 18788 26525 18816
rect 25556 18776 25562 18788
rect 26513 18785 26525 18788
rect 26559 18785 26571 18819
rect 28350 18816 28356 18828
rect 28311 18788 28356 18816
rect 26513 18779 26571 18785
rect 28350 18776 28356 18788
rect 28408 18776 28414 18828
rect 25958 18748 25964 18760
rect 24044 18720 25964 18748
rect 23937 18711 23995 18717
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 28721 18751 28779 18757
rect 28721 18717 28733 18751
rect 28767 18748 28779 18751
rect 29288 18748 29316 18847
rect 29914 18816 29920 18828
rect 29875 18788 29920 18816
rect 29914 18776 29920 18788
rect 29972 18776 29978 18828
rect 30006 18776 30012 18828
rect 30064 18816 30070 18828
rect 32140 18816 32168 18856
rect 32306 18816 32312 18828
rect 30064 18788 30109 18816
rect 31864 18788 32168 18816
rect 32267 18788 32312 18816
rect 30064 18776 30070 18788
rect 28767 18720 29316 18748
rect 29932 18748 29960 18776
rect 31864 18757 31892 18788
rect 32306 18776 32312 18788
rect 32364 18776 32370 18828
rect 32398 18776 32404 18828
rect 32456 18816 32462 18828
rect 32784 18825 32812 18856
rect 32876 18856 33508 18884
rect 32876 18825 32904 18856
rect 33502 18844 33508 18856
rect 33560 18844 33566 18896
rect 33612 18884 33640 18924
rect 33686 18912 33692 18964
rect 33744 18952 33750 18964
rect 36170 18952 36176 18964
rect 33744 18924 33789 18952
rect 36131 18924 36176 18952
rect 33744 18912 33750 18924
rect 36170 18912 36176 18924
rect 36228 18912 36234 18964
rect 36262 18912 36268 18964
rect 36320 18952 36326 18964
rect 37642 18952 37648 18964
rect 36320 18924 37648 18952
rect 36320 18912 36326 18924
rect 37642 18912 37648 18924
rect 37700 18952 37706 18964
rect 41506 18952 41512 18964
rect 37700 18924 41512 18952
rect 37700 18912 37706 18924
rect 41506 18912 41512 18924
rect 41564 18912 41570 18964
rect 41690 18952 41696 18964
rect 41651 18924 41696 18952
rect 41690 18912 41696 18924
rect 41748 18912 41754 18964
rect 48590 18912 48596 18964
rect 48648 18952 48654 18964
rect 53374 18952 53380 18964
rect 48648 18924 53380 18952
rect 48648 18912 48654 18924
rect 33612 18856 39712 18884
rect 32769 18819 32827 18825
rect 32456 18788 32501 18816
rect 32456 18776 32462 18788
rect 32769 18785 32781 18819
rect 32815 18785 32827 18819
rect 32769 18779 32827 18785
rect 32861 18819 32919 18825
rect 32861 18785 32873 18819
rect 32907 18785 32919 18819
rect 32861 18779 32919 18785
rect 36170 18776 36176 18828
rect 36228 18816 36234 18828
rect 36541 18819 36599 18825
rect 36541 18816 36553 18819
rect 36228 18788 36553 18816
rect 36228 18776 36234 18788
rect 36541 18785 36553 18788
rect 36587 18785 36599 18819
rect 36541 18779 36599 18785
rect 36722 18776 36728 18828
rect 36780 18816 36786 18828
rect 38749 18819 38807 18825
rect 36780 18788 38700 18816
rect 36780 18776 36786 18788
rect 31849 18751 31907 18757
rect 31849 18748 31861 18751
rect 29932 18720 31861 18748
rect 28767 18717 28779 18720
rect 28721 18711 28779 18717
rect 31849 18717 31861 18720
rect 31895 18717 31907 18751
rect 31849 18711 31907 18717
rect 33413 18751 33471 18757
rect 33413 18717 33425 18751
rect 33459 18748 33471 18751
rect 33594 18748 33600 18760
rect 33459 18720 33600 18748
rect 33459 18717 33471 18720
rect 33413 18711 33471 18717
rect 33594 18708 33600 18720
rect 33652 18708 33658 18760
rect 33686 18708 33692 18760
rect 33744 18748 33750 18760
rect 34330 18748 34336 18760
rect 33744 18720 34336 18748
rect 33744 18708 33750 18720
rect 34330 18708 34336 18720
rect 34388 18748 34394 18760
rect 38197 18751 38255 18757
rect 38197 18748 38209 18751
rect 34388 18720 38209 18748
rect 34388 18708 34394 18720
rect 38197 18717 38209 18720
rect 38243 18717 38255 18751
rect 38197 18711 38255 18717
rect 38565 18751 38623 18757
rect 38565 18717 38577 18751
rect 38611 18717 38623 18751
rect 38672 18748 38700 18788
rect 38749 18785 38761 18819
rect 38795 18816 38807 18819
rect 38838 18816 38844 18828
rect 38795 18788 38844 18816
rect 38795 18785 38807 18788
rect 38749 18779 38807 18785
rect 38838 18776 38844 18788
rect 38896 18776 38902 18828
rect 39298 18816 39304 18828
rect 39259 18788 39304 18816
rect 39298 18776 39304 18788
rect 39356 18776 39362 18828
rect 39482 18816 39488 18828
rect 39443 18788 39488 18816
rect 39482 18776 39488 18788
rect 39540 18776 39546 18828
rect 39684 18748 39712 18856
rect 39850 18844 39856 18896
rect 39908 18884 39914 18896
rect 39908 18856 39953 18884
rect 39908 18844 39914 18856
rect 40034 18844 40040 18896
rect 40092 18884 40098 18896
rect 41969 18887 42027 18893
rect 41969 18884 41981 18887
rect 40092 18856 41981 18884
rect 40092 18844 40098 18856
rect 41969 18853 41981 18856
rect 42015 18884 42027 18887
rect 49602 18884 49608 18896
rect 42015 18856 44588 18884
rect 49563 18856 49608 18884
rect 42015 18853 42027 18856
rect 41969 18847 42027 18853
rect 41690 18776 41696 18828
rect 41748 18816 41754 18828
rect 41877 18819 41935 18825
rect 41877 18816 41889 18819
rect 41748 18788 41889 18816
rect 41748 18776 41754 18788
rect 41877 18785 41889 18788
rect 41923 18785 41935 18819
rect 41877 18779 41935 18785
rect 44085 18819 44143 18825
rect 44085 18785 44097 18819
rect 44131 18816 44143 18819
rect 44450 18816 44456 18828
rect 44131 18788 44456 18816
rect 44131 18785 44143 18788
rect 44085 18779 44143 18785
rect 44450 18776 44456 18788
rect 44508 18776 44514 18828
rect 44560 18825 44588 18856
rect 49602 18844 49608 18856
rect 49660 18844 49666 18896
rect 44545 18819 44603 18825
rect 44545 18785 44557 18819
rect 44591 18785 44603 18819
rect 44545 18779 44603 18785
rect 44634 18776 44640 18828
rect 44692 18816 44698 18828
rect 47854 18816 47860 18828
rect 44692 18788 44737 18816
rect 47815 18788 47860 18816
rect 44692 18776 44698 18788
rect 47854 18776 47860 18788
rect 47912 18816 47918 18828
rect 48133 18819 48191 18825
rect 48133 18816 48145 18819
rect 47912 18788 48145 18816
rect 47912 18776 47918 18788
rect 48133 18785 48145 18788
rect 48179 18816 48191 18819
rect 48866 18816 48872 18828
rect 48179 18788 48872 18816
rect 48179 18785 48191 18788
rect 48133 18779 48191 18785
rect 48866 18776 48872 18788
rect 48924 18776 48930 18828
rect 49050 18816 49056 18828
rect 49011 18788 49056 18816
rect 49050 18776 49056 18788
rect 49108 18776 49114 18828
rect 49234 18816 49240 18828
rect 49195 18788 49240 18816
rect 49234 18776 49240 18788
rect 49292 18776 49298 18828
rect 49970 18776 49976 18828
rect 50028 18816 50034 18828
rect 50617 18819 50675 18825
rect 50617 18816 50629 18819
rect 50028 18788 50629 18816
rect 50028 18776 50034 18788
rect 50617 18785 50629 18788
rect 50663 18816 50675 18819
rect 50709 18819 50767 18825
rect 50709 18816 50721 18819
rect 50663 18788 50721 18816
rect 50663 18785 50675 18788
rect 50617 18779 50675 18785
rect 50709 18785 50721 18788
rect 50755 18785 50767 18819
rect 50709 18779 50767 18785
rect 50893 18819 50951 18825
rect 50893 18785 50905 18819
rect 50939 18785 50951 18819
rect 51350 18816 51356 18828
rect 51311 18788 51356 18816
rect 50893 18779 50951 18785
rect 43993 18751 44051 18757
rect 38672 18720 38746 18748
rect 39684 18720 39804 18748
rect 38565 18711 38623 18717
rect 18322 18680 18328 18692
rect 15795 18652 18328 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 18322 18640 18328 18652
rect 18380 18680 18386 18692
rect 18380 18652 23060 18680
rect 18380 18640 18386 18652
rect 16025 18615 16083 18621
rect 16025 18612 16037 18615
rect 15120 18584 16037 18612
rect 16025 18581 16037 18584
rect 16071 18581 16083 18615
rect 16025 18575 16083 18581
rect 21358 18572 21364 18624
rect 21416 18612 21422 18624
rect 21821 18615 21879 18621
rect 21821 18612 21833 18615
rect 21416 18584 21833 18612
rect 21416 18572 21422 18584
rect 21821 18581 21833 18584
rect 21867 18581 21879 18615
rect 23032 18612 23060 18652
rect 25222 18640 25228 18692
rect 25280 18680 25286 18692
rect 26605 18683 26663 18689
rect 26605 18680 26617 18683
rect 25280 18652 26617 18680
rect 25280 18640 25286 18652
rect 26605 18649 26617 18652
rect 26651 18649 26663 18683
rect 26605 18643 26663 18649
rect 28629 18683 28687 18689
rect 28629 18649 28641 18683
rect 28675 18680 28687 18683
rect 36446 18680 36452 18692
rect 28675 18652 36452 18680
rect 28675 18649 28687 18652
rect 28629 18643 28687 18649
rect 36446 18640 36452 18652
rect 36504 18640 36510 18692
rect 26694 18612 26700 18624
rect 23032 18584 26700 18612
rect 21821 18575 21879 18581
rect 26694 18572 26700 18584
rect 26752 18572 26758 18624
rect 27338 18572 27344 18624
rect 27396 18612 27402 18624
rect 28491 18615 28549 18621
rect 28491 18612 28503 18615
rect 27396 18584 28503 18612
rect 27396 18572 27402 18584
rect 28491 18581 28503 18584
rect 28537 18581 28549 18615
rect 28994 18612 29000 18624
rect 28955 18584 29000 18612
rect 28491 18575 28549 18581
rect 28994 18572 29000 18584
rect 29052 18572 29058 18624
rect 29270 18572 29276 18624
rect 29328 18612 29334 18624
rect 33686 18612 33692 18624
rect 29328 18584 33692 18612
rect 29328 18572 29334 18584
rect 33686 18572 33692 18584
rect 33744 18572 33750 18624
rect 33870 18612 33876 18624
rect 33831 18584 33876 18612
rect 33870 18572 33876 18584
rect 33928 18572 33934 18624
rect 36357 18615 36415 18621
rect 36357 18581 36369 18615
rect 36403 18612 36415 18615
rect 37366 18612 37372 18624
rect 36403 18584 37372 18612
rect 36403 18581 36415 18584
rect 36357 18575 36415 18581
rect 37366 18572 37372 18584
rect 37424 18572 37430 18624
rect 38212 18612 38240 18711
rect 38286 18640 38292 18692
rect 38344 18680 38350 18692
rect 38381 18683 38439 18689
rect 38381 18680 38393 18683
rect 38344 18652 38393 18680
rect 38344 18640 38350 18652
rect 38381 18649 38393 18652
rect 38427 18680 38439 18683
rect 38580 18680 38608 18711
rect 38427 18652 38608 18680
rect 38718 18680 38746 18720
rect 39776 18680 39804 18720
rect 43993 18717 44005 18751
rect 44039 18748 44051 18751
rect 44174 18748 44180 18760
rect 44039 18720 44180 18748
rect 44039 18717 44051 18720
rect 43993 18711 44051 18717
rect 44174 18708 44180 18720
rect 44232 18708 44238 18760
rect 46934 18708 46940 18760
rect 46992 18748 46998 18760
rect 50908 18748 50936 18779
rect 51350 18776 51356 18788
rect 51408 18776 51414 18828
rect 51445 18819 51503 18825
rect 51445 18785 51457 18819
rect 51491 18816 51503 18819
rect 52454 18816 52460 18828
rect 51491 18788 52460 18816
rect 51491 18785 51503 18788
rect 51445 18779 51503 18785
rect 52454 18776 52460 18788
rect 52512 18776 52518 18828
rect 52932 18825 52960 18924
rect 53374 18912 53380 18924
rect 53432 18912 53438 18964
rect 52917 18819 52975 18825
rect 52917 18785 52929 18819
rect 52963 18785 52975 18819
rect 52917 18779 52975 18785
rect 53101 18819 53159 18825
rect 53101 18785 53113 18819
rect 53147 18816 53159 18819
rect 53282 18816 53288 18828
rect 53147 18788 53288 18816
rect 53147 18785 53159 18788
rect 53101 18779 53159 18785
rect 53282 18776 53288 18788
rect 53340 18776 53346 18828
rect 46992 18720 50936 18748
rect 46992 18708 46998 18720
rect 44450 18680 44456 18692
rect 38718 18652 39712 18680
rect 39776 18652 44456 18680
rect 38427 18649 38439 18652
rect 38381 18643 38439 18649
rect 38838 18612 38844 18624
rect 38212 18584 38844 18612
rect 38838 18572 38844 18584
rect 38896 18572 38902 18624
rect 39114 18572 39120 18624
rect 39172 18612 39178 18624
rect 39574 18612 39580 18624
rect 39172 18584 39580 18612
rect 39172 18572 39178 18584
rect 39574 18572 39580 18584
rect 39632 18572 39638 18624
rect 39684 18612 39712 18652
rect 44450 18640 44456 18652
rect 44508 18640 44514 18692
rect 45002 18680 45008 18692
rect 44963 18652 45008 18680
rect 45002 18640 45008 18652
rect 45060 18640 45066 18692
rect 45646 18640 45652 18692
rect 45704 18680 45710 18692
rect 51813 18683 51871 18689
rect 51813 18680 51825 18683
rect 45704 18652 51825 18680
rect 45704 18640 45710 18652
rect 51813 18649 51825 18652
rect 51859 18649 51871 18683
rect 51813 18643 51871 18649
rect 40218 18612 40224 18624
rect 39684 18584 40224 18612
rect 40218 18572 40224 18584
rect 40276 18572 40282 18624
rect 41506 18572 41512 18624
rect 41564 18612 41570 18624
rect 47946 18612 47952 18624
rect 41564 18584 47952 18612
rect 41564 18572 41570 18584
rect 47946 18572 47952 18584
rect 48004 18572 48010 18624
rect 52546 18572 52552 18624
rect 52604 18612 52610 18624
rect 53193 18615 53251 18621
rect 53193 18612 53205 18615
rect 52604 18584 53205 18612
rect 52604 18572 52610 18584
rect 53193 18581 53205 18584
rect 53239 18581 53251 18615
rect 53193 18575 53251 18581
rect 1104 18522 54832 18544
rect 1104 18470 9947 18522
rect 9999 18470 10011 18522
rect 10063 18470 10075 18522
rect 10127 18470 10139 18522
rect 10191 18470 27878 18522
rect 27930 18470 27942 18522
rect 27994 18470 28006 18522
rect 28058 18470 28070 18522
rect 28122 18470 45808 18522
rect 45860 18470 45872 18522
rect 45924 18470 45936 18522
rect 45988 18470 46000 18522
rect 46052 18470 54832 18522
rect 1104 18448 54832 18470
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 8110 18408 8116 18420
rect 6972 18380 8116 18408
rect 6972 18368 6978 18380
rect 8110 18368 8116 18380
rect 8168 18408 8174 18420
rect 8168 18380 9352 18408
rect 8168 18368 8174 18380
rect 4154 18340 4160 18352
rect 4115 18312 4160 18340
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 9324 18340 9352 18380
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10376 18380 10977 18408
rect 10376 18368 10382 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 13078 18368 13084 18420
rect 13136 18408 13142 18420
rect 13136 18380 17724 18408
rect 13136 18368 13142 18380
rect 12253 18343 12311 18349
rect 12253 18340 12265 18343
rect 9324 18312 12265 18340
rect 12253 18309 12265 18312
rect 12299 18340 12311 18343
rect 17696 18340 17724 18380
rect 17770 18368 17776 18420
rect 17828 18408 17834 18420
rect 17828 18380 22048 18408
rect 17828 18368 17834 18380
rect 18046 18340 18052 18352
rect 12299 18312 12480 18340
rect 17696 18312 18052 18340
rect 12299 18309 12311 18312
rect 12253 18303 12311 18309
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 7374 18272 7380 18284
rect 1903 18244 7380 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 8662 18272 8668 18284
rect 8623 18244 8668 18272
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 12452 18281 12480 18312
rect 18046 18300 18052 18312
rect 18104 18300 18110 18352
rect 19889 18343 19947 18349
rect 19889 18309 19901 18343
rect 19935 18340 19947 18343
rect 20990 18340 20996 18352
rect 19935 18312 20996 18340
rect 19935 18309 19947 18312
rect 19889 18303 19947 18309
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 13725 18275 13783 18281
rect 13725 18241 13737 18275
rect 13771 18272 13783 18275
rect 15010 18272 15016 18284
rect 13771 18244 14872 18272
rect 14971 18244 15016 18272
rect 13771 18241 13783 18244
rect 13725 18235 13783 18241
rect 1581 18207 1639 18213
rect 1581 18173 1593 18207
rect 1627 18204 1639 18207
rect 2866 18204 2872 18216
rect 1627 18176 2872 18204
rect 1627 18173 1639 18176
rect 1581 18167 1639 18173
rect 2866 18164 2872 18176
rect 2924 18204 2930 18216
rect 3329 18207 3387 18213
rect 3329 18204 3341 18207
rect 2924 18176 3341 18204
rect 2924 18164 2930 18176
rect 3329 18173 3341 18176
rect 3375 18173 3387 18207
rect 4338 18204 4344 18216
rect 4299 18176 4344 18204
rect 3329 18167 3387 18173
rect 4338 18164 4344 18176
rect 4396 18164 4402 18216
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18173 4675 18207
rect 5074 18204 5080 18216
rect 5035 18176 5080 18204
rect 4617 18167 4675 18173
rect 3237 18139 3295 18145
rect 3237 18105 3249 18139
rect 3283 18136 3295 18139
rect 4246 18136 4252 18148
rect 3283 18108 4252 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 4246 18096 4252 18108
rect 4304 18136 4310 18148
rect 4632 18136 4660 18167
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5258 18204 5264 18216
rect 5219 18176 5264 18204
rect 5258 18164 5264 18176
rect 5316 18164 5322 18216
rect 6822 18204 6828 18216
rect 6783 18176 6828 18204
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 8386 18204 8392 18216
rect 8347 18176 8392 18204
rect 8386 18164 8392 18176
rect 8444 18204 8450 18216
rect 8444 18176 9352 18204
rect 8444 18164 8450 18176
rect 4304 18108 4660 18136
rect 9324 18136 9352 18176
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 9732 18176 10057 18204
rect 9732 18164 9738 18176
rect 10045 18173 10057 18176
rect 10091 18204 10103 18207
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 10091 18176 10885 18204
rect 10091 18173 10103 18176
rect 10045 18167 10103 18173
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18173 12679 18207
rect 13078 18204 13084 18216
rect 13039 18176 13084 18204
rect 12621 18167 12679 18173
rect 10137 18139 10195 18145
rect 10137 18136 10149 18139
rect 9324 18108 10149 18136
rect 4304 18096 4310 18108
rect 10137 18105 10149 18108
rect 10183 18105 10195 18139
rect 10137 18099 10195 18105
rect 11974 18096 11980 18148
rect 12032 18136 12038 18148
rect 12636 18136 12664 18167
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18204 13231 18207
rect 13262 18204 13268 18216
rect 13219 18176 13268 18204
rect 13219 18173 13231 18176
rect 13173 18167 13231 18173
rect 13188 18136 13216 18167
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 14568 18176 14749 18204
rect 12032 18108 13216 18136
rect 12032 18096 12038 18108
rect 6362 18028 6368 18080
rect 6420 18068 6426 18080
rect 7009 18071 7067 18077
rect 7009 18068 7021 18071
rect 6420 18040 7021 18068
rect 6420 18028 6426 18040
rect 7009 18037 7021 18040
rect 7055 18037 7067 18071
rect 7009 18031 7067 18037
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 14568 18077 14596 18176
rect 14737 18173 14749 18176
rect 14783 18173 14795 18207
rect 14844 18204 14872 18244
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 16040 18244 18337 18272
rect 16040 18204 16068 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 14844 18176 16068 18204
rect 18049 18207 18107 18213
rect 14737 18167 14795 18173
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18782 18204 18788 18216
rect 18095 18176 18788 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18782 18164 18788 18176
rect 18840 18204 18846 18216
rect 19904 18204 19932 18303
rect 20990 18300 20996 18312
rect 21048 18340 21054 18352
rect 22020 18340 22048 18380
rect 23014 18368 23020 18420
rect 23072 18408 23078 18420
rect 29362 18408 29368 18420
rect 23072 18380 29368 18408
rect 23072 18368 23078 18380
rect 29362 18368 29368 18380
rect 29420 18368 29426 18420
rect 31386 18408 31392 18420
rect 29472 18380 31392 18408
rect 28077 18343 28135 18349
rect 28077 18340 28089 18343
rect 21048 18312 21128 18340
rect 22020 18312 28089 18340
rect 21048 18300 21054 18312
rect 21100 18281 21128 18312
rect 28077 18309 28089 18312
rect 28123 18340 28135 18343
rect 29472 18340 29500 18380
rect 31386 18368 31392 18380
rect 31444 18368 31450 18420
rect 32398 18368 32404 18420
rect 32456 18408 32462 18420
rect 32493 18411 32551 18417
rect 32493 18408 32505 18411
rect 32456 18380 32505 18408
rect 32456 18368 32462 18380
rect 32493 18377 32505 18380
rect 32539 18377 32551 18411
rect 33505 18411 33563 18417
rect 33505 18408 33517 18411
rect 32493 18371 32551 18377
rect 32876 18380 33517 18408
rect 28123 18312 29500 18340
rect 29549 18343 29607 18349
rect 28123 18309 28135 18312
rect 28077 18303 28135 18309
rect 29549 18309 29561 18343
rect 29595 18340 29607 18343
rect 32122 18340 32128 18352
rect 29595 18312 32128 18340
rect 29595 18309 29607 18312
rect 29549 18303 29607 18309
rect 32122 18300 32128 18312
rect 32180 18300 32186 18352
rect 32217 18343 32275 18349
rect 32217 18309 32229 18343
rect 32263 18340 32275 18343
rect 32876 18340 32904 18380
rect 33505 18377 33517 18380
rect 33551 18377 33563 18411
rect 33505 18371 33563 18377
rect 34974 18368 34980 18420
rect 35032 18408 35038 18420
rect 36541 18411 36599 18417
rect 36541 18408 36553 18411
rect 35032 18380 36553 18408
rect 35032 18368 35038 18380
rect 36541 18377 36553 18380
rect 36587 18408 36599 18411
rect 39006 18411 39064 18417
rect 36587 18380 37688 18408
rect 36587 18377 36599 18380
rect 36541 18371 36599 18377
rect 32263 18312 32904 18340
rect 32263 18309 32275 18312
rect 32217 18303 32275 18309
rect 32950 18300 32956 18352
rect 33008 18340 33014 18352
rect 33394 18343 33452 18349
rect 33008 18312 33053 18340
rect 33008 18300 33014 18312
rect 33394 18309 33406 18343
rect 33440 18340 33452 18343
rect 37274 18340 37280 18352
rect 33440 18312 36124 18340
rect 33440 18309 33452 18312
rect 33394 18303 33452 18309
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18241 21143 18275
rect 21358 18272 21364 18284
rect 21319 18244 21364 18272
rect 21085 18235 21143 18241
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 25222 18272 25228 18284
rect 25183 18244 25228 18272
rect 25222 18232 25228 18244
rect 25280 18232 25286 18284
rect 25498 18232 25504 18284
rect 25556 18272 25562 18284
rect 25685 18275 25743 18281
rect 25685 18272 25697 18275
rect 25556 18244 25697 18272
rect 25556 18232 25562 18244
rect 25685 18241 25697 18244
rect 25731 18241 25743 18275
rect 25685 18235 25743 18241
rect 28994 18232 29000 18284
rect 29052 18272 29058 18284
rect 29420 18275 29478 18281
rect 29420 18272 29432 18275
rect 29052 18244 29432 18272
rect 29052 18232 29058 18244
rect 29420 18241 29432 18244
rect 29466 18241 29478 18275
rect 29638 18272 29644 18284
rect 29599 18244 29644 18272
rect 29420 18235 29478 18241
rect 29638 18232 29644 18244
rect 29696 18232 29702 18284
rect 29733 18275 29791 18281
rect 29733 18241 29745 18275
rect 29779 18241 29791 18275
rect 32398 18272 32404 18284
rect 29733 18235 29791 18241
rect 32232 18244 32404 18272
rect 18840 18176 19932 18204
rect 25409 18207 25467 18213
rect 18840 18164 18846 18176
rect 25409 18173 25421 18207
rect 25455 18173 25467 18207
rect 25409 18167 25467 18173
rect 25777 18207 25835 18213
rect 25777 18173 25789 18207
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 16393 18139 16451 18145
rect 16393 18105 16405 18139
rect 16439 18136 16451 18139
rect 16482 18136 16488 18148
rect 16439 18108 16488 18136
rect 16439 18105 16451 18108
rect 16393 18099 16451 18105
rect 16482 18096 16488 18108
rect 16540 18096 16546 18148
rect 19702 18136 19708 18148
rect 19663 18108 19708 18136
rect 19702 18096 19708 18108
rect 19760 18096 19766 18148
rect 22741 18139 22799 18145
rect 22741 18105 22753 18139
rect 22787 18136 22799 18139
rect 23474 18136 23480 18148
rect 22787 18108 23480 18136
rect 22787 18105 22799 18108
rect 22741 18099 22799 18105
rect 23474 18096 23480 18108
rect 23532 18136 23538 18148
rect 23934 18136 23940 18148
rect 23532 18108 23940 18136
rect 23532 18096 23538 18108
rect 23934 18096 23940 18108
rect 23992 18096 23998 18148
rect 14553 18071 14611 18077
rect 14553 18068 14565 18071
rect 14424 18040 14565 18068
rect 14424 18028 14430 18040
rect 14553 18037 14565 18040
rect 14599 18037 14611 18071
rect 14553 18031 14611 18037
rect 22002 18028 22008 18080
rect 22060 18068 22066 18080
rect 23014 18068 23020 18080
rect 22060 18040 23020 18068
rect 22060 18028 22066 18040
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 25041 18071 25099 18077
rect 25041 18037 25053 18071
rect 25087 18068 25099 18071
rect 25222 18068 25228 18080
rect 25087 18040 25228 18068
rect 25087 18037 25099 18040
rect 25041 18031 25099 18037
rect 25222 18028 25228 18040
rect 25280 18028 25286 18080
rect 25424 18068 25452 18167
rect 25792 18136 25820 18167
rect 25958 18164 25964 18216
rect 26016 18204 26022 18216
rect 29748 18204 29776 18235
rect 26016 18176 29776 18204
rect 31021 18207 31079 18213
rect 26016 18164 26022 18176
rect 31021 18173 31033 18207
rect 31067 18173 31079 18207
rect 31202 18204 31208 18216
rect 31115 18176 31208 18204
rect 31021 18167 31079 18173
rect 26602 18136 26608 18148
rect 25792 18108 26608 18136
rect 26602 18096 26608 18108
rect 26660 18096 26666 18148
rect 26697 18139 26755 18145
rect 26697 18105 26709 18139
rect 26743 18136 26755 18139
rect 26789 18139 26847 18145
rect 26789 18136 26801 18139
rect 26743 18108 26801 18136
rect 26743 18105 26755 18108
rect 26697 18099 26755 18105
rect 26789 18105 26801 18108
rect 26835 18136 26847 18139
rect 26970 18136 26976 18148
rect 26835 18108 26976 18136
rect 26835 18105 26847 18108
rect 26789 18099 26847 18105
rect 26970 18096 26976 18108
rect 27028 18096 27034 18148
rect 28258 18096 28264 18148
rect 28316 18136 28322 18148
rect 28902 18136 28908 18148
rect 28316 18108 28908 18136
rect 28316 18096 28322 18108
rect 28902 18096 28908 18108
rect 28960 18096 28966 18148
rect 28994 18096 29000 18148
rect 29052 18136 29058 18148
rect 29273 18139 29331 18145
rect 29273 18136 29285 18139
rect 29052 18108 29285 18136
rect 29052 18096 29058 18108
rect 29273 18105 29285 18108
rect 29319 18105 29331 18139
rect 29273 18099 29331 18105
rect 27430 18068 27436 18080
rect 25424 18040 27436 18068
rect 27430 18028 27436 18040
rect 27488 18028 27494 18080
rect 28810 18028 28816 18080
rect 28868 18068 28874 18080
rect 31036 18068 31064 18167
rect 31202 18164 31208 18176
rect 31260 18204 31266 18216
rect 31260 18176 31708 18204
rect 31260 18164 31266 18176
rect 28868 18040 31064 18068
rect 31680 18068 31708 18176
rect 31754 18164 31760 18216
rect 31812 18204 31818 18216
rect 31941 18207 31999 18213
rect 31812 18176 31857 18204
rect 31812 18164 31818 18176
rect 31941 18173 31953 18207
rect 31987 18204 31999 18207
rect 32232 18204 32260 18244
rect 32398 18232 32404 18244
rect 32456 18232 32462 18284
rect 33594 18272 33600 18284
rect 33555 18244 33600 18272
rect 33594 18232 33600 18244
rect 33652 18232 33658 18284
rect 33689 18275 33747 18281
rect 33689 18241 33701 18275
rect 33735 18241 33747 18275
rect 33689 18235 33747 18241
rect 31987 18176 32260 18204
rect 31987 18173 31999 18176
rect 31941 18167 31999 18173
rect 32306 18164 32312 18216
rect 32364 18204 32370 18216
rect 33704 18204 33732 18235
rect 34974 18204 34980 18216
rect 32364 18176 33732 18204
rect 34935 18176 34980 18204
rect 32364 18164 32370 18176
rect 34974 18164 34980 18176
rect 35032 18164 35038 18216
rect 35158 18204 35164 18216
rect 35119 18176 35164 18204
rect 35158 18164 35164 18176
rect 35216 18164 35222 18216
rect 35618 18204 35624 18216
rect 35579 18176 35624 18204
rect 35618 18164 35624 18176
rect 35676 18164 35682 18216
rect 35710 18164 35716 18216
rect 35768 18204 35774 18216
rect 36096 18204 36124 18312
rect 36648 18312 37280 18340
rect 36648 18204 36676 18312
rect 37274 18300 37280 18312
rect 37332 18300 37338 18352
rect 37660 18272 37688 18380
rect 39006 18377 39018 18411
rect 39052 18408 39064 18411
rect 39666 18408 39672 18420
rect 39052 18380 39672 18408
rect 39052 18377 39064 18380
rect 39006 18371 39064 18377
rect 39666 18368 39672 18380
rect 39724 18368 39730 18420
rect 39758 18368 39764 18420
rect 39816 18408 39822 18420
rect 39816 18380 39861 18408
rect 39816 18368 39822 18380
rect 39942 18368 39948 18420
rect 40000 18408 40006 18420
rect 41598 18408 41604 18420
rect 40000 18380 41604 18408
rect 40000 18368 40006 18380
rect 41598 18368 41604 18380
rect 41656 18368 41662 18420
rect 44158 18411 44216 18417
rect 44158 18377 44170 18411
rect 44204 18408 44216 18411
rect 45002 18408 45008 18420
rect 44204 18380 45008 18408
rect 44204 18377 44216 18380
rect 44158 18371 44216 18377
rect 45002 18368 45008 18380
rect 45060 18368 45066 18420
rect 47946 18368 47952 18420
rect 48004 18408 48010 18420
rect 48133 18411 48191 18417
rect 48133 18408 48145 18411
rect 48004 18380 48145 18408
rect 48004 18368 48010 18380
rect 48133 18377 48145 18380
rect 48179 18377 48191 18411
rect 48133 18371 48191 18377
rect 39114 18340 39120 18352
rect 39075 18312 39120 18340
rect 39114 18300 39120 18312
rect 39172 18300 39178 18352
rect 39298 18300 39304 18352
rect 39356 18340 39362 18352
rect 43349 18343 43407 18349
rect 43349 18340 43361 18343
rect 39356 18312 42012 18340
rect 39356 18300 39362 18312
rect 39022 18272 39028 18284
rect 37660 18244 39028 18272
rect 39022 18232 39028 18244
rect 39080 18232 39086 18284
rect 39209 18275 39267 18281
rect 39209 18241 39221 18275
rect 39255 18272 39267 18275
rect 40126 18272 40132 18284
rect 39255 18244 40132 18272
rect 39255 18241 39267 18244
rect 39209 18235 39267 18241
rect 40126 18232 40132 18244
rect 40184 18232 40190 18284
rect 41785 18275 41843 18281
rect 41785 18272 41797 18275
rect 40236 18244 41797 18272
rect 35768 18176 35813 18204
rect 36096 18176 36676 18204
rect 36725 18207 36783 18213
rect 35768 18164 35774 18176
rect 36725 18173 36737 18207
rect 36771 18204 36783 18207
rect 38930 18204 38936 18216
rect 36771 18176 38936 18204
rect 36771 18173 36783 18176
rect 36725 18167 36783 18173
rect 33229 18139 33287 18145
rect 33229 18105 33241 18139
rect 33275 18136 33287 18139
rect 36265 18139 36323 18145
rect 36265 18136 36277 18139
rect 33275 18108 36277 18136
rect 33275 18105 33287 18108
rect 33229 18099 33287 18105
rect 36265 18105 36277 18108
rect 36311 18105 36323 18139
rect 36740 18136 36768 18167
rect 38930 18164 38936 18176
rect 38988 18164 38994 18216
rect 39942 18164 39948 18216
rect 40000 18204 40006 18216
rect 40236 18204 40264 18244
rect 41785 18241 41797 18244
rect 41831 18241 41843 18275
rect 41785 18235 41843 18241
rect 40770 18204 40776 18216
rect 40000 18176 40264 18204
rect 40731 18176 40776 18204
rect 40000 18164 40006 18176
rect 40770 18164 40776 18176
rect 40828 18164 40834 18216
rect 41984 18213 42012 18312
rect 42996 18312 43361 18340
rect 41969 18207 42027 18213
rect 41969 18173 41981 18207
rect 42015 18173 42027 18207
rect 42518 18204 42524 18216
rect 42479 18176 42524 18204
rect 41969 18167 42027 18173
rect 38838 18136 38844 18148
rect 36265 18099 36323 18105
rect 36372 18108 36768 18136
rect 38799 18108 38844 18136
rect 32769 18071 32827 18077
rect 32769 18068 32781 18071
rect 31680 18040 32781 18068
rect 28868 18028 28874 18040
rect 32769 18037 32781 18040
rect 32815 18068 32827 18071
rect 33042 18068 33048 18080
rect 32815 18040 33048 18068
rect 32815 18037 32827 18040
rect 32769 18031 32827 18037
rect 33042 18028 33048 18040
rect 33100 18028 33106 18080
rect 35158 18028 35164 18080
rect 35216 18068 35222 18080
rect 36372 18068 36400 18108
rect 38838 18096 38844 18108
rect 38896 18096 38902 18148
rect 41984 18136 42012 18167
rect 42518 18164 42524 18176
rect 42576 18164 42582 18216
rect 42610 18164 42616 18216
rect 42668 18204 42674 18216
rect 42705 18207 42763 18213
rect 42705 18204 42717 18207
rect 42668 18176 42717 18204
rect 42668 18164 42674 18176
rect 42705 18173 42717 18176
rect 42751 18204 42763 18207
rect 42996 18204 43024 18312
rect 43349 18309 43361 18312
rect 43395 18340 43407 18343
rect 48148 18340 48176 18371
rect 52730 18368 52736 18420
rect 52788 18408 52794 18420
rect 52825 18411 52883 18417
rect 52825 18408 52837 18411
rect 52788 18380 52837 18408
rect 52788 18368 52794 18380
rect 52825 18377 52837 18380
rect 52871 18377 52883 18411
rect 52825 18371 52883 18377
rect 48409 18343 48467 18349
rect 48409 18340 48421 18343
rect 43395 18312 47256 18340
rect 48148 18312 48421 18340
rect 43395 18309 43407 18312
rect 43349 18303 43407 18309
rect 43073 18275 43131 18281
rect 43073 18241 43085 18275
rect 43119 18272 43131 18275
rect 44361 18275 44419 18281
rect 44361 18272 44373 18275
rect 43119 18244 44373 18272
rect 43119 18241 43131 18244
rect 43073 18235 43131 18241
rect 44361 18241 44373 18244
rect 44407 18241 44419 18275
rect 44361 18235 44419 18241
rect 44450 18232 44456 18284
rect 44508 18272 44514 18284
rect 46106 18272 46112 18284
rect 44508 18244 44553 18272
rect 46067 18244 46112 18272
rect 44508 18232 44514 18244
rect 46106 18232 46112 18244
rect 46164 18232 46170 18284
rect 47228 18272 47256 18312
rect 48409 18309 48421 18312
rect 48455 18340 48467 18343
rect 49697 18343 49755 18349
rect 49697 18340 49709 18343
rect 48455 18312 49709 18340
rect 48455 18309 48467 18312
rect 48409 18303 48467 18309
rect 49697 18309 49709 18312
rect 49743 18309 49755 18343
rect 49697 18303 49755 18309
rect 49050 18272 49056 18284
rect 47228 18244 48728 18272
rect 49011 18244 49056 18272
rect 44266 18213 44272 18216
rect 42751 18176 43024 18204
rect 44223 18207 44272 18213
rect 42751 18173 42763 18176
rect 42705 18167 42763 18173
rect 44223 18173 44235 18207
rect 44269 18173 44272 18207
rect 44223 18167 44272 18173
rect 44266 18164 44272 18167
rect 44324 18164 44330 18216
rect 44726 18164 44732 18216
rect 44784 18204 44790 18216
rect 46290 18204 46296 18216
rect 44784 18176 45968 18204
rect 46251 18176 46296 18204
rect 44784 18164 44790 18176
rect 42978 18136 42984 18148
rect 41984 18108 42984 18136
rect 42978 18096 42984 18108
rect 43036 18096 43042 18148
rect 43993 18139 44051 18145
rect 43993 18105 44005 18139
rect 44039 18136 44051 18139
rect 45646 18136 45652 18148
rect 44039 18108 45652 18136
rect 44039 18105 44051 18108
rect 43993 18099 44051 18105
rect 45646 18096 45652 18108
rect 45704 18096 45710 18148
rect 45940 18145 45968 18176
rect 46290 18164 46296 18176
rect 46348 18164 46354 18216
rect 46753 18207 46811 18213
rect 46753 18173 46765 18207
rect 46799 18173 46811 18207
rect 46753 18167 46811 18173
rect 46845 18207 46903 18213
rect 46845 18173 46857 18207
rect 46891 18173 46903 18207
rect 48314 18204 48320 18216
rect 48275 18176 48320 18204
rect 46845 18167 46903 18173
rect 45925 18139 45983 18145
rect 45925 18105 45937 18139
rect 45971 18136 45983 18139
rect 46768 18136 46796 18167
rect 45971 18108 46796 18136
rect 46860 18136 46888 18167
rect 48314 18164 48320 18176
rect 48372 18164 48378 18216
rect 48590 18204 48596 18216
rect 48551 18176 48596 18204
rect 48590 18164 48596 18176
rect 48648 18164 48654 18216
rect 48700 18204 48728 18244
rect 49050 18232 49056 18244
rect 49108 18232 49114 18284
rect 49712 18204 49740 18303
rect 50065 18207 50123 18213
rect 50065 18204 50077 18207
rect 48700 18176 49188 18204
rect 49712 18176 50077 18204
rect 49050 18136 49056 18148
rect 46860 18108 49056 18136
rect 45971 18105 45983 18108
rect 45925 18099 45983 18105
rect 49050 18096 49056 18108
rect 49108 18096 49114 18148
rect 35216 18040 36400 18068
rect 35216 18028 35222 18040
rect 36446 18028 36452 18080
rect 36504 18068 36510 18080
rect 39485 18071 39543 18077
rect 39485 18068 39497 18071
rect 36504 18040 39497 18068
rect 36504 18028 36510 18040
rect 39485 18037 39497 18040
rect 39531 18037 39543 18071
rect 39485 18031 39543 18037
rect 40034 18028 40040 18080
rect 40092 18068 40098 18080
rect 40865 18071 40923 18077
rect 40865 18068 40877 18071
rect 40092 18040 40877 18068
rect 40092 18028 40098 18040
rect 40865 18037 40877 18040
rect 40911 18068 40923 18071
rect 41966 18068 41972 18080
rect 40911 18040 41972 18068
rect 40911 18037 40923 18040
rect 40865 18031 40923 18037
rect 41966 18028 41972 18040
rect 42024 18028 42030 18080
rect 47302 18068 47308 18080
rect 47263 18040 47308 18068
rect 47302 18028 47308 18040
rect 47360 18028 47366 18080
rect 49160 18068 49188 18176
rect 50065 18173 50077 18176
rect 50111 18173 50123 18207
rect 50065 18167 50123 18173
rect 51350 18164 51356 18216
rect 51408 18204 51414 18216
rect 52365 18207 52423 18213
rect 52365 18204 52377 18207
rect 51408 18176 52377 18204
rect 51408 18164 51414 18176
rect 52365 18173 52377 18176
rect 52411 18173 52423 18207
rect 52638 18204 52644 18216
rect 52599 18176 52644 18204
rect 52365 18167 52423 18173
rect 52638 18164 52644 18176
rect 52696 18164 52702 18216
rect 49878 18136 49884 18148
rect 49839 18108 49884 18136
rect 49878 18096 49884 18108
rect 49936 18096 49942 18148
rect 50433 18139 50491 18145
rect 50433 18105 50445 18139
rect 50479 18136 50491 18139
rect 51626 18136 51632 18148
rect 50479 18108 51632 18136
rect 50479 18105 50491 18108
rect 50433 18099 50491 18105
rect 51626 18096 51632 18108
rect 51684 18096 51690 18148
rect 52546 18136 52552 18148
rect 52507 18108 52552 18136
rect 52546 18096 52552 18108
rect 52604 18096 52610 18148
rect 49970 18068 49976 18080
rect 49160 18040 49976 18068
rect 49970 18028 49976 18040
rect 50028 18028 50034 18080
rect 1104 17978 54832 18000
rect 1104 17926 18912 17978
rect 18964 17926 18976 17978
rect 19028 17926 19040 17978
rect 19092 17926 19104 17978
rect 19156 17926 36843 17978
rect 36895 17926 36907 17978
rect 36959 17926 36971 17978
rect 37023 17926 37035 17978
rect 37087 17926 54832 17978
rect 1104 17904 54832 17926
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17833 3019 17867
rect 2961 17827 3019 17833
rect 2976 17796 3004 17827
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4801 17867 4859 17873
rect 4801 17864 4813 17867
rect 4396 17836 4813 17864
rect 4396 17824 4402 17836
rect 4801 17833 4813 17836
rect 4847 17833 4859 17867
rect 4801 17827 4859 17833
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 11609 17867 11667 17873
rect 11609 17864 11621 17867
rect 11296 17836 11621 17864
rect 11296 17824 11302 17836
rect 11609 17833 11621 17836
rect 11655 17864 11667 17867
rect 11790 17864 11796 17876
rect 11655 17836 11796 17864
rect 11655 17833 11667 17836
rect 11609 17827 11667 17833
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 12618 17864 12624 17876
rect 12544 17836 12624 17864
rect 2976 17768 6040 17796
rect 2130 17688 2136 17740
rect 2188 17728 2194 17740
rect 6012 17737 6040 17768
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 12342 17796 12348 17808
rect 8352 17768 12348 17796
rect 8352 17756 8358 17768
rect 12342 17756 12348 17768
rect 12400 17796 12406 17808
rect 12400 17768 12480 17796
rect 12400 17756 12406 17768
rect 3145 17731 3203 17737
rect 3145 17728 3157 17731
rect 2188 17700 3157 17728
rect 2188 17688 2194 17700
rect 3145 17697 3157 17700
rect 3191 17697 3203 17731
rect 3145 17691 3203 17697
rect 4985 17731 5043 17737
rect 4985 17697 4997 17731
rect 5031 17728 5043 17731
rect 5997 17731 6055 17737
rect 5031 17700 5856 17728
rect 5031 17697 5043 17700
rect 4985 17691 5043 17697
rect 5828 17601 5856 17700
rect 5997 17697 6009 17731
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17728 6699 17731
rect 6822 17728 6828 17740
rect 6687 17700 6828 17728
rect 6687 17697 6699 17700
rect 6641 17691 6699 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 7837 17731 7895 17737
rect 7837 17697 7849 17731
rect 7883 17728 7895 17731
rect 8570 17728 8576 17740
rect 7883 17700 8576 17728
rect 7883 17697 7895 17700
rect 7837 17691 7895 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 10962 17728 10968 17740
rect 10551 17700 10968 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11790 17728 11796 17740
rect 11751 17700 11796 17728
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 11974 17728 11980 17740
rect 11935 17700 11980 17728
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12452 17737 12480 17768
rect 12544 17737 12572 17836
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 15930 17864 15936 17876
rect 14231 17836 15936 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 19242 17864 19248 17876
rect 18104 17836 19248 17864
rect 18104 17824 18110 17836
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 21177 17867 21235 17873
rect 21177 17864 21189 17867
rect 19392 17836 21189 17864
rect 19392 17824 19398 17836
rect 21177 17833 21189 17836
rect 21223 17864 21235 17867
rect 23661 17867 23719 17873
rect 21223 17836 22508 17864
rect 21223 17833 21235 17836
rect 21177 17827 21235 17833
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 16117 17799 16175 17805
rect 16117 17796 16129 17799
rect 13872 17768 16129 17796
rect 13872 17756 13878 17768
rect 16117 17765 16129 17768
rect 16163 17796 16175 17799
rect 16163 17768 22140 17796
rect 16163 17765 16175 17768
rect 16117 17759 16175 17765
rect 12437 17731 12495 17737
rect 12437 17697 12449 17731
rect 12483 17697 12495 17731
rect 12437 17691 12495 17697
rect 12529 17731 12587 17737
rect 12529 17697 12541 17731
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 14369 17731 14427 17737
rect 14369 17697 14381 17731
rect 14415 17728 14427 17731
rect 16025 17731 16083 17737
rect 14415 17700 14596 17728
rect 14415 17697 14427 17700
rect 14369 17691 14427 17697
rect 5813 17595 5871 17601
rect 5813 17561 5825 17595
rect 5859 17561 5871 17595
rect 5813 17555 5871 17561
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 6825 17527 6883 17533
rect 6825 17524 6837 17527
rect 6788 17496 6837 17524
rect 6788 17484 6794 17496
rect 6825 17493 6837 17496
rect 6871 17493 6883 17527
rect 8018 17524 8024 17536
rect 7979 17496 8024 17524
rect 6825 17487 6883 17493
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 10686 17524 10692 17536
rect 10647 17496 10692 17524
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 12986 17524 12992 17536
rect 12947 17496 12992 17524
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 14568 17533 14596 17700
rect 16025 17697 16037 17731
rect 16071 17728 16083 17731
rect 16482 17728 16488 17740
rect 16071 17700 16488 17728
rect 16071 17697 16083 17700
rect 16025 17691 16083 17697
rect 16482 17688 16488 17700
rect 16540 17688 16546 17740
rect 17037 17731 17095 17737
rect 17037 17697 17049 17731
rect 17083 17728 17095 17731
rect 17218 17728 17224 17740
rect 17083 17700 17224 17728
rect 17083 17697 17095 17700
rect 17037 17691 17095 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 18230 17728 18236 17740
rect 18191 17700 18236 17728
rect 18230 17688 18236 17700
rect 18288 17688 18294 17740
rect 19153 17731 19211 17737
rect 19153 17697 19165 17731
rect 19199 17728 19211 17731
rect 19702 17728 19708 17740
rect 19199 17700 19708 17728
rect 19199 17697 19211 17700
rect 19153 17691 19211 17697
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 21082 17728 21088 17740
rect 21043 17700 21088 17728
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 22002 17728 22008 17740
rect 21963 17700 22008 17728
rect 22002 17688 22008 17700
rect 22060 17688 22066 17740
rect 22112 17737 22140 17768
rect 22097 17731 22155 17737
rect 22097 17697 22109 17731
rect 22143 17697 22155 17731
rect 22097 17691 22155 17697
rect 22281 17731 22339 17737
rect 22281 17697 22293 17731
rect 22327 17728 22339 17731
rect 22370 17728 22376 17740
rect 22327 17700 22376 17728
rect 22327 17697 22339 17700
rect 22281 17691 22339 17697
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 22480 17592 22508 17836
rect 23661 17833 23673 17867
rect 23707 17864 23719 17867
rect 29270 17864 29276 17876
rect 23707 17836 29276 17864
rect 23707 17833 23719 17836
rect 23661 17827 23719 17833
rect 23676 17796 23704 17827
rect 29270 17824 29276 17836
rect 29328 17824 29334 17876
rect 30006 17824 30012 17876
rect 30064 17864 30070 17876
rect 30064 17836 37872 17864
rect 30064 17824 30070 17836
rect 22848 17768 23704 17796
rect 24857 17799 24915 17805
rect 22848 17737 22876 17768
rect 24857 17765 24869 17799
rect 24903 17796 24915 17799
rect 25774 17796 25780 17808
rect 24903 17768 25780 17796
rect 24903 17765 24915 17768
rect 24857 17759 24915 17765
rect 25774 17756 25780 17768
rect 25832 17756 25838 17808
rect 29638 17756 29644 17808
rect 29696 17796 29702 17808
rect 29733 17799 29791 17805
rect 29733 17796 29745 17799
rect 29696 17768 29745 17796
rect 29696 17756 29702 17768
rect 29733 17765 29745 17768
rect 29779 17765 29791 17799
rect 29733 17759 29791 17765
rect 29917 17799 29975 17805
rect 29917 17765 29929 17799
rect 29963 17796 29975 17799
rect 31202 17796 31208 17808
rect 29963 17768 31208 17796
rect 29963 17765 29975 17768
rect 29917 17759 29975 17765
rect 22833 17731 22891 17737
rect 22833 17697 22845 17731
rect 22879 17697 22891 17731
rect 23014 17728 23020 17740
rect 22975 17700 23020 17728
rect 22833 17691 22891 17697
rect 23014 17688 23020 17700
rect 23072 17688 23078 17740
rect 28718 17728 28724 17740
rect 28679 17700 28724 17728
rect 28718 17688 28724 17700
rect 28776 17688 28782 17740
rect 29089 17731 29147 17737
rect 29089 17697 29101 17731
rect 29135 17697 29147 17731
rect 29454 17728 29460 17740
rect 29415 17700 29460 17728
rect 29089 17691 29147 17697
rect 24946 17620 24952 17672
rect 25004 17669 25010 17672
rect 25004 17663 25062 17669
rect 25004 17629 25016 17663
rect 25050 17629 25062 17663
rect 25222 17660 25228 17672
rect 25183 17632 25228 17660
rect 25004 17623 25062 17629
rect 25004 17620 25010 17623
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 29104 17660 29132 17691
rect 29454 17688 29460 17700
rect 29512 17688 29518 17740
rect 29932 17660 29960 17759
rect 31202 17756 31208 17768
rect 31260 17756 31266 17808
rect 36265 17799 36323 17805
rect 32876 17768 36216 17796
rect 32306 17688 32312 17740
rect 32364 17728 32370 17740
rect 32766 17728 32772 17740
rect 32364 17700 32409 17728
rect 32727 17700 32772 17728
rect 32364 17688 32370 17700
rect 32766 17688 32772 17700
rect 32824 17688 32830 17740
rect 32876 17737 32904 17768
rect 32861 17731 32919 17737
rect 32861 17697 32873 17731
rect 32907 17697 32919 17731
rect 32861 17691 32919 17697
rect 34333 17731 34391 17737
rect 34333 17697 34345 17731
rect 34379 17728 34391 17731
rect 34606 17728 34612 17740
rect 34379 17700 34612 17728
rect 34379 17697 34391 17700
rect 34333 17691 34391 17697
rect 34606 17688 34612 17700
rect 34664 17728 34670 17740
rect 35710 17728 35716 17740
rect 34664 17700 35716 17728
rect 34664 17688 34670 17700
rect 35710 17688 35716 17700
rect 35768 17688 35774 17740
rect 36188 17737 36216 17768
rect 36265 17765 36277 17799
rect 36311 17796 36323 17799
rect 36630 17796 36636 17808
rect 36311 17768 36636 17796
rect 36311 17765 36323 17768
rect 36265 17759 36323 17765
rect 36630 17756 36636 17768
rect 36688 17756 36694 17808
rect 37182 17756 37188 17808
rect 37240 17796 37246 17808
rect 37240 17768 37780 17796
rect 37240 17756 37246 17768
rect 36081 17731 36139 17737
rect 36081 17697 36093 17731
rect 36127 17697 36139 17731
rect 36081 17691 36139 17697
rect 36173 17731 36231 17737
rect 36173 17697 36185 17731
rect 36219 17728 36231 17731
rect 36354 17728 36360 17740
rect 36219 17700 36360 17728
rect 36219 17697 36231 17700
rect 36173 17691 36231 17697
rect 29104 17632 29960 17660
rect 30374 17620 30380 17672
rect 30432 17660 30438 17672
rect 31941 17663 31999 17669
rect 31941 17660 31953 17663
rect 30432 17632 31953 17660
rect 30432 17620 30438 17632
rect 31941 17629 31953 17632
rect 31987 17660 31999 17663
rect 32125 17663 32183 17669
rect 32125 17660 32137 17663
rect 31987 17632 32137 17660
rect 31987 17629 31999 17632
rect 31941 17623 31999 17629
rect 32125 17629 32137 17632
rect 32171 17629 32183 17663
rect 32125 17623 32183 17629
rect 33502 17620 33508 17672
rect 33560 17660 33566 17672
rect 34425 17663 34483 17669
rect 34425 17660 34437 17663
rect 33560 17632 34437 17660
rect 33560 17620 33566 17632
rect 34425 17629 34437 17632
rect 34471 17629 34483 17663
rect 36096 17660 36124 17691
rect 36354 17688 36360 17700
rect 36412 17688 36418 17740
rect 37366 17688 37372 17740
rect 37424 17728 37430 17740
rect 37752 17737 37780 17768
rect 37553 17731 37611 17737
rect 37553 17728 37565 17731
rect 37424 17700 37565 17728
rect 37424 17688 37430 17700
rect 37553 17697 37565 17700
rect 37599 17697 37611 17731
rect 37553 17691 37611 17697
rect 37737 17731 37795 17737
rect 37737 17697 37749 17731
rect 37783 17697 37795 17731
rect 37737 17691 37795 17697
rect 36096 17632 37780 17660
rect 34425 17623 34483 17629
rect 25133 17595 25191 17601
rect 22480 17564 24624 17592
rect 14553 17527 14611 17533
rect 14553 17493 14565 17527
rect 14599 17524 14611 17527
rect 14734 17524 14740 17536
rect 14599 17496 14740 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 17126 17524 17132 17536
rect 17087 17496 17132 17524
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 18046 17524 18052 17536
rect 18007 17496 18052 17524
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 23290 17524 23296 17536
rect 23251 17496 23296 17524
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 24596 17524 24624 17564
rect 25133 17561 25145 17595
rect 25179 17592 25191 17595
rect 25406 17592 25412 17604
rect 25179 17564 25412 17592
rect 25179 17561 25191 17564
rect 25133 17555 25191 17561
rect 25406 17552 25412 17564
rect 25464 17552 25470 17604
rect 25501 17595 25559 17601
rect 25501 17561 25513 17595
rect 25547 17592 25559 17595
rect 28994 17592 29000 17604
rect 25547 17564 29000 17592
rect 25547 17561 25559 17564
rect 25501 17555 25559 17561
rect 28994 17552 29000 17564
rect 29052 17552 29058 17604
rect 35894 17592 35900 17604
rect 35855 17564 35900 17592
rect 35894 17552 35900 17564
rect 35952 17552 35958 17604
rect 37384 17601 37412 17632
rect 37369 17595 37427 17601
rect 37369 17561 37381 17595
rect 37415 17561 37427 17595
rect 37369 17555 37427 17561
rect 28626 17524 28632 17536
rect 24596 17496 28632 17524
rect 28626 17484 28632 17496
rect 28684 17484 28690 17536
rect 28902 17484 28908 17536
rect 28960 17524 28966 17536
rect 29730 17524 29736 17536
rect 28960 17496 29736 17524
rect 28960 17484 28966 17496
rect 29730 17484 29736 17496
rect 29788 17484 29794 17536
rect 33318 17524 33324 17536
rect 33279 17496 33324 17524
rect 33318 17484 33324 17496
rect 33376 17484 33382 17536
rect 37752 17524 37780 17632
rect 37844 17592 37872 17836
rect 37918 17824 37924 17876
rect 37976 17864 37982 17876
rect 37976 17836 38792 17864
rect 37976 17824 37982 17836
rect 38654 17796 38660 17808
rect 38488 17768 38660 17796
rect 37921 17731 37979 17737
rect 37921 17697 37933 17731
rect 37967 17728 37979 17731
rect 38102 17728 38108 17740
rect 37967 17700 38108 17728
rect 37967 17697 37979 17700
rect 37921 17691 37979 17697
rect 38102 17688 38108 17700
rect 38160 17688 38166 17740
rect 38378 17728 38384 17740
rect 38339 17700 38384 17728
rect 38378 17688 38384 17700
rect 38436 17688 38442 17740
rect 38488 17737 38516 17768
rect 38654 17756 38660 17768
rect 38712 17756 38718 17808
rect 38764 17796 38792 17836
rect 38838 17824 38844 17876
rect 38896 17864 38902 17876
rect 38933 17867 38991 17873
rect 38933 17864 38945 17867
rect 38896 17836 38945 17864
rect 38896 17824 38902 17836
rect 38933 17833 38945 17836
rect 38979 17833 38991 17867
rect 38933 17827 38991 17833
rect 39022 17824 39028 17876
rect 39080 17864 39086 17876
rect 44174 17864 44180 17876
rect 39080 17836 44180 17864
rect 39080 17824 39086 17836
rect 44174 17824 44180 17836
rect 44232 17824 44238 17876
rect 44542 17824 44548 17876
rect 44600 17864 44606 17876
rect 48590 17864 48596 17876
rect 44600 17836 48596 17864
rect 44600 17824 44606 17836
rect 40037 17799 40095 17805
rect 40037 17796 40049 17799
rect 38764 17768 40049 17796
rect 40037 17765 40049 17768
rect 40083 17765 40095 17799
rect 45465 17799 45523 17805
rect 40037 17759 40095 17765
rect 40328 17768 43944 17796
rect 38473 17731 38531 17737
rect 38473 17697 38485 17731
rect 38519 17697 38531 17731
rect 38473 17691 38531 17697
rect 38562 17688 38568 17740
rect 38620 17728 38626 17740
rect 39209 17731 39267 17737
rect 39209 17728 39221 17731
rect 38620 17700 39221 17728
rect 38620 17688 38626 17700
rect 39209 17697 39221 17700
rect 39255 17697 39267 17731
rect 39209 17691 39267 17697
rect 39942 17592 39948 17604
rect 37844 17564 39948 17592
rect 39942 17552 39948 17564
rect 40000 17552 40006 17604
rect 39298 17524 39304 17536
rect 37752 17496 39304 17524
rect 39298 17484 39304 17496
rect 39356 17484 39362 17536
rect 40052 17524 40080 17759
rect 40328 17737 40356 17768
rect 40313 17731 40371 17737
rect 40313 17697 40325 17731
rect 40359 17697 40371 17731
rect 40313 17691 40371 17697
rect 40405 17731 40463 17737
rect 40405 17697 40417 17731
rect 40451 17728 40463 17731
rect 40770 17728 40776 17740
rect 40451 17700 40776 17728
rect 40451 17697 40463 17700
rect 40405 17691 40463 17697
rect 40770 17688 40776 17700
rect 40828 17688 40834 17740
rect 40862 17688 40868 17740
rect 40920 17728 40926 17740
rect 41049 17731 41107 17737
rect 40920 17700 40965 17728
rect 40920 17688 40926 17700
rect 41049 17697 41061 17731
rect 41095 17728 41107 17731
rect 41095 17700 41276 17728
rect 41095 17697 41107 17700
rect 41049 17691 41107 17697
rect 41248 17660 41276 17700
rect 41322 17688 41328 17740
rect 41380 17728 41386 17740
rect 41601 17731 41659 17737
rect 41601 17728 41613 17731
rect 41380 17700 41613 17728
rect 41380 17688 41386 17700
rect 41601 17697 41613 17700
rect 41647 17697 41659 17731
rect 43916 17728 43944 17768
rect 45465 17765 45477 17799
rect 45511 17796 45523 17799
rect 45554 17796 45560 17808
rect 45511 17768 45560 17796
rect 45511 17765 45523 17768
rect 45465 17759 45523 17765
rect 45554 17756 45560 17768
rect 45612 17796 45618 17808
rect 46290 17796 46296 17808
rect 45612 17768 46296 17796
rect 45612 17756 45618 17768
rect 46290 17756 46296 17768
rect 46348 17756 46354 17808
rect 45646 17728 45652 17740
rect 43916 17700 45652 17728
rect 41601 17691 41659 17697
rect 45646 17688 45652 17700
rect 45704 17688 45710 17740
rect 47412 17737 47440 17836
rect 48590 17824 48596 17836
rect 48648 17824 48654 17876
rect 52454 17824 52460 17876
rect 52512 17864 52518 17876
rect 53009 17867 53067 17873
rect 53009 17864 53021 17867
rect 52512 17836 53021 17864
rect 52512 17824 52518 17836
rect 53009 17833 53021 17836
rect 53055 17833 53067 17867
rect 53009 17827 53067 17833
rect 48608 17796 48636 17824
rect 49513 17799 49571 17805
rect 48608 17768 49188 17796
rect 47029 17731 47087 17737
rect 47029 17697 47041 17731
rect 47075 17697 47087 17731
rect 47029 17691 47087 17697
rect 47397 17731 47455 17737
rect 47397 17697 47409 17731
rect 47443 17697 47455 17731
rect 47397 17691 47455 17697
rect 47581 17731 47639 17737
rect 47581 17697 47593 17731
rect 47627 17728 47639 17731
rect 48314 17728 48320 17740
rect 47627 17700 48320 17728
rect 47627 17697 47639 17700
rect 47581 17691 47639 17697
rect 43809 17663 43867 17669
rect 41248 17632 41368 17660
rect 40770 17552 40776 17604
rect 40828 17592 40834 17604
rect 41233 17595 41291 17601
rect 41233 17592 41245 17595
rect 40828 17564 41245 17592
rect 40828 17552 40834 17564
rect 41233 17561 41245 17564
rect 41279 17561 41291 17595
rect 41233 17555 41291 17561
rect 41340 17524 41368 17632
rect 43809 17629 43821 17663
rect 43855 17629 43867 17663
rect 44082 17660 44088 17672
rect 44043 17632 44088 17660
rect 43809 17623 43867 17629
rect 40052 17496 41368 17524
rect 43717 17527 43775 17533
rect 43717 17493 43729 17527
rect 43763 17524 43775 17527
rect 43824 17524 43852 17623
rect 44082 17620 44088 17632
rect 44140 17620 44146 17672
rect 47044 17592 47072 17691
rect 48314 17688 48320 17700
rect 48372 17728 48378 17740
rect 49160 17737 49188 17768
rect 49513 17765 49525 17799
rect 49559 17796 49571 17799
rect 49878 17796 49884 17808
rect 49559 17768 49884 17796
rect 49559 17765 49571 17768
rect 49513 17759 49571 17765
rect 49878 17756 49884 17768
rect 49936 17756 49942 17808
rect 48961 17731 49019 17737
rect 48961 17728 48973 17731
rect 48372 17700 48973 17728
rect 48372 17688 48378 17700
rect 48961 17697 48973 17700
rect 49007 17697 49019 17731
rect 48961 17691 49019 17697
rect 49145 17731 49203 17737
rect 49145 17697 49157 17731
rect 49191 17697 49203 17731
rect 49896 17728 49924 17756
rect 50341 17731 50399 17737
rect 50341 17728 50353 17731
rect 49896 17700 50353 17728
rect 49145 17691 49203 17697
rect 50341 17697 50353 17700
rect 50387 17697 50399 17731
rect 50341 17691 50399 17697
rect 50798 17688 50804 17740
rect 50856 17728 50862 17740
rect 51537 17731 51595 17737
rect 51537 17728 51549 17731
rect 50856 17700 51549 17728
rect 50856 17688 50862 17700
rect 51537 17697 51549 17700
rect 51583 17697 51595 17731
rect 51537 17691 51595 17697
rect 51626 17688 51632 17740
rect 51684 17728 51690 17740
rect 52917 17731 52975 17737
rect 51684 17700 51729 17728
rect 51684 17688 51690 17700
rect 52917 17697 52929 17731
rect 52963 17728 52975 17731
rect 53282 17728 53288 17740
rect 52963 17700 53288 17728
rect 52963 17697 52975 17700
rect 52917 17691 52975 17697
rect 53282 17688 53288 17700
rect 53340 17688 53346 17740
rect 47118 17620 47124 17672
rect 47176 17660 47182 17672
rect 51350 17660 51356 17672
rect 47176 17632 47221 17660
rect 51311 17632 51356 17660
rect 47176 17620 47182 17632
rect 51350 17620 51356 17632
rect 51408 17620 51414 17672
rect 52089 17663 52147 17669
rect 52089 17629 52101 17663
rect 52135 17660 52147 17663
rect 52362 17660 52368 17672
rect 52135 17632 52368 17660
rect 52135 17629 52147 17632
rect 52089 17623 52147 17629
rect 52362 17620 52368 17632
rect 52420 17620 52426 17672
rect 50246 17592 50252 17604
rect 47044 17564 50252 17592
rect 50246 17552 50252 17564
rect 50304 17592 50310 17604
rect 50433 17595 50491 17601
rect 50433 17592 50445 17595
rect 50304 17564 50445 17592
rect 50304 17552 50310 17564
rect 50433 17561 50445 17564
rect 50479 17561 50491 17595
rect 50433 17555 50491 17561
rect 43990 17524 43996 17536
rect 43763 17496 43996 17524
rect 43763 17493 43775 17496
rect 43717 17487 43775 17493
rect 43990 17484 43996 17496
rect 44048 17524 44054 17536
rect 45186 17524 45192 17536
rect 44048 17496 45192 17524
rect 44048 17484 44054 17496
rect 45186 17484 45192 17496
rect 45244 17484 45250 17536
rect 46474 17524 46480 17536
rect 46435 17496 46480 17524
rect 46474 17484 46480 17496
rect 46532 17484 46538 17536
rect 1104 17434 54832 17456
rect 1104 17382 9947 17434
rect 9999 17382 10011 17434
rect 10063 17382 10075 17434
rect 10127 17382 10139 17434
rect 10191 17382 27878 17434
rect 27930 17382 27942 17434
rect 27994 17382 28006 17434
rect 28058 17382 28070 17434
rect 28122 17382 45808 17434
rect 45860 17382 45872 17434
rect 45924 17382 45936 17434
rect 45988 17382 46000 17434
rect 46052 17382 54832 17434
rect 1104 17360 54832 17382
rect 2130 17320 2136 17332
rect 2091 17292 2136 17320
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 4801 17323 4859 17329
rect 4801 17320 4813 17323
rect 2332 17292 4813 17320
rect 2332 17125 2360 17292
rect 4801 17289 4813 17292
rect 4847 17320 4859 17323
rect 5258 17320 5264 17332
rect 4847 17292 5264 17320
rect 4847 17289 4859 17292
rect 4801 17283 4859 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 15013 17323 15071 17329
rect 15013 17320 15025 17323
rect 10888 17292 15025 17320
rect 8018 17212 8024 17264
rect 8076 17252 8082 17264
rect 8076 17224 10456 17252
rect 8076 17212 8082 17224
rect 7190 17184 7196 17196
rect 7151 17156 7196 17184
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 9582 17184 9588 17196
rect 7300 17156 9588 17184
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2590 17076 2596 17128
rect 2648 17116 2654 17128
rect 3329 17119 3387 17125
rect 3329 17116 3341 17119
rect 2648 17088 3341 17116
rect 2648 17076 2654 17088
rect 3329 17085 3341 17088
rect 3375 17085 3387 17119
rect 3329 17079 3387 17085
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 3881 17119 3939 17125
rect 3881 17085 3893 17119
rect 3927 17085 3939 17119
rect 3881 17079 3939 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17085 4399 17119
rect 4341 17079 4399 17085
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 7300 17116 7328 17156
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 9766 17184 9772 17196
rect 9727 17156 9772 17184
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10428 17128 10456 17224
rect 7558 17116 7564 17128
rect 4571 17088 7328 17116
rect 7519 17088 7564 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 3804 17048 3832 17079
rect 3160 17020 3832 17048
rect 3160 16989 3188 17020
rect 3145 16983 3203 16989
rect 3145 16949 3157 16983
rect 3191 16949 3203 16983
rect 3896 16980 3924 17079
rect 4062 17008 4068 17060
rect 4120 17048 4126 17060
rect 4356 17048 4384 17079
rect 4120 17020 4384 17048
rect 4120 17008 4126 17020
rect 4540 16980 4568 17079
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 7745 17119 7803 17125
rect 7745 17085 7757 17119
rect 7791 17116 7803 17119
rect 8018 17116 8024 17128
rect 7791 17088 8024 17116
rect 7791 17085 7803 17088
rect 7745 17079 7803 17085
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8294 17116 8300 17128
rect 8255 17088 8300 17116
rect 8113 17079 8171 17085
rect 8128 17048 8156 17079
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 10229 17119 10287 17125
rect 10229 17116 10241 17119
rect 9732 17088 10241 17116
rect 9732 17076 9738 17088
rect 10229 17085 10241 17088
rect 10275 17085 10287 17119
rect 10410 17116 10416 17128
rect 10323 17088 10416 17116
rect 10229 17079 10287 17085
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 10888 17125 10916 17292
rect 15013 17289 15025 17292
rect 15059 17289 15071 17323
rect 15013 17283 15071 17289
rect 16022 17280 16028 17332
rect 16080 17320 16086 17332
rect 16574 17320 16580 17332
rect 16080 17292 16580 17320
rect 16080 17280 16086 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 24946 17320 24952 17332
rect 24903 17292 24952 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 24946 17280 24952 17292
rect 25004 17280 25010 17332
rect 28261 17323 28319 17329
rect 27632 17292 28120 17320
rect 14274 17252 14280 17264
rect 14187 17224 14280 17252
rect 14274 17212 14280 17224
rect 14332 17252 14338 17264
rect 18690 17252 18696 17264
rect 14332 17224 18696 17252
rect 14332 17212 14338 17224
rect 18690 17212 18696 17224
rect 18748 17212 18754 17264
rect 19794 17252 19800 17264
rect 19260 17224 19800 17252
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 18877 17187 18935 17193
rect 18877 17184 18889 17187
rect 16540 17156 18889 17184
rect 16540 17144 16546 17156
rect 18877 17153 18889 17156
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 10781 17119 10839 17125
rect 10781 17116 10793 17119
rect 10744 17088 10793 17116
rect 10744 17076 10750 17088
rect 10781 17085 10793 17088
rect 10827 17085 10839 17119
rect 10781 17079 10839 17085
rect 10873 17119 10931 17125
rect 10873 17085 10885 17119
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 12713 17119 12771 17125
rect 12713 17085 12725 17119
rect 12759 17116 12771 17119
rect 14366 17116 14372 17128
rect 12759 17088 14372 17116
rect 12759 17085 12771 17088
rect 12713 17079 12771 17085
rect 8570 17048 8576 17060
rect 8128 17020 8576 17048
rect 8570 17008 8576 17020
rect 8628 17048 8634 17060
rect 10796 17048 10824 17079
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 15102 17076 15108 17128
rect 15160 17116 15166 17128
rect 15286 17116 15292 17128
rect 15160 17088 15292 17116
rect 15160 17076 15166 17088
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 16022 17116 16028 17128
rect 15519 17088 16028 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 16209 17119 16267 17125
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 17126 17116 17132 17128
rect 16255 17088 17132 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 8628 17020 10824 17048
rect 15013 17051 15071 17057
rect 8628 17008 8634 17020
rect 15013 17017 15025 17051
rect 15059 17048 15071 17051
rect 16224 17048 16252 17079
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 19061 17119 19119 17125
rect 19061 17085 19073 17119
rect 19107 17116 19119 17119
rect 19260 17116 19288 17224
rect 19794 17212 19800 17224
rect 19852 17252 19858 17264
rect 21177 17255 21235 17261
rect 21177 17252 21189 17255
rect 19852 17224 21189 17252
rect 19852 17212 19858 17224
rect 21177 17221 21189 17224
rect 21223 17221 21235 17255
rect 21177 17215 21235 17221
rect 24489 17255 24547 17261
rect 24489 17221 24501 17255
rect 24535 17252 24547 17255
rect 27632 17252 27660 17292
rect 24535 17224 27660 17252
rect 27893 17255 27951 17261
rect 24535 17221 24547 17224
rect 24489 17215 24547 17221
rect 27893 17221 27905 17255
rect 27939 17221 27951 17255
rect 28092 17252 28120 17292
rect 28261 17289 28273 17323
rect 28307 17320 28319 17323
rect 28350 17320 28356 17332
rect 28307 17292 28356 17320
rect 28307 17289 28319 17292
rect 28261 17283 28319 17289
rect 28350 17280 28356 17292
rect 28408 17280 28414 17332
rect 28442 17280 28448 17332
rect 28500 17320 28506 17332
rect 28537 17323 28595 17329
rect 28537 17320 28549 17323
rect 28500 17292 28549 17320
rect 28500 17280 28506 17292
rect 28537 17289 28549 17292
rect 28583 17320 28595 17323
rect 29822 17320 29828 17332
rect 28583 17292 29828 17320
rect 28583 17289 28595 17292
rect 28537 17283 28595 17289
rect 29822 17280 29828 17292
rect 29880 17280 29886 17332
rect 29914 17280 29920 17332
rect 29972 17320 29978 17332
rect 30745 17323 30803 17329
rect 30745 17320 30757 17323
rect 29972 17292 30757 17320
rect 29972 17280 29978 17292
rect 30745 17289 30757 17292
rect 30791 17289 30803 17323
rect 30745 17283 30803 17289
rect 31849 17323 31907 17329
rect 31849 17289 31861 17323
rect 31895 17320 31907 17323
rect 31938 17320 31944 17332
rect 31895 17292 31944 17320
rect 31895 17289 31907 17292
rect 31849 17283 31907 17289
rect 31938 17280 31944 17292
rect 31996 17280 32002 17332
rect 33318 17280 33324 17332
rect 33376 17320 33382 17332
rect 39022 17320 39028 17332
rect 33376 17292 39028 17320
rect 33376 17280 33382 17292
rect 39022 17280 39028 17292
rect 39080 17280 39086 17332
rect 41233 17323 41291 17329
rect 41233 17320 41245 17323
rect 39132 17292 41245 17320
rect 35989 17255 36047 17261
rect 35989 17252 36001 17255
rect 28092 17224 36001 17252
rect 27893 17215 27951 17221
rect 35989 17221 36001 17224
rect 36035 17221 36047 17255
rect 35989 17215 36047 17221
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17184 20223 17187
rect 24581 17187 24639 17193
rect 24581 17184 24593 17187
rect 20211 17156 24593 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 24581 17153 24593 17156
rect 24627 17153 24639 17187
rect 24581 17147 24639 17153
rect 19107 17088 19288 17116
rect 19521 17119 19579 17125
rect 19107 17085 19119 17088
rect 19061 17079 19119 17085
rect 19521 17085 19533 17119
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 15059 17020 16252 17048
rect 15059 17017 15071 17020
rect 15013 17011 15071 17017
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 19536 17048 19564 17079
rect 19610 17076 19616 17128
rect 19668 17116 19674 17128
rect 21085 17119 21143 17125
rect 19668 17088 19713 17116
rect 19668 17076 19674 17088
rect 21085 17085 21097 17119
rect 21131 17116 21143 17119
rect 22370 17116 22376 17128
rect 21131 17088 22376 17116
rect 21131 17085 21143 17088
rect 21085 17079 21143 17085
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 23290 17076 23296 17128
rect 23348 17116 23354 17128
rect 24213 17119 24271 17125
rect 24213 17116 24225 17119
rect 23348 17088 24225 17116
rect 23348 17076 23354 17088
rect 24213 17085 24225 17088
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 24360 17119 24418 17125
rect 24360 17085 24372 17119
rect 24406 17116 24418 17119
rect 25314 17116 25320 17128
rect 24406 17088 25320 17116
rect 24406 17085 24418 17088
rect 24360 17079 24418 17085
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 26234 17076 26240 17128
rect 26292 17116 26298 17128
rect 27764 17119 27822 17125
rect 27764 17116 27776 17119
rect 26292 17088 27776 17116
rect 26292 17076 26298 17088
rect 27764 17085 27776 17088
rect 27810 17085 27822 17119
rect 27908 17116 27936 17215
rect 36078 17212 36084 17264
rect 36136 17252 36142 17264
rect 39132 17252 39160 17292
rect 41233 17289 41245 17292
rect 41279 17289 41291 17323
rect 41233 17283 41291 17289
rect 41509 17323 41567 17329
rect 41509 17289 41521 17323
rect 41555 17320 41567 17323
rect 41690 17320 41696 17332
rect 41555 17292 41696 17320
rect 41555 17289 41567 17292
rect 41509 17283 41567 17289
rect 41690 17280 41696 17292
rect 41748 17320 41754 17332
rect 42242 17320 42248 17332
rect 41748 17292 42248 17320
rect 41748 17280 41754 17292
rect 42242 17280 42248 17292
rect 42300 17280 42306 17332
rect 44082 17320 44088 17332
rect 44043 17292 44088 17320
rect 44082 17280 44088 17292
rect 44140 17280 44146 17332
rect 44542 17280 44548 17332
rect 44600 17320 44606 17332
rect 45097 17323 45155 17329
rect 45097 17320 45109 17323
rect 44600 17292 45109 17320
rect 44600 17280 44606 17292
rect 45097 17289 45109 17292
rect 45143 17289 45155 17323
rect 45097 17283 45155 17289
rect 45186 17280 45192 17332
rect 45244 17320 45250 17332
rect 46845 17323 46903 17329
rect 46845 17320 46857 17323
rect 45244 17292 46857 17320
rect 45244 17280 45250 17292
rect 46845 17289 46857 17292
rect 46891 17320 46903 17323
rect 50890 17320 50896 17332
rect 46891 17292 50896 17320
rect 46891 17289 46903 17292
rect 46845 17283 46903 17289
rect 36136 17224 39160 17252
rect 36136 17212 36142 17224
rect 39206 17212 39212 17264
rect 39264 17252 39270 17264
rect 39853 17255 39911 17261
rect 39853 17252 39865 17255
rect 39264 17224 39865 17252
rect 39264 17212 39270 17224
rect 39853 17221 39865 17224
rect 39899 17252 39911 17255
rect 39942 17252 39948 17264
rect 39899 17224 39948 17252
rect 39899 17221 39911 17224
rect 39853 17215 39911 17221
rect 39942 17212 39948 17224
rect 40000 17252 40006 17264
rect 43990 17252 43996 17264
rect 40000 17224 43996 17252
rect 40000 17212 40006 17224
rect 43990 17212 43996 17224
rect 44048 17212 44054 17264
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17184 28043 17187
rect 29270 17184 29276 17196
rect 28031 17156 29276 17184
rect 28031 17153 28043 17156
rect 27985 17147 28043 17153
rect 29270 17144 29276 17156
rect 29328 17144 29334 17196
rect 29454 17184 29460 17196
rect 29415 17156 29460 17184
rect 29454 17144 29460 17156
rect 29512 17144 29518 17196
rect 30006 17184 30012 17196
rect 29564 17156 30012 17184
rect 28442 17116 28448 17128
rect 27908 17088 28448 17116
rect 27764 17079 27822 17085
rect 28442 17076 28448 17088
rect 28500 17076 28506 17128
rect 28534 17076 28540 17128
rect 28592 17116 28598 17128
rect 29564 17116 29592 17156
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 30374 17184 30380 17196
rect 30287 17156 30380 17184
rect 30374 17144 30380 17156
rect 30432 17144 30438 17196
rect 34514 17144 34520 17196
rect 34572 17184 34578 17196
rect 34609 17187 34667 17193
rect 34609 17184 34621 17187
rect 34572 17156 34621 17184
rect 34572 17144 34578 17156
rect 34609 17153 34621 17156
rect 34655 17184 34667 17187
rect 34885 17187 34943 17193
rect 34885 17184 34897 17187
rect 34655 17156 34897 17184
rect 34655 17153 34667 17156
rect 34609 17147 34667 17153
rect 34885 17153 34897 17156
rect 34931 17153 34943 17187
rect 34885 17147 34943 17153
rect 37553 17187 37611 17193
rect 37553 17153 37565 17187
rect 37599 17184 37611 17187
rect 37645 17187 37703 17193
rect 37645 17184 37657 17187
rect 37599 17156 37657 17184
rect 37599 17153 37611 17156
rect 37553 17147 37611 17153
rect 37645 17153 37657 17156
rect 37691 17184 37703 17187
rect 38010 17184 38016 17196
rect 37691 17156 38016 17184
rect 37691 17153 37703 17156
rect 37645 17147 37703 17153
rect 38010 17144 38016 17156
rect 38068 17144 38074 17196
rect 39298 17144 39304 17196
rect 39356 17184 39362 17196
rect 41598 17184 41604 17196
rect 39356 17156 40080 17184
rect 41559 17156 41604 17184
rect 39356 17144 39362 17156
rect 28592 17088 29592 17116
rect 28592 17076 28598 17088
rect 29638 17076 29644 17128
rect 29696 17116 29702 17128
rect 29914 17116 29920 17128
rect 29696 17088 29920 17116
rect 29696 17076 29702 17088
rect 29914 17076 29920 17088
rect 29972 17076 29978 17128
rect 30101 17119 30159 17125
rect 30101 17085 30113 17119
rect 30147 17085 30159 17119
rect 30101 17079 30159 17085
rect 27154 17048 27160 17060
rect 19300 17020 19564 17048
rect 21100 17020 27160 17048
rect 19300 17008 19306 17020
rect 21100 16992 21128 17020
rect 27154 17008 27160 17020
rect 27212 17008 27218 17060
rect 27614 17048 27620 17060
rect 27575 17020 27620 17048
rect 27614 17008 27620 17020
rect 27672 17008 27678 17060
rect 28994 17008 29000 17060
rect 29052 17048 29058 17060
rect 30116 17048 30144 17079
rect 29052 17020 30144 17048
rect 29052 17008 29058 17020
rect 3896 16952 4568 16980
rect 3145 16943 3203 16949
rect 5626 16940 5632 16992
rect 5684 16980 5690 16992
rect 11238 16980 11244 16992
rect 5684 16952 11244 16980
rect 5684 16940 5690 16952
rect 11238 16940 11244 16952
rect 11296 16940 11302 16992
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 14461 16983 14519 16989
rect 14461 16980 14473 16983
rect 14424 16952 14473 16980
rect 14424 16940 14430 16952
rect 14461 16949 14473 16952
rect 14507 16949 14519 16983
rect 15102 16980 15108 16992
rect 15063 16952 15108 16980
rect 14461 16943 14519 16949
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 16482 16980 16488 16992
rect 16443 16952 16488 16980
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 21082 16940 21088 16992
rect 21140 16940 21146 16992
rect 21266 16940 21272 16992
rect 21324 16980 21330 16992
rect 24578 16980 24584 16992
rect 21324 16952 24584 16980
rect 21324 16940 21330 16952
rect 24578 16940 24584 16952
rect 24636 16940 24642 16992
rect 28258 16940 28264 16992
rect 28316 16980 28322 16992
rect 29273 16983 29331 16989
rect 29273 16980 29285 16983
rect 28316 16952 29285 16980
rect 28316 16940 28322 16952
rect 29273 16949 29285 16952
rect 29319 16980 29331 16983
rect 30392 16980 30420 17144
rect 30469 17119 30527 17125
rect 30469 17085 30481 17119
rect 30515 17085 30527 17119
rect 30469 17079 30527 17085
rect 30484 17048 30512 17079
rect 31110 17076 31116 17128
rect 31168 17116 31174 17128
rect 31757 17119 31815 17125
rect 31757 17116 31769 17119
rect 31168 17088 31769 17116
rect 31168 17076 31174 17088
rect 31757 17085 31769 17088
rect 31803 17116 31815 17119
rect 33594 17116 33600 17128
rect 31803 17088 33600 17116
rect 31803 17085 31815 17088
rect 31757 17079 31815 17085
rect 33594 17076 33600 17088
rect 33652 17076 33658 17128
rect 35069 17119 35127 17125
rect 35069 17085 35081 17119
rect 35115 17085 35127 17119
rect 35618 17116 35624 17128
rect 35579 17088 35624 17116
rect 35069 17079 35127 17085
rect 32214 17048 32220 17060
rect 30484 17020 32220 17048
rect 32214 17008 32220 17020
rect 32272 17008 32278 17060
rect 33226 17008 33232 17060
rect 33284 17048 33290 17060
rect 35084 17048 35112 17079
rect 35618 17076 35624 17088
rect 35676 17076 35682 17128
rect 35805 17119 35863 17125
rect 35805 17085 35817 17119
rect 35851 17116 35863 17119
rect 35851 17088 36032 17116
rect 35851 17085 35863 17088
rect 35805 17079 35863 17085
rect 35894 17048 35900 17060
rect 33284 17020 35900 17048
rect 33284 17008 33290 17020
rect 35894 17008 35900 17020
rect 35952 17008 35958 17060
rect 36004 17048 36032 17088
rect 36078 17076 36084 17128
rect 36136 17116 36142 17128
rect 36357 17119 36415 17125
rect 36357 17116 36369 17119
rect 36136 17088 36369 17116
rect 36136 17076 36142 17088
rect 36357 17085 36369 17088
rect 36403 17116 36415 17119
rect 36446 17116 36452 17128
rect 36403 17088 36452 17116
rect 36403 17085 36415 17088
rect 36357 17079 36415 17085
rect 36446 17076 36452 17088
rect 36504 17076 36510 17128
rect 37826 17116 37832 17128
rect 37787 17088 37832 17116
rect 37826 17076 37832 17088
rect 37884 17076 37890 17128
rect 38289 17119 38347 17125
rect 38289 17085 38301 17119
rect 38335 17085 38347 17119
rect 38289 17079 38347 17085
rect 38381 17119 38439 17125
rect 38381 17085 38393 17119
rect 38427 17116 38439 17119
rect 39209 17119 39267 17125
rect 39209 17116 39221 17119
rect 38427 17088 39221 17116
rect 38427 17085 38439 17088
rect 38381 17079 38439 17085
rect 39209 17085 39221 17088
rect 39255 17116 39267 17119
rect 39482 17116 39488 17128
rect 39255 17088 39488 17116
rect 39255 17085 39267 17088
rect 39209 17079 39267 17085
rect 37182 17048 37188 17060
rect 36004 17020 37188 17048
rect 37182 17008 37188 17020
rect 37240 17008 37246 17060
rect 38304 17048 38332 17079
rect 39482 17076 39488 17088
rect 39540 17076 39546 17128
rect 40052 17125 40080 17156
rect 41598 17144 41604 17156
rect 41656 17144 41662 17196
rect 46474 17184 46480 17196
rect 41708 17156 41920 17184
rect 40037 17119 40095 17125
rect 40037 17085 40049 17119
rect 40083 17085 40095 17119
rect 40037 17079 40095 17085
rect 41233 17119 41291 17125
rect 41233 17085 41245 17119
rect 41279 17116 41291 17119
rect 41708 17116 41736 17156
rect 41279 17088 41736 17116
rect 41785 17119 41843 17125
rect 41279 17085 41291 17088
rect 41233 17079 41291 17085
rect 41785 17085 41797 17119
rect 41831 17085 41843 17119
rect 41892 17116 41920 17156
rect 44008 17156 46480 17184
rect 42242 17116 42248 17128
rect 41892 17088 42104 17116
rect 42203 17088 42248 17116
rect 41785 17079 41843 17085
rect 38746 17048 38752 17060
rect 38304 17020 38752 17048
rect 38746 17008 38752 17020
rect 38804 17008 38810 17060
rect 38933 17051 38991 17057
rect 38933 17017 38945 17051
rect 38979 17048 38991 17051
rect 39666 17048 39672 17060
rect 38979 17020 39672 17048
rect 38979 17017 38991 17020
rect 38933 17011 38991 17017
rect 39666 17008 39672 17020
rect 39724 17008 39730 17060
rect 29319 16952 30420 16980
rect 29319 16949 29331 16952
rect 29273 16943 29331 16949
rect 35618 16940 35624 16992
rect 35676 16980 35682 16992
rect 38102 16980 38108 16992
rect 35676 16952 38108 16980
rect 35676 16940 35682 16952
rect 38102 16940 38108 16952
rect 38160 16980 38166 16992
rect 39758 16980 39764 16992
rect 38160 16952 39764 16980
rect 38160 16940 38166 16952
rect 39758 16940 39764 16952
rect 39816 16940 39822 16992
rect 41800 16980 41828 17079
rect 42076 17048 42104 17088
rect 42242 17076 42248 17088
rect 42300 17076 42306 17128
rect 42337 17119 42395 17125
rect 42337 17085 42349 17119
rect 42383 17116 42395 17119
rect 42702 17116 42708 17128
rect 42383 17088 42708 17116
rect 42383 17085 42395 17088
rect 42337 17079 42395 17085
rect 42702 17076 42708 17088
rect 42760 17076 42766 17128
rect 44008 17125 44036 17156
rect 46474 17144 46480 17156
rect 46532 17144 46538 17196
rect 46952 17193 46980 17292
rect 50890 17280 50896 17292
rect 50948 17280 50954 17332
rect 48866 17212 48872 17264
rect 48924 17252 48930 17264
rect 50430 17252 50436 17264
rect 48924 17224 50436 17252
rect 48924 17212 48930 17224
rect 50430 17212 50436 17224
rect 50488 17252 50494 17264
rect 50488 17224 50936 17252
rect 50488 17212 50494 17224
rect 46937 17187 46995 17193
rect 46937 17153 46949 17187
rect 46983 17153 46995 17187
rect 50798 17184 50804 17196
rect 50759 17156 50804 17184
rect 46937 17147 46995 17153
rect 50798 17144 50804 17156
rect 50856 17144 50862 17196
rect 50908 17193 50936 17224
rect 50893 17187 50951 17193
rect 50893 17153 50905 17187
rect 50939 17184 50951 17187
rect 50982 17184 50988 17196
rect 50939 17156 50988 17184
rect 50939 17153 50951 17156
rect 50893 17147 50951 17153
rect 50982 17144 50988 17156
rect 51040 17144 51046 17196
rect 51074 17144 51080 17196
rect 51132 17184 51138 17196
rect 52362 17184 52368 17196
rect 51132 17156 52224 17184
rect 52323 17156 52368 17184
rect 51132 17144 51138 17156
rect 43993 17119 44051 17125
rect 43993 17085 44005 17119
rect 44039 17085 44051 17119
rect 43993 17079 44051 17085
rect 45005 17119 45063 17125
rect 45005 17085 45017 17119
rect 45051 17116 45063 17119
rect 45554 17116 45560 17128
rect 45051 17088 45560 17116
rect 45051 17085 45063 17088
rect 45005 17079 45063 17085
rect 45554 17076 45560 17088
rect 45612 17076 45618 17128
rect 47213 17119 47271 17125
rect 47213 17085 47225 17119
rect 47259 17116 47271 17119
rect 47486 17116 47492 17128
rect 47259 17088 47492 17116
rect 47259 17085 47271 17088
rect 47213 17079 47271 17085
rect 47486 17076 47492 17088
rect 47544 17076 47550 17128
rect 50246 17116 50252 17128
rect 50207 17088 50252 17116
rect 50246 17076 50252 17088
rect 50304 17076 50310 17128
rect 50430 17125 50436 17128
rect 50413 17119 50436 17125
rect 50413 17085 50425 17119
rect 50413 17079 50436 17085
rect 50430 17076 50436 17079
rect 50488 17076 50494 17128
rect 52089 17119 52147 17125
rect 52089 17116 52101 17119
rect 51920 17088 52101 17116
rect 42889 17051 42947 17057
rect 42889 17048 42901 17051
rect 42076 17020 42901 17048
rect 42889 17017 42901 17020
rect 42935 17017 42947 17051
rect 42889 17011 42947 17017
rect 42978 17008 42984 17060
rect 43036 17048 43042 17060
rect 43036 17020 44312 17048
rect 43036 17008 43042 17020
rect 44174 16980 44180 16992
rect 41800 16952 44180 16980
rect 44174 16940 44180 16952
rect 44232 16940 44238 16992
rect 44284 16980 44312 17020
rect 47946 17008 47952 17060
rect 48004 17048 48010 17060
rect 51350 17048 51356 17060
rect 48004 17020 51356 17048
rect 48004 17008 48010 17020
rect 51350 17008 51356 17020
rect 51408 17008 51414 17060
rect 48498 16980 48504 16992
rect 44284 16952 48504 16980
rect 48498 16940 48504 16952
rect 48556 16940 48562 16992
rect 51258 16940 51264 16992
rect 51316 16980 51322 16992
rect 51920 16989 51948 17088
rect 52089 17085 52101 17088
rect 52135 17085 52147 17119
rect 52196 17116 52224 17156
rect 52362 17144 52368 17156
rect 52420 17144 52426 17196
rect 53469 17187 53527 17193
rect 53469 17153 53481 17187
rect 53515 17153 53527 17187
rect 53469 17147 53527 17153
rect 53484 17116 53512 17147
rect 52196 17088 53512 17116
rect 52089 17079 52147 17085
rect 51905 16983 51963 16989
rect 51905 16980 51917 16983
rect 51316 16952 51917 16980
rect 51316 16940 51322 16952
rect 51905 16949 51917 16952
rect 51951 16949 51963 16983
rect 51905 16943 51963 16949
rect 1104 16890 54832 16912
rect 1104 16838 18912 16890
rect 18964 16838 18976 16890
rect 19028 16838 19040 16890
rect 19092 16838 19104 16890
rect 19156 16838 36843 16890
rect 36895 16838 36907 16890
rect 36959 16838 36971 16890
rect 37023 16838 37035 16890
rect 37087 16838 54832 16890
rect 1104 16816 54832 16838
rect 2590 16776 2596 16788
rect 2551 16748 2596 16776
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 4157 16779 4215 16785
rect 4157 16745 4169 16779
rect 4203 16776 4215 16779
rect 10781 16779 10839 16785
rect 4203 16748 8064 16776
rect 4203 16745 4215 16748
rect 4157 16739 4215 16745
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 3786 16640 3792 16652
rect 2832 16612 2877 16640
rect 3747 16612 3792 16640
rect 2832 16600 2838 16612
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 4062 16640 4068 16652
rect 4023 16612 4068 16640
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16640 5595 16643
rect 5626 16640 5632 16652
rect 5583 16612 5632 16640
rect 5583 16609 5595 16612
rect 5537 16603 5595 16609
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 5813 16643 5871 16649
rect 5813 16609 5825 16643
rect 5859 16640 5871 16643
rect 6362 16640 6368 16652
rect 5859 16612 6368 16640
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 6546 16640 6552 16652
rect 6459 16612 6552 16640
rect 6546 16600 6552 16612
rect 6604 16640 6610 16652
rect 7558 16640 7564 16652
rect 6604 16612 7564 16640
rect 6604 16600 6610 16612
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8036 16649 8064 16748
rect 10781 16745 10793 16779
rect 10827 16776 10839 16779
rect 11422 16776 11428 16788
rect 10827 16748 11428 16776
rect 10827 16745 10839 16748
rect 10781 16739 10839 16745
rect 11422 16736 11428 16748
rect 11480 16736 11486 16788
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 12400 16748 13461 16776
rect 12400 16736 12406 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13449 16739 13507 16745
rect 14568 16748 17172 16776
rect 10686 16668 10692 16720
rect 10744 16708 10750 16720
rect 10744 16680 11560 16708
rect 10744 16668 10750 16680
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 11532 16649 11560 16680
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 10468 16612 11161 16640
rect 10468 16600 10474 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16640 11759 16643
rect 13170 16640 13176 16652
rect 11747 16612 13176 16640
rect 11747 16609 11759 16612
rect 11701 16603 11759 16609
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16640 13415 16643
rect 14274 16640 14280 16652
rect 13403 16612 14280 16640
rect 13403 16609 13415 16612
rect 13357 16603 13415 16609
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 14568 16649 14596 16748
rect 14553 16643 14611 16649
rect 14553 16609 14565 16643
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 14918 16600 14924 16652
rect 14976 16640 14982 16652
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 14976 16612 16037 16640
rect 14976 16600 14982 16612
rect 16025 16609 16037 16612
rect 16071 16640 16083 16643
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 16071 16612 16221 16640
rect 16071 16609 16083 16612
rect 16025 16603 16083 16609
rect 16209 16609 16221 16612
rect 16255 16609 16267 16643
rect 16482 16640 16488 16652
rect 16443 16612 16488 16640
rect 16209 16603 16267 16609
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 17144 16640 17172 16748
rect 17218 16736 17224 16788
rect 17276 16776 17282 16788
rect 17773 16779 17831 16785
rect 17773 16776 17785 16779
rect 17276 16748 17785 16776
rect 17276 16736 17282 16748
rect 17773 16745 17785 16748
rect 17819 16776 17831 16779
rect 21266 16776 21272 16788
rect 17819 16748 21272 16776
rect 17819 16745 17831 16748
rect 17773 16739 17831 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 25777 16779 25835 16785
rect 25777 16776 25789 16779
rect 24504 16748 25789 16776
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 21637 16711 21695 16717
rect 21637 16708 21649 16711
rect 17920 16680 21649 16708
rect 17920 16668 17926 16680
rect 21637 16677 21649 16680
rect 21683 16708 21695 16711
rect 21821 16711 21879 16717
rect 21821 16708 21833 16711
rect 21683 16680 21833 16708
rect 21683 16677 21695 16680
rect 21637 16671 21695 16677
rect 21821 16677 21833 16680
rect 21867 16708 21879 16711
rect 21867 16680 22692 16708
rect 21867 16677 21879 16680
rect 21821 16671 21879 16677
rect 18046 16640 18052 16652
rect 17144 16612 18052 16640
rect 18046 16600 18052 16612
rect 18104 16640 18110 16652
rect 18877 16643 18935 16649
rect 18877 16640 18889 16643
rect 18104 16612 18889 16640
rect 18104 16600 18110 16612
rect 18877 16609 18889 16612
rect 18923 16609 18935 16643
rect 19334 16640 19340 16652
rect 19295 16612 19340 16640
rect 18877 16603 18935 16609
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 22020 16649 22048 16680
rect 22005 16643 22063 16649
rect 22005 16609 22017 16643
rect 22051 16640 22063 16643
rect 22189 16643 22247 16649
rect 22051 16612 22085 16640
rect 22051 16609 22063 16612
rect 22005 16603 22063 16609
rect 22189 16609 22201 16643
rect 22235 16640 22247 16643
rect 22554 16640 22560 16652
rect 22235 16612 22560 16640
rect 22235 16609 22247 16612
rect 22189 16603 22247 16609
rect 22554 16600 22560 16612
rect 22612 16600 22618 16652
rect 22664 16649 22692 16680
rect 22649 16643 22707 16649
rect 22649 16609 22661 16643
rect 22695 16609 22707 16643
rect 22649 16603 22707 16609
rect 22738 16600 22744 16652
rect 22796 16640 22802 16652
rect 23382 16640 23388 16652
rect 22796 16612 23388 16640
rect 22796 16600 22802 16612
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 24394 16640 24400 16652
rect 24355 16612 24400 16640
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 24504 16649 24532 16748
rect 25777 16745 25789 16748
rect 25823 16776 25835 16779
rect 28534 16776 28540 16788
rect 25823 16748 28540 16776
rect 25823 16745 25835 16748
rect 25777 16739 25835 16745
rect 28534 16736 28540 16748
rect 28592 16736 28598 16788
rect 28626 16736 28632 16788
rect 28684 16776 28690 16788
rect 28721 16779 28779 16785
rect 28721 16776 28733 16779
rect 28684 16748 28733 16776
rect 28684 16736 28690 16748
rect 28721 16745 28733 16748
rect 28767 16745 28779 16779
rect 30653 16779 30711 16785
rect 30653 16776 30665 16779
rect 28721 16739 28779 16745
rect 29104 16748 30665 16776
rect 24670 16668 24676 16720
rect 24728 16708 24734 16720
rect 28994 16708 29000 16720
rect 24728 16680 24992 16708
rect 24728 16668 24734 16680
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16609 24547 16643
rect 24489 16603 24547 16609
rect 24578 16600 24584 16652
rect 24636 16640 24642 16652
rect 24964 16649 24992 16680
rect 26712 16680 29000 16708
rect 24857 16643 24915 16649
rect 24857 16640 24869 16643
rect 24636 16612 24869 16640
rect 24636 16600 24642 16612
rect 24857 16609 24869 16612
rect 24903 16609 24915 16643
rect 24857 16603 24915 16609
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16609 25007 16643
rect 26510 16640 26516 16652
rect 26471 16612 26516 16640
rect 24949 16603 25007 16609
rect 26510 16600 26516 16612
rect 26568 16640 26574 16652
rect 26712 16649 26740 16680
rect 28994 16668 29000 16680
rect 29052 16668 29058 16720
rect 26697 16643 26755 16649
rect 26568 16612 26648 16640
rect 26568 16600 26574 16612
rect 11241 16575 11299 16581
rect 11241 16541 11253 16575
rect 11287 16541 11299 16575
rect 11241 16535 11299 16541
rect 11256 16504 11284 16535
rect 12342 16532 12348 16584
rect 12400 16572 12406 16584
rect 15102 16572 15108 16584
rect 12400 16544 15108 16572
rect 12400 16532 12406 16544
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 11698 16504 11704 16516
rect 11256 16476 11704 16504
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 18506 16464 18512 16516
rect 18564 16504 18570 16516
rect 18693 16507 18751 16513
rect 18693 16504 18705 16507
rect 18564 16476 18705 16504
rect 18564 16464 18570 16476
rect 18693 16473 18705 16476
rect 18739 16504 18751 16507
rect 18782 16504 18788 16516
rect 18739 16476 18788 16504
rect 18739 16473 18751 16476
rect 18693 16467 18751 16473
rect 18782 16464 18788 16476
rect 18840 16464 18846 16516
rect 25314 16504 25320 16516
rect 25275 16476 25320 16504
rect 25314 16464 25320 16476
rect 25372 16464 25378 16516
rect 26234 16504 26240 16516
rect 25516 16476 26240 16504
rect 3142 16396 3148 16448
rect 3200 16436 3206 16448
rect 3605 16439 3663 16445
rect 3605 16436 3617 16439
rect 3200 16408 3617 16436
rect 3200 16396 3206 16408
rect 3605 16405 3617 16408
rect 3651 16405 3663 16439
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 3605 16399 3663 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7837 16439 7895 16445
rect 7837 16436 7849 16439
rect 6972 16408 7849 16436
rect 6972 16396 6978 16408
rect 7837 16405 7849 16408
rect 7883 16405 7895 16439
rect 14366 16436 14372 16448
rect 14327 16408 14372 16436
rect 7837 16399 7895 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 19426 16436 19432 16448
rect 19387 16408 19432 16436
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 23201 16439 23259 16445
rect 23201 16405 23213 16439
rect 23247 16436 23259 16439
rect 25516 16436 25544 16476
rect 26234 16464 26240 16476
rect 26292 16464 26298 16516
rect 26620 16504 26648 16612
rect 26697 16609 26709 16643
rect 26743 16609 26755 16643
rect 27154 16640 27160 16652
rect 27115 16612 27160 16640
rect 26697 16603 26755 16609
rect 27154 16600 27160 16612
rect 27212 16600 27218 16652
rect 27249 16643 27307 16649
rect 27249 16609 27261 16643
rect 27295 16640 27307 16643
rect 27706 16640 27712 16652
rect 27295 16612 27712 16640
rect 27295 16609 27307 16612
rect 27249 16603 27307 16609
rect 27706 16600 27712 16612
rect 27764 16640 27770 16652
rect 28902 16640 28908 16652
rect 27764 16612 28908 16640
rect 27764 16600 27770 16612
rect 28902 16600 28908 16612
rect 28960 16600 28966 16652
rect 29104 16649 29132 16748
rect 30653 16745 30665 16748
rect 30699 16776 30711 16779
rect 33594 16776 33600 16788
rect 30699 16748 33180 16776
rect 33555 16748 33600 16776
rect 30699 16745 30711 16748
rect 30653 16739 30711 16745
rect 33152 16708 33180 16748
rect 33594 16736 33600 16748
rect 33652 16736 33658 16788
rect 33704 16748 36124 16776
rect 33704 16708 33732 16748
rect 29196 16680 30512 16708
rect 33152 16680 33732 16708
rect 29196 16649 29224 16680
rect 30484 16652 30512 16680
rect 29089 16643 29147 16649
rect 29089 16609 29101 16643
rect 29135 16609 29147 16643
rect 29089 16603 29147 16609
rect 29181 16643 29239 16649
rect 29181 16609 29193 16643
rect 29227 16609 29239 16643
rect 29454 16640 29460 16652
rect 29181 16603 29239 16609
rect 29288 16612 29460 16640
rect 29288 16572 29316 16612
rect 29454 16600 29460 16612
rect 29512 16600 29518 16652
rect 29546 16600 29552 16652
rect 29604 16640 29610 16652
rect 29641 16643 29699 16649
rect 29641 16640 29653 16643
rect 29604 16612 29653 16640
rect 29604 16600 29610 16612
rect 29641 16609 29653 16612
rect 29687 16609 29699 16643
rect 29641 16603 29699 16609
rect 29730 16600 29736 16652
rect 29788 16640 29794 16652
rect 29825 16643 29883 16649
rect 29825 16640 29837 16643
rect 29788 16612 29837 16640
rect 29788 16600 29794 16612
rect 29825 16609 29837 16612
rect 29871 16609 29883 16643
rect 30466 16640 30472 16652
rect 30427 16612 30472 16640
rect 29825 16603 29883 16609
rect 30466 16600 30472 16612
rect 30524 16600 30530 16652
rect 32217 16643 32275 16649
rect 32217 16609 32229 16643
rect 32263 16640 32275 16643
rect 32950 16640 32956 16652
rect 32263 16612 32956 16640
rect 32263 16609 32275 16612
rect 32217 16603 32275 16609
rect 32950 16600 32956 16612
rect 33008 16640 33014 16652
rect 34057 16643 34115 16649
rect 34057 16640 34069 16643
rect 33008 16612 34069 16640
rect 33008 16600 33014 16612
rect 34057 16609 34069 16612
rect 34103 16640 34115 16643
rect 35161 16643 35219 16649
rect 35161 16640 35173 16643
rect 34103 16612 35173 16640
rect 34103 16609 34115 16612
rect 34057 16603 34115 16609
rect 35161 16609 35173 16612
rect 35207 16640 35219 16643
rect 35802 16640 35808 16652
rect 35207 16612 35808 16640
rect 35207 16609 35219 16612
rect 35161 16603 35219 16609
rect 35802 16600 35808 16612
rect 35860 16600 35866 16652
rect 28000 16544 29316 16572
rect 32493 16575 32551 16581
rect 28000 16513 28028 16544
rect 32493 16541 32505 16575
rect 32539 16572 32551 16575
rect 32858 16572 32864 16584
rect 32539 16544 32864 16572
rect 32539 16541 32551 16544
rect 32493 16535 32551 16541
rect 32858 16532 32864 16544
rect 32916 16532 32922 16584
rect 35437 16575 35495 16581
rect 35437 16541 35449 16575
rect 35483 16572 35495 16575
rect 35894 16572 35900 16584
rect 35483 16544 35900 16572
rect 35483 16541 35495 16544
rect 35437 16535 35495 16541
rect 35894 16532 35900 16544
rect 35952 16532 35958 16584
rect 36096 16572 36124 16748
rect 37182 16736 37188 16788
rect 37240 16776 37246 16788
rect 42245 16779 42303 16785
rect 42245 16776 42257 16779
rect 37240 16748 42257 16776
rect 37240 16736 37246 16748
rect 42245 16745 42257 16748
rect 42291 16776 42303 16779
rect 42334 16776 42340 16788
rect 42291 16748 42340 16776
rect 42291 16745 42303 16748
rect 42245 16739 42303 16745
rect 42334 16736 42340 16748
rect 42392 16736 42398 16788
rect 47486 16776 47492 16788
rect 47447 16748 47492 16776
rect 47486 16736 47492 16748
rect 47544 16736 47550 16788
rect 39942 16708 39948 16720
rect 39903 16680 39948 16708
rect 39942 16668 39948 16680
rect 40000 16668 40006 16720
rect 40494 16668 40500 16720
rect 40552 16708 40558 16720
rect 40589 16711 40647 16717
rect 40589 16708 40601 16711
rect 40552 16680 40601 16708
rect 40552 16668 40558 16680
rect 40589 16677 40601 16680
rect 40635 16677 40647 16711
rect 47302 16708 47308 16720
rect 40589 16671 40647 16677
rect 40972 16680 47308 16708
rect 40770 16649 40776 16652
rect 40736 16643 40776 16649
rect 36648 16612 40632 16640
rect 36648 16572 36676 16612
rect 36096 16544 36676 16572
rect 38105 16575 38163 16581
rect 38105 16541 38117 16575
rect 38151 16541 38163 16575
rect 38378 16572 38384 16584
rect 38339 16544 38384 16572
rect 38105 16535 38163 16541
rect 27985 16507 28043 16513
rect 27985 16504 27997 16507
rect 26620 16476 27997 16504
rect 27985 16473 27997 16476
rect 28031 16473 28043 16507
rect 27985 16467 28043 16473
rect 29270 16464 29276 16516
rect 29328 16504 29334 16516
rect 30009 16507 30067 16513
rect 30009 16504 30021 16507
rect 29328 16476 30021 16504
rect 29328 16464 29334 16476
rect 30009 16473 30021 16476
rect 30055 16473 30067 16507
rect 30009 16467 30067 16473
rect 36354 16464 36360 16516
rect 36412 16504 36418 16516
rect 36541 16507 36599 16513
rect 36541 16504 36553 16507
rect 36412 16476 36553 16504
rect 36412 16464 36418 16476
rect 36541 16473 36553 16476
rect 36587 16473 36599 16507
rect 36541 16467 36599 16473
rect 25958 16436 25964 16448
rect 23247 16408 25544 16436
rect 25871 16408 25964 16436
rect 23247 16405 23259 16408
rect 23201 16399 23259 16405
rect 25958 16396 25964 16408
rect 26016 16436 26022 16448
rect 26878 16436 26884 16448
rect 26016 16408 26884 16436
rect 26016 16396 26022 16408
rect 26878 16396 26884 16408
rect 26936 16396 26942 16448
rect 27062 16396 27068 16448
rect 27120 16436 27126 16448
rect 27709 16439 27767 16445
rect 27709 16436 27721 16439
rect 27120 16408 27721 16436
rect 27120 16396 27126 16408
rect 27709 16405 27721 16408
rect 27755 16405 27767 16439
rect 27709 16399 27767 16405
rect 35802 16396 35808 16448
rect 35860 16436 35866 16448
rect 36446 16436 36452 16448
rect 35860 16408 36452 16436
rect 35860 16396 35866 16408
rect 36446 16396 36452 16408
rect 36504 16436 36510 16448
rect 36909 16439 36967 16445
rect 36909 16436 36921 16439
rect 36504 16408 36921 16436
rect 36504 16396 36510 16408
rect 36909 16405 36921 16408
rect 36955 16405 36967 16439
rect 38120 16436 38148 16535
rect 38378 16532 38384 16544
rect 38436 16532 38442 16584
rect 38746 16532 38752 16584
rect 38804 16572 38810 16584
rect 39114 16572 39120 16584
rect 38804 16544 39120 16572
rect 38804 16532 38810 16544
rect 39114 16532 39120 16544
rect 39172 16572 39178 16584
rect 39485 16575 39543 16581
rect 39485 16572 39497 16575
rect 39172 16544 39497 16572
rect 39172 16532 39178 16544
rect 39485 16541 39497 16544
rect 39531 16541 39543 16575
rect 39485 16535 39543 16541
rect 39666 16532 39672 16584
rect 39724 16572 39730 16584
rect 40494 16572 40500 16584
rect 39724 16544 40500 16572
rect 39724 16532 39730 16544
rect 40494 16532 40500 16544
rect 40552 16532 40558 16584
rect 40604 16504 40632 16612
rect 40736 16609 40748 16643
rect 40736 16603 40776 16609
rect 40770 16600 40776 16603
rect 40828 16600 40834 16652
rect 40972 16581 41000 16680
rect 47302 16668 47308 16680
rect 47360 16668 47366 16720
rect 49050 16668 49056 16720
rect 49108 16708 49114 16720
rect 53285 16711 53343 16717
rect 53285 16708 53297 16711
rect 49108 16680 53297 16708
rect 49108 16668 49114 16680
rect 41046 16600 41052 16652
rect 41104 16640 41110 16652
rect 41325 16643 41383 16649
rect 41325 16640 41337 16643
rect 41104 16612 41337 16640
rect 41104 16600 41110 16612
rect 41325 16609 41337 16612
rect 41371 16609 41383 16643
rect 41325 16603 41383 16609
rect 41782 16600 41788 16652
rect 41840 16640 41846 16652
rect 42153 16643 42211 16649
rect 42153 16640 42165 16643
rect 41840 16612 42165 16640
rect 41840 16600 41846 16612
rect 42153 16609 42165 16612
rect 42199 16609 42211 16643
rect 42153 16603 42211 16609
rect 43349 16643 43407 16649
rect 43349 16609 43361 16643
rect 43395 16640 43407 16643
rect 44634 16640 44640 16652
rect 43395 16612 44640 16640
rect 43395 16609 43407 16612
rect 43349 16603 43407 16609
rect 40957 16575 41015 16581
rect 40957 16541 40969 16575
rect 41003 16541 41015 16575
rect 40957 16535 41015 16541
rect 42058 16532 42064 16584
rect 42116 16572 42122 16584
rect 43364 16572 43392 16603
rect 44634 16600 44640 16612
rect 44692 16640 44698 16652
rect 45462 16640 45468 16652
rect 44692 16612 45468 16640
rect 44692 16600 44698 16612
rect 45462 16600 45468 16612
rect 45520 16600 45526 16652
rect 47394 16640 47400 16652
rect 47355 16612 47400 16640
rect 47394 16600 47400 16612
rect 47452 16600 47458 16652
rect 48498 16600 48504 16652
rect 48556 16640 48562 16652
rect 48961 16643 49019 16649
rect 48961 16640 48973 16643
rect 48556 16612 48973 16640
rect 48556 16600 48562 16612
rect 48961 16609 48973 16612
rect 49007 16609 49019 16643
rect 48961 16603 49019 16609
rect 50154 16600 50160 16652
rect 50212 16640 50218 16652
rect 50448 16649 50476 16680
rect 53285 16677 53297 16680
rect 53331 16677 53343 16711
rect 53285 16671 53343 16677
rect 50249 16643 50307 16649
rect 50249 16640 50261 16643
rect 50212 16612 50261 16640
rect 50212 16600 50218 16612
rect 50249 16609 50261 16612
rect 50295 16609 50307 16643
rect 50249 16603 50307 16609
rect 50433 16643 50491 16649
rect 50433 16609 50445 16643
rect 50479 16609 50491 16643
rect 50433 16603 50491 16609
rect 51442 16600 51448 16652
rect 51500 16640 51506 16652
rect 51629 16643 51687 16649
rect 51629 16640 51641 16643
rect 51500 16612 51641 16640
rect 51500 16600 51506 16612
rect 51629 16609 51641 16612
rect 51675 16609 51687 16643
rect 51629 16603 51687 16609
rect 51718 16600 51724 16652
rect 51776 16640 51782 16652
rect 51813 16643 51871 16649
rect 51813 16640 51825 16643
rect 51776 16612 51825 16640
rect 51776 16600 51782 16612
rect 51813 16609 51825 16612
rect 51859 16609 51871 16643
rect 51813 16603 51871 16609
rect 51905 16643 51963 16649
rect 51905 16609 51917 16643
rect 51951 16609 51963 16643
rect 51905 16603 51963 16609
rect 53193 16643 53251 16649
rect 53193 16609 53205 16643
rect 53239 16609 53251 16643
rect 53193 16603 53251 16609
rect 42116 16544 43392 16572
rect 50801 16575 50859 16581
rect 42116 16532 42122 16544
rect 50801 16541 50813 16575
rect 50847 16572 50859 16575
rect 51920 16572 51948 16603
rect 52362 16572 52368 16584
rect 50847 16544 51948 16572
rect 52323 16544 52368 16572
rect 50847 16541 50859 16544
rect 50801 16535 50859 16541
rect 52362 16532 52368 16544
rect 52420 16532 52426 16584
rect 42886 16504 42892 16516
rect 40604 16476 42892 16504
rect 42886 16464 42892 16476
rect 42944 16464 42950 16516
rect 50890 16464 50896 16516
rect 50948 16504 50954 16516
rect 51258 16504 51264 16516
rect 50948 16476 51264 16504
rect 50948 16464 50954 16476
rect 51258 16464 51264 16476
rect 51316 16464 51322 16516
rect 51350 16464 51356 16516
rect 51408 16504 51414 16516
rect 53208 16504 53236 16603
rect 53466 16504 53472 16516
rect 51408 16476 53472 16504
rect 51408 16464 51414 16476
rect 53466 16464 53472 16476
rect 53524 16464 53530 16516
rect 39942 16436 39948 16448
rect 38120 16408 39948 16436
rect 36909 16399 36967 16405
rect 39942 16396 39948 16408
rect 40000 16396 40006 16448
rect 40310 16396 40316 16448
rect 40368 16436 40374 16448
rect 40405 16439 40463 16445
rect 40405 16436 40417 16439
rect 40368 16408 40417 16436
rect 40368 16396 40374 16408
rect 40405 16405 40417 16408
rect 40451 16436 40463 16439
rect 40865 16439 40923 16445
rect 40865 16436 40877 16439
rect 40451 16408 40877 16436
rect 40451 16405 40463 16408
rect 40405 16399 40463 16405
rect 40865 16405 40877 16408
rect 40911 16405 40923 16439
rect 40865 16399 40923 16405
rect 42702 16396 42708 16448
rect 42760 16436 42766 16448
rect 43441 16439 43499 16445
rect 43441 16436 43453 16439
rect 42760 16408 43453 16436
rect 42760 16396 42766 16408
rect 43441 16405 43453 16408
rect 43487 16405 43499 16439
rect 43441 16399 43499 16405
rect 48590 16396 48596 16448
rect 48648 16436 48654 16448
rect 49053 16439 49111 16445
rect 49053 16436 49065 16439
rect 48648 16408 49065 16436
rect 48648 16396 48654 16408
rect 49053 16405 49065 16408
rect 49099 16405 49111 16439
rect 49053 16399 49111 16405
rect 1104 16346 54832 16368
rect 1104 16294 9947 16346
rect 9999 16294 10011 16346
rect 10063 16294 10075 16346
rect 10127 16294 10139 16346
rect 10191 16294 27878 16346
rect 27930 16294 27942 16346
rect 27994 16294 28006 16346
rect 28058 16294 28070 16346
rect 28122 16294 45808 16346
rect 45860 16294 45872 16346
rect 45924 16294 45936 16346
rect 45988 16294 46000 16346
rect 46052 16294 54832 16346
rect 1104 16272 54832 16294
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 4709 16235 4767 16241
rect 4709 16232 4721 16235
rect 4212 16204 4721 16232
rect 4212 16192 4218 16204
rect 4709 16201 4721 16204
rect 4755 16232 4767 16235
rect 6546 16232 6552 16244
rect 4755 16204 6552 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 8754 16192 8760 16244
rect 8812 16232 8818 16244
rect 8849 16235 8907 16241
rect 8849 16232 8861 16235
rect 8812 16204 8861 16232
rect 8812 16192 8818 16204
rect 8849 16201 8861 16204
rect 8895 16201 8907 16235
rect 8849 16195 8907 16201
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 13906 16232 13912 16244
rect 12032 16204 13912 16232
rect 12032 16192 12038 16204
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 15286 16232 15292 16244
rect 14875 16204 15292 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 15286 16192 15292 16204
rect 15344 16232 15350 16244
rect 25685 16235 25743 16241
rect 15344 16204 24900 16232
rect 15344 16192 15350 16204
rect 6730 16124 6736 16176
rect 6788 16164 6794 16176
rect 6788 16136 7144 16164
rect 6788 16124 6794 16136
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 6822 16096 6828 16108
rect 2455 16068 6828 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 2866 16028 2872 16040
rect 2179 16000 2872 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2866 15988 2872 16000
rect 2924 16028 2930 16040
rect 3789 16031 3847 16037
rect 2924 16000 3740 16028
rect 2924 15988 2930 16000
rect 3712 15960 3740 16000
rect 3789 15997 3801 16031
rect 3835 16028 3847 16031
rect 3878 16028 3884 16040
rect 3835 16000 3884 16028
rect 3835 15997 3847 16000
rect 3789 15991 3847 15997
rect 3878 15988 3884 16000
rect 3936 16028 3942 16040
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 3936 16000 4629 16028
rect 3936 15988 3942 16000
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 6914 16028 6920 16040
rect 5859 16000 6920 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 7116 16037 7144 16136
rect 8018 16124 8024 16176
rect 8076 16164 8082 16176
rect 19426 16164 19432 16176
rect 8076 16136 9260 16164
rect 8076 16124 8082 16136
rect 7101 16031 7159 16037
rect 7101 15997 7113 16031
rect 7147 15997 7159 16031
rect 9030 16028 9036 16040
rect 8991 16000 9036 16028
rect 7101 15991 7159 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 9232 16037 9260 16136
rect 16132 16136 19432 16164
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 16132 16096 16160 16136
rect 19426 16124 19432 16136
rect 19484 16164 19490 16176
rect 19484 16136 21496 16164
rect 19484 16124 19490 16136
rect 19518 16096 19524 16108
rect 13228 16068 16160 16096
rect 13228 16056 13234 16068
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 15997 9643 16031
rect 9585 15991 9643 15997
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 16028 9827 16031
rect 10781 16031 10839 16037
rect 10781 16028 10793 16031
rect 9815 16000 9996 16028
rect 9815 15997 9827 16000
rect 9769 15991 9827 15997
rect 3970 15960 3976 15972
rect 3712 15932 3976 15960
rect 3970 15920 3976 15932
rect 4028 15920 4034 15972
rect 8570 15920 8576 15972
rect 8628 15960 8634 15972
rect 9600 15960 9628 15991
rect 8628 15932 9628 15960
rect 8628 15920 8634 15932
rect 9968 15904 9996 16000
rect 10428 16000 10793 16028
rect 10428 15904 10456 16000
rect 10781 15997 10793 16000
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 15997 13323 16031
rect 13538 16028 13544 16040
rect 13499 16000 13544 16028
rect 13265 15991 13323 15997
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5629 15895 5687 15901
rect 5629 15892 5641 15895
rect 5040 15864 5641 15892
rect 5040 15852 5046 15864
rect 5629 15861 5641 15864
rect 5675 15861 5687 15895
rect 5629 15855 5687 15861
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7558 15892 7564 15904
rect 7331 15864 7564 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7558 15852 7564 15864
rect 7616 15852 7622 15904
rect 9950 15892 9956 15904
rect 9911 15864 9956 15892
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10410 15892 10416 15904
rect 10371 15864 10416 15892
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 10597 15895 10655 15901
rect 10597 15892 10609 15895
rect 10560 15864 10609 15892
rect 10560 15852 10566 15864
rect 10597 15861 10609 15864
rect 10643 15861 10655 15895
rect 13280 15892 13308 15991
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 15997 15991 16031
rect 16132 16028 16160 16068
rect 19352 16068 19524 16096
rect 16393 16031 16451 16037
rect 16393 16028 16405 16031
rect 16132 16000 16405 16028
rect 15933 15991 15991 15997
rect 16393 15997 16405 16000
rect 16439 15997 16451 16031
rect 16393 15991 16451 15997
rect 16485 16031 16543 16037
rect 16485 15997 16497 16031
rect 16531 16028 16543 16031
rect 16574 16028 16580 16040
rect 16531 16000 16580 16028
rect 16531 15997 16543 16000
rect 16485 15991 16543 15997
rect 14366 15892 14372 15904
rect 13280 15864 14372 15892
rect 10597 15855 10655 15861
rect 14366 15852 14372 15864
rect 14424 15892 14430 15904
rect 14918 15892 14924 15904
rect 14424 15864 14924 15892
rect 14424 15852 14430 15864
rect 14918 15852 14924 15864
rect 14976 15892 14982 15904
rect 15013 15895 15071 15901
rect 15013 15892 15025 15895
rect 14976 15864 15025 15892
rect 14976 15852 14982 15864
rect 15013 15861 15025 15864
rect 15059 15861 15071 15895
rect 15013 15855 15071 15861
rect 15470 15852 15476 15904
rect 15528 15892 15534 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15528 15864 15669 15892
rect 15528 15852 15534 15864
rect 15657 15861 15669 15864
rect 15703 15892 15715 15895
rect 15764 15892 15792 15991
rect 15948 15960 15976 15991
rect 16500 15960 16528 15991
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 19352 16037 19380 16068
rect 19518 16056 19524 16068
rect 19576 16056 19582 16108
rect 21468 16105 21496 16136
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16065 21511 16099
rect 24578 16096 24584 16108
rect 24539 16068 24584 16096
rect 21453 16059 21511 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 18969 16031 19027 16037
rect 18969 16028 18981 16031
rect 18616 16000 18981 16028
rect 17034 15960 17040 15972
rect 15948 15932 16528 15960
rect 16995 15932 17040 15960
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 18616 15904 18644 16000
rect 18969 15997 18981 16000
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 19337 16031 19395 16037
rect 19337 15997 19349 16031
rect 19383 15997 19395 16031
rect 19337 15991 19395 15997
rect 19429 16031 19487 16037
rect 19429 15997 19441 16031
rect 19475 16028 19487 16031
rect 19475 16000 19656 16028
rect 19475 15997 19487 16000
rect 19429 15991 19487 15997
rect 18690 15920 18696 15972
rect 18748 15960 18754 15972
rect 19628 15960 19656 16000
rect 19702 15988 19708 16040
rect 19760 16028 19766 16040
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 19760 16000 19809 16028
rect 19760 15988 19766 16000
rect 19797 15997 19809 16000
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 19886 15988 19892 16040
rect 19944 16028 19950 16040
rect 21542 16028 21548 16040
rect 19944 16000 19989 16028
rect 21503 16000 21548 16028
rect 19944 15988 19950 16000
rect 21542 15988 21548 16000
rect 21600 15988 21606 16040
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 21692 16000 22017 16028
rect 21692 15988 21698 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 24670 16028 24676 16040
rect 22152 16000 22197 16028
rect 24631 16000 24676 16028
rect 22152 15988 22158 16000
rect 24670 15988 24676 16000
rect 24728 15988 24734 16040
rect 24872 16028 24900 16204
rect 25685 16201 25697 16235
rect 25731 16232 25743 16235
rect 26973 16235 27031 16241
rect 26973 16232 26985 16235
rect 25731 16204 26985 16232
rect 25731 16201 25743 16204
rect 25685 16195 25743 16201
rect 26973 16201 26985 16204
rect 27019 16201 27031 16235
rect 27338 16232 27344 16244
rect 27299 16204 27344 16232
rect 26973 16195 27031 16201
rect 27338 16192 27344 16204
rect 27396 16192 27402 16244
rect 28902 16192 28908 16244
rect 28960 16232 28966 16244
rect 29365 16235 29423 16241
rect 29365 16232 29377 16235
rect 28960 16204 29377 16232
rect 28960 16192 28966 16204
rect 29365 16201 29377 16204
rect 29411 16201 29423 16235
rect 32858 16232 32864 16244
rect 32819 16204 32864 16232
rect 29365 16195 29423 16201
rect 32858 16192 32864 16204
rect 32916 16192 32922 16244
rect 35894 16232 35900 16244
rect 35855 16204 35900 16232
rect 35894 16192 35900 16204
rect 35952 16192 35958 16244
rect 39209 16235 39267 16241
rect 39209 16201 39221 16235
rect 39255 16232 39267 16235
rect 39390 16232 39396 16244
rect 39255 16204 39396 16232
rect 39255 16201 39267 16204
rect 39209 16195 39267 16201
rect 39390 16192 39396 16204
rect 39448 16192 39454 16244
rect 47394 16192 47400 16244
rect 47452 16232 47458 16244
rect 47673 16235 47731 16241
rect 47673 16232 47685 16235
rect 47452 16204 47685 16232
rect 47452 16192 47458 16204
rect 47673 16201 47685 16204
rect 47719 16201 47731 16235
rect 53466 16232 53472 16244
rect 53427 16204 53472 16232
rect 47673 16195 47731 16201
rect 53466 16192 53472 16204
rect 53524 16192 53530 16244
rect 32401 16167 32459 16173
rect 32401 16133 32413 16167
rect 32447 16164 32459 16167
rect 50614 16164 50620 16176
rect 32447 16136 35572 16164
rect 32447 16133 32459 16136
rect 32401 16127 32459 16133
rect 27062 16096 27068 16108
rect 27023 16068 27068 16096
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 31573 16099 31631 16105
rect 31573 16065 31585 16099
rect 31619 16096 31631 16099
rect 31619 16068 32720 16096
rect 31619 16065 31631 16068
rect 31573 16059 31631 16065
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24872 16000 25145 16028
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 25225 16031 25283 16037
rect 25225 15997 25237 16031
rect 25271 16028 25283 16031
rect 26234 16028 26240 16040
rect 25271 16000 26240 16028
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 26234 15988 26240 16000
rect 26292 15988 26298 16040
rect 26418 15988 26424 16040
rect 26476 16028 26482 16040
rect 26844 16031 26902 16037
rect 26844 16028 26856 16031
rect 26476 16000 26856 16028
rect 26476 15988 26482 16000
rect 26844 15997 26856 16000
rect 26890 15997 26902 16031
rect 26844 15991 26902 15997
rect 29273 16031 29331 16037
rect 29273 15997 29285 16031
rect 29319 16028 29331 16031
rect 29546 16028 29552 16040
rect 29319 16000 29552 16028
rect 29319 15997 29331 16000
rect 29273 15991 29331 15997
rect 29546 15988 29552 16000
rect 29604 15988 29610 16040
rect 31110 15988 31116 16040
rect 31168 16028 31174 16040
rect 32692 16037 32720 16068
rect 35544 16040 35572 16136
rect 48240 16136 50620 16164
rect 41782 16056 41788 16108
rect 41840 16096 41846 16108
rect 42702 16096 42708 16108
rect 41840 16068 42708 16096
rect 41840 16056 41846 16068
rect 42702 16056 42708 16068
rect 42760 16096 42766 16108
rect 43349 16099 43407 16105
rect 43349 16096 43361 16099
rect 42760 16068 43361 16096
rect 42760 16056 42766 16068
rect 43349 16065 43361 16068
rect 43395 16065 43407 16099
rect 43349 16059 43407 16065
rect 47026 16056 47032 16108
rect 47084 16096 47090 16108
rect 48130 16096 48136 16108
rect 47084 16068 48136 16096
rect 47084 16056 47090 16068
rect 48130 16056 48136 16068
rect 48188 16056 48194 16108
rect 31205 16031 31263 16037
rect 31205 16028 31217 16031
rect 31168 16000 31217 16028
rect 31168 15988 31174 16000
rect 31205 15997 31217 16000
rect 31251 15997 31263 16031
rect 31205 15991 31263 15997
rect 32677 16031 32735 16037
rect 32677 15997 32689 16031
rect 32723 15997 32735 16031
rect 35526 16028 35532 16040
rect 35487 16000 35532 16028
rect 32677 15991 32735 15997
rect 35526 15988 35532 16000
rect 35584 15988 35590 16040
rect 35713 16031 35771 16037
rect 35713 15997 35725 16031
rect 35759 16028 35771 16031
rect 35802 16028 35808 16040
rect 35759 16000 35808 16028
rect 35759 15997 35771 16000
rect 35713 15991 35771 15997
rect 35802 15988 35808 16000
rect 35860 15988 35866 16040
rect 39114 16028 39120 16040
rect 39075 16000 39120 16028
rect 39114 15988 39120 16000
rect 39172 15988 39178 16040
rect 42058 16028 42064 16040
rect 42019 16000 42064 16028
rect 42058 15988 42064 16000
rect 42116 15988 42122 16040
rect 42794 15988 42800 16040
rect 42852 16028 42858 16040
rect 43257 16031 43315 16037
rect 43257 16028 43269 16031
rect 42852 16000 43269 16028
rect 42852 15988 42858 16000
rect 43257 15997 43269 16000
rect 43303 15997 43315 16031
rect 43530 16028 43536 16040
rect 43491 16000 43536 16028
rect 43257 15991 43315 15997
rect 43530 15988 43536 16000
rect 43588 15988 43594 16040
rect 48240 16037 48268 16136
rect 50614 16124 50620 16136
rect 50672 16124 50678 16176
rect 52362 16096 52368 16108
rect 48608 16068 49832 16096
rect 52323 16068 52368 16096
rect 48608 16040 48636 16068
rect 48225 16031 48283 16037
rect 48225 15997 48237 16031
rect 48271 15997 48283 16031
rect 48590 16028 48596 16040
rect 48551 16000 48596 16028
rect 48225 15991 48283 15997
rect 48590 15988 48596 16000
rect 48648 15988 48654 16040
rect 49804 16037 49832 16068
rect 52362 16056 52368 16068
rect 52420 16056 52426 16108
rect 48685 16031 48743 16037
rect 48685 15997 48697 16031
rect 48731 15997 48743 16031
rect 48685 15991 48743 15997
rect 49789 16031 49847 16037
rect 49789 15997 49801 16031
rect 49835 15997 49847 16031
rect 49789 15991 49847 15997
rect 18748 15932 19656 15960
rect 18748 15920 18754 15932
rect 16758 15892 16764 15904
rect 15703 15864 16764 15892
rect 15703 15861 15715 15864
rect 15657 15855 15715 15861
rect 16758 15852 16764 15864
rect 16816 15852 16822 15904
rect 18598 15892 18604 15904
rect 18559 15864 18604 15892
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 18782 15892 18788 15904
rect 18743 15864 18788 15892
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 19628 15892 19656 15932
rect 20441 15963 20499 15969
rect 20441 15929 20453 15963
rect 20487 15960 20499 15963
rect 26697 15963 26755 15969
rect 26697 15960 26709 15963
rect 20487 15932 26709 15960
rect 20487 15929 20499 15932
rect 20441 15923 20499 15929
rect 26697 15929 26709 15932
rect 26743 15929 26755 15963
rect 26697 15923 26755 15929
rect 30742 15920 30748 15972
rect 30800 15960 30806 15972
rect 31021 15963 31079 15969
rect 31021 15960 31033 15963
rect 30800 15932 31033 15960
rect 30800 15920 30806 15932
rect 31021 15929 31033 15932
rect 31067 15929 31079 15963
rect 31021 15923 31079 15929
rect 32585 15963 32643 15969
rect 32585 15929 32597 15963
rect 32631 15960 32643 15963
rect 33962 15960 33968 15972
rect 32631 15932 33968 15960
rect 32631 15929 32643 15932
rect 32585 15923 32643 15929
rect 33962 15920 33968 15932
rect 34020 15920 34026 15972
rect 35618 15960 35624 15972
rect 35579 15932 35624 15960
rect 35618 15920 35624 15932
rect 35676 15920 35682 15972
rect 41874 15960 41880 15972
rect 41835 15932 41880 15960
rect 41874 15920 41880 15932
rect 41932 15920 41938 15972
rect 43993 15963 44051 15969
rect 43993 15929 44005 15963
rect 44039 15960 44051 15963
rect 48700 15960 48728 15991
rect 51258 15988 51264 16040
rect 51316 16028 51322 16040
rect 52089 16031 52147 16037
rect 52089 16028 52101 16031
rect 51316 16000 52101 16028
rect 51316 15988 51322 16000
rect 48958 15960 48964 15972
rect 44039 15932 48964 15960
rect 44039 15929 44051 15932
rect 43993 15923 44051 15929
rect 48958 15920 48964 15932
rect 49016 15960 49022 15972
rect 49605 15963 49663 15969
rect 49605 15960 49617 15963
rect 49016 15932 49617 15960
rect 49016 15920 49022 15932
rect 49605 15929 49617 15932
rect 49651 15929 49663 15963
rect 50154 15960 50160 15972
rect 50115 15932 50160 15960
rect 49605 15923 49663 15929
rect 50154 15920 50160 15932
rect 50212 15920 50218 15972
rect 21634 15892 21640 15904
rect 19628 15864 21640 15892
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 22557 15895 22615 15901
rect 22557 15861 22569 15895
rect 22603 15892 22615 15895
rect 29730 15892 29736 15904
rect 22603 15864 29736 15892
rect 22603 15861 22615 15864
rect 22557 15855 22615 15861
rect 29730 15852 29736 15864
rect 29788 15852 29794 15904
rect 42150 15892 42156 15904
rect 42111 15864 42156 15892
rect 42150 15852 42156 15864
rect 42208 15852 42214 15904
rect 51810 15852 51816 15904
rect 51868 15892 51874 15904
rect 51920 15901 51948 16000
rect 52089 15997 52101 16000
rect 52135 15997 52147 16031
rect 52089 15991 52147 15997
rect 51905 15895 51963 15901
rect 51905 15892 51917 15895
rect 51868 15864 51917 15892
rect 51868 15852 51874 15864
rect 51905 15861 51917 15864
rect 51951 15861 51963 15895
rect 51905 15855 51963 15861
rect 1104 15802 54832 15824
rect 1104 15750 18912 15802
rect 18964 15750 18976 15802
rect 19028 15750 19040 15802
rect 19092 15750 19104 15802
rect 19156 15750 36843 15802
rect 36895 15750 36907 15802
rect 36959 15750 36971 15802
rect 37023 15750 37035 15802
rect 37087 15750 54832 15802
rect 1104 15728 54832 15750
rect 2133 15691 2191 15697
rect 2133 15657 2145 15691
rect 2179 15688 2191 15691
rect 2774 15688 2780 15700
rect 2179 15660 2780 15688
rect 2179 15657 2191 15660
rect 2133 15651 2191 15657
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 3145 15691 3203 15697
rect 3145 15657 3157 15691
rect 3191 15688 3203 15691
rect 3786 15688 3792 15700
rect 3191 15660 3792 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 3786 15648 3792 15660
rect 3844 15648 3850 15700
rect 7650 15688 7656 15700
rect 6012 15660 7512 15688
rect 7611 15660 7656 15688
rect 2498 15580 2504 15632
rect 2556 15620 2562 15632
rect 6012 15620 6040 15660
rect 6362 15620 6368 15632
rect 2556 15592 6040 15620
rect 6104 15592 6368 15620
rect 2556 15580 2562 15592
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15552 2375 15555
rect 3142 15552 3148 15564
rect 2363 15524 3148 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 3329 15555 3387 15561
rect 3329 15521 3341 15555
rect 3375 15552 3387 15555
rect 4982 15552 4988 15564
rect 3375 15524 4844 15552
rect 4943 15524 4988 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 4816 15425 4844 15524
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 6104 15561 6132 15592
rect 6362 15580 6368 15592
rect 6420 15580 6426 15632
rect 7484 15620 7512 15660
rect 7650 15648 7656 15660
rect 7708 15648 7714 15700
rect 10410 15688 10416 15700
rect 7944 15660 10416 15688
rect 7944 15620 7972 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 11425 15691 11483 15697
rect 11425 15657 11437 15691
rect 11471 15688 11483 15691
rect 14182 15688 14188 15700
rect 11471 15660 14188 15688
rect 11471 15657 11483 15660
rect 11425 15651 11483 15657
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 18506 15688 18512 15700
rect 16776 15660 18512 15688
rect 7484 15592 7972 15620
rect 8018 15580 8024 15632
rect 8076 15620 8082 15632
rect 8076 15592 8248 15620
rect 8076 15580 8082 15592
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15552 5595 15555
rect 6089 15555 6147 15561
rect 6089 15552 6101 15555
rect 5583 15524 6101 15552
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 6089 15521 6101 15524
rect 6135 15521 6147 15555
rect 6270 15552 6276 15564
rect 6183 15524 6276 15552
rect 6089 15515 6147 15521
rect 6270 15512 6276 15524
rect 6328 15552 6334 15564
rect 8220 15561 8248 15592
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 13173 15623 13231 15629
rect 10008 15592 12848 15620
rect 10008 15580 10014 15592
rect 8205 15555 8263 15561
rect 6328 15524 8064 15552
rect 6328 15512 6334 15524
rect 8036 15493 8064 15524
rect 8205 15521 8217 15555
rect 8251 15521 8263 15555
rect 8570 15552 8576 15564
rect 8531 15524 8576 15552
rect 8205 15515 8263 15521
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15552 8815 15555
rect 10318 15552 10324 15564
rect 8803 15524 10324 15552
rect 8803 15521 8815 15524
rect 8757 15515 8815 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 10594 15552 10600 15564
rect 10555 15524 10600 15552
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 11572 15524 11621 15552
rect 11572 15512 11578 15524
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15552 12127 15555
rect 12618 15552 12624 15564
rect 12115 15524 12624 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 12820 15561 12848 15592
rect 13173 15589 13185 15623
rect 13219 15620 13231 15623
rect 13538 15620 13544 15632
rect 13219 15592 13544 15620
rect 13219 15589 13231 15592
rect 13173 15583 13231 15589
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 12805 15555 12863 15561
rect 12805 15521 12817 15555
rect 12851 15552 12863 15555
rect 14274 15552 14280 15564
rect 12851 15524 13400 15552
rect 14235 15524 14280 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15484 5319 15487
rect 5353 15487 5411 15493
rect 5353 15484 5365 15487
rect 5307 15456 5365 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 5353 15453 5365 15456
rect 5399 15453 5411 15487
rect 5353 15447 5411 15453
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 4801 15419 4859 15425
rect 4801 15385 4813 15419
rect 4847 15385 4859 15419
rect 4801 15379 4859 15385
rect 5368 15348 5396 15447
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11296 15456 11805 15484
rect 11296 15444 11302 15456
rect 11793 15453 11805 15456
rect 11839 15484 11851 15487
rect 11974 15484 11980 15496
rect 11839 15456 11980 15484
rect 11839 15453 11851 15456
rect 11793 15447 11851 15453
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 13372 15484 13400 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16776 15561 16804 15660
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 19886 15648 19892 15700
rect 19944 15688 19950 15700
rect 20993 15691 21051 15697
rect 20993 15688 21005 15691
rect 19944 15660 21005 15688
rect 19944 15648 19950 15660
rect 20993 15657 21005 15660
rect 21039 15657 21051 15691
rect 20993 15651 21051 15657
rect 28994 15648 29000 15700
rect 29052 15688 29058 15700
rect 29273 15691 29331 15697
rect 29273 15688 29285 15691
rect 29052 15660 29285 15688
rect 29052 15648 29058 15660
rect 29273 15657 29285 15660
rect 29319 15657 29331 15691
rect 33962 15688 33968 15700
rect 33923 15660 33968 15688
rect 29273 15651 29331 15657
rect 19337 15623 19395 15629
rect 19337 15589 19349 15623
rect 19383 15620 19395 15623
rect 20806 15620 20812 15632
rect 19383 15592 20812 15620
rect 19383 15589 19395 15592
rect 19337 15583 19395 15589
rect 20806 15580 20812 15592
rect 20864 15580 20870 15632
rect 29288 15620 29316 15651
rect 33962 15648 33968 15660
rect 34020 15648 34026 15700
rect 43990 15688 43996 15700
rect 43951 15660 43996 15688
rect 43990 15648 43996 15660
rect 44048 15648 44054 15700
rect 45462 15688 45468 15700
rect 45423 15660 45468 15688
rect 45462 15648 45468 15660
rect 45520 15648 45526 15700
rect 29288 15592 30420 15620
rect 16761 15555 16819 15561
rect 16761 15521 16773 15555
rect 16807 15521 16819 15555
rect 17034 15552 17040 15564
rect 16995 15524 17040 15552
rect 16761 15515 16819 15521
rect 17034 15512 17040 15524
rect 17092 15512 17098 15564
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15552 19579 15555
rect 19610 15552 19616 15564
rect 19567 15524 19616 15552
rect 19567 15521 19579 15524
rect 19521 15515 19579 15521
rect 19610 15512 19616 15524
rect 19668 15552 19674 15564
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 19668 15524 20913 15552
rect 19668 15512 19674 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 30392 15561 30420 15592
rect 31938 15580 31944 15632
rect 31996 15620 32002 15632
rect 32309 15623 32367 15629
rect 32309 15620 32321 15623
rect 31996 15592 32321 15620
rect 31996 15580 32002 15592
rect 32309 15589 32321 15592
rect 32355 15620 32367 15623
rect 32355 15592 33916 15620
rect 32355 15589 32367 15592
rect 32309 15583 32367 15589
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 23992 15524 24593 15552
rect 23992 15512 23998 15524
rect 24581 15521 24593 15524
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 30377 15555 30435 15561
rect 30377 15521 30389 15555
rect 30423 15521 30435 15555
rect 32490 15552 32496 15564
rect 32451 15524 32496 15552
rect 30377 15515 30435 15521
rect 32490 15512 32496 15524
rect 32548 15512 32554 15564
rect 32674 15512 32680 15564
rect 32732 15552 32738 15564
rect 33888 15561 33916 15592
rect 33689 15555 33747 15561
rect 33689 15552 33701 15555
rect 32732 15524 33701 15552
rect 32732 15512 32738 15524
rect 33689 15521 33701 15524
rect 33735 15521 33747 15555
rect 33689 15515 33747 15521
rect 33873 15555 33931 15561
rect 33873 15521 33885 15555
rect 33919 15521 33931 15555
rect 33980 15552 34008 15648
rect 38197 15623 38255 15629
rect 38197 15589 38209 15623
rect 38243 15620 38255 15623
rect 38378 15620 38384 15632
rect 38243 15592 38384 15620
rect 38243 15589 38255 15592
rect 38197 15583 38255 15589
rect 38378 15580 38384 15592
rect 38436 15580 38442 15632
rect 41782 15620 41788 15632
rect 40512 15592 41788 15620
rect 34974 15552 34980 15564
rect 33980 15524 34980 15552
rect 33873 15515 33931 15521
rect 34974 15512 34980 15524
rect 35032 15552 35038 15564
rect 35437 15555 35495 15561
rect 35437 15552 35449 15555
rect 35032 15524 35449 15552
rect 35032 15512 35038 15524
rect 35437 15521 35449 15524
rect 35483 15521 35495 15555
rect 35802 15552 35808 15564
rect 35763 15524 35808 15552
rect 35437 15515 35495 15521
rect 35802 15512 35808 15524
rect 35860 15512 35866 15564
rect 36173 15555 36231 15561
rect 36173 15521 36185 15555
rect 36219 15552 36231 15555
rect 36630 15552 36636 15564
rect 36219 15524 36636 15552
rect 36219 15521 36231 15524
rect 36173 15515 36231 15521
rect 36630 15512 36636 15524
rect 36688 15512 36694 15564
rect 39022 15552 39028 15564
rect 38983 15524 39028 15552
rect 39022 15512 39028 15524
rect 39080 15512 39086 15564
rect 39209 15555 39267 15561
rect 39209 15521 39221 15555
rect 39255 15552 39267 15555
rect 39390 15552 39396 15564
rect 39255 15524 39396 15552
rect 39255 15521 39267 15524
rect 39209 15515 39267 15521
rect 39390 15512 39396 15524
rect 39448 15512 39454 15564
rect 40313 15555 40371 15561
rect 40313 15521 40325 15555
rect 40359 15552 40371 15555
rect 40402 15552 40408 15564
rect 40359 15524 40408 15552
rect 40359 15521 40371 15524
rect 40313 15515 40371 15521
rect 40402 15512 40408 15524
rect 40460 15512 40466 15564
rect 40512 15561 40540 15592
rect 41782 15580 41788 15592
rect 41840 15580 41846 15632
rect 41877 15623 41935 15629
rect 41877 15589 41889 15623
rect 41923 15620 41935 15623
rect 42150 15620 42156 15632
rect 41923 15592 42156 15620
rect 41923 15589 41935 15592
rect 41877 15583 41935 15589
rect 42150 15580 42156 15592
rect 42208 15580 42214 15632
rect 48590 15580 48596 15632
rect 48648 15620 48654 15632
rect 51718 15620 51724 15632
rect 48648 15592 49280 15620
rect 51679 15592 51724 15620
rect 48648 15580 48654 15592
rect 40497 15555 40555 15561
rect 40497 15521 40509 15555
rect 40543 15521 40555 15555
rect 40497 15515 40555 15521
rect 40865 15555 40923 15561
rect 40865 15521 40877 15555
rect 40911 15552 40923 15555
rect 41969 15555 42027 15561
rect 41969 15552 41981 15555
rect 40911 15524 41981 15552
rect 40911 15521 40923 15524
rect 40865 15515 40923 15521
rect 41969 15521 41981 15524
rect 42015 15521 42027 15555
rect 41969 15515 42027 15521
rect 42429 15555 42487 15561
rect 42429 15521 42441 15555
rect 42475 15552 42487 15555
rect 44361 15555 44419 15561
rect 44361 15552 44373 15555
rect 42475 15524 44373 15552
rect 42475 15521 42487 15524
rect 42429 15515 42487 15521
rect 44361 15521 44373 15524
rect 44407 15521 44419 15555
rect 46750 15552 46756 15564
rect 46711 15524 46756 15552
rect 44361 15515 44419 15521
rect 46750 15512 46756 15524
rect 46808 15512 46814 15564
rect 46934 15552 46940 15564
rect 46895 15524 46940 15552
rect 46934 15512 46940 15524
rect 46992 15552 46998 15564
rect 47210 15552 47216 15564
rect 46992 15524 47216 15552
rect 46992 15512 46998 15524
rect 47210 15512 47216 15524
rect 47268 15512 47274 15564
rect 48958 15552 48964 15564
rect 48919 15524 48964 15552
rect 48958 15512 48964 15524
rect 49016 15512 49022 15564
rect 49050 15512 49056 15564
rect 49108 15552 49114 15564
rect 49252 15561 49280 15592
rect 51718 15580 51724 15592
rect 51776 15580 51782 15632
rect 49237 15555 49295 15561
rect 49108 15524 49153 15552
rect 49108 15512 49114 15524
rect 49237 15521 49249 15555
rect 49283 15521 49295 15555
rect 49237 15515 49295 15521
rect 50614 15512 50620 15564
rect 50672 15552 50678 15564
rect 51169 15555 51227 15561
rect 51169 15552 51181 15555
rect 50672 15524 51181 15552
rect 50672 15512 50678 15524
rect 51169 15521 51181 15524
rect 51215 15521 51227 15555
rect 51350 15552 51356 15564
rect 51311 15524 51356 15552
rect 51169 15515 51227 15521
rect 51350 15512 51356 15524
rect 51408 15552 51414 15564
rect 51813 15555 51871 15561
rect 51813 15552 51825 15555
rect 51408 15524 51825 15552
rect 51408 15512 51414 15524
rect 51813 15521 51825 15524
rect 51859 15521 51871 15555
rect 51813 15515 51871 15521
rect 18417 15487 18475 15493
rect 13372 15456 14228 15484
rect 6454 15416 6460 15428
rect 6415 15388 6460 15416
rect 6454 15376 6460 15388
rect 6512 15376 6518 15428
rect 12434 15376 12440 15428
rect 12492 15416 12498 15428
rect 14093 15419 14151 15425
rect 14093 15416 14105 15419
rect 12492 15388 14105 15416
rect 12492 15376 12498 15388
rect 14093 15385 14105 15388
rect 14139 15385 14151 15419
rect 14093 15379 14151 15385
rect 9766 15348 9772 15360
rect 5368 15320 9772 15348
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 10410 15348 10416 15360
rect 10371 15320 10416 15348
rect 10410 15308 10416 15320
rect 10468 15308 10474 15360
rect 13449 15351 13507 15357
rect 13449 15317 13461 15351
rect 13495 15348 13507 15351
rect 14200 15348 14228 15456
rect 18417 15453 18429 15487
rect 18463 15484 18475 15487
rect 19334 15484 19340 15496
rect 18463 15456 19340 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 21726 15444 21732 15496
rect 21784 15484 21790 15496
rect 21913 15487 21971 15493
rect 21913 15484 21925 15487
rect 21784 15456 21925 15484
rect 21784 15444 21790 15456
rect 21913 15453 21925 15456
rect 21959 15453 21971 15487
rect 22186 15484 22192 15496
rect 22147 15456 22192 15484
rect 21913 15447 21971 15453
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 27614 15444 27620 15496
rect 27672 15484 27678 15496
rect 27893 15487 27951 15493
rect 27893 15484 27905 15487
rect 27672 15456 27905 15484
rect 27672 15444 27678 15456
rect 27893 15453 27905 15456
rect 27939 15453 27951 15487
rect 27893 15447 27951 15453
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15484 28227 15487
rect 29362 15484 29368 15496
rect 28215 15456 29368 15484
rect 28215 15453 28227 15456
rect 28169 15447 28227 15453
rect 29362 15444 29368 15456
rect 29420 15444 29426 15496
rect 31202 15484 31208 15496
rect 29564 15456 31208 15484
rect 24762 15416 24768 15428
rect 17696 15388 21864 15416
rect 15381 15351 15439 15357
rect 15381 15348 15393 15351
rect 13495 15320 15393 15348
rect 13495 15317 13507 15320
rect 13449 15311 13507 15317
rect 15381 15317 15393 15320
rect 15427 15348 15439 15351
rect 17696 15348 17724 15388
rect 15427 15320 17724 15348
rect 19613 15351 19671 15357
rect 15427 15317 15439 15320
rect 15381 15311 15439 15317
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 19702 15348 19708 15360
rect 19659 15320 19708 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 21726 15348 21732 15360
rect 21687 15320 21732 15348
rect 21726 15308 21732 15320
rect 21784 15308 21790 15360
rect 21836 15348 21864 15388
rect 23308 15388 24768 15416
rect 23308 15348 23336 15388
rect 24762 15376 24768 15388
rect 24820 15376 24826 15428
rect 21836 15320 23336 15348
rect 23382 15308 23388 15360
rect 23440 15348 23446 15360
rect 23477 15351 23535 15357
rect 23477 15348 23489 15351
rect 23440 15320 23489 15348
rect 23440 15308 23446 15320
rect 23477 15317 23489 15320
rect 23523 15317 23535 15351
rect 23477 15311 23535 15317
rect 23934 15308 23940 15360
rect 23992 15348 23998 15360
rect 24213 15351 24271 15357
rect 24213 15348 24225 15351
rect 23992 15320 24225 15348
rect 23992 15308 23998 15320
rect 24213 15317 24225 15320
rect 24259 15317 24271 15351
rect 24213 15311 24271 15317
rect 24397 15351 24455 15357
rect 24397 15317 24409 15351
rect 24443 15348 24455 15351
rect 29564 15348 29592 15456
rect 31202 15444 31208 15456
rect 31260 15444 31266 15496
rect 32861 15487 32919 15493
rect 32861 15453 32873 15487
rect 32907 15484 32919 15487
rect 34422 15484 34428 15496
rect 32907 15456 34428 15484
rect 32907 15453 32919 15456
rect 32861 15447 32919 15453
rect 34422 15444 34428 15456
rect 34480 15444 34486 15496
rect 38746 15484 38752 15496
rect 38707 15456 38752 15484
rect 38746 15444 38752 15456
rect 38804 15444 38810 15496
rect 43990 15444 43996 15496
rect 44048 15484 44054 15496
rect 44085 15487 44143 15493
rect 44085 15484 44097 15487
rect 44048 15456 44097 15484
rect 44048 15444 44054 15456
rect 44085 15453 44097 15456
rect 44131 15453 44143 15487
rect 49602 15484 49608 15496
rect 49563 15456 49608 15484
rect 44085 15447 44143 15453
rect 49602 15444 49608 15456
rect 49660 15444 49666 15496
rect 29730 15376 29736 15428
rect 29788 15416 29794 15428
rect 40310 15416 40316 15428
rect 29788 15388 40316 15416
rect 29788 15376 29794 15388
rect 40310 15376 40316 15388
rect 40368 15376 40374 15428
rect 24443 15320 29592 15348
rect 29641 15351 29699 15357
rect 24443 15317 24455 15320
rect 24397 15311 24455 15317
rect 29641 15317 29653 15351
rect 29687 15348 29699 15351
rect 30098 15348 30104 15360
rect 29687 15320 30104 15348
rect 29687 15317 29699 15320
rect 29641 15311 29699 15317
rect 30098 15308 30104 15320
rect 30156 15308 30162 15360
rect 30469 15351 30527 15357
rect 30469 15317 30481 15351
rect 30515 15348 30527 15351
rect 31110 15348 31116 15360
rect 30515 15320 31116 15348
rect 30515 15317 30527 15320
rect 30469 15311 30527 15317
rect 31110 15308 31116 15320
rect 31168 15308 31174 15360
rect 41690 15348 41696 15360
rect 41651 15320 41696 15348
rect 41690 15308 41696 15320
rect 41748 15308 41754 15360
rect 47026 15348 47032 15360
rect 46987 15320 47032 15348
rect 47026 15308 47032 15320
rect 47084 15308 47090 15360
rect 1104 15258 54832 15280
rect 1104 15206 9947 15258
rect 9999 15206 10011 15258
rect 10063 15206 10075 15258
rect 10127 15206 10139 15258
rect 10191 15206 27878 15258
rect 27930 15206 27942 15258
rect 27994 15206 28006 15258
rect 28058 15206 28070 15258
rect 28122 15206 45808 15258
rect 45860 15206 45872 15258
rect 45924 15206 45936 15258
rect 45988 15206 46000 15258
rect 46052 15206 54832 15258
rect 1104 15184 54832 15206
rect 11238 15144 11244 15156
rect 7208 15116 11244 15144
rect 2133 15079 2191 15085
rect 2133 15045 2145 15079
rect 2179 15076 2191 15079
rect 2179 15048 3280 15076
rect 2179 15045 2191 15048
rect 2133 15039 2191 15045
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 3252 14949 3280 15048
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 15008 3755 15011
rect 4062 15008 4068 15020
rect 3743 14980 4068 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 6362 14968 6368 15020
rect 6420 15008 6426 15020
rect 6420 14980 7052 15008
rect 6420 14968 6426 14980
rect 2317 14943 2375 14949
rect 2317 14940 2329 14943
rect 2280 14912 2329 14940
rect 2280 14900 2286 14912
rect 2317 14909 2329 14912
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14909 3295 14943
rect 3878 14940 3884 14952
rect 3839 14912 3884 14940
rect 3237 14903 3295 14909
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 4154 14940 4160 14952
rect 4115 14912 4160 14940
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 4430 14940 4436 14952
rect 4391 14912 4436 14940
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 5629 14943 5687 14949
rect 5629 14909 5641 14943
rect 5675 14940 5687 14943
rect 6546 14940 6552 14952
rect 5675 14912 6552 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 7024 14949 7052 14980
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6687 14912 6837 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 6840 14872 6868 14903
rect 7208 14872 7236 15116
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 11333 15147 11391 15153
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 11379 15116 13308 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 12342 15076 12348 15088
rect 9140 15048 12348 15076
rect 9140 15017 9168 15048
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 13170 15076 13176 15088
rect 12676 15048 13176 15076
rect 12676 15036 12682 15048
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 13280 15076 13308 15116
rect 14274 15104 14280 15156
rect 14332 15144 14338 15156
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 14332 15116 14657 15144
rect 14332 15104 14338 15116
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 20806 15104 20812 15156
rect 20864 15144 20870 15156
rect 22465 15147 22523 15153
rect 22465 15144 22477 15147
rect 20864 15116 22477 15144
rect 20864 15104 20870 15116
rect 22465 15113 22477 15116
rect 22511 15113 22523 15147
rect 22465 15107 22523 15113
rect 24026 15104 24032 15156
rect 24084 15144 24090 15156
rect 27522 15144 27528 15156
rect 24084 15116 27528 15144
rect 24084 15104 24090 15116
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 32582 15104 32588 15156
rect 32640 15144 32646 15156
rect 33321 15147 33379 15153
rect 33321 15144 33333 15147
rect 32640 15116 33333 15144
rect 32640 15104 32646 15116
rect 33321 15113 33333 15116
rect 33367 15113 33379 15147
rect 33321 15107 33379 15113
rect 17954 15076 17960 15088
rect 13280 15048 17960 15076
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 18506 15036 18512 15088
rect 18564 15076 18570 15088
rect 20714 15076 20720 15088
rect 18564 15048 20720 15076
rect 18564 15036 18570 15048
rect 20714 15036 20720 15048
rect 20772 15076 20778 15088
rect 21726 15076 21732 15088
rect 20772 15048 21732 15076
rect 20772 15036 20778 15048
rect 21726 15036 21732 15048
rect 21784 15076 21790 15088
rect 24673 15079 24731 15085
rect 24673 15076 24685 15079
rect 21784 15048 24685 15076
rect 21784 15036 21790 15048
rect 24673 15045 24685 15048
rect 24719 15076 24731 15079
rect 24719 15048 24900 15076
rect 24719 15045 24731 15048
rect 24673 15039 24731 15045
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 15008 8999 15011
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 8987 14980 9137 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 9125 14977 9137 14980
rect 9171 14977 9183 15011
rect 9125 14971 9183 14977
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 15008 12311 15011
rect 12526 15008 12532 15020
rect 12299 14980 12532 15008
rect 12299 14977 12311 14980
rect 12253 14971 12311 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 13630 15008 13636 15020
rect 13591 14980 13636 15008
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 18230 15008 18236 15020
rect 14752 14980 18236 15008
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 6840 14844 7236 14872
rect 7484 14872 7512 14903
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 7616 14912 9229 14940
rect 7616 14900 7622 14912
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9674 14940 9680 14952
rect 9635 14912 9680 14940
rect 9217 14903 9275 14909
rect 8294 14872 8300 14884
rect 7484 14844 8300 14872
rect 8294 14832 8300 14844
rect 8352 14872 8358 14884
rect 9030 14872 9036 14884
rect 8352 14844 9036 14872
rect 8352 14832 8358 14844
rect 9030 14832 9036 14844
rect 9088 14832 9094 14884
rect 9232 14872 9260 14903
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 11146 14940 11152 14952
rect 9815 14912 11152 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 9784 14872 9812 14903
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 11517 14943 11575 14949
rect 11517 14909 11529 14943
rect 11563 14940 11575 14943
rect 12342 14940 12348 14952
rect 11563 14912 12348 14940
rect 11563 14909 11575 14912
rect 11517 14903 11575 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12618 14940 12624 14952
rect 12579 14912 12624 14940
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 13078 14940 13084 14952
rect 13039 14912 13084 14940
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13228 14912 13273 14940
rect 13228 14900 13234 14912
rect 10318 14872 10324 14884
rect 9232 14844 9812 14872
rect 10279 14844 10324 14872
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 12802 14832 12808 14884
rect 12860 14872 12866 14884
rect 14752 14872 14780 14980
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 24872 15017 24900 15048
rect 25866 15036 25872 15088
rect 25924 15076 25930 15088
rect 33226 15076 33232 15088
rect 25924 15048 33232 15076
rect 25924 15036 25930 15048
rect 33226 15036 33232 15048
rect 33284 15036 33290 15088
rect 24857 15011 24915 15017
rect 19392 14980 24716 15008
rect 19392 14968 19398 14980
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14909 14887 14943
rect 15838 14940 15844 14952
rect 15799 14912 15844 14940
rect 14829 14903 14887 14909
rect 12860 14844 14780 14872
rect 14844 14872 14872 14903
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 18782 14940 18788 14952
rect 16899 14912 18788 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14940 19763 14943
rect 19886 14940 19892 14952
rect 19751 14912 19892 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 16482 14872 16488 14884
rect 14844 14844 16488 14872
rect 12860 14832 12866 14844
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 18984 14872 19012 14903
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 20806 14900 20812 14952
rect 20864 14940 20870 14952
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20864 14912 20913 14940
rect 20864 14900 20870 14912
rect 20901 14909 20913 14912
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 22189 14943 22247 14949
rect 22189 14909 22201 14943
rect 22235 14909 22247 14943
rect 22189 14903 22247 14909
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14940 22339 14943
rect 23382 14940 23388 14952
rect 22327 14912 23388 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 18380 14844 19012 14872
rect 19521 14875 19579 14881
rect 18380 14832 18386 14844
rect 19521 14841 19533 14875
rect 19567 14872 19579 14875
rect 20993 14875 21051 14881
rect 20993 14872 21005 14875
rect 19567 14844 21005 14872
rect 19567 14841 19579 14844
rect 19521 14835 19579 14841
rect 20993 14841 21005 14844
rect 21039 14872 21051 14875
rect 22002 14872 22008 14884
rect 21039 14844 22008 14872
rect 21039 14841 21051 14844
rect 20993 14835 21051 14841
rect 22002 14832 22008 14844
rect 22060 14832 22066 14884
rect 22204 14872 22232 14903
rect 23382 14900 23388 14912
rect 23440 14900 23446 14952
rect 24581 14943 24639 14949
rect 24581 14909 24593 14943
rect 24627 14909 24639 14943
rect 24688 14940 24716 14980
rect 24857 14977 24869 15011
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 27430 14968 27436 15020
rect 27488 15008 27494 15020
rect 27617 15011 27675 15017
rect 27617 15008 27629 15011
rect 27488 14980 27629 15008
rect 27488 14968 27494 14980
rect 27617 14977 27629 14980
rect 27663 15008 27675 15011
rect 28902 15008 28908 15020
rect 27663 14980 28908 15008
rect 27663 14977 27675 14980
rect 27617 14971 27675 14977
rect 28902 14968 28908 14980
rect 28960 14968 28966 15020
rect 32490 15008 32496 15020
rect 31128 14980 32496 15008
rect 31128 14952 31156 14980
rect 24946 14940 24952 14952
rect 24688 14912 24952 14940
rect 24581 14903 24639 14909
rect 22204 14844 22968 14872
rect 22940 14816 22968 14844
rect 3418 14764 3424 14816
rect 3476 14804 3482 14816
rect 5445 14807 5503 14813
rect 5445 14804 5457 14807
rect 3476 14776 5457 14804
rect 3476 14764 3482 14776
rect 5445 14773 5457 14776
rect 5491 14773 5503 14807
rect 5445 14767 5503 14773
rect 7190 14764 7196 14816
rect 7248 14804 7254 14816
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7248 14776 8033 14804
rect 7248 14764 7254 14776
rect 8021 14773 8033 14776
rect 8067 14773 8079 14807
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 8021 14767 8079 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 16666 14804 16672 14816
rect 16627 14776 16672 14804
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 18506 14764 18512 14816
rect 18564 14804 18570 14816
rect 18785 14807 18843 14813
rect 18785 14804 18797 14807
rect 18564 14776 18797 14804
rect 18564 14764 18570 14776
rect 18785 14773 18797 14776
rect 18831 14773 18843 14807
rect 18785 14767 18843 14773
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19484 14776 19809 14804
rect 19484 14764 19490 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 22922 14804 22928 14816
rect 22883 14776 22928 14804
rect 19797 14767 19855 14773
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 24394 14804 24400 14816
rect 24355 14776 24400 14804
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 24596 14804 24624 14903
rect 24946 14900 24952 14912
rect 25004 14900 25010 14952
rect 25130 14940 25136 14952
rect 25091 14912 25136 14940
rect 25130 14900 25136 14912
rect 25188 14900 25194 14952
rect 26602 14900 26608 14952
rect 26660 14940 26666 14952
rect 27522 14940 27528 14952
rect 26660 14912 27528 14940
rect 26660 14900 26666 14912
rect 27522 14900 27528 14912
rect 27580 14900 27586 14952
rect 30742 14940 30748 14952
rect 30703 14912 30748 14940
rect 30742 14900 30748 14912
rect 30800 14900 30806 14952
rect 30837 14943 30895 14949
rect 30837 14909 30849 14943
rect 30883 14909 30895 14943
rect 31110 14940 31116 14952
rect 31071 14912 31116 14940
rect 30837 14903 30895 14909
rect 26344 14844 29224 14872
rect 26344 14804 26372 14844
rect 24596 14776 26372 14804
rect 26421 14807 26479 14813
rect 26421 14773 26433 14807
rect 26467 14804 26479 14807
rect 26510 14804 26516 14816
rect 26467 14776 26516 14804
rect 26467 14773 26479 14776
rect 26421 14767 26479 14773
rect 26510 14764 26516 14776
rect 26568 14764 26574 14816
rect 29196 14804 29224 14844
rect 29270 14832 29276 14884
rect 29328 14872 29334 14884
rect 30101 14875 30159 14881
rect 30101 14872 30113 14875
rect 29328 14844 30113 14872
rect 29328 14832 29334 14844
rect 30101 14841 30113 14844
rect 30147 14841 30159 14875
rect 30852 14872 30880 14903
rect 31110 14900 31116 14912
rect 31168 14900 31174 14952
rect 32324 14949 32352 14980
rect 32490 14968 32496 14980
rect 32548 14968 32554 15020
rect 32674 15008 32680 15020
rect 32635 14980 32680 15008
rect 32674 14968 32680 14980
rect 32732 14968 32738 15020
rect 31297 14943 31355 14949
rect 31297 14909 31309 14943
rect 31343 14940 31355 14943
rect 32125 14943 32183 14949
rect 32125 14940 32137 14943
rect 31343 14912 32137 14940
rect 31343 14909 31355 14912
rect 31297 14903 31355 14909
rect 32125 14909 32137 14912
rect 32171 14909 32183 14943
rect 32125 14903 32183 14909
rect 32309 14943 32367 14949
rect 32309 14909 32321 14943
rect 32355 14909 32367 14943
rect 33336 14940 33364 15107
rect 34422 15104 34428 15156
rect 34480 15144 34486 15156
rect 36495 15147 36553 15153
rect 36495 15144 36507 15147
rect 34480 15116 36507 15144
rect 34480 15104 34486 15116
rect 36495 15113 36507 15116
rect 36541 15113 36553 15147
rect 36495 15107 36553 15113
rect 36633 15147 36691 15153
rect 36633 15113 36645 15147
rect 36679 15144 36691 15147
rect 39390 15144 39396 15156
rect 36679 15116 39396 15144
rect 36679 15113 36691 15116
rect 36633 15107 36691 15113
rect 39390 15104 39396 15116
rect 39448 15104 39454 15156
rect 46934 15144 46940 15156
rect 42076 15116 46940 15144
rect 38565 15079 38623 15085
rect 35176 15048 35756 15076
rect 33505 14943 33563 14949
rect 33505 14940 33517 14943
rect 33336 14912 33517 14940
rect 32309 14903 32367 14909
rect 33505 14909 33517 14912
rect 33551 14909 33563 14943
rect 34974 14940 34980 14952
rect 34935 14912 34980 14940
rect 33505 14903 33563 14909
rect 32140 14872 32168 14903
rect 34974 14900 34980 14912
rect 35032 14900 35038 14952
rect 35176 14949 35204 15048
rect 35529 15011 35587 15017
rect 35529 14977 35541 15011
rect 35575 15008 35587 15011
rect 35618 15008 35624 15020
rect 35575 14980 35624 15008
rect 35575 14977 35587 14980
rect 35529 14971 35587 14977
rect 35618 14968 35624 14980
rect 35676 14968 35682 15020
rect 35728 15008 35756 15048
rect 38565 15045 38577 15079
rect 38611 15076 38623 15079
rect 38746 15076 38752 15088
rect 38611 15048 38752 15076
rect 38611 15045 38623 15048
rect 38565 15039 38623 15045
rect 38746 15036 38752 15048
rect 38804 15036 38810 15088
rect 36722 15008 36728 15020
rect 35728 14980 36728 15008
rect 36722 14968 36728 14980
rect 36780 14968 36786 15020
rect 39022 15008 39028 15020
rect 38212 14980 39028 15008
rect 35161 14943 35219 14949
rect 35161 14909 35173 14943
rect 35207 14909 35219 14943
rect 35636 14940 35664 14968
rect 38212 14940 38240 14980
rect 39022 14968 39028 14980
rect 39080 15008 39086 15020
rect 39117 15011 39175 15017
rect 39117 15008 39129 15011
rect 39080 14980 39129 15008
rect 39080 14968 39086 14980
rect 39117 14977 39129 14980
rect 39163 14977 39175 15011
rect 39117 14971 39175 14977
rect 41506 14968 41512 15020
rect 41564 15008 41570 15020
rect 42076 15017 42104 15116
rect 46934 15104 46940 15116
rect 46992 15104 46998 15156
rect 47026 15104 47032 15156
rect 47084 15153 47090 15156
rect 47084 15147 47133 15153
rect 47084 15113 47087 15147
rect 47121 15113 47133 15147
rect 47084 15107 47133 15113
rect 47581 15147 47639 15153
rect 47581 15113 47593 15147
rect 47627 15144 47639 15147
rect 48314 15144 48320 15156
rect 47627 15116 48320 15144
rect 47627 15113 47639 15116
rect 47581 15107 47639 15113
rect 47084 15104 47090 15107
rect 48314 15104 48320 15116
rect 48372 15104 48378 15156
rect 50614 15144 50620 15156
rect 50575 15116 50620 15144
rect 50614 15104 50620 15116
rect 50672 15104 50678 15156
rect 51442 15104 51448 15156
rect 51500 15144 51506 15156
rect 51721 15147 51779 15153
rect 51721 15144 51733 15147
rect 51500 15116 51733 15144
rect 51500 15104 51506 15116
rect 51721 15113 51733 15116
rect 51767 15113 51779 15147
rect 51721 15107 51779 15113
rect 44174 15036 44180 15088
rect 44232 15076 44238 15088
rect 47213 15079 47271 15085
rect 47213 15076 47225 15079
rect 44232 15048 47225 15076
rect 44232 15036 44238 15048
rect 47213 15045 47225 15048
rect 47259 15045 47271 15079
rect 47213 15039 47271 15045
rect 42061 15011 42119 15017
rect 42061 15008 42073 15011
rect 41564 14980 42073 15008
rect 41564 14968 41570 14980
rect 42061 14977 42073 14980
rect 42107 14977 42119 15011
rect 43530 15008 43536 15020
rect 42061 14971 42119 14977
rect 42536 14980 43536 15008
rect 42536 14952 42564 14980
rect 43530 14968 43536 14980
rect 43588 15008 43594 15020
rect 43809 15011 43867 15017
rect 43809 15008 43821 15011
rect 43588 14980 43821 15008
rect 43588 14968 43594 14980
rect 43809 14977 43821 14980
rect 43855 14977 43867 15011
rect 45278 15008 45284 15020
rect 43809 14971 43867 14977
rect 45020 14980 45284 15008
rect 35636 14912 38240 14940
rect 38473 14943 38531 14949
rect 35161 14903 35219 14909
rect 38473 14909 38485 14943
rect 38519 14909 38531 14943
rect 38473 14903 38531 14909
rect 38933 14943 38991 14949
rect 38933 14909 38945 14943
rect 38979 14940 38991 14943
rect 39390 14940 39396 14952
rect 38979 14912 39396 14940
rect 38979 14909 38991 14912
rect 38933 14903 38991 14909
rect 35710 14872 35716 14884
rect 30852 14844 31524 14872
rect 32140 14844 35716 14872
rect 30101 14835 30159 14841
rect 31496 14816 31524 14844
rect 35710 14832 35716 14844
rect 35768 14872 35774 14884
rect 36357 14875 36415 14881
rect 36357 14872 36369 14875
rect 35768 14844 36369 14872
rect 35768 14832 35774 14844
rect 36357 14841 36369 14844
rect 36403 14841 36415 14875
rect 38488 14872 38516 14903
rect 39390 14900 39396 14912
rect 39448 14900 39454 14952
rect 40494 14940 40500 14952
rect 40455 14912 40500 14940
rect 40494 14900 40500 14912
rect 40552 14900 40558 14952
rect 40589 14943 40647 14949
rect 40589 14909 40601 14943
rect 40635 14940 40647 14943
rect 41874 14940 41880 14952
rect 40635 14912 41880 14940
rect 40635 14909 40647 14912
rect 40589 14903 40647 14909
rect 41874 14900 41880 14912
rect 41932 14940 41938 14952
rect 42153 14943 42211 14949
rect 42153 14940 42165 14943
rect 41932 14912 42165 14940
rect 41932 14900 41938 14912
rect 42153 14909 42165 14912
rect 42199 14909 42211 14943
rect 42518 14940 42524 14952
rect 42479 14912 42524 14940
rect 42153 14903 42211 14909
rect 42518 14900 42524 14912
rect 42576 14900 42582 14952
rect 42705 14943 42763 14949
rect 42705 14909 42717 14943
rect 42751 14940 42763 14943
rect 42794 14940 42800 14952
rect 42751 14912 42800 14940
rect 42751 14909 42763 14912
rect 42705 14903 42763 14909
rect 42794 14900 42800 14912
rect 42852 14900 42858 14952
rect 43714 14940 43720 14952
rect 43675 14912 43720 14940
rect 43714 14900 43720 14912
rect 43772 14900 43778 14952
rect 44358 14900 44364 14952
rect 44416 14940 44422 14952
rect 45020 14949 45048 14980
rect 45278 14968 45284 14980
rect 45336 14968 45342 15020
rect 45646 14968 45652 15020
rect 45704 15008 45710 15020
rect 47305 15011 47363 15017
rect 47305 15008 47317 15011
rect 45704 14980 47317 15008
rect 45704 14968 45710 14980
rect 47305 14977 47317 14980
rect 47351 14977 47363 15011
rect 55582 15008 55588 15020
rect 47305 14971 47363 14977
rect 47412 14980 55588 15008
rect 45005 14943 45063 14949
rect 45005 14940 45017 14943
rect 44416 14912 45017 14940
rect 44416 14900 44422 14912
rect 45005 14909 45017 14912
rect 45051 14909 45063 14943
rect 45005 14903 45063 14909
rect 45186 14900 45192 14952
rect 45244 14940 45250 14952
rect 47412 14940 47440 14980
rect 55582 14968 55588 14980
rect 55640 14968 55646 15020
rect 45244 14912 47440 14940
rect 45244 14900 45250 14912
rect 47578 14900 47584 14952
rect 47636 14940 47642 14952
rect 49237 14943 49295 14949
rect 49237 14940 49249 14943
rect 47636 14912 49249 14940
rect 47636 14900 47642 14912
rect 49237 14909 49249 14912
rect 49283 14909 49295 14943
rect 49237 14903 49295 14909
rect 50154 14900 50160 14952
rect 50212 14940 50218 14952
rect 50525 14943 50583 14949
rect 50525 14940 50537 14943
rect 50212 14912 50537 14940
rect 50212 14900 50218 14912
rect 50525 14909 50537 14912
rect 50571 14909 50583 14943
rect 51994 14940 52000 14952
rect 51955 14912 52000 14940
rect 50525 14903 50583 14909
rect 51994 14900 52000 14912
rect 52052 14900 52058 14952
rect 38488 14844 39620 14872
rect 36357 14835 36415 14841
rect 30006 14804 30012 14816
rect 29196 14776 30012 14804
rect 30006 14764 30012 14776
rect 30064 14764 30070 14816
rect 31478 14804 31484 14816
rect 31439 14776 31484 14804
rect 31478 14764 31484 14776
rect 31536 14764 31542 14816
rect 33597 14807 33655 14813
rect 33597 14773 33609 14807
rect 33643 14804 33655 14807
rect 34054 14804 34060 14816
rect 33643 14776 34060 14804
rect 33643 14773 33655 14776
rect 33597 14767 33655 14773
rect 34054 14764 34060 14776
rect 34112 14764 34118 14816
rect 37001 14807 37059 14813
rect 37001 14773 37013 14807
rect 37047 14804 37059 14807
rect 39390 14804 39396 14816
rect 37047 14776 39396 14804
rect 37047 14773 37059 14776
rect 37001 14767 37059 14773
rect 39390 14764 39396 14776
rect 39448 14764 39454 14816
rect 39592 14813 39620 14844
rect 40126 14832 40132 14884
rect 40184 14872 40190 14884
rect 41509 14875 41567 14881
rect 41509 14872 41521 14875
rect 40184 14844 41521 14872
rect 40184 14832 40190 14844
rect 41509 14841 41521 14844
rect 41555 14841 41567 14875
rect 41509 14835 41567 14841
rect 45097 14875 45155 14881
rect 45097 14841 45109 14875
rect 45143 14872 45155 14875
rect 45830 14872 45836 14884
rect 45143 14844 45836 14872
rect 45143 14841 45155 14844
rect 45097 14835 45155 14841
rect 45830 14832 45836 14844
rect 45888 14832 45894 14884
rect 46934 14872 46940 14884
rect 46895 14844 46940 14872
rect 46934 14832 46940 14844
rect 46992 14832 46998 14884
rect 51905 14875 51963 14881
rect 51905 14872 51917 14875
rect 47044 14844 51917 14872
rect 39577 14807 39635 14813
rect 39577 14773 39589 14807
rect 39623 14804 39635 14807
rect 39666 14804 39672 14816
rect 39623 14776 39672 14804
rect 39623 14773 39635 14776
rect 39577 14767 39635 14773
rect 39666 14764 39672 14776
rect 39724 14764 39730 14816
rect 46198 14764 46204 14816
rect 46256 14804 46262 14816
rect 47044 14804 47072 14844
rect 51905 14841 51917 14844
rect 51951 14841 51963 14875
rect 51905 14835 51963 14841
rect 52270 14832 52276 14884
rect 52328 14872 52334 14884
rect 52457 14875 52515 14881
rect 52457 14872 52469 14875
rect 52328 14844 52469 14872
rect 52328 14832 52334 14844
rect 52457 14841 52469 14844
rect 52503 14841 52515 14875
rect 52457 14835 52515 14841
rect 46256 14776 47072 14804
rect 49329 14807 49387 14813
rect 46256 14764 46262 14776
rect 49329 14773 49341 14807
rect 49375 14804 49387 14807
rect 49694 14804 49700 14816
rect 49375 14776 49700 14804
rect 49375 14773 49387 14776
rect 49329 14767 49387 14773
rect 49694 14764 49700 14776
rect 49752 14764 49758 14816
rect 1104 14714 54832 14736
rect 1104 14662 18912 14714
rect 18964 14662 18976 14714
rect 19028 14662 19040 14714
rect 19092 14662 19104 14714
rect 19156 14662 36843 14714
rect 36895 14662 36907 14714
rect 36959 14662 36971 14714
rect 37023 14662 37035 14714
rect 37087 14662 54832 14714
rect 1104 14640 54832 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14569 3295 14603
rect 5813 14603 5871 14609
rect 5813 14600 5825 14603
rect 3237 14563 3295 14569
rect 4080 14572 5825 14600
rect 3252 14532 3280 14563
rect 2424 14504 3280 14532
rect 2424 14473 2452 14504
rect 2409 14467 2467 14473
rect 2409 14433 2421 14467
rect 2455 14433 2467 14467
rect 3418 14464 3424 14476
rect 3379 14436 3424 14464
rect 2409 14427 2467 14433
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4080 14473 4108 14572
rect 5813 14569 5825 14572
rect 5859 14569 5871 14603
rect 6546 14600 6552 14612
rect 6507 14572 6552 14600
rect 5813 14563 5871 14569
rect 5828 14532 5856 14563
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 12802 14600 12808 14612
rect 12763 14572 12808 14600
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13814 14600 13820 14612
rect 13775 14572 13820 14600
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 15378 14600 15384 14612
rect 15339 14572 15384 14600
rect 15378 14560 15384 14572
rect 15436 14600 15442 14612
rect 15746 14600 15752 14612
rect 15436 14572 15752 14600
rect 15436 14560 15442 14572
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 24026 14600 24032 14612
rect 17000 14572 24032 14600
rect 17000 14560 17006 14572
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 24121 14603 24179 14609
rect 24121 14569 24133 14603
rect 24167 14600 24179 14603
rect 25866 14600 25872 14612
rect 24167 14572 25872 14600
rect 24167 14569 24179 14572
rect 24121 14563 24179 14569
rect 6914 14532 6920 14544
rect 5828 14504 6920 14532
rect 6914 14492 6920 14504
rect 6972 14532 6978 14544
rect 8386 14532 8392 14544
rect 6972 14504 8392 14532
rect 6972 14492 6978 14504
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 10505 14535 10563 14541
rect 10505 14501 10517 14535
rect 10551 14532 10563 14535
rect 13722 14532 13728 14544
rect 10551 14504 13728 14532
rect 10551 14501 10563 14504
rect 10505 14495 10563 14501
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 4028 14436 4077 14464
rect 4028 14424 4034 14436
rect 4065 14433 4077 14436
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14464 4399 14467
rect 6454 14464 6460 14476
rect 4387 14436 6460 14464
rect 4387 14433 4399 14436
rect 4341 14427 4399 14433
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 6748 14396 6776 14427
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7340 14436 7757 14464
rect 7340 14424 7346 14436
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 8757 14467 8815 14473
rect 8757 14433 8769 14467
rect 8803 14464 8815 14467
rect 10410 14464 10416 14476
rect 8803 14436 10416 14464
rect 8803 14433 8815 14436
rect 8757 14427 8815 14433
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 10888 14473 10916 14504
rect 13722 14492 13728 14504
rect 13780 14492 13786 14544
rect 18414 14532 18420 14544
rect 18375 14504 18420 14532
rect 18414 14492 18420 14504
rect 18472 14492 18478 14544
rect 20073 14535 20131 14541
rect 20073 14532 20085 14535
rect 19352 14504 20085 14532
rect 10781 14467 10839 14473
rect 10781 14433 10793 14467
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 10873 14467 10931 14473
rect 10873 14433 10885 14467
rect 10919 14433 10931 14467
rect 11146 14464 11152 14476
rect 10873 14427 10931 14433
rect 10980 14436 11152 14464
rect 4580 14368 6776 14396
rect 10796 14396 10824 14427
rect 10980 14396 11008 14436
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 11517 14467 11575 14473
rect 11388 14436 11433 14464
rect 11388 14424 11394 14436
rect 11517 14433 11529 14467
rect 11563 14464 11575 14467
rect 11698 14464 11704 14476
rect 11563 14436 11704 14464
rect 11563 14433 11575 14436
rect 11517 14427 11575 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 12768 14436 13001 14464
rect 12768 14424 12774 14436
rect 12989 14433 13001 14436
rect 13035 14433 13047 14467
rect 12989 14427 13047 14433
rect 14001 14467 14059 14473
rect 14001 14433 14013 14467
rect 14047 14433 14059 14467
rect 14001 14427 14059 14433
rect 10796 14368 11008 14396
rect 14016 14396 14044 14427
rect 14826 14424 14832 14476
rect 14884 14464 14890 14476
rect 19352 14473 19380 14504
rect 20073 14501 20085 14504
rect 20119 14532 20131 14535
rect 20806 14532 20812 14544
rect 20119 14504 20812 14532
rect 20119 14501 20131 14504
rect 20073 14495 20131 14501
rect 20806 14492 20812 14504
rect 20864 14532 20870 14544
rect 22002 14532 22008 14544
rect 20864 14504 21864 14532
rect 21963 14504 22008 14532
rect 20864 14492 20870 14504
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 14884 14436 15301 14464
rect 14884 14424 14890 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 19337 14467 19395 14473
rect 19337 14433 19349 14467
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19562 14467 19620 14473
rect 19484 14436 19529 14464
rect 19484 14424 19490 14436
rect 19562 14433 19574 14467
rect 19608 14464 19620 14467
rect 19702 14464 19708 14476
rect 19608 14436 19708 14464
rect 19608 14433 19620 14436
rect 19562 14427 19620 14433
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 21836 14473 21864 14504
rect 22002 14492 22008 14504
rect 22060 14492 22066 14544
rect 23382 14532 23388 14544
rect 23343 14504 23388 14532
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 21821 14467 21879 14473
rect 21821 14433 21833 14467
rect 21867 14433 21879 14467
rect 21821 14427 21879 14433
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14433 22155 14467
rect 22097 14427 22155 14433
rect 16022 14396 16028 14408
rect 14016 14368 16028 14396
rect 4580 14356 4586 14368
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14396 16911 14399
rect 19981 14399 20039 14405
rect 19981 14396 19993 14399
rect 16899 14368 19993 14396
rect 16899 14365 16911 14368
rect 16853 14359 16911 14365
rect 19981 14365 19993 14368
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 8573 14331 8631 14337
rect 8573 14297 8585 14331
rect 8619 14328 8631 14331
rect 8619 14300 12940 14328
rect 8619 14297 8631 14300
rect 8573 14291 8631 14297
rect 5442 14260 5448 14272
rect 5403 14232 5448 14260
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 6638 14220 6644 14272
rect 6696 14260 6702 14272
rect 7561 14263 7619 14269
rect 7561 14260 7573 14263
rect 6696 14232 7573 14260
rect 6696 14220 6702 14232
rect 7561 14229 7573 14232
rect 7607 14229 7619 14263
rect 7561 14223 7619 14229
rect 11793 14263 11851 14269
rect 11793 14229 11805 14263
rect 11839 14260 11851 14263
rect 12434 14260 12440 14272
rect 11839 14232 12440 14260
rect 11839 14229 11851 14232
rect 11793 14223 11851 14229
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 12912 14260 12940 14300
rect 12986 14288 12992 14340
rect 13044 14328 13050 14340
rect 15194 14328 15200 14340
rect 13044 14300 15200 14328
rect 13044 14288 13050 14300
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15378 14260 15384 14272
rect 12912 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 16592 14260 16620 14359
rect 18141 14331 18199 14337
rect 18141 14297 18153 14331
rect 18187 14328 18199 14331
rect 19610 14328 19616 14340
rect 18187 14300 19616 14328
rect 18187 14297 18199 14300
rect 18141 14291 18199 14297
rect 19610 14288 19616 14300
rect 19668 14288 19674 14340
rect 21836 14328 21864 14427
rect 22112 14396 22140 14427
rect 22922 14424 22928 14476
rect 22980 14464 22986 14476
rect 23569 14467 23627 14473
rect 23569 14464 23581 14467
rect 22980 14436 23581 14464
rect 22980 14424 22986 14436
rect 23569 14433 23581 14436
rect 23615 14464 23627 14467
rect 24136 14464 24164 14563
rect 25866 14560 25872 14572
rect 25924 14560 25930 14612
rect 27522 14560 27528 14612
rect 27580 14600 27586 14612
rect 29181 14603 29239 14609
rect 29181 14600 29193 14603
rect 27580 14572 29193 14600
rect 27580 14560 27586 14572
rect 29181 14569 29193 14572
rect 29227 14569 29239 14603
rect 29181 14563 29239 14569
rect 30742 14560 30748 14612
rect 30800 14600 30806 14612
rect 31113 14603 31171 14609
rect 31113 14600 31125 14603
rect 30800 14572 31125 14600
rect 30800 14560 30806 14572
rect 31113 14569 31125 14572
rect 31159 14569 31171 14603
rect 35710 14600 35716 14612
rect 35671 14572 35716 14600
rect 31113 14563 31171 14569
rect 35710 14560 35716 14572
rect 35768 14560 35774 14612
rect 40494 14560 40500 14612
rect 40552 14600 40558 14612
rect 41417 14603 41475 14609
rect 41417 14600 41429 14603
rect 40552 14572 41429 14600
rect 40552 14560 40558 14572
rect 41417 14569 41429 14572
rect 41463 14569 41475 14603
rect 41417 14563 41475 14569
rect 44085 14603 44143 14609
rect 44085 14569 44097 14603
rect 44131 14600 44143 14603
rect 44174 14600 44180 14612
rect 44131 14572 44180 14600
rect 44131 14569 44143 14572
rect 44085 14563 44143 14569
rect 44174 14560 44180 14572
rect 44232 14560 44238 14612
rect 48130 14560 48136 14612
rect 48188 14600 48194 14612
rect 48961 14603 49019 14609
rect 48961 14600 48973 14603
rect 48188 14572 48973 14600
rect 48188 14560 48194 14572
rect 48961 14569 48973 14572
rect 49007 14569 49019 14603
rect 48961 14563 49019 14569
rect 37734 14532 37740 14544
rect 33704 14504 37740 14532
rect 23615 14436 24164 14464
rect 23615 14433 23627 14436
rect 23569 14427 23627 14433
rect 25038 14424 25044 14476
rect 25096 14464 25102 14476
rect 25133 14467 25191 14473
rect 25133 14464 25145 14467
rect 25096 14436 25145 14464
rect 25096 14424 25102 14436
rect 25133 14433 25145 14436
rect 25179 14433 25191 14467
rect 26510 14464 26516 14476
rect 26471 14436 26516 14464
rect 25133 14427 25191 14433
rect 26510 14424 26516 14436
rect 26568 14424 26574 14476
rect 27614 14424 27620 14476
rect 27672 14464 27678 14476
rect 27801 14467 27859 14473
rect 27801 14464 27813 14467
rect 27672 14436 27813 14464
rect 27672 14424 27678 14436
rect 27801 14433 27813 14436
rect 27847 14464 27859 14467
rect 30098 14464 30104 14476
rect 27847 14436 30104 14464
rect 27847 14433 27859 14436
rect 27801 14427 27859 14433
rect 30098 14424 30104 14436
rect 30156 14424 30162 14476
rect 31021 14467 31079 14473
rect 31021 14433 31033 14467
rect 31067 14464 31079 14467
rect 32674 14464 32680 14476
rect 31067 14436 32680 14464
rect 31067 14433 31079 14436
rect 31021 14427 31079 14433
rect 32674 14424 32680 14436
rect 32732 14424 32738 14476
rect 33704 14473 33732 14504
rect 37734 14492 37740 14504
rect 37792 14492 37798 14544
rect 39390 14492 39396 14544
rect 39448 14532 39454 14544
rect 41141 14535 41199 14541
rect 41141 14532 41153 14535
rect 39448 14504 41153 14532
rect 39448 14492 39454 14504
rect 41141 14501 41153 14504
rect 41187 14532 41199 14535
rect 42794 14532 42800 14544
rect 41187 14504 42800 14532
rect 41187 14501 41199 14504
rect 41141 14495 41199 14501
rect 42794 14492 42800 14504
rect 42852 14492 42858 14544
rect 45649 14535 45707 14541
rect 45649 14501 45661 14535
rect 45695 14532 45707 14535
rect 47578 14532 47584 14544
rect 45695 14504 47584 14532
rect 45695 14501 45707 14504
rect 45649 14495 45707 14501
rect 47578 14492 47584 14504
rect 47636 14492 47642 14544
rect 49602 14532 49608 14544
rect 48424 14504 49608 14532
rect 33689 14467 33747 14473
rect 33689 14433 33701 14467
rect 33735 14433 33747 14467
rect 34054 14464 34060 14476
rect 33967 14436 34060 14464
rect 33689 14427 33747 14433
rect 34054 14424 34060 14436
rect 34112 14464 34118 14476
rect 35158 14464 35164 14476
rect 34112 14436 35164 14464
rect 34112 14424 34118 14436
rect 35158 14424 35164 14436
rect 35216 14424 35222 14476
rect 35253 14467 35311 14473
rect 35253 14433 35265 14467
rect 35299 14433 35311 14467
rect 35253 14427 35311 14433
rect 23845 14399 23903 14405
rect 23845 14396 23857 14399
rect 22112 14368 23857 14396
rect 23845 14365 23857 14368
rect 23891 14365 23903 14399
rect 23845 14359 23903 14365
rect 28077 14399 28135 14405
rect 28077 14365 28089 14399
rect 28123 14396 28135 14399
rect 28258 14396 28264 14408
rect 28123 14368 28264 14396
rect 28123 14365 28135 14368
rect 28077 14359 28135 14365
rect 28258 14356 28264 14368
rect 28316 14356 28322 14408
rect 31478 14356 31484 14408
rect 31536 14396 31542 14408
rect 33781 14399 33839 14405
rect 33781 14396 33793 14399
rect 31536 14368 33793 14396
rect 31536 14356 31542 14368
rect 33781 14365 33793 14368
rect 33827 14365 33839 14399
rect 34146 14396 34152 14408
rect 34107 14368 34152 14396
rect 33781 14359 33839 14365
rect 33796 14328 33824 14359
rect 34146 14356 34152 14368
rect 34204 14396 34210 14408
rect 35268 14396 35296 14427
rect 35434 14424 35440 14476
rect 35492 14464 35498 14476
rect 35529 14467 35587 14473
rect 35529 14464 35541 14467
rect 35492 14436 35541 14464
rect 35492 14424 35498 14436
rect 35529 14433 35541 14436
rect 35575 14464 35587 14467
rect 37826 14464 37832 14476
rect 35575 14436 37832 14464
rect 35575 14433 35587 14436
rect 35529 14427 35587 14433
rect 37826 14424 37832 14436
rect 37884 14424 37890 14476
rect 37921 14467 37979 14473
rect 37921 14433 37933 14467
rect 37967 14464 37979 14467
rect 38562 14464 38568 14476
rect 37967 14436 38568 14464
rect 37967 14433 37979 14436
rect 37921 14427 37979 14433
rect 38562 14424 38568 14436
rect 38620 14424 38626 14476
rect 40126 14464 40132 14476
rect 40087 14436 40132 14464
rect 40126 14424 40132 14436
rect 40184 14424 40190 14476
rect 41325 14467 41383 14473
rect 41325 14433 41337 14467
rect 41371 14464 41383 14467
rect 42518 14464 42524 14476
rect 41371 14436 42524 14464
rect 41371 14433 41383 14436
rect 41325 14427 41383 14433
rect 34204 14368 35296 14396
rect 34204 14356 34210 14368
rect 39758 14356 39764 14408
rect 39816 14396 39822 14408
rect 41340 14396 41368 14427
rect 42518 14424 42524 14436
rect 42576 14424 42582 14476
rect 42886 14424 42892 14476
rect 42944 14464 42950 14476
rect 43993 14467 44051 14473
rect 43993 14464 44005 14467
rect 42944 14436 44005 14464
rect 42944 14424 42950 14436
rect 43993 14433 44005 14436
rect 44039 14464 44051 14467
rect 44269 14467 44327 14473
rect 44269 14464 44281 14467
rect 44039 14436 44281 14464
rect 44039 14433 44051 14436
rect 43993 14427 44051 14433
rect 44269 14433 44281 14436
rect 44315 14464 44327 14467
rect 44726 14464 44732 14476
rect 44315 14436 44732 14464
rect 44315 14433 44327 14436
rect 44269 14427 44327 14433
rect 44726 14424 44732 14436
rect 44784 14424 44790 14476
rect 45830 14464 45836 14476
rect 45743 14436 45836 14464
rect 45830 14424 45836 14436
rect 45888 14464 45894 14476
rect 46750 14464 46756 14476
rect 45888 14436 46756 14464
rect 45888 14424 45894 14436
rect 46750 14424 46756 14436
rect 46808 14424 46814 14476
rect 46934 14424 46940 14476
rect 46992 14464 46998 14476
rect 47029 14467 47087 14473
rect 47029 14464 47041 14467
rect 46992 14436 47041 14464
rect 46992 14424 46998 14436
rect 47029 14433 47041 14436
rect 47075 14433 47087 14467
rect 47210 14464 47216 14476
rect 47171 14436 47216 14464
rect 47029 14427 47087 14433
rect 46198 14396 46204 14408
rect 39816 14368 41368 14396
rect 46159 14368 46204 14396
rect 39816 14356 39822 14368
rect 46198 14356 46204 14368
rect 46256 14356 46262 14408
rect 47044 14396 47072 14427
rect 47210 14424 47216 14436
rect 47268 14424 47274 14476
rect 48424 14396 48452 14504
rect 49602 14492 49608 14504
rect 49660 14532 49666 14544
rect 49660 14504 50200 14532
rect 49660 14492 49666 14504
rect 49694 14464 49700 14476
rect 49655 14436 49700 14464
rect 49694 14424 49700 14436
rect 49752 14424 49758 14476
rect 50172 14473 50200 14504
rect 50065 14467 50123 14473
rect 50065 14433 50077 14467
rect 50111 14433 50123 14467
rect 50065 14427 50123 14433
rect 50157 14467 50215 14473
rect 50157 14433 50169 14467
rect 50203 14433 50215 14467
rect 52270 14464 52276 14476
rect 52231 14436 52276 14464
rect 50157 14427 50215 14433
rect 47044 14368 48452 14396
rect 48961 14399 49019 14405
rect 48961 14365 48973 14399
rect 49007 14396 49019 14399
rect 49605 14399 49663 14405
rect 49605 14396 49617 14399
rect 49007 14368 49617 14396
rect 49007 14365 49019 14368
rect 48961 14359 49019 14365
rect 49605 14365 49617 14368
rect 49651 14365 49663 14399
rect 49605 14359 49663 14365
rect 34422 14328 34428 14340
rect 21836 14300 22784 14328
rect 33796 14300 34428 14328
rect 22756 14272 22784 14300
rect 34422 14288 34428 14300
rect 34480 14288 34486 14340
rect 35342 14328 35348 14340
rect 35303 14300 35348 14328
rect 35342 14288 35348 14300
rect 35400 14288 35406 14340
rect 35526 14288 35532 14340
rect 35584 14328 35590 14340
rect 37366 14328 37372 14340
rect 35584 14300 37372 14328
rect 35584 14288 35590 14300
rect 37366 14288 37372 14300
rect 37424 14328 37430 14340
rect 41690 14328 41696 14340
rect 37424 14300 41696 14328
rect 37424 14288 37430 14300
rect 41690 14288 41696 14300
rect 41748 14328 41754 14340
rect 42150 14328 42156 14340
rect 41748 14300 42156 14328
rect 41748 14288 41754 14300
rect 42150 14288 42156 14300
rect 42208 14288 42214 14340
rect 47210 14288 47216 14340
rect 47268 14328 47274 14340
rect 50080 14328 50108 14427
rect 52270 14424 52276 14436
rect 52328 14424 52334 14476
rect 51997 14399 52055 14405
rect 51997 14396 52009 14399
rect 51828 14368 52009 14396
rect 50706 14328 50712 14340
rect 47268 14300 50712 14328
rect 47268 14288 47274 14300
rect 50706 14288 50712 14300
rect 50764 14288 50770 14340
rect 51828 14272 51856 14368
rect 51997 14365 52009 14368
rect 52043 14365 52055 14399
rect 51997 14359 52055 14365
rect 18414 14260 18420 14272
rect 16592 14232 18420 14260
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 22186 14220 22192 14272
rect 22244 14260 22250 14272
rect 22281 14263 22339 14269
rect 22281 14260 22293 14263
rect 22244 14232 22293 14260
rect 22244 14220 22250 14232
rect 22281 14229 22293 14232
rect 22327 14229 22339 14263
rect 22738 14260 22744 14272
rect 22699 14232 22744 14260
rect 22281 14223 22339 14229
rect 22738 14220 22744 14232
rect 22796 14220 22802 14272
rect 25222 14260 25228 14272
rect 25183 14232 25228 14260
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 26234 14220 26240 14272
rect 26292 14260 26298 14272
rect 26605 14263 26663 14269
rect 26605 14260 26617 14263
rect 26292 14232 26617 14260
rect 26292 14220 26298 14232
rect 26605 14229 26617 14232
rect 26651 14229 26663 14263
rect 26605 14223 26663 14229
rect 29641 14263 29699 14269
rect 29641 14229 29653 14263
rect 29687 14260 29699 14263
rect 30098 14260 30104 14272
rect 29687 14232 30104 14260
rect 29687 14229 29699 14232
rect 29641 14223 29699 14229
rect 30098 14220 30104 14232
rect 30156 14220 30162 14272
rect 32030 14220 32036 14272
rect 32088 14260 32094 14272
rect 33137 14263 33195 14269
rect 33137 14260 33149 14263
rect 32088 14232 33149 14260
rect 32088 14220 32094 14232
rect 33137 14229 33149 14232
rect 33183 14229 33195 14263
rect 33137 14223 33195 14229
rect 37550 14220 37556 14272
rect 37608 14260 37614 14272
rect 38013 14263 38071 14269
rect 38013 14260 38025 14263
rect 37608 14232 38025 14260
rect 37608 14220 37614 14232
rect 38013 14229 38025 14232
rect 38059 14229 38071 14263
rect 38013 14223 38071 14229
rect 38473 14263 38531 14269
rect 38473 14229 38485 14263
rect 38519 14260 38531 14263
rect 38562 14260 38568 14272
rect 38519 14232 38568 14260
rect 38519 14229 38531 14232
rect 38473 14223 38531 14229
rect 38562 14220 38568 14232
rect 38620 14220 38626 14272
rect 40218 14260 40224 14272
rect 40179 14232 40224 14260
rect 40218 14220 40224 14232
rect 40276 14220 40282 14272
rect 49145 14263 49203 14269
rect 49145 14229 49157 14263
rect 49191 14260 49203 14263
rect 49602 14260 49608 14272
rect 49191 14232 49608 14260
rect 49191 14229 49203 14232
rect 49145 14223 49203 14229
rect 49602 14220 49608 14232
rect 49660 14220 49666 14272
rect 49786 14220 49792 14272
rect 49844 14260 49850 14272
rect 51442 14260 51448 14272
rect 49844 14232 51448 14260
rect 49844 14220 49850 14232
rect 51442 14220 51448 14232
rect 51500 14220 51506 14272
rect 51810 14260 51816 14272
rect 51771 14232 51816 14260
rect 51810 14220 51816 14232
rect 51868 14220 51874 14272
rect 52454 14220 52460 14272
rect 52512 14260 52518 14272
rect 53377 14263 53435 14269
rect 53377 14260 53389 14263
rect 52512 14232 53389 14260
rect 52512 14220 52518 14232
rect 53377 14229 53389 14232
rect 53423 14229 53435 14263
rect 53377 14223 53435 14229
rect 1104 14170 54832 14192
rect 1104 14118 9947 14170
rect 9999 14118 10011 14170
rect 10063 14118 10075 14170
rect 10127 14118 10139 14170
rect 10191 14118 27878 14170
rect 27930 14118 27942 14170
rect 27994 14118 28006 14170
rect 28058 14118 28070 14170
rect 28122 14118 45808 14170
rect 45860 14118 45872 14170
rect 45924 14118 45936 14170
rect 45988 14118 46000 14170
rect 46052 14118 54832 14170
rect 1104 14096 54832 14118
rect 5445 14059 5503 14065
rect 5445 14025 5457 14059
rect 5491 14056 5503 14059
rect 5534 14056 5540 14068
rect 5491 14028 5540 14056
rect 5491 14025 5503 14028
rect 5445 14019 5503 14025
rect 5534 14016 5540 14028
rect 5592 14056 5598 14068
rect 6270 14056 6276 14068
rect 5592 14028 6276 14056
rect 5592 14016 5598 14028
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8294 14056 8300 14068
rect 8159 14028 8300 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 14274 14056 14280 14068
rect 10827 14028 14280 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14826 14056 14832 14068
rect 14787 14028 14832 14056
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 18785 14059 18843 14065
rect 18785 14056 18797 14059
rect 15896 14028 18797 14056
rect 15896 14016 15902 14028
rect 18785 14025 18797 14028
rect 18831 14025 18843 14059
rect 20806 14056 20812 14068
rect 20767 14028 20812 14056
rect 18785 14019 18843 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 24305 14059 24363 14065
rect 24305 14025 24317 14059
rect 24351 14056 24363 14059
rect 25130 14056 25136 14068
rect 24351 14028 25136 14056
rect 24351 14025 24363 14028
rect 24305 14019 24363 14025
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 26418 14056 26424 14068
rect 26379 14028 26424 14056
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 28258 14056 28264 14068
rect 28219 14028 28264 14056
rect 28258 14016 28264 14028
rect 28316 14016 28322 14068
rect 29362 14056 29368 14068
rect 29323 14028 29368 14056
rect 29362 14016 29368 14028
rect 29420 14016 29426 14068
rect 41230 14056 41236 14068
rect 29472 14028 41236 14056
rect 4249 13991 4307 13997
rect 4249 13957 4261 13991
rect 4295 13957 4307 13991
rect 4249 13951 4307 13957
rect 7561 13991 7619 13997
rect 7561 13957 7573 13991
rect 7607 13988 7619 13991
rect 8754 13988 8760 14000
rect 7607 13960 8760 13988
rect 7607 13957 7619 13960
rect 7561 13951 7619 13957
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2317 13855 2375 13861
rect 2317 13852 2329 13855
rect 2280 13824 2329 13852
rect 2280 13812 2286 13824
rect 2317 13821 2329 13824
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 4264 13852 4292 13951
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 9769 13991 9827 13997
rect 9769 13957 9781 13991
rect 9815 13988 9827 13991
rect 11514 13988 11520 14000
rect 9815 13960 11520 13988
rect 9815 13957 9827 13960
rect 9769 13951 9827 13957
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 16942 13988 16948 14000
rect 16903 13960 16948 13988
rect 16942 13948 16948 13960
rect 17000 13948 17006 14000
rect 20824 13988 20852 14016
rect 21637 13991 21695 13997
rect 21637 13988 21649 13991
rect 20824 13960 21649 13988
rect 21637 13957 21649 13960
rect 21683 13957 21695 13991
rect 21637 13951 21695 13957
rect 22557 13991 22615 13997
rect 22557 13957 22569 13991
rect 22603 13957 22615 13991
rect 22557 13951 22615 13957
rect 12986 13920 12992 13932
rect 11256 13892 12992 13920
rect 4430 13852 4436 13864
rect 3467 13824 4292 13852
rect 4391 13824 4436 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 4430 13812 4436 13824
rect 4488 13812 4494 13864
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 5442 13852 5448 13864
rect 5399 13824 5448 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7156 13824 7757 13852
rect 7156 13812 7162 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 8018 13852 8024 13864
rect 7979 13824 8024 13852
rect 7745 13815 7803 13821
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 10965 13855 11023 13861
rect 9999 13824 10916 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 2133 13719 2191 13725
rect 2133 13685 2145 13719
rect 2179 13716 2191 13719
rect 2314 13716 2320 13728
rect 2179 13688 2320 13716
rect 2179 13685 2191 13688
rect 2133 13679 2191 13685
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 3234 13716 3240 13728
rect 3195 13688 3240 13716
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 10888 13716 10916 13824
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 11011 13824 11100 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11072 13784 11100 13824
rect 11256 13784 11284 13892
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13541 13923 13599 13929
rect 13096 13892 13400 13920
rect 13096 13852 13124 13892
rect 13262 13852 13268 13864
rect 11072 13756 11284 13784
rect 11348 13824 13124 13852
rect 13223 13824 13268 13852
rect 11348 13716 11376 13824
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13372 13852 13400 13892
rect 13541 13889 13553 13923
rect 13587 13920 13599 13923
rect 13630 13920 13636 13932
rect 13587 13892 13636 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 15470 13920 15476 13932
rect 13780 13892 15476 13920
rect 13780 13880 13786 13892
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15746 13920 15752 13932
rect 15707 13892 15752 13920
rect 15746 13880 15752 13892
rect 15804 13920 15810 13932
rect 19613 13923 19671 13929
rect 15804 13892 16068 13920
rect 15804 13880 15810 13892
rect 13814 13852 13820 13864
rect 13372 13824 13820 13852
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13821 15991 13855
rect 16040 13852 16068 13892
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 22572 13920 22600 13951
rect 22738 13948 22744 14000
rect 22796 13988 22802 14000
rect 29472 13988 29500 14028
rect 41230 14016 41236 14028
rect 41288 14016 41294 14068
rect 43714 14056 43720 14068
rect 43675 14028 43720 14056
rect 43714 14016 43720 14028
rect 43772 14016 43778 14068
rect 44729 14059 44787 14065
rect 44729 14025 44741 14059
rect 44775 14056 44787 14059
rect 44818 14056 44824 14068
rect 44775 14028 44824 14056
rect 44775 14025 44787 14028
rect 44729 14019 44787 14025
rect 44818 14016 44824 14028
rect 44876 14056 44882 14068
rect 45186 14056 45192 14068
rect 44876 14028 45192 14056
rect 44876 14016 44882 14028
rect 45186 14016 45192 14028
rect 45244 14016 45250 14068
rect 46293 14059 46351 14065
rect 46293 14025 46305 14059
rect 46339 14056 46351 14059
rect 47213 14059 47271 14065
rect 47213 14056 47225 14059
rect 46339 14028 47225 14056
rect 46339 14025 46351 14028
rect 46293 14019 46351 14025
rect 47213 14025 47225 14028
rect 47259 14056 47271 14059
rect 49786 14056 49792 14068
rect 47259 14028 49792 14056
rect 47259 14025 47271 14028
rect 47213 14019 47271 14025
rect 49786 14016 49792 14028
rect 49844 14016 49850 14068
rect 50706 14056 50712 14068
rect 50667 14028 50712 14056
rect 50706 14016 50712 14028
rect 50764 14016 50770 14068
rect 51994 14056 52000 14068
rect 51955 14028 52000 14056
rect 51994 14016 52000 14028
rect 52052 14016 52058 14068
rect 52454 14056 52460 14068
rect 52415 14028 52460 14056
rect 52454 14016 52460 14028
rect 52512 14016 52518 14068
rect 32582 13988 32588 14000
rect 22796 13960 29500 13988
rect 32543 13960 32588 13988
rect 22796 13948 22802 13960
rect 32582 13948 32588 13960
rect 32640 13948 32646 14000
rect 32950 13988 32956 14000
rect 32911 13960 32956 13988
rect 32950 13948 32956 13960
rect 33008 13948 33014 14000
rect 33873 13991 33931 13997
rect 33873 13957 33885 13991
rect 33919 13988 33931 13991
rect 35342 13988 35348 14000
rect 33919 13960 35348 13988
rect 33919 13957 33931 13960
rect 33873 13951 33931 13957
rect 35342 13948 35348 13960
rect 35400 13948 35406 14000
rect 37366 13988 37372 14000
rect 37327 13960 37372 13988
rect 37366 13948 37372 13960
rect 37424 13948 37430 14000
rect 45005 13991 45063 13997
rect 45005 13957 45017 13991
rect 45051 13957 45063 13991
rect 45005 13951 45063 13957
rect 24854 13920 24860 13932
rect 19659 13892 21128 13920
rect 22572 13892 24860 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 16040 13824 16405 13852
rect 15933 13815 15991 13821
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13852 16543 13855
rect 16574 13852 16580 13864
rect 16531 13824 16580 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 15948 13784 15976 13815
rect 16500 13784 16528 13815
rect 16574 13812 16580 13824
rect 16632 13812 16638 13864
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 18969 13855 19027 13861
rect 18969 13852 18981 13855
rect 16724 13824 18981 13852
rect 16724 13812 16730 13824
rect 18969 13821 18981 13824
rect 19015 13821 19027 13855
rect 19426 13852 19432 13864
rect 19387 13824 19432 13852
rect 18969 13815 19027 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19794 13852 19800 13864
rect 19755 13824 19800 13852
rect 19794 13812 19800 13824
rect 19852 13812 19858 13864
rect 21100 13861 21128 13892
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 24946 13880 24952 13932
rect 25004 13920 25010 13932
rect 25225 13923 25283 13929
rect 25225 13920 25237 13923
rect 25004 13892 25237 13920
rect 25004 13880 25010 13892
rect 25225 13889 25237 13892
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 30098 13880 30104 13932
rect 30156 13920 30162 13932
rect 31205 13923 31263 13929
rect 31205 13920 31217 13923
rect 30156 13892 31217 13920
rect 30156 13880 30162 13892
rect 31205 13889 31217 13892
rect 31251 13920 31263 13923
rect 32968 13920 32996 13948
rect 38562 13920 38568 13932
rect 31251 13892 32996 13920
rect 34072 13892 38568 13920
rect 31251 13889 31263 13892
rect 31205 13883 31263 13889
rect 21085 13855 21143 13861
rect 21085 13821 21097 13855
rect 21131 13821 21143 13855
rect 22738 13852 22744 13864
rect 22699 13824 22744 13852
rect 21085 13815 21143 13821
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 24210 13852 24216 13864
rect 24171 13824 24216 13852
rect 24210 13812 24216 13824
rect 24268 13812 24274 13864
rect 24762 13812 24768 13864
rect 24820 13852 24826 13864
rect 25041 13855 25099 13861
rect 25041 13852 25053 13855
rect 24820 13824 25053 13852
rect 24820 13812 24826 13824
rect 25041 13821 25053 13824
rect 25087 13852 25099 13855
rect 25406 13852 25412 13864
rect 25087 13824 25268 13852
rect 25367 13824 25412 13852
rect 25087 13821 25099 13824
rect 25041 13815 25099 13821
rect 20990 13784 20996 13796
rect 15948 13756 16528 13784
rect 20951 13756 20996 13784
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 25240 13784 25268 13824
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 25869 13855 25927 13861
rect 25869 13852 25881 13855
rect 25516 13824 25881 13852
rect 25516 13784 25544 13824
rect 25869 13821 25881 13824
rect 25915 13821 25927 13855
rect 25869 13815 25927 13821
rect 25961 13855 26019 13861
rect 25961 13821 25973 13855
rect 26007 13852 26019 13855
rect 26510 13852 26516 13864
rect 26007 13824 26516 13852
rect 26007 13821 26019 13824
rect 25961 13815 26019 13821
rect 26510 13812 26516 13824
rect 26568 13812 26574 13864
rect 28169 13855 28227 13861
rect 28169 13821 28181 13855
rect 28215 13852 28227 13855
rect 29086 13852 29092 13864
rect 28215 13824 29092 13852
rect 28215 13821 28227 13824
rect 28169 13815 28227 13821
rect 29086 13812 29092 13824
rect 29144 13812 29150 13864
rect 29270 13852 29276 13864
rect 29231 13824 29276 13852
rect 29270 13812 29276 13824
rect 29328 13812 29334 13864
rect 31478 13852 31484 13864
rect 31439 13824 31484 13852
rect 31478 13812 31484 13824
rect 31536 13812 31542 13864
rect 33042 13812 33048 13864
rect 33100 13852 33106 13864
rect 34072 13861 34100 13892
rect 38562 13880 38568 13892
rect 38620 13880 38626 13932
rect 40218 13880 40224 13932
rect 40276 13920 40282 13932
rect 42613 13923 42671 13929
rect 42613 13920 42625 13923
rect 40276 13892 42625 13920
rect 40276 13880 40282 13892
rect 42613 13889 42625 13892
rect 42659 13889 42671 13923
rect 42613 13883 42671 13889
rect 42702 13880 42708 13932
rect 42760 13920 42766 13932
rect 45020 13920 45048 13951
rect 45278 13948 45284 14000
rect 45336 13988 45342 14000
rect 45336 13960 51948 13988
rect 45336 13948 45342 13960
rect 42760 13892 46152 13920
rect 42760 13880 42766 13892
rect 33781 13855 33839 13861
rect 33781 13852 33793 13855
rect 33100 13824 33793 13852
rect 33100 13812 33106 13824
rect 33781 13821 33793 13824
rect 33827 13852 33839 13855
rect 34057 13855 34115 13861
rect 34057 13852 34069 13855
rect 33827 13824 34069 13852
rect 33827 13821 33839 13824
rect 33781 13815 33839 13821
rect 34057 13821 34069 13824
rect 34103 13821 34115 13855
rect 34057 13815 34115 13821
rect 34146 13812 34152 13864
rect 34204 13852 34210 13864
rect 35253 13855 35311 13861
rect 35253 13852 35265 13855
rect 34204 13824 35265 13852
rect 34204 13812 34210 13824
rect 35253 13821 35265 13824
rect 35299 13821 35311 13855
rect 35434 13852 35440 13864
rect 35395 13824 35440 13852
rect 35253 13815 35311 13821
rect 35434 13812 35440 13824
rect 35492 13812 35498 13864
rect 35805 13855 35863 13861
rect 35805 13821 35817 13855
rect 35851 13852 35863 13855
rect 35986 13852 35992 13864
rect 35851 13824 35992 13852
rect 35851 13821 35863 13824
rect 35805 13815 35863 13821
rect 35986 13812 35992 13824
rect 36044 13812 36050 13864
rect 37550 13852 37556 13864
rect 37511 13824 37556 13852
rect 37550 13812 37556 13824
rect 37608 13812 37614 13864
rect 37642 13812 37648 13864
rect 37700 13852 37706 13864
rect 39393 13855 39451 13861
rect 37700 13824 37745 13852
rect 37700 13812 37706 13824
rect 39393 13821 39405 13855
rect 39439 13821 39451 13855
rect 39393 13815 39451 13821
rect 39485 13855 39543 13861
rect 39485 13821 39497 13855
rect 39531 13852 39543 13855
rect 40862 13852 40868 13864
rect 39531 13824 40868 13852
rect 39531 13821 39543 13824
rect 39485 13815 39543 13821
rect 25240 13756 25544 13784
rect 38105 13787 38163 13793
rect 38105 13753 38117 13787
rect 38151 13784 38163 13787
rect 38194 13784 38200 13796
rect 38151 13756 38200 13784
rect 38151 13753 38163 13756
rect 38105 13747 38163 13753
rect 38194 13744 38200 13756
rect 38252 13744 38258 13796
rect 39301 13787 39359 13793
rect 39301 13753 39313 13787
rect 39347 13784 39359 13787
rect 39408 13784 39436 13815
rect 40862 13812 40868 13824
rect 40920 13852 40926 13864
rect 41233 13855 41291 13861
rect 41233 13852 41245 13855
rect 40920 13824 41245 13852
rect 40920 13812 40926 13824
rect 41233 13821 41245 13824
rect 41279 13821 41291 13855
rect 41233 13815 41291 13821
rect 42245 13855 42303 13861
rect 42245 13821 42257 13855
rect 42291 13852 42303 13855
rect 42337 13855 42395 13861
rect 42337 13852 42349 13855
rect 42291 13824 42349 13852
rect 42291 13821 42303 13824
rect 42245 13815 42303 13821
rect 42337 13821 42349 13824
rect 42383 13852 42395 13855
rect 43070 13852 43076 13864
rect 42383 13824 43076 13852
rect 42383 13821 42395 13824
rect 42337 13815 42395 13821
rect 43070 13812 43076 13824
rect 43128 13852 43134 13864
rect 43990 13852 43996 13864
rect 43128 13824 43996 13852
rect 43128 13812 43134 13824
rect 43990 13812 43996 13824
rect 44048 13812 44054 13864
rect 44818 13852 44824 13864
rect 44779 13824 44824 13852
rect 44818 13812 44824 13824
rect 44876 13812 44882 13864
rect 46124 13861 46152 13892
rect 49694 13880 49700 13932
rect 49752 13920 49758 13932
rect 49752 13892 51764 13920
rect 49752 13880 49758 13892
rect 46109 13855 46167 13861
rect 46109 13821 46121 13855
rect 46155 13852 46167 13855
rect 46477 13855 46535 13861
rect 46477 13852 46489 13855
rect 46155 13824 46489 13852
rect 46155 13821 46167 13824
rect 46109 13815 46167 13821
rect 46477 13821 46489 13824
rect 46523 13821 46535 13855
rect 46477 13815 46535 13821
rect 47302 13812 47308 13864
rect 47360 13852 47366 13864
rect 47489 13855 47547 13861
rect 47489 13852 47501 13855
rect 47360 13824 47501 13852
rect 47360 13812 47366 13824
rect 47489 13821 47501 13824
rect 47535 13821 47547 13855
rect 49602 13852 49608 13864
rect 49563 13824 49608 13852
rect 47489 13815 47547 13821
rect 49602 13812 49608 13824
rect 49660 13812 49666 13864
rect 50617 13855 50675 13861
rect 50617 13821 50629 13855
rect 50663 13852 50675 13855
rect 51442 13852 51448 13864
rect 50663 13824 51448 13852
rect 50663 13821 50675 13824
rect 50617 13815 50675 13821
rect 51442 13812 51448 13824
rect 51500 13812 51506 13864
rect 51736 13861 51764 13892
rect 51920 13861 51948 13960
rect 51721 13855 51779 13861
rect 51721 13821 51733 13855
rect 51767 13821 51779 13855
rect 51721 13815 51779 13821
rect 51905 13855 51963 13861
rect 51905 13821 51917 13855
rect 51951 13852 51963 13855
rect 52472 13852 52500 14016
rect 51951 13824 52500 13852
rect 51951 13821 51963 13824
rect 51905 13815 51963 13821
rect 41690 13784 41696 13796
rect 39347 13756 41696 13784
rect 39347 13753 39359 13756
rect 39301 13747 39359 13753
rect 41690 13744 41696 13756
rect 41748 13744 41754 13796
rect 47118 13744 47124 13796
rect 47176 13784 47182 13796
rect 47397 13787 47455 13793
rect 47397 13784 47409 13787
rect 47176 13756 47409 13784
rect 47176 13744 47182 13756
rect 47397 13753 47409 13756
rect 47443 13753 47455 13787
rect 47397 13747 47455 13753
rect 47949 13787 48007 13793
rect 47949 13753 47961 13787
rect 47995 13784 48007 13787
rect 48222 13784 48228 13796
rect 47995 13756 48228 13784
rect 47995 13753 48007 13756
rect 47949 13747 48007 13753
rect 48222 13744 48228 13756
rect 48280 13744 48286 13796
rect 10888 13688 11376 13716
rect 13262 13676 13268 13728
rect 13320 13716 13326 13728
rect 14918 13716 14924 13728
rect 13320 13688 14924 13716
rect 13320 13676 13326 13688
rect 14918 13676 14924 13688
rect 14976 13716 14982 13728
rect 15013 13719 15071 13725
rect 15013 13716 15025 13719
rect 14976 13688 15025 13716
rect 14976 13676 14982 13688
rect 15013 13685 15025 13688
rect 15059 13685 15071 13719
rect 15013 13679 15071 13685
rect 30926 13676 30932 13728
rect 30984 13716 30990 13728
rect 41322 13716 41328 13728
rect 30984 13688 41328 13716
rect 30984 13676 30990 13688
rect 41322 13676 41328 13688
rect 41380 13676 41386 13728
rect 41417 13719 41475 13725
rect 41417 13685 41429 13719
rect 41463 13716 41475 13719
rect 41506 13716 41512 13728
rect 41463 13688 41512 13716
rect 41463 13685 41475 13688
rect 41417 13679 41475 13685
rect 41506 13676 41512 13688
rect 41564 13676 41570 13728
rect 49694 13716 49700 13728
rect 49655 13688 49700 13716
rect 49694 13676 49700 13688
rect 49752 13676 49758 13728
rect 1104 13626 54832 13648
rect 1104 13574 18912 13626
rect 18964 13574 18976 13626
rect 19028 13574 19040 13626
rect 19092 13574 19104 13626
rect 19156 13574 36843 13626
rect 36895 13574 36907 13626
rect 36959 13574 36971 13626
rect 37023 13574 37035 13626
rect 37087 13574 54832 13626
rect 1104 13552 54832 13574
rect 4430 13512 4436 13524
rect 4391 13484 4436 13512
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 8386 13472 8392 13524
rect 8444 13512 8450 13524
rect 8665 13515 8723 13521
rect 8665 13512 8677 13515
rect 8444 13484 8677 13512
rect 8444 13472 8450 13484
rect 8665 13481 8677 13484
rect 8711 13481 8723 13515
rect 16022 13512 16028 13524
rect 15983 13484 16028 13512
rect 8665 13475 8723 13481
rect 7006 13444 7012 13456
rect 5368 13416 7012 13444
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 5368 13385 5396 13416
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 4985 13379 5043 13385
rect 4985 13376 4997 13379
rect 4948 13348 4997 13376
rect 4948 13336 4954 13348
rect 4985 13345 4997 13348
rect 5031 13345 5043 13379
rect 4985 13339 5043 13345
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 6914 13376 6920 13388
rect 5500 13348 5545 13376
rect 6875 13348 6920 13376
rect 5500 13336 5506 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7190 13376 7196 13388
rect 7151 13348 7196 13376
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 8680 13376 8708 13475
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 22370 13512 22376 13524
rect 22331 13484 22376 13512
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 24946 13472 24952 13524
rect 25004 13512 25010 13524
rect 26789 13515 26847 13521
rect 26789 13512 26801 13515
rect 25004 13484 26801 13512
rect 25004 13472 25010 13484
rect 26789 13481 26801 13484
rect 26835 13481 26847 13515
rect 29546 13512 29552 13524
rect 29507 13484 29552 13512
rect 26789 13475 26847 13481
rect 29546 13472 29552 13484
rect 29604 13472 29610 13524
rect 30009 13515 30067 13521
rect 30009 13481 30021 13515
rect 30055 13512 30067 13515
rect 30098 13512 30104 13524
rect 30055 13484 30104 13512
rect 30055 13481 30067 13484
rect 30009 13475 30067 13481
rect 30098 13472 30104 13484
rect 30156 13472 30162 13524
rect 31113 13515 31171 13521
rect 31113 13481 31125 13515
rect 31159 13512 31171 13515
rect 31478 13512 31484 13524
rect 31159 13484 31484 13512
rect 31159 13481 31171 13484
rect 31113 13475 31171 13481
rect 31478 13472 31484 13484
rect 31536 13472 31542 13524
rect 42150 13512 42156 13524
rect 42111 13484 42156 13512
rect 42150 13472 42156 13484
rect 42208 13472 42214 13524
rect 45557 13515 45615 13521
rect 45557 13481 45569 13515
rect 45603 13512 45615 13515
rect 45646 13512 45652 13524
rect 45603 13484 45652 13512
rect 45603 13481 45615 13484
rect 45557 13475 45615 13481
rect 45646 13472 45652 13484
rect 45704 13472 45710 13524
rect 51442 13512 51448 13524
rect 51403 13484 51448 13512
rect 51442 13472 51448 13484
rect 51500 13472 51506 13524
rect 16761 13447 16819 13453
rect 16761 13413 16773 13447
rect 16807 13444 16819 13447
rect 17218 13444 17224 13456
rect 16807 13416 17224 13444
rect 16807 13413 16819 13416
rect 16761 13407 16819 13413
rect 17218 13404 17224 13416
rect 17276 13444 17282 13456
rect 19245 13447 19303 13453
rect 19245 13444 19257 13447
rect 17276 13416 19257 13444
rect 17276 13404 17282 13416
rect 19245 13413 19257 13416
rect 19291 13413 19303 13447
rect 19245 13407 19303 13413
rect 24210 13404 24216 13456
rect 24268 13444 24274 13456
rect 24397 13447 24455 13453
rect 24397 13444 24409 13447
rect 24268 13416 24409 13444
rect 24268 13404 24274 13416
rect 24397 13413 24409 13416
rect 24443 13413 24455 13447
rect 25682 13444 25688 13456
rect 24397 13407 24455 13413
rect 25332 13416 25688 13444
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 8680 13348 9689 13376
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13376 10011 13379
rect 10318 13376 10324 13388
rect 9999 13348 10324 13376
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 5534 13308 5540 13320
rect 5123 13280 5540 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 9692 13308 9720 13339
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 16209 13379 16267 13385
rect 12492 13348 12537 13376
rect 12492 13336 12498 13348
rect 16209 13345 16221 13379
rect 16255 13345 16267 13379
rect 16666 13376 16672 13388
rect 16627 13348 16672 13376
rect 16209 13339 16267 13345
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 9692 13280 11437 13308
rect 11425 13277 11437 13280
rect 11471 13308 11483 13311
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 11471 13280 12173 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 12161 13277 12173 13280
rect 12207 13308 12219 13311
rect 13262 13308 13268 13320
rect 12207 13280 13268 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 13262 13268 13268 13280
rect 13320 13308 13326 13320
rect 13909 13311 13967 13317
rect 13909 13308 13921 13311
rect 13320 13280 13921 13308
rect 13320 13268 13326 13280
rect 13909 13277 13921 13280
rect 13955 13277 13967 13311
rect 16224 13308 16252 13339
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13345 17923 13379
rect 17865 13339 17923 13345
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 21266 13376 21272 13388
rect 18095 13348 19656 13376
rect 21227 13348 21272 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 17678 13308 17684 13320
rect 16224 13280 17684 13308
rect 13909 13271 13967 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 17880 13240 17908 13339
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13308 18475 13311
rect 19334 13308 19340 13320
rect 18463 13280 19340 13308
rect 18463 13277 18475 13280
rect 18417 13271 18475 13277
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19628 13317 19656 13348
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 25038 13376 25044 13388
rect 24951 13348 25044 13376
rect 25038 13336 25044 13348
rect 25096 13376 25102 13388
rect 25222 13376 25228 13388
rect 25096 13348 25228 13376
rect 25096 13336 25102 13348
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 19613 13311 19671 13317
rect 19484 13280 19564 13308
rect 19484 13268 19490 13280
rect 19536 13249 19564 13280
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 19794 13308 19800 13320
rect 19659 13280 19800 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 19794 13268 19800 13280
rect 19852 13268 19858 13320
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 20993 13311 21051 13317
rect 20993 13308 21005 13311
rect 20772 13280 21005 13308
rect 20772 13268 20778 13280
rect 20993 13277 21005 13280
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13308 25191 13311
rect 25332 13308 25360 13416
rect 25682 13404 25688 13416
rect 25740 13404 25746 13456
rect 26252 13416 26740 13444
rect 26252 13388 26280 13416
rect 25409 13379 25467 13385
rect 25409 13345 25421 13379
rect 25455 13376 25467 13379
rect 26234 13376 26240 13388
rect 25455 13348 26240 13376
rect 25455 13345 25467 13348
rect 25409 13339 25467 13345
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 26712 13385 26740 13416
rect 26878 13404 26884 13456
rect 26936 13444 26942 13456
rect 32861 13447 32919 13453
rect 26936 13416 28304 13444
rect 26936 13404 26942 13416
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13345 26571 13379
rect 26513 13339 26571 13345
rect 26697 13379 26755 13385
rect 26697 13345 26709 13379
rect 26743 13345 26755 13379
rect 26697 13339 26755 13345
rect 25179 13280 25360 13308
rect 25501 13311 25559 13317
rect 25179 13277 25191 13280
rect 25133 13271 25191 13277
rect 25501 13277 25513 13311
rect 25547 13308 25559 13311
rect 26528 13308 26556 13339
rect 27614 13336 27620 13388
rect 27672 13376 27678 13388
rect 28169 13379 28227 13385
rect 28169 13376 28181 13379
rect 27672 13348 28181 13376
rect 27672 13336 27678 13348
rect 28169 13345 28181 13348
rect 28215 13345 28227 13379
rect 28276 13376 28304 13416
rect 32861 13413 32873 13447
rect 32907 13444 32919 13447
rect 34146 13444 34152 13456
rect 32907 13416 34152 13444
rect 32907 13413 32919 13416
rect 32861 13407 32919 13413
rect 34146 13404 34152 13416
rect 34204 13404 34210 13456
rect 35342 13404 35348 13456
rect 35400 13444 35406 13456
rect 36541 13447 36599 13453
rect 35400 13416 36216 13444
rect 35400 13404 35406 13416
rect 30926 13376 30932 13388
rect 28276 13348 30932 13376
rect 28169 13339 28227 13345
rect 30926 13336 30932 13348
rect 30984 13336 30990 13388
rect 31021 13379 31079 13385
rect 31021 13345 31033 13379
rect 31067 13376 31079 13379
rect 32030 13376 32036 13388
rect 31067 13348 32036 13376
rect 31067 13345 31079 13348
rect 31021 13339 31079 13345
rect 32030 13336 32036 13348
rect 32088 13336 32094 13388
rect 32125 13379 32183 13385
rect 32125 13345 32137 13379
rect 32171 13345 32183 13379
rect 32398 13376 32404 13388
rect 32359 13348 32404 13376
rect 32125 13339 32183 13345
rect 28442 13308 28448 13320
rect 25547 13280 26556 13308
rect 28403 13280 28448 13308
rect 25547 13277 25559 13280
rect 25501 13271 25559 13277
rect 19521 13243 19579 13249
rect 19521 13240 19533 13243
rect 17880 13212 19533 13240
rect 19521 13209 19533 13212
rect 19567 13209 19579 13243
rect 19521 13203 19579 13209
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 2314 13172 2320 13184
rect 2179 13144 2320 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8297 13175 8355 13181
rect 8297 13172 8309 13175
rect 8076 13144 8309 13172
rect 8076 13132 8082 13144
rect 8297 13141 8309 13144
rect 8343 13141 8355 13175
rect 8297 13135 8355 13141
rect 10318 13132 10324 13184
rect 10376 13172 10382 13184
rect 10870 13172 10876 13184
rect 10376 13144 10876 13172
rect 10376 13132 10382 13144
rect 10870 13132 10876 13144
rect 10928 13172 10934 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10928 13144 11069 13172
rect 10928 13132 10934 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 13538 13172 13544 13184
rect 13499 13144 13544 13172
rect 11057 13135 11115 13141
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 19426 13181 19432 13184
rect 19410 13175 19432 13181
rect 19410 13141 19422 13175
rect 19484 13172 19490 13184
rect 19794 13172 19800 13184
rect 19484 13144 19800 13172
rect 19410 13135 19432 13141
rect 19426 13132 19432 13135
rect 19484 13132 19490 13144
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 19889 13175 19947 13181
rect 19889 13141 19901 13175
rect 19935 13172 19947 13175
rect 25608 13172 25636 13280
rect 28442 13268 28448 13280
rect 28500 13268 28506 13320
rect 31662 13268 31668 13320
rect 31720 13308 31726 13320
rect 32140 13308 32168 13339
rect 32398 13336 32404 13348
rect 32456 13336 32462 13388
rect 33962 13336 33968 13388
rect 34020 13376 34026 13388
rect 34425 13379 34483 13385
rect 34425 13376 34437 13379
rect 34020 13348 34437 13376
rect 34020 13336 34026 13348
rect 34425 13345 34437 13348
rect 34471 13345 34483 13379
rect 34425 13339 34483 13345
rect 34514 13336 34520 13388
rect 34572 13376 34578 13388
rect 35986 13376 35992 13388
rect 34572 13348 34617 13376
rect 35947 13348 35992 13376
rect 34572 13336 34578 13348
rect 35986 13336 35992 13348
rect 36044 13336 36050 13388
rect 36188 13385 36216 13416
rect 36541 13413 36553 13447
rect 36587 13444 36599 13447
rect 37642 13444 37648 13456
rect 36587 13416 37648 13444
rect 36587 13413 36599 13416
rect 36541 13407 36599 13413
rect 37642 13404 37648 13416
rect 37700 13404 37706 13456
rect 41322 13404 41328 13456
rect 41380 13444 41386 13456
rect 45664 13444 45692 13472
rect 46750 13444 46756 13456
rect 41380 13416 45508 13444
rect 45664 13416 46756 13444
rect 41380 13404 41386 13416
rect 36173 13379 36231 13385
rect 36173 13345 36185 13379
rect 36219 13345 36231 13379
rect 38194 13376 38200 13388
rect 38155 13348 38200 13376
rect 36173 13339 36231 13345
rect 38194 13336 38200 13348
rect 38252 13336 38258 13388
rect 40862 13376 40868 13388
rect 38304 13348 39804 13376
rect 40823 13348 40868 13376
rect 31720 13280 32168 13308
rect 32217 13311 32275 13317
rect 31720 13268 31726 13280
rect 32217 13277 32229 13311
rect 32263 13308 32275 13311
rect 33226 13308 33232 13320
rect 32263 13280 33232 13308
rect 32263 13277 32275 13280
rect 32217 13271 32275 13277
rect 33226 13268 33232 13280
rect 33284 13308 33290 13320
rect 33502 13308 33508 13320
rect 33284 13280 33508 13308
rect 33284 13268 33290 13280
rect 33502 13268 33508 13280
rect 33560 13268 33566 13320
rect 34974 13308 34980 13320
rect 34935 13280 34980 13308
rect 34974 13268 34980 13280
rect 35032 13268 35038 13320
rect 37921 13311 37979 13317
rect 37921 13277 37933 13311
rect 37967 13308 37979 13311
rect 38304 13308 38332 13348
rect 37967 13280 38332 13308
rect 37967 13277 37979 13280
rect 37921 13271 37979 13277
rect 38562 13268 38568 13320
rect 38620 13308 38626 13320
rect 39301 13311 39359 13317
rect 39301 13308 39313 13311
rect 38620 13280 39313 13308
rect 38620 13268 38626 13280
rect 39301 13277 39313 13280
rect 39347 13277 39359 13311
rect 39301 13271 39359 13277
rect 34241 13243 34299 13249
rect 34241 13209 34253 13243
rect 34287 13240 34299 13243
rect 35526 13240 35532 13252
rect 34287 13212 35532 13240
rect 34287 13209 34299 13212
rect 34241 13203 34299 13209
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 39776 13181 39804 13348
rect 40862 13336 40868 13348
rect 40920 13336 40926 13388
rect 41414 13336 41420 13388
rect 41472 13376 41478 13388
rect 41969 13379 42027 13385
rect 41969 13376 41981 13379
rect 41472 13348 41981 13376
rect 41472 13336 41478 13348
rect 41969 13345 41981 13348
rect 42015 13376 42027 13379
rect 42337 13379 42395 13385
rect 42337 13376 42349 13379
rect 42015 13348 42349 13376
rect 42015 13345 42027 13348
rect 41969 13339 42027 13345
rect 42337 13345 42349 13348
rect 42383 13376 42395 13379
rect 42702 13376 42708 13388
rect 42383 13348 42708 13376
rect 42383 13345 42395 13348
rect 42337 13339 42395 13345
rect 42702 13336 42708 13348
rect 42760 13336 42766 13388
rect 44450 13376 44456 13388
rect 44411 13348 44456 13376
rect 44450 13336 44456 13348
rect 44508 13336 44514 13388
rect 45480 13385 45508 13416
rect 46750 13404 46756 13416
rect 46808 13444 46814 13456
rect 46808 13416 47532 13444
rect 46808 13404 46814 13416
rect 45465 13379 45523 13385
rect 45465 13345 45477 13379
rect 45511 13376 45523 13379
rect 45741 13379 45799 13385
rect 45741 13376 45753 13379
rect 45511 13348 45753 13376
rect 45511 13345 45523 13348
rect 45465 13339 45523 13345
rect 45741 13345 45753 13348
rect 45787 13345 45799 13379
rect 45741 13339 45799 13345
rect 43622 13308 43628 13320
rect 43583 13280 43628 13308
rect 43622 13268 43628 13280
rect 43680 13268 43686 13320
rect 44082 13268 44088 13320
rect 44140 13308 44146 13320
rect 44177 13311 44235 13317
rect 44177 13308 44189 13311
rect 44140 13280 44189 13308
rect 44140 13268 44146 13280
rect 44177 13277 44189 13280
rect 44223 13277 44235 13311
rect 44177 13271 44235 13277
rect 44266 13268 44272 13320
rect 44324 13308 44330 13320
rect 44637 13311 44695 13317
rect 44637 13308 44649 13311
rect 44324 13280 44649 13308
rect 44324 13268 44330 13280
rect 44637 13277 44649 13280
rect 44683 13277 44695 13311
rect 44637 13271 44695 13277
rect 19935 13144 25636 13172
rect 39761 13175 39819 13181
rect 19935 13141 19947 13144
rect 19889 13135 19947 13141
rect 39761 13141 39773 13175
rect 39807 13172 39819 13175
rect 40862 13172 40868 13184
rect 39807 13144 40868 13172
rect 39807 13141 39819 13144
rect 39761 13135 39819 13141
rect 40862 13132 40868 13144
rect 40920 13132 40926 13184
rect 41046 13172 41052 13184
rect 41007 13144 41052 13172
rect 41046 13132 41052 13144
rect 41104 13132 41110 13184
rect 45756 13172 45784 13339
rect 46198 13336 46204 13388
rect 46256 13376 46262 13388
rect 46566 13376 46572 13388
rect 46256 13348 46572 13376
rect 46256 13336 46262 13348
rect 46566 13336 46572 13348
rect 46624 13376 46630 13388
rect 46937 13379 46995 13385
rect 46937 13376 46949 13379
rect 46624 13348 46949 13376
rect 46624 13336 46630 13348
rect 46937 13345 46949 13348
rect 46983 13345 46995 13379
rect 47302 13376 47308 13388
rect 47263 13348 47308 13376
rect 46937 13339 46995 13345
rect 47302 13336 47308 13348
rect 47360 13336 47366 13388
rect 47504 13385 47532 13416
rect 47489 13379 47547 13385
rect 47489 13345 47501 13379
rect 47535 13345 47547 13379
rect 47489 13339 47547 13345
rect 49694 13336 49700 13388
rect 49752 13376 49758 13388
rect 50341 13379 50399 13385
rect 50341 13376 50353 13379
rect 49752 13348 50353 13376
rect 49752 13336 49758 13348
rect 50341 13345 50353 13348
rect 50387 13345 50399 13379
rect 50341 13339 50399 13345
rect 47854 13268 47860 13320
rect 47912 13308 47918 13320
rect 49973 13311 50031 13317
rect 49973 13308 49985 13311
rect 47912 13280 49985 13308
rect 47912 13268 47918 13280
rect 49973 13277 49985 13280
rect 50019 13308 50031 13311
rect 50065 13311 50123 13317
rect 50065 13308 50077 13311
rect 50019 13280 50077 13308
rect 50019 13277 50031 13280
rect 49973 13271 50031 13277
rect 50065 13277 50077 13280
rect 50111 13308 50123 13311
rect 51810 13308 51816 13320
rect 50111 13280 51816 13308
rect 50111 13277 50123 13280
rect 50065 13271 50123 13277
rect 51810 13268 51816 13280
rect 51868 13268 51874 13320
rect 49326 13172 49332 13184
rect 45756 13144 49332 13172
rect 49326 13132 49332 13144
rect 49384 13132 49390 13184
rect 1104 13082 54832 13104
rect 1104 13030 9947 13082
rect 9999 13030 10011 13082
rect 10063 13030 10075 13082
rect 10127 13030 10139 13082
rect 10191 13030 27878 13082
rect 27930 13030 27942 13082
rect 27994 13030 28006 13082
rect 28058 13030 28070 13082
rect 28122 13030 45808 13082
rect 45860 13030 45872 13082
rect 45924 13030 45936 13082
rect 45988 13030 46000 13082
rect 46052 13030 54832 13082
rect 1104 13008 54832 13030
rect 2222 12968 2228 12980
rect 2183 12940 2228 12968
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 7098 12968 7104 12980
rect 7059 12940 7104 12968
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10410 12968 10416 12980
rect 9732 12940 10416 12968
rect 9732 12928 9738 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 11756 12940 13093 12968
rect 11756 12928 11762 12940
rect 13081 12937 13093 12940
rect 13127 12968 13139 12971
rect 13354 12968 13360 12980
rect 13127 12940 13360 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 14918 12968 14924 12980
rect 14879 12940 14924 12968
rect 14918 12928 14924 12940
rect 14976 12928 14982 12980
rect 16666 12968 16672 12980
rect 16627 12940 16672 12968
rect 16666 12928 16672 12940
rect 16724 12928 16730 12980
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 19797 12971 19855 12977
rect 19797 12968 19809 12971
rect 19576 12940 19809 12968
rect 19576 12928 19582 12940
rect 19797 12937 19809 12940
rect 19843 12937 19855 12971
rect 19797 12931 19855 12937
rect 21361 12971 21419 12977
rect 21361 12937 21373 12971
rect 21407 12968 21419 12971
rect 22738 12968 22744 12980
rect 21407 12940 22744 12968
rect 21407 12937 21419 12940
rect 21361 12931 21419 12937
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 25685 12971 25743 12977
rect 25685 12968 25697 12971
rect 23532 12940 25697 12968
rect 23532 12928 23538 12940
rect 25685 12937 25697 12940
rect 25731 12937 25743 12971
rect 25685 12931 25743 12937
rect 29086 12928 29092 12980
rect 29144 12968 29150 12980
rect 29641 12971 29699 12977
rect 29641 12968 29653 12971
rect 29144 12940 29653 12968
rect 29144 12928 29150 12940
rect 29641 12937 29653 12940
rect 29687 12937 29699 12971
rect 29641 12931 29699 12937
rect 30929 12971 30987 12977
rect 30929 12937 30941 12971
rect 30975 12968 30987 12971
rect 31386 12968 31392 12980
rect 30975 12940 31392 12968
rect 30975 12937 30987 12940
rect 30929 12931 30987 12937
rect 8294 12900 8300 12912
rect 7392 12872 8300 12900
rect 7392 12841 7420 12872
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 8849 12903 8907 12909
rect 8849 12869 8861 12903
rect 8895 12869 8907 12903
rect 8849 12863 8907 12869
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 8864 12832 8892 12863
rect 7377 12795 7435 12801
rect 7484 12804 8892 12832
rect 14936 12832 14964 12928
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 18785 12903 18843 12909
rect 18785 12900 18797 12903
rect 16540 12872 18797 12900
rect 16540 12860 16546 12872
rect 18785 12869 18797 12872
rect 18831 12869 18843 12903
rect 18785 12863 18843 12869
rect 19337 12903 19395 12909
rect 19337 12869 19349 12903
rect 19383 12900 19395 12903
rect 20257 12903 20315 12909
rect 20257 12900 20269 12903
rect 19383 12872 20269 12900
rect 19383 12869 19395 12872
rect 19337 12863 19395 12869
rect 20257 12869 20269 12872
rect 20303 12900 20315 12903
rect 25225 12903 25283 12909
rect 25225 12900 25237 12903
rect 20303 12872 25237 12900
rect 20303 12869 20315 12872
rect 20257 12863 20315 12869
rect 25225 12869 25237 12872
rect 25271 12900 25283 12903
rect 26050 12900 26056 12912
rect 25271 12872 26056 12900
rect 25271 12869 25283 12872
rect 25225 12863 25283 12869
rect 26050 12860 26056 12872
rect 26108 12860 26114 12912
rect 30944 12900 30972 12931
rect 31386 12928 31392 12940
rect 31444 12928 31450 12980
rect 34422 12928 34428 12980
rect 34480 12968 34486 12980
rect 41690 12968 41696 12980
rect 34480 12940 36952 12968
rect 41603 12940 41696 12968
rect 34480 12928 34486 12940
rect 30116 12872 30972 12900
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14936 12804 15117 12832
rect 2406 12773 2412 12776
rect 2401 12764 2412 12773
rect 2367 12736 2412 12764
rect 2401 12727 2412 12736
rect 2406 12724 2412 12727
rect 2464 12724 2470 12776
rect 3418 12764 3424 12776
rect 3379 12736 3424 12764
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 4430 12764 4436 12776
rect 4391 12736 4436 12764
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12764 5503 12767
rect 6178 12764 6184 12776
rect 5491 12736 6184 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 7484 12773 7512 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 25682 12792 25688 12844
rect 25740 12832 25746 12844
rect 30116 12841 30144 12872
rect 36446 12860 36452 12912
rect 36504 12900 36510 12912
rect 36817 12903 36875 12909
rect 36817 12900 36829 12903
rect 36504 12872 36829 12900
rect 36504 12860 36510 12872
rect 36817 12869 36829 12872
rect 36863 12869 36875 12903
rect 36817 12863 36875 12869
rect 30101 12835 30159 12841
rect 30101 12832 30113 12835
rect 25740 12804 30113 12832
rect 25740 12792 25746 12804
rect 30101 12801 30113 12804
rect 30147 12801 30159 12835
rect 33962 12832 33968 12844
rect 30101 12795 30159 12801
rect 30208 12804 33456 12832
rect 33923 12804 33968 12832
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 8018 12764 8024 12776
rect 7979 12736 8024 12764
rect 7837 12727 7895 12733
rect 7852 12696 7880 12727
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8904 12736 9045 12764
rect 8904 12724 8910 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 10318 12764 10324 12776
rect 10279 12736 10324 12764
rect 9033 12727 9091 12733
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 11514 12764 11520 12776
rect 11475 12736 11520 12764
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12764 13047 12767
rect 13170 12764 13176 12776
rect 13035 12736 13176 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 13170 12724 13176 12736
rect 13228 12764 13234 12776
rect 13538 12764 13544 12776
rect 13228 12736 13544 12764
rect 13228 12724 13234 12736
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14182 12764 14188 12776
rect 14143 12736 14188 12764
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 15381 12767 15439 12773
rect 15381 12733 15393 12767
rect 15427 12764 15439 12767
rect 16022 12764 16028 12776
rect 15427 12736 16028 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 16022 12724 16028 12736
rect 16080 12724 16086 12776
rect 17586 12724 17592 12776
rect 17644 12764 17650 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 17644 12736 18981 12764
rect 17644 12724 17650 12736
rect 18969 12733 18981 12736
rect 19015 12733 19027 12767
rect 19610 12764 19616 12776
rect 19571 12736 19616 12764
rect 18969 12727 19027 12733
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 21542 12764 21548 12776
rect 21600 12773 21606 12776
rect 21511 12736 21548 12764
rect 21542 12724 21548 12736
rect 21600 12727 21611 12773
rect 21600 12724 21606 12727
rect 22462 12724 22468 12776
rect 22520 12764 22526 12776
rect 22557 12767 22615 12773
rect 22557 12764 22569 12767
rect 22520 12736 22569 12764
rect 22520 12724 22526 12736
rect 22557 12733 22569 12736
rect 22603 12733 22615 12767
rect 24026 12764 24032 12776
rect 23987 12736 24032 12764
rect 22557 12727 22615 12733
rect 24026 12724 24032 12736
rect 24084 12724 24090 12776
rect 24946 12764 24952 12776
rect 24320 12736 24952 12764
rect 9950 12696 9956 12708
rect 7852 12668 9956 12696
rect 9950 12656 9956 12668
rect 10008 12656 10014 12708
rect 19521 12699 19579 12705
rect 19521 12665 19533 12699
rect 19567 12696 19579 12699
rect 19702 12696 19708 12708
rect 19567 12668 19708 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 19702 12656 19708 12668
rect 19760 12656 19766 12708
rect 23845 12699 23903 12705
rect 23845 12665 23857 12699
rect 23891 12696 23903 12699
rect 24320 12696 24348 12736
rect 24946 12724 24952 12736
rect 25004 12724 25010 12776
rect 25501 12767 25559 12773
rect 25501 12733 25513 12767
rect 25547 12764 25559 12767
rect 26418 12764 26424 12776
rect 25547 12736 26424 12764
rect 25547 12733 25559 12736
rect 25501 12727 25559 12733
rect 26418 12724 26424 12736
rect 26476 12724 26482 12776
rect 26786 12764 26792 12776
rect 26747 12736 26792 12764
rect 26786 12724 26792 12736
rect 26844 12724 26850 12776
rect 27246 12724 27252 12776
rect 27304 12764 27310 12776
rect 27985 12767 28043 12773
rect 27985 12764 27997 12767
rect 27304 12736 27997 12764
rect 27304 12724 27310 12736
rect 27985 12733 27997 12736
rect 28031 12733 28043 12767
rect 27985 12727 28043 12733
rect 28902 12724 28908 12776
rect 28960 12764 28966 12776
rect 30208 12773 30236 12804
rect 33428 12776 33456 12804
rect 33962 12792 33968 12804
rect 34020 12792 34026 12844
rect 34974 12792 34980 12844
rect 35032 12832 35038 12844
rect 35345 12835 35403 12841
rect 35345 12832 35357 12835
rect 35032 12804 35357 12832
rect 35032 12792 35038 12804
rect 35345 12801 35357 12804
rect 35391 12801 35403 12835
rect 36464 12832 36492 12860
rect 35345 12795 35403 12801
rect 35452 12804 36492 12832
rect 36924 12832 36952 12940
rect 41690 12928 41696 12940
rect 41748 12968 41754 12980
rect 44818 12968 44824 12980
rect 41748 12940 44824 12968
rect 41748 12928 41754 12940
rect 37645 12903 37703 12909
rect 37645 12869 37657 12903
rect 37691 12900 37703 12903
rect 37734 12900 37740 12912
rect 37691 12872 37740 12900
rect 37691 12869 37703 12872
rect 37645 12863 37703 12869
rect 37734 12860 37740 12872
rect 37792 12860 37798 12912
rect 39945 12903 40003 12909
rect 39040 12872 39896 12900
rect 39040 12832 39068 12872
rect 39666 12832 39672 12844
rect 36924 12804 39068 12832
rect 39132 12804 39672 12832
rect 30193 12767 30251 12773
rect 28960 12736 30144 12764
rect 28960 12724 28966 12736
rect 23891 12668 24348 12696
rect 24397 12699 24455 12705
rect 23891 12665 23903 12668
rect 23845 12659 23903 12665
rect 24397 12665 24409 12699
rect 24443 12696 24455 12699
rect 25130 12696 25136 12708
rect 24443 12668 25136 12696
rect 24443 12665 24455 12668
rect 24397 12659 24455 12665
rect 25130 12656 25136 12668
rect 25188 12696 25194 12708
rect 25409 12699 25467 12705
rect 25409 12696 25421 12699
rect 25188 12668 25421 12696
rect 25188 12656 25194 12668
rect 25409 12665 25421 12668
rect 25455 12665 25467 12699
rect 25409 12659 25467 12665
rect 27706 12656 27712 12708
rect 27764 12696 27770 12708
rect 27801 12699 27859 12705
rect 27801 12696 27813 12699
rect 27764 12668 27813 12696
rect 27764 12656 27770 12668
rect 27801 12665 27813 12668
rect 27847 12696 27859 12699
rect 28166 12696 28172 12708
rect 27847 12668 28172 12696
rect 27847 12665 27859 12668
rect 27801 12659 27859 12665
rect 28166 12656 28172 12668
rect 28224 12656 28230 12708
rect 28353 12699 28411 12705
rect 28353 12665 28365 12699
rect 28399 12696 28411 12699
rect 29454 12696 29460 12708
rect 28399 12668 29460 12696
rect 28399 12665 28411 12668
rect 28353 12659 28411 12665
rect 29454 12656 29460 12668
rect 29512 12656 29518 12708
rect 30116 12696 30144 12736
rect 30193 12733 30205 12767
rect 30239 12733 30251 12767
rect 30193 12727 30251 12733
rect 30561 12767 30619 12773
rect 30561 12733 30573 12767
rect 30607 12733 30619 12767
rect 30561 12727 30619 12733
rect 30745 12767 30803 12773
rect 30745 12733 30757 12767
rect 30791 12764 30803 12767
rect 31662 12764 31668 12776
rect 30791 12736 31668 12764
rect 30791 12733 30803 12736
rect 30745 12727 30803 12733
rect 30576 12696 30604 12727
rect 31662 12724 31668 12736
rect 31720 12764 31726 12776
rect 31757 12767 31815 12773
rect 31757 12764 31769 12767
rect 31720 12736 31769 12764
rect 31720 12724 31726 12736
rect 31757 12733 31769 12736
rect 31803 12733 31815 12767
rect 31757 12727 31815 12733
rect 31941 12767 31999 12773
rect 31941 12733 31953 12767
rect 31987 12764 31999 12767
rect 32398 12764 32404 12776
rect 31987 12736 32404 12764
rect 31987 12733 31999 12736
rect 31941 12727 31999 12733
rect 31956 12696 31984 12727
rect 32398 12724 32404 12736
rect 32456 12724 32462 12776
rect 33410 12764 33416 12776
rect 33323 12736 33416 12764
rect 33410 12724 33416 12736
rect 33468 12724 33474 12776
rect 33597 12767 33655 12773
rect 33597 12733 33609 12767
rect 33643 12733 33655 12767
rect 33597 12727 33655 12733
rect 35069 12767 35127 12773
rect 35069 12733 35081 12767
rect 35115 12764 35127 12767
rect 35452 12764 35480 12804
rect 39132 12776 39160 12804
rect 39666 12792 39672 12804
rect 39724 12792 39730 12844
rect 35115 12736 35480 12764
rect 35115 12733 35127 12736
rect 35069 12727 35127 12733
rect 30116 12668 31984 12696
rect 32309 12699 32367 12705
rect 32309 12665 32321 12699
rect 32355 12696 32367 12699
rect 33318 12696 33324 12708
rect 32355 12668 33324 12696
rect 32355 12665 32367 12668
rect 32309 12659 32367 12665
rect 33318 12656 33324 12668
rect 33376 12656 33382 12708
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 3237 12631 3295 12637
rect 3237 12628 3249 12631
rect 2464 12600 3249 12628
rect 2464 12588 2470 12600
rect 3237 12597 3249 12600
rect 3283 12597 3295 12631
rect 4246 12628 4252 12640
rect 4207 12600 4252 12628
rect 3237 12591 3295 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4982 12588 4988 12640
rect 5040 12628 5046 12640
rect 5261 12631 5319 12637
rect 5261 12628 5273 12631
rect 5040 12600 5273 12628
rect 5040 12588 5046 12600
rect 5261 12597 5273 12600
rect 5307 12597 5319 12631
rect 5261 12591 5319 12597
rect 11333 12631 11391 12637
rect 11333 12597 11345 12631
rect 11379 12628 11391 12631
rect 12986 12628 12992 12640
rect 11379 12600 12992 12628
rect 11379 12597 11391 12600
rect 11333 12591 11391 12597
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 13964 12600 14013 12628
rect 13964 12588 13970 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 14001 12591 14059 12597
rect 22373 12631 22431 12637
rect 22373 12597 22385 12631
rect 22419 12628 22431 12631
rect 23750 12628 23756 12640
rect 22419 12600 23756 12628
rect 22419 12597 22431 12600
rect 22373 12591 22431 12597
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 24026 12588 24032 12640
rect 24084 12628 24090 12640
rect 24670 12628 24676 12640
rect 24084 12600 24676 12628
rect 24084 12588 24090 12600
rect 24670 12588 24676 12600
rect 24728 12628 24734 12640
rect 26881 12631 26939 12637
rect 26881 12628 26893 12631
rect 24728 12600 26893 12628
rect 24728 12588 24734 12600
rect 26881 12597 26893 12600
rect 26927 12597 26939 12631
rect 33612 12628 33640 12727
rect 35986 12724 35992 12776
rect 36044 12764 36050 12776
rect 37553 12767 37611 12773
rect 37553 12764 37565 12767
rect 36044 12736 37565 12764
rect 36044 12724 36050 12736
rect 37553 12733 37565 12736
rect 37599 12733 37611 12767
rect 39114 12764 39120 12776
rect 39027 12736 39120 12764
rect 37553 12727 37611 12733
rect 39114 12724 39120 12736
rect 39172 12724 39178 12776
rect 39393 12767 39451 12773
rect 39393 12733 39405 12767
rect 39439 12733 39451 12767
rect 39868 12764 39896 12872
rect 39945 12869 39957 12903
rect 39991 12900 40003 12903
rect 40034 12900 40040 12912
rect 39991 12872 40040 12900
rect 39991 12869 40003 12872
rect 39945 12863 40003 12869
rect 40034 12860 40040 12872
rect 40092 12860 40098 12912
rect 40681 12767 40739 12773
rect 40681 12764 40693 12767
rect 39868 12736 40693 12764
rect 39393 12727 39451 12733
rect 40681 12733 40693 12736
rect 40727 12764 40739 12767
rect 41046 12764 41052 12776
rect 40727 12736 41052 12764
rect 40727 12733 40739 12736
rect 40681 12727 40739 12733
rect 34606 12628 34612 12640
rect 33612 12600 34612 12628
rect 26881 12591 26939 12597
rect 34606 12588 34612 12600
rect 34664 12628 34670 12640
rect 36449 12631 36507 12637
rect 36449 12628 36461 12631
rect 34664 12600 36461 12628
rect 34664 12588 34670 12600
rect 36449 12597 36461 12600
rect 36495 12597 36507 12631
rect 39408 12628 39436 12727
rect 41046 12724 41052 12736
rect 41104 12724 41110 12776
rect 41800 12773 41828 12940
rect 44818 12928 44824 12940
rect 44876 12928 44882 12980
rect 47854 12968 47860 12980
rect 47815 12940 47860 12968
rect 47854 12928 47860 12940
rect 47912 12928 47918 12980
rect 49326 12968 49332 12980
rect 49287 12940 49332 12968
rect 49326 12928 49332 12940
rect 49384 12928 49390 12980
rect 44082 12900 44088 12912
rect 44043 12872 44088 12900
rect 44082 12860 44088 12872
rect 44140 12860 44146 12912
rect 44450 12792 44456 12844
rect 44508 12832 44514 12844
rect 44821 12835 44879 12841
rect 44821 12832 44833 12835
rect 44508 12804 44833 12832
rect 44508 12792 44514 12804
rect 44821 12801 44833 12804
rect 44867 12832 44879 12835
rect 47118 12832 47124 12844
rect 44867 12804 47124 12832
rect 44867 12801 44879 12804
rect 44821 12795 44879 12801
rect 47118 12792 47124 12804
rect 47176 12792 47182 12844
rect 47872 12832 47900 12928
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47872 12804 47961 12832
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 48222 12832 48228 12844
rect 48183 12804 48228 12832
rect 47949 12795 48007 12801
rect 48222 12792 48228 12804
rect 48280 12792 48286 12844
rect 41785 12767 41843 12773
rect 41785 12733 41797 12767
rect 41831 12733 41843 12767
rect 41785 12727 41843 12733
rect 43717 12767 43775 12773
rect 43717 12733 43729 12767
rect 43763 12764 43775 12767
rect 43809 12767 43867 12773
rect 43809 12764 43821 12767
rect 43763 12736 43821 12764
rect 43763 12733 43775 12736
rect 43717 12727 43775 12733
rect 43809 12733 43821 12736
rect 43855 12733 43867 12767
rect 43809 12727 43867 12733
rect 39574 12696 39580 12708
rect 39535 12668 39580 12696
rect 39574 12656 39580 12668
rect 39632 12656 39638 12708
rect 39666 12656 39672 12708
rect 39724 12696 39730 12708
rect 39761 12699 39819 12705
rect 39761 12696 39773 12699
rect 39724 12668 39773 12696
rect 39724 12656 39730 12668
rect 39761 12665 39773 12668
rect 39807 12696 39819 12699
rect 43732 12696 43760 12727
rect 44266 12724 44272 12776
rect 44324 12764 44330 12776
rect 44361 12767 44419 12773
rect 44361 12764 44373 12767
rect 44324 12736 44373 12764
rect 44324 12724 44330 12736
rect 44361 12733 44373 12736
rect 44407 12733 44419 12767
rect 46566 12764 46572 12776
rect 46527 12736 46572 12764
rect 44361 12727 44419 12733
rect 46566 12724 46572 12736
rect 46624 12724 46630 12776
rect 46750 12764 46756 12776
rect 46711 12736 46756 12764
rect 46750 12724 46756 12736
rect 46808 12724 46814 12776
rect 39807 12668 43760 12696
rect 39807 12665 39819 12668
rect 39761 12659 39819 12665
rect 40034 12628 40040 12640
rect 39408 12600 40040 12628
rect 36449 12591 36507 12597
rect 40034 12588 40040 12600
rect 40092 12628 40098 12640
rect 40310 12628 40316 12640
rect 40092 12600 40316 12628
rect 40092 12588 40098 12600
rect 40310 12588 40316 12600
rect 40368 12588 40374 12640
rect 40880 12637 40908 12668
rect 40865 12631 40923 12637
rect 40865 12597 40877 12631
rect 40911 12597 40923 12631
rect 41966 12628 41972 12640
rect 41927 12600 41972 12628
rect 40865 12591 40923 12597
rect 41966 12588 41972 12600
rect 42024 12588 42030 12640
rect 1104 12538 54832 12560
rect 1104 12486 18912 12538
rect 18964 12486 18976 12538
rect 19028 12486 19040 12538
rect 19092 12486 19104 12538
rect 19156 12486 36843 12538
rect 36895 12486 36907 12538
rect 36959 12486 36971 12538
rect 37023 12486 37035 12538
rect 37087 12486 54832 12538
rect 1104 12464 54832 12486
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3418 12424 3424 12436
rect 2915 12396 3424 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 4801 12427 4859 12433
rect 4801 12393 4813 12427
rect 4847 12424 4859 12427
rect 4890 12424 4896 12436
rect 4847 12396 4896 12424
rect 4847 12393 4859 12396
rect 4801 12387 4859 12393
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 6178 12384 6184 12436
rect 6236 12424 6242 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 6236 12396 7849 12424
rect 6236 12384 6242 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 9950 12424 9956 12436
rect 9911 12396 9956 12424
rect 7837 12387 7895 12393
rect 9950 12384 9956 12396
rect 10008 12424 10014 12436
rect 10594 12424 10600 12436
rect 10008 12396 10600 12424
rect 10008 12384 10014 12396
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 19702 12424 19708 12436
rect 18800 12396 19708 12424
rect 13817 12359 13875 12365
rect 13817 12356 13829 12359
rect 10704 12328 12388 12356
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3234 12288 3240 12300
rect 3099 12260 3240 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 3234 12248 3240 12260
rect 3292 12248 3298 12300
rect 4982 12288 4988 12300
rect 4943 12260 4988 12288
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12288 6055 12291
rect 6914 12288 6920 12300
rect 6043 12260 6920 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 7558 12288 7564 12300
rect 7055 12260 7564 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 10704 12297 10732 12328
rect 9033 12291 9091 12297
rect 9033 12288 9045 12291
rect 8628 12260 9045 12288
rect 8628 12248 8634 12260
rect 9033 12257 9045 12260
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10689 12291 10747 12297
rect 10367 12260 10548 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 5813 12087 5871 12093
rect 5813 12084 5825 12087
rect 5592 12056 5825 12084
rect 5592 12044 5598 12056
rect 5813 12053 5825 12056
rect 5859 12053 5871 12087
rect 6822 12084 6828 12096
rect 6783 12056 6828 12084
rect 5813 12047 5871 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 8849 12087 8907 12093
rect 8849 12084 8861 12087
rect 7984 12056 8861 12084
rect 7984 12044 7990 12056
rect 8849 12053 8861 12056
rect 8895 12053 8907 12087
rect 10520 12084 10548 12260
rect 10689 12257 10701 12291
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10870 12220 10876 12232
rect 10643 12192 10876 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 12360 12220 12388 12328
rect 13096 12328 13829 12356
rect 13096 12297 13124 12328
rect 13817 12325 13829 12328
rect 13863 12356 13875 12359
rect 13863 12328 16804 12356
rect 13863 12325 13875 12328
rect 13817 12319 13875 12325
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12257 13139 12291
rect 13081 12251 13139 12257
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 15654 12288 15660 12300
rect 13495 12260 15660 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 16209 12291 16267 12297
rect 16209 12257 16221 12291
rect 16255 12288 16267 12291
rect 16574 12288 16580 12300
rect 16255 12260 16580 12288
rect 16255 12257 16267 12260
rect 16209 12251 16267 12257
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 13170 12220 13176 12232
rect 12360 12192 12756 12220
rect 13131 12192 13176 12220
rect 12728 12161 12756 12192
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 13354 12220 13360 12232
rect 13315 12192 13360 12220
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 12713 12155 12771 12161
rect 12713 12121 12725 12155
rect 12759 12152 12771 12155
rect 15286 12152 15292 12164
rect 12759 12124 15292 12152
rect 12759 12121 12771 12124
rect 12713 12115 12771 12121
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 16574 12152 16580 12164
rect 16535 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 13906 12084 13912 12096
rect 10520 12056 13912 12084
rect 8849 12047 8907 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 14700 12056 16037 12084
rect 14700 12044 14706 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16684 12084 16712 12251
rect 16776 12152 16804 12328
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17494 12288 17500 12300
rect 17407 12260 17500 12288
rect 17494 12248 17500 12260
rect 17552 12288 17558 12300
rect 18800 12288 18828 12396
rect 19702 12384 19708 12396
rect 19760 12424 19766 12436
rect 21177 12427 21235 12433
rect 21177 12424 21189 12427
rect 19760 12396 21189 12424
rect 19760 12384 19766 12396
rect 21177 12393 21189 12396
rect 21223 12393 21235 12427
rect 21177 12387 21235 12393
rect 26418 12384 26424 12436
rect 26476 12424 26482 12436
rect 26789 12427 26847 12433
rect 26789 12424 26801 12427
rect 26476 12396 26801 12424
rect 26476 12384 26482 12396
rect 26789 12393 26801 12396
rect 26835 12393 26847 12427
rect 29086 12424 29092 12436
rect 28999 12396 29092 12424
rect 26789 12387 26847 12393
rect 29086 12384 29092 12396
rect 29144 12424 29150 12436
rect 30742 12424 30748 12436
rect 29144 12396 30748 12424
rect 29144 12384 29150 12396
rect 30742 12384 30748 12396
rect 30800 12384 30806 12436
rect 34241 12427 34299 12433
rect 34241 12424 34253 12427
rect 30852 12396 34253 12424
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 20901 12359 20959 12365
rect 20901 12356 20913 12359
rect 19392 12328 20913 12356
rect 19392 12316 19398 12328
rect 19444 12297 19472 12328
rect 20901 12325 20913 12328
rect 20947 12356 20959 12359
rect 20990 12356 20996 12368
rect 20947 12328 20996 12356
rect 20947 12325 20959 12328
rect 20901 12319 20959 12325
rect 20990 12316 20996 12328
rect 21048 12316 21054 12368
rect 25038 12316 25044 12368
rect 25096 12356 25102 12368
rect 26513 12359 26571 12365
rect 26513 12356 26525 12359
rect 25096 12328 26525 12356
rect 25096 12316 25102 12328
rect 26513 12325 26525 12328
rect 26559 12325 26571 12359
rect 26513 12319 26571 12325
rect 28353 12359 28411 12365
rect 28353 12325 28365 12359
rect 28399 12356 28411 12359
rect 30098 12356 30104 12368
rect 28399 12328 30104 12356
rect 28399 12325 28411 12328
rect 28353 12319 28411 12325
rect 30098 12316 30104 12328
rect 30156 12316 30162 12368
rect 17552 12260 18828 12288
rect 19429 12291 19487 12297
rect 17552 12248 17558 12260
rect 19429 12257 19441 12291
rect 19475 12257 19487 12291
rect 19610 12288 19616 12300
rect 19571 12260 19616 12288
rect 19429 12251 19487 12257
rect 19610 12248 19616 12260
rect 19668 12248 19674 12300
rect 19794 12288 19800 12300
rect 19755 12260 19800 12288
rect 19794 12248 19800 12260
rect 19852 12288 19858 12300
rect 21082 12288 21088 12300
rect 19852 12260 21088 12288
rect 19852 12248 19858 12260
rect 21082 12248 21088 12260
rect 21140 12248 21146 12300
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 23474 12288 23480 12300
rect 22603 12260 23480 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 25130 12288 25136 12300
rect 25091 12260 25136 12288
rect 25130 12248 25136 12260
rect 25188 12248 25194 12300
rect 25406 12248 25412 12300
rect 25464 12288 25470 12300
rect 25593 12291 25651 12297
rect 25593 12288 25605 12291
rect 25464 12260 25605 12288
rect 25464 12248 25470 12260
rect 25593 12257 25605 12260
rect 25639 12288 25651 12291
rect 26234 12288 26240 12300
rect 25639 12260 26240 12288
rect 25639 12257 25651 12260
rect 25593 12251 25651 12257
rect 26234 12248 26240 12260
rect 26292 12248 26298 12300
rect 26697 12291 26755 12297
rect 26697 12257 26709 12291
rect 26743 12288 26755 12291
rect 26786 12288 26792 12300
rect 26743 12260 26792 12288
rect 26743 12257 26755 12260
rect 26697 12251 26755 12257
rect 22002 12180 22008 12232
rect 22060 12220 22066 12232
rect 22189 12223 22247 12229
rect 22189 12220 22201 12223
rect 22060 12192 22201 12220
rect 22060 12180 22066 12192
rect 22189 12189 22201 12192
rect 22235 12220 22247 12223
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22235 12192 22293 12220
rect 22235 12189 22247 12192
rect 22189 12183 22247 12189
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12220 23903 12223
rect 26712 12220 26740 12251
rect 26786 12248 26792 12260
rect 26844 12248 26850 12300
rect 28258 12248 28264 12300
rect 28316 12288 28322 12300
rect 28445 12291 28503 12297
rect 28445 12288 28457 12291
rect 28316 12260 28457 12288
rect 28316 12248 28322 12260
rect 28445 12257 28457 12260
rect 28491 12257 28503 12291
rect 30466 12288 30472 12300
rect 30427 12260 30472 12288
rect 28445 12251 28503 12257
rect 30466 12248 30472 12260
rect 30524 12248 30530 12300
rect 23891 12192 26740 12220
rect 23891 12189 23903 12192
rect 23845 12183 23903 12189
rect 29454 12180 29460 12232
rect 29512 12220 29518 12232
rect 30852 12229 30880 12396
rect 34241 12393 34253 12396
rect 34287 12424 34299 12427
rect 34698 12424 34704 12436
rect 34287 12396 34704 12424
rect 34287 12393 34299 12396
rect 34241 12387 34299 12393
rect 34698 12384 34704 12396
rect 34756 12384 34762 12436
rect 40310 12384 40316 12436
rect 40368 12424 40374 12436
rect 40773 12427 40831 12433
rect 40773 12424 40785 12427
rect 40368 12396 40785 12424
rect 40368 12384 40374 12396
rect 40773 12393 40785 12396
rect 40819 12393 40831 12427
rect 40773 12387 40831 12393
rect 40862 12384 40868 12436
rect 40920 12424 40926 12436
rect 41233 12427 41291 12433
rect 41233 12424 41245 12427
rect 40920 12396 41245 12424
rect 40920 12384 40926 12396
rect 41233 12393 41245 12396
rect 41279 12424 41291 12427
rect 43070 12424 43076 12436
rect 41279 12396 43076 12424
rect 41279 12393 41291 12396
rect 41233 12387 41291 12393
rect 43070 12384 43076 12396
rect 43128 12384 43134 12436
rect 44726 12424 44732 12436
rect 44687 12396 44732 12424
rect 44726 12384 44732 12396
rect 44784 12384 44790 12436
rect 31205 12359 31263 12365
rect 31205 12325 31217 12359
rect 31251 12356 31263 12359
rect 31662 12356 31668 12368
rect 31251 12328 31668 12356
rect 31251 12325 31263 12328
rect 31205 12319 31263 12325
rect 31662 12316 31668 12328
rect 31720 12316 31726 12368
rect 32968 12328 35112 12356
rect 32582 12248 32588 12300
rect 32640 12288 32646 12300
rect 32968 12297 32996 12328
rect 35084 12300 35112 12328
rect 32953 12291 33011 12297
rect 32953 12288 32965 12291
rect 32640 12260 32965 12288
rect 32640 12248 32646 12260
rect 32953 12257 32965 12260
rect 32999 12257 33011 12291
rect 32953 12251 33011 12257
rect 34149 12291 34207 12297
rect 34149 12257 34161 12291
rect 34195 12288 34207 12291
rect 34330 12288 34336 12300
rect 34195 12260 34336 12288
rect 34195 12257 34207 12260
rect 34149 12251 34207 12257
rect 34330 12248 34336 12260
rect 34388 12288 34394 12300
rect 34425 12291 34483 12297
rect 34425 12288 34437 12291
rect 34388 12260 34437 12288
rect 34388 12248 34394 12260
rect 34425 12257 34437 12260
rect 34471 12257 34483 12291
rect 34425 12251 34483 12257
rect 35066 12248 35072 12300
rect 35124 12288 35130 12300
rect 35345 12291 35403 12297
rect 35345 12288 35357 12291
rect 35124 12260 35357 12288
rect 35124 12248 35130 12260
rect 35345 12257 35357 12260
rect 35391 12257 35403 12291
rect 35345 12251 35403 12257
rect 35434 12248 35440 12300
rect 35492 12288 35498 12300
rect 39393 12291 39451 12297
rect 35492 12260 35537 12288
rect 35492 12248 35498 12260
rect 39393 12257 39405 12291
rect 39439 12288 39451 12291
rect 40880 12288 40908 12384
rect 39439 12260 40908 12288
rect 43088 12288 43116 12384
rect 43349 12291 43407 12297
rect 43349 12288 43361 12291
rect 43088 12260 43361 12288
rect 39439 12257 39451 12260
rect 39393 12251 39451 12257
rect 43349 12257 43361 12260
rect 43395 12257 43407 12291
rect 43622 12288 43628 12300
rect 43583 12260 43628 12288
rect 43349 12251 43407 12257
rect 43622 12248 43628 12260
rect 43680 12248 43686 12300
rect 30616 12223 30674 12229
rect 30616 12220 30628 12223
rect 29512 12192 30628 12220
rect 29512 12180 29518 12192
rect 30616 12189 30628 12192
rect 30662 12189 30674 12223
rect 30616 12183 30674 12189
rect 30837 12223 30895 12229
rect 30837 12189 30849 12223
rect 30883 12189 30895 12223
rect 30837 12183 30895 12189
rect 31110 12180 31116 12232
rect 31168 12220 31174 12232
rect 32125 12223 32183 12229
rect 32125 12220 32137 12223
rect 31168 12192 32137 12220
rect 31168 12180 31174 12192
rect 32125 12189 32137 12192
rect 32171 12189 32183 12223
rect 32674 12220 32680 12232
rect 32635 12192 32680 12220
rect 32125 12183 32183 12189
rect 32674 12180 32680 12192
rect 32732 12180 32738 12232
rect 32766 12180 32772 12232
rect 32824 12229 32830 12232
rect 32824 12223 32873 12229
rect 32824 12189 32827 12223
rect 32861 12189 32873 12223
rect 32824 12183 32873 12189
rect 32824 12180 32830 12183
rect 39574 12180 39580 12232
rect 39632 12220 39638 12232
rect 39669 12223 39727 12229
rect 39669 12220 39681 12223
rect 39632 12192 39681 12220
rect 39632 12180 39638 12192
rect 39669 12189 39681 12192
rect 39715 12189 39727 12223
rect 39669 12183 39727 12189
rect 16776 12124 22324 12152
rect 17773 12087 17831 12093
rect 17773 12084 17785 12087
rect 16684 12056 17785 12084
rect 16025 12047 16083 12053
rect 17773 12053 17785 12056
rect 17819 12084 17831 12087
rect 18874 12084 18880 12096
rect 17819 12056 18880 12084
rect 17819 12053 17831 12056
rect 17773 12047 17831 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 22296 12084 22324 12124
rect 26050 12112 26056 12164
rect 26108 12152 26114 12164
rect 28169 12155 28227 12161
rect 28169 12152 28181 12155
rect 26108 12124 28181 12152
rect 26108 12112 26114 12124
rect 28169 12121 28181 12124
rect 28215 12152 28227 12155
rect 29086 12152 29092 12164
rect 28215 12124 29092 12152
rect 28215 12121 28227 12124
rect 28169 12115 28227 12121
rect 29086 12112 29092 12124
rect 29144 12112 29150 12164
rect 30745 12155 30803 12161
rect 30745 12121 30757 12155
rect 30791 12152 30803 12155
rect 30791 12124 30880 12152
rect 30791 12121 30803 12124
rect 30745 12115 30803 12121
rect 23934 12084 23940 12096
rect 22296 12056 23940 12084
rect 23934 12044 23940 12056
rect 23992 12044 23998 12096
rect 24946 12084 24952 12096
rect 24907 12056 24952 12084
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 28442 12044 28448 12096
rect 28500 12084 28506 12096
rect 28629 12087 28687 12093
rect 28629 12084 28641 12087
rect 28500 12056 28641 12084
rect 28500 12044 28506 12056
rect 28629 12053 28641 12056
rect 28675 12053 28687 12087
rect 30852 12084 30880 12124
rect 30926 12112 30932 12164
rect 30984 12152 30990 12164
rect 35161 12155 35219 12161
rect 35161 12152 35173 12155
rect 30984 12124 35173 12152
rect 30984 12112 30990 12124
rect 35161 12121 35173 12124
rect 35207 12152 35219 12155
rect 35207 12124 36124 12152
rect 35207 12121 35219 12124
rect 35161 12115 35219 12121
rect 32766 12084 32772 12096
rect 30852 12056 32772 12084
rect 28629 12047 28687 12053
rect 32766 12044 32772 12056
rect 32824 12044 32830 12096
rect 35618 12084 35624 12096
rect 35579 12056 35624 12084
rect 35618 12044 35624 12056
rect 35676 12044 35682 12096
rect 36096 12093 36124 12124
rect 36081 12087 36139 12093
rect 36081 12053 36093 12087
rect 36127 12084 36139 12087
rect 41966 12084 41972 12096
rect 36127 12056 41972 12084
rect 36127 12053 36139 12056
rect 36081 12047 36139 12053
rect 41966 12044 41972 12056
rect 42024 12044 42030 12096
rect 1104 11994 54832 12016
rect 1104 11942 9947 11994
rect 9999 11942 10011 11994
rect 10063 11942 10075 11994
rect 10127 11942 10139 11994
rect 10191 11942 27878 11994
rect 27930 11942 27942 11994
rect 27994 11942 28006 11994
rect 28058 11942 28070 11994
rect 28122 11942 45808 11994
rect 45860 11942 45872 11994
rect 45924 11942 45936 11994
rect 45988 11942 46000 11994
rect 46052 11942 54832 11994
rect 1104 11920 54832 11942
rect 2133 11883 2191 11889
rect 2133 11849 2145 11883
rect 2179 11880 2191 11883
rect 4522 11880 4528 11892
rect 2179 11852 4528 11880
rect 2179 11849 2191 11852
rect 2133 11843 2191 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 7558 11880 7564 11892
rect 7519 11852 7564 11880
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 8570 11880 8576 11892
rect 8531 11852 8576 11880
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14185 11883 14243 11889
rect 14185 11880 14197 11883
rect 13872 11852 14197 11880
rect 13872 11840 13878 11852
rect 14185 11849 14197 11852
rect 14231 11849 14243 11883
rect 15194 11880 15200 11892
rect 15155 11852 15200 11880
rect 14185 11843 14243 11849
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 17586 11880 17592 11892
rect 15344 11852 17592 11880
rect 15344 11840 15350 11852
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 17678 11840 17684 11892
rect 17736 11880 17742 11892
rect 18785 11883 18843 11889
rect 18785 11880 18797 11883
rect 17736 11852 18797 11880
rect 17736 11840 17742 11852
rect 18785 11849 18797 11852
rect 18831 11849 18843 11883
rect 18785 11843 18843 11849
rect 18874 11840 18880 11892
rect 18932 11880 18938 11892
rect 30006 11880 30012 11892
rect 18932 11852 25728 11880
rect 29967 11852 30012 11880
rect 18932 11840 18938 11852
rect 11609 11815 11667 11821
rect 11609 11781 11621 11815
rect 11655 11812 11667 11815
rect 13906 11812 13912 11824
rect 11655 11784 13912 11812
rect 11655 11781 11667 11784
rect 11609 11775 11667 11781
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 22002 11812 22008 11824
rect 20772 11784 22008 11812
rect 20772 11772 20778 11784
rect 22002 11772 22008 11784
rect 22060 11812 22066 11824
rect 24305 11815 24363 11821
rect 24305 11812 24317 11815
rect 22060 11784 24317 11812
rect 22060 11772 22066 11784
rect 24305 11781 24317 11784
rect 24351 11812 24363 11815
rect 25700 11812 25728 11852
rect 30006 11840 30012 11852
rect 30064 11840 30070 11892
rect 30116 11852 32904 11880
rect 30116 11812 30144 11852
rect 24351 11784 24532 11812
rect 25700 11784 30144 11812
rect 31021 11815 31079 11821
rect 24351 11781 24363 11784
rect 24305 11775 24363 11781
rect 6822 11744 6828 11756
rect 3528 11716 6828 11744
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 3528 11685 3556 11716
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 16022 11744 16028 11756
rect 15983 11716 16028 11744
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16574 11744 16580 11756
rect 16535 11716 16580 11744
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17126 11744 17132 11756
rect 17083 11716 17132 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 19153 11747 19211 11753
rect 19153 11713 19165 11747
rect 19199 11744 19211 11747
rect 19245 11747 19303 11753
rect 19245 11744 19257 11747
rect 19199 11716 19257 11744
rect 19199 11713 19211 11716
rect 19153 11707 19211 11713
rect 19245 11713 19257 11716
rect 19291 11713 19303 11747
rect 19518 11744 19524 11756
rect 19479 11716 19524 11744
rect 19245 11707 19303 11713
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 2188 11648 2329 11676
rect 2188 11636 2194 11648
rect 2317 11645 2329 11648
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11645 3571 11679
rect 4522 11676 4528 11688
rect 4483 11648 4528 11676
rect 3513 11639 3571 11645
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 5534 11676 5540 11688
rect 5495 11648 5540 11676
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 7745 11679 7803 11685
rect 7745 11645 7757 11679
rect 7791 11676 7803 11679
rect 7926 11676 7932 11688
rect 7791 11648 7932 11676
rect 7791 11645 7803 11648
rect 7745 11639 7803 11645
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 8754 11676 8760 11688
rect 8715 11648 8760 11676
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 9766 11676 9772 11688
rect 9727 11648 9772 11676
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 10778 11676 10784 11688
rect 10739 11648 10784 11676
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11480 11648 11805 11676
rect 11480 11636 11486 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 13446 11676 13452 11688
rect 13403 11648 13452 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 14332 11648 14381 11676
rect 14332 11636 14338 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 15378 11676 15384 11688
rect 15339 11648 15384 11676
rect 14369 11639 14427 11645
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11676 16911 11679
rect 17494 11676 17500 11688
rect 16899 11648 17500 11676
rect 16899 11645 16911 11648
rect 16853 11639 16911 11645
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18012 11648 18981 11676
rect 18012 11636 18018 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 19260 11676 19288 11707
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 24504 11753 24532 11784
rect 31021 11781 31033 11815
rect 31067 11781 31079 11815
rect 31021 11775 31079 11781
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 20714 11676 20720 11688
rect 19260 11648 20720 11676
rect 18969 11639 19027 11645
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 21910 11676 21916 11688
rect 21871 11648 21916 11676
rect 21910 11636 21916 11648
rect 21968 11636 21974 11688
rect 24762 11676 24768 11688
rect 24723 11648 24768 11676
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 25130 11636 25136 11688
rect 25188 11676 25194 11688
rect 25188 11648 25452 11676
rect 25188 11636 25194 11648
rect 20898 11608 20904 11620
rect 20859 11580 20904 11608
rect 20898 11568 20904 11580
rect 20956 11568 20962 11620
rect 21634 11568 21640 11620
rect 21692 11608 21698 11620
rect 25424 11608 25452 11648
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 27157 11679 27215 11685
rect 27157 11676 27169 11679
rect 26292 11648 27169 11676
rect 26292 11636 26298 11648
rect 27157 11645 27169 11648
rect 27203 11676 27215 11679
rect 27246 11676 27252 11688
rect 27203 11648 27252 11676
rect 27203 11645 27215 11648
rect 27157 11639 27215 11645
rect 27246 11636 27252 11648
rect 27304 11636 27310 11688
rect 30193 11679 30251 11685
rect 30193 11645 30205 11679
rect 30239 11676 30251 11679
rect 31036 11676 31064 11775
rect 31202 11676 31208 11688
rect 30239 11648 31064 11676
rect 31163 11648 31208 11676
rect 30239 11645 30251 11648
rect 30193 11639 30251 11645
rect 31202 11636 31208 11648
rect 31260 11636 31266 11688
rect 31588 11685 31616 11852
rect 31849 11815 31907 11821
rect 31849 11781 31861 11815
rect 31895 11812 31907 11815
rect 32674 11812 32680 11824
rect 31895 11784 32680 11812
rect 31895 11781 31907 11784
rect 31849 11775 31907 11781
rect 32674 11772 32680 11784
rect 32732 11772 32738 11824
rect 32876 11821 32904 11852
rect 33410 11840 33416 11892
rect 33468 11880 33474 11892
rect 33597 11883 33655 11889
rect 33597 11880 33609 11883
rect 33468 11852 33609 11880
rect 33468 11840 33474 11852
rect 33597 11849 33609 11852
rect 33643 11849 33655 11883
rect 33597 11843 33655 11849
rect 34440 11852 35572 11880
rect 32861 11815 32919 11821
rect 32861 11781 32873 11815
rect 32907 11812 32919 11815
rect 34440 11812 34468 11852
rect 35434 11812 35440 11824
rect 32907 11784 34468 11812
rect 35268 11784 35440 11812
rect 32907 11781 32919 11784
rect 32861 11775 32919 11781
rect 32766 11744 32772 11756
rect 32324 11716 32772 11744
rect 32324 11685 32352 11716
rect 32766 11704 32772 11716
rect 32824 11704 32830 11756
rect 35268 11753 35296 11784
rect 35434 11772 35440 11784
rect 35492 11772 35498 11824
rect 35544 11812 35572 11852
rect 36446 11840 36452 11892
rect 36504 11880 36510 11892
rect 36814 11880 36820 11892
rect 36504 11852 36820 11880
rect 36504 11840 36510 11852
rect 36814 11840 36820 11852
rect 36872 11840 36878 11892
rect 39114 11880 39120 11892
rect 36924 11852 39120 11880
rect 36924 11812 36952 11852
rect 39114 11840 39120 11852
rect 39172 11840 39178 11892
rect 35544 11784 36952 11812
rect 35253 11747 35311 11753
rect 35253 11713 35265 11747
rect 35299 11713 35311 11747
rect 35253 11707 35311 11713
rect 36814 11704 36820 11756
rect 36872 11744 36878 11756
rect 37001 11747 37059 11753
rect 37001 11744 37013 11747
rect 36872 11716 37013 11744
rect 36872 11704 36878 11716
rect 37001 11713 37013 11716
rect 37047 11713 37059 11747
rect 37001 11707 37059 11713
rect 31573 11679 31631 11685
rect 31573 11645 31585 11679
rect 31619 11645 31631 11679
rect 31573 11639 31631 11645
rect 32309 11679 32367 11685
rect 32309 11645 32321 11679
rect 32355 11645 32367 11679
rect 32582 11676 32588 11688
rect 32543 11648 32588 11676
rect 32309 11639 32367 11645
rect 32582 11636 32588 11648
rect 32640 11636 32646 11688
rect 33318 11636 33324 11688
rect 33376 11676 33382 11688
rect 33505 11679 33563 11685
rect 33505 11676 33517 11679
rect 33376 11648 33517 11676
rect 33376 11636 33382 11648
rect 33505 11645 33517 11648
rect 33551 11645 33563 11679
rect 33505 11639 33563 11645
rect 34606 11636 34612 11688
rect 34664 11676 34670 11688
rect 34885 11679 34943 11685
rect 34885 11676 34897 11679
rect 34664 11648 34897 11676
rect 34664 11636 34670 11648
rect 34885 11645 34897 11648
rect 34931 11645 34943 11679
rect 34885 11639 34943 11645
rect 35437 11679 35495 11685
rect 35437 11645 35449 11679
rect 35483 11645 35495 11679
rect 35437 11639 35495 11645
rect 26973 11611 27031 11617
rect 26973 11608 26985 11611
rect 21692 11580 24403 11608
rect 25424 11580 26985 11608
rect 21692 11568 21698 11580
rect 3326 11540 3332 11552
rect 3287 11512 3332 11540
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 4341 11543 4399 11549
rect 4341 11509 4353 11543
rect 4387 11540 4399 11543
rect 5258 11540 5264 11552
rect 4387 11512 5264 11540
rect 4387 11509 4399 11512
rect 4341 11503 4399 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5353 11543 5411 11549
rect 5353 11509 5365 11543
rect 5399 11540 5411 11543
rect 7006 11540 7012 11552
rect 5399 11512 7012 11540
rect 5399 11509 5411 11512
rect 5353 11503 5411 11509
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9088 11512 9597 11540
rect 9088 11500 9094 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 9732 11512 10609 11540
rect 9732 11500 9738 11512
rect 10597 11509 10609 11512
rect 10643 11509 10655 11543
rect 10597 11503 10655 11509
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 14366 11540 14372 11552
rect 13219 11512 14372 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 21726 11540 21732 11552
rect 21687 11512 21732 11540
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 24375 11540 24403 11580
rect 26973 11577 26985 11580
rect 27019 11608 27031 11611
rect 30466 11608 30472 11620
rect 27019 11580 30472 11608
rect 27019 11577 27031 11580
rect 26973 11571 27031 11577
rect 30466 11568 30472 11580
rect 30524 11568 30530 11620
rect 34698 11568 34704 11620
rect 34756 11608 34762 11620
rect 35452 11608 35480 11639
rect 35618 11636 35624 11688
rect 35676 11676 35682 11688
rect 37277 11679 37335 11685
rect 37277 11676 37289 11679
rect 35676 11648 37289 11676
rect 35676 11636 35682 11648
rect 37277 11645 37289 11648
rect 37323 11645 37335 11679
rect 37277 11639 37335 11645
rect 34756 11580 35480 11608
rect 34756 11568 34762 11580
rect 25590 11540 25596 11552
rect 24375 11512 25596 11540
rect 25590 11500 25596 11512
rect 25648 11540 25654 11552
rect 25869 11543 25927 11549
rect 25869 11540 25881 11543
rect 25648 11512 25881 11540
rect 25648 11500 25654 11512
rect 25869 11509 25881 11512
rect 25915 11509 25927 11543
rect 27246 11540 27252 11552
rect 27207 11512 27252 11540
rect 25869 11503 25927 11509
rect 27246 11500 27252 11512
rect 27304 11500 27310 11552
rect 34330 11500 34336 11552
rect 34388 11540 34394 11552
rect 38381 11543 38439 11549
rect 38381 11540 38393 11543
rect 34388 11512 38393 11540
rect 34388 11500 34394 11512
rect 38381 11509 38393 11512
rect 38427 11509 38439 11543
rect 38381 11503 38439 11509
rect 1104 11450 54832 11472
rect 1104 11398 18912 11450
rect 18964 11398 18976 11450
rect 19028 11398 19040 11450
rect 19092 11398 19104 11450
rect 19156 11398 36843 11450
rect 36895 11398 36907 11450
rect 36959 11398 36971 11450
rect 37023 11398 37035 11450
rect 37087 11398 54832 11450
rect 1104 11376 54832 11398
rect 2130 11336 2136 11348
rect 2091 11308 2136 11336
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 4580 11308 6837 11336
rect 4580 11296 4586 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 6972 11308 7849 11336
rect 6972 11296 6978 11308
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 8846 11336 8852 11348
rect 8807 11308 8852 11336
rect 7837 11299 7895 11305
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 11422 11336 11428 11348
rect 11383 11308 11428 11336
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 13446 11336 13452 11348
rect 13407 11308 13452 11336
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 20993 11339 21051 11345
rect 20993 11305 21005 11339
rect 21039 11336 21051 11339
rect 21082 11336 21088 11348
rect 21039 11308 21088 11336
rect 21039 11305 21051 11308
rect 20993 11299 21051 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 24688 11308 25636 11336
rect 3326 11228 3332 11280
rect 3384 11268 3390 11280
rect 3384 11240 8064 11268
rect 3384 11228 3390 11240
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 4246 11200 4252 11212
rect 2363 11172 4252 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5000 11132 5028 11163
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5316 11172 6009 11200
rect 5316 11160 5322 11172
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 7006 11200 7012 11212
rect 6967 11172 7012 11200
rect 5997 11163 6055 11169
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 8036 11209 8064 11240
rect 13998 11228 14004 11280
rect 14056 11268 14062 11280
rect 14056 11240 19288 11268
rect 14056 11228 14062 11240
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 9030 11200 9036 11212
rect 8991 11172 9036 11200
rect 8021 11163 8079 11169
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 11422 11200 11428 11212
rect 10643 11172 11428 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 12526 11200 12532 11212
rect 11655 11172 12532 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 6178 11132 6184 11144
rect 5000 11104 6184 11132
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 12636 11132 12664 11163
rect 12986 11160 12992 11212
rect 13044 11200 13050 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 13044 11172 13645 11200
rect 13044 11160 13050 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 17126 11200 17132 11212
rect 16255 11172 17132 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17221 11203 17279 11209
rect 17221 11169 17233 11203
rect 17267 11200 17279 11203
rect 18046 11200 18052 11212
rect 17267 11172 18052 11200
rect 17267 11169 17279 11172
rect 17221 11163 17279 11169
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 18230 11200 18236 11212
rect 18191 11172 18236 11200
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 19260 11209 19288 11240
rect 19245 11203 19303 11209
rect 19245 11169 19257 11203
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 20070 11160 20076 11212
rect 20128 11200 20134 11212
rect 20257 11203 20315 11209
rect 20257 11200 20269 11203
rect 20128 11172 20269 11200
rect 20128 11160 20134 11172
rect 20257 11169 20269 11172
rect 20303 11169 20315 11203
rect 20898 11200 20904 11212
rect 20859 11172 20904 11200
rect 20257 11163 20315 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 22094 11160 22100 11212
rect 22152 11200 22158 11212
rect 22152 11172 22197 11200
rect 22152 11160 22158 11172
rect 22370 11160 22376 11212
rect 22428 11200 22434 11212
rect 23109 11203 23167 11209
rect 23109 11200 23121 11203
rect 22428 11172 23121 11200
rect 22428 11160 22434 11172
rect 23109 11169 23121 11172
rect 23155 11169 23167 11203
rect 24118 11200 24124 11212
rect 24079 11172 24124 11200
rect 23109 11163 23167 11169
rect 24118 11160 24124 11172
rect 24176 11160 24182 11212
rect 24688 11209 24716 11308
rect 24762 11228 24768 11280
rect 24820 11268 24826 11280
rect 25608 11277 25636 11308
rect 25682 11296 25688 11348
rect 25740 11336 25746 11348
rect 27249 11339 27307 11345
rect 27249 11336 27261 11339
rect 25740 11308 27261 11336
rect 25740 11296 25746 11308
rect 27249 11305 27261 11308
rect 27295 11305 27307 11339
rect 27249 11299 27307 11305
rect 32217 11339 32275 11345
rect 32217 11305 32229 11339
rect 32263 11336 32275 11339
rect 32766 11336 32772 11348
rect 32263 11308 32772 11336
rect 32263 11305 32275 11308
rect 32217 11299 32275 11305
rect 32766 11296 32772 11308
rect 32824 11296 32830 11348
rect 33318 11336 33324 11348
rect 33152 11308 33324 11336
rect 25409 11271 25467 11277
rect 25409 11268 25421 11271
rect 24820 11240 25421 11268
rect 24820 11228 24826 11240
rect 25409 11237 25421 11240
rect 25455 11237 25467 11271
rect 25409 11231 25467 11237
rect 25593 11271 25651 11277
rect 25593 11237 25605 11271
rect 25639 11268 25651 11271
rect 26050 11268 26056 11280
rect 25639 11240 26056 11268
rect 25639 11237 25651 11240
rect 25593 11231 25651 11237
rect 26050 11228 26056 11240
rect 26108 11228 26114 11280
rect 29549 11271 29607 11277
rect 29549 11268 29561 11271
rect 28000 11240 29561 11268
rect 24673 11203 24731 11209
rect 24673 11169 24685 11203
rect 24719 11169 24731 11203
rect 24673 11163 24731 11169
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 14182 11132 14188 11144
rect 12636 11104 14188 11132
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 24872 11132 24900 11163
rect 24946 11160 24952 11212
rect 25004 11200 25010 11212
rect 27430 11200 27436 11212
rect 25004 11172 25049 11200
rect 27391 11172 27436 11200
rect 25004 11160 25010 11172
rect 27430 11160 27436 11172
rect 27488 11160 27494 11212
rect 28000 11209 28028 11240
rect 29549 11237 29561 11240
rect 29595 11237 29607 11271
rect 30098 11268 30104 11280
rect 30059 11240 30104 11268
rect 29549 11231 29607 11237
rect 30098 11228 30104 11240
rect 30156 11228 30162 11280
rect 33152 11277 33180 11308
rect 33318 11296 33324 11308
rect 33376 11296 33382 11348
rect 34514 11336 34520 11348
rect 33704 11308 34520 11336
rect 33704 11277 33732 11308
rect 34514 11296 34520 11308
rect 34572 11296 34578 11348
rect 33137 11271 33195 11277
rect 33137 11237 33149 11271
rect 33183 11237 33195 11271
rect 33137 11231 33195 11237
rect 33689 11271 33747 11277
rect 33689 11237 33701 11271
rect 33735 11237 33747 11271
rect 35066 11268 35072 11280
rect 35027 11240 35072 11268
rect 33689 11231 33747 11237
rect 35066 11228 35072 11240
rect 35124 11228 35130 11280
rect 27985 11203 28043 11209
rect 27985 11169 27997 11203
rect 28031 11169 28043 11203
rect 27985 11163 28043 11169
rect 27246 11132 27252 11144
rect 24872 11104 27252 11132
rect 27246 11092 27252 11104
rect 27304 11132 27310 11144
rect 28000 11132 28028 11163
rect 28258 11160 28264 11212
rect 28316 11200 28322 11212
rect 28353 11203 28411 11209
rect 28353 11200 28365 11203
rect 28316 11172 28365 11200
rect 28316 11160 28322 11172
rect 28353 11169 28365 11172
rect 28399 11169 28411 11203
rect 28353 11163 28411 11169
rect 28537 11203 28595 11209
rect 28537 11169 28549 11203
rect 28583 11200 28595 11203
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 28583 11172 29745 11200
rect 28583 11169 28595 11172
rect 28537 11163 28595 11169
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 27304 11104 28028 11132
rect 27304 11092 27310 11104
rect 28166 11092 28172 11144
rect 28224 11132 28230 11144
rect 28552 11132 28580 11163
rect 28224 11104 28580 11132
rect 30116 11132 30144 11228
rect 32125 11203 32183 11209
rect 32125 11169 32137 11203
rect 32171 11200 32183 11203
rect 32214 11200 32220 11212
rect 32171 11172 32220 11200
rect 32171 11169 32183 11172
rect 32125 11163 32183 11169
rect 32214 11160 32220 11172
rect 32272 11160 32278 11212
rect 33226 11160 33232 11212
rect 33284 11200 33290 11212
rect 33321 11203 33379 11209
rect 33321 11200 33333 11203
rect 33284 11172 33333 11200
rect 33284 11160 33290 11172
rect 33321 11169 33333 11172
rect 33367 11169 33379 11203
rect 33321 11163 33379 11169
rect 34517 11203 34575 11209
rect 34517 11169 34529 11203
rect 34563 11200 34575 11203
rect 34606 11200 34612 11212
rect 34563 11172 34612 11200
rect 34563 11169 34575 11172
rect 34517 11163 34575 11169
rect 34532 11132 34560 11163
rect 34606 11160 34612 11172
rect 34664 11160 34670 11212
rect 34698 11160 34704 11212
rect 34756 11200 34762 11212
rect 34756 11172 34801 11200
rect 34756 11160 34762 11172
rect 30116 11104 34560 11132
rect 28224 11092 28230 11104
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 4801 11067 4859 11073
rect 4801 11064 4813 11067
rect 4672 11036 4813 11064
rect 4672 11024 4678 11036
rect 4801 11033 4813 11036
rect 4847 11033 4859 11067
rect 4801 11027 4859 11033
rect 10413 11067 10471 11073
rect 10413 11033 10425 11067
rect 10459 11064 10471 11067
rect 13630 11064 13636 11076
rect 10459 11036 13636 11064
rect 10459 11033 10471 11036
rect 10413 11027 10471 11033
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 15378 11024 15384 11076
rect 15436 11064 15442 11076
rect 16025 11067 16083 11073
rect 16025 11064 16037 11067
rect 15436 11036 16037 11064
rect 15436 11024 15442 11036
rect 16025 11033 16037 11036
rect 16071 11033 16083 11067
rect 16025 11027 16083 11033
rect 18414 11024 18420 11076
rect 18472 11064 18478 11076
rect 19061 11067 19119 11073
rect 19061 11064 19073 11067
rect 18472 11036 19073 11064
rect 18472 11024 18478 11036
rect 19061 11033 19073 11036
rect 19107 11033 19119 11067
rect 19061 11027 19119 11033
rect 21913 11067 21971 11073
rect 21913 11033 21925 11067
rect 21959 11064 21971 11067
rect 22554 11064 22560 11076
rect 21959 11036 22560 11064
rect 21959 11033 21971 11036
rect 21913 11027 21971 11033
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 22925 11067 22983 11073
rect 22925 11033 22937 11067
rect 22971 11064 22983 11067
rect 23014 11064 23020 11076
rect 22971 11036 23020 11064
rect 22971 11033 22983 11036
rect 22925 11027 22983 11033
rect 23014 11024 23020 11036
rect 23072 11024 23078 11076
rect 5813 10999 5871 11005
rect 5813 10965 5825 10999
rect 5859 10996 5871 10999
rect 6362 10996 6368 11008
rect 5859 10968 6368 10996
rect 5859 10965 5871 10968
rect 5813 10959 5871 10965
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 12437 10999 12495 11005
rect 12437 10965 12449 10999
rect 12483 10996 12495 10999
rect 13722 10996 13728 11008
rect 12483 10968 13728 10996
rect 12483 10965 12495 10968
rect 12437 10959 12495 10965
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 17037 10999 17095 11005
rect 17037 10965 17049 10999
rect 17083 10996 17095 10999
rect 17402 10996 17408 11008
rect 17083 10968 17408 10996
rect 17083 10965 17095 10968
rect 17037 10959 17095 10965
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 18049 10999 18107 11005
rect 18049 10965 18061 10999
rect 18095 10996 18107 10999
rect 18966 10996 18972 11008
rect 18095 10968 18972 10996
rect 18095 10965 18107 10968
rect 18049 10959 18107 10965
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 20073 10999 20131 11005
rect 20073 10996 20085 10999
rect 20036 10968 20085 10996
rect 20036 10956 20042 10968
rect 20073 10965 20085 10968
rect 20119 10965 20131 10999
rect 23934 10996 23940 11008
rect 23895 10968 23940 10996
rect 20073 10959 20131 10965
rect 23934 10956 23940 10968
rect 23992 10956 23998 11008
rect 1104 10906 54832 10928
rect 1104 10854 9947 10906
rect 9999 10854 10011 10906
rect 10063 10854 10075 10906
rect 10127 10854 10139 10906
rect 10191 10854 27878 10906
rect 27930 10854 27942 10906
rect 27994 10854 28006 10906
rect 28058 10854 28070 10906
rect 28122 10854 45808 10906
rect 45860 10854 45872 10906
rect 45924 10854 45936 10906
rect 45988 10854 46000 10906
rect 46052 10854 54832 10906
rect 1104 10832 54832 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 4430 10792 4436 10804
rect 2179 10764 4436 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 4430 10752 4436 10764
rect 4488 10752 4494 10804
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 8573 10795 8631 10801
rect 8573 10761 8585 10795
rect 8619 10792 8631 10795
rect 9766 10792 9772 10804
rect 8619 10764 9772 10792
rect 8619 10761 8631 10764
rect 8573 10755 8631 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 11422 10792 11428 10804
rect 11383 10764 11428 10792
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12584 10764 13185 10792
rect 12584 10752 12590 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 14182 10792 14188 10804
rect 14143 10764 14188 10792
rect 13173 10755 13231 10761
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 17184 10764 17233 10792
rect 17184 10752 17190 10764
rect 17221 10761 17233 10764
rect 17267 10761 17279 10795
rect 17221 10755 17279 10761
rect 21542 10752 21548 10804
rect 21600 10792 21606 10804
rect 25222 10792 25228 10804
rect 21600 10764 25228 10792
rect 21600 10752 21606 10764
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 25685 10795 25743 10801
rect 25685 10761 25697 10795
rect 25731 10792 25743 10795
rect 26234 10792 26240 10804
rect 25731 10764 26240 10792
rect 25731 10761 25743 10764
rect 25685 10755 25743 10761
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 32125 10795 32183 10801
rect 32125 10761 32137 10795
rect 32171 10792 32183 10795
rect 32214 10792 32220 10804
rect 32171 10764 32220 10792
rect 32171 10761 32183 10764
rect 32125 10755 32183 10761
rect 32214 10752 32220 10764
rect 32272 10752 32278 10804
rect 32585 10795 32643 10801
rect 32585 10761 32597 10795
rect 32631 10792 32643 10795
rect 32950 10792 32956 10804
rect 32631 10764 32956 10792
rect 32631 10761 32643 10764
rect 32585 10755 32643 10761
rect 16666 10684 16672 10736
rect 16724 10724 16730 10736
rect 18785 10727 18843 10733
rect 18785 10724 18797 10727
rect 16724 10696 18797 10724
rect 16724 10684 16730 10696
rect 18785 10693 18797 10696
rect 18831 10693 18843 10727
rect 18785 10687 18843 10693
rect 21821 10727 21879 10733
rect 21821 10693 21833 10727
rect 21867 10693 21879 10727
rect 21821 10687 21879 10693
rect 2314 10588 2320 10600
rect 2275 10560 2320 10588
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 3326 10588 3332 10600
rect 3287 10560 3332 10588
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 4338 10588 4344 10600
rect 4299 10560 4344 10588
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 5350 10588 5356 10600
rect 5311 10560 5356 10588
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 6362 10588 6368 10600
rect 6323 10560 6368 10588
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 9674 10588 9680 10600
rect 8803 10560 9680 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 7760 10520 7788 10551
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10588 10655 10591
rect 11514 10588 11520 10600
rect 10643 10560 11520 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11609 10591 11667 10597
rect 11609 10557 11621 10591
rect 11655 10588 11667 10591
rect 12526 10588 12532 10600
rect 11655 10560 12532 10588
rect 11655 10557 11667 10560
rect 11609 10551 11667 10557
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13538 10588 13544 10600
rect 13403 10560 13544 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13538 10548 13544 10560
rect 13596 10548 13602 10600
rect 14366 10588 14372 10600
rect 14327 10560 14372 10588
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10588 15439 10591
rect 16022 10588 16028 10600
rect 15427 10560 16028 10588
rect 15427 10557 15439 10560
rect 15381 10551 15439 10557
rect 16022 10548 16028 10560
rect 16080 10548 16086 10600
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 17034 10588 17040 10600
rect 16439 10560 17040 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 17402 10588 17408 10600
rect 17363 10560 17408 10588
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 18966 10588 18972 10600
rect 18927 10560 18972 10588
rect 18966 10548 18972 10560
rect 19024 10548 19030 10600
rect 19978 10588 19984 10600
rect 19939 10560 19984 10588
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10588 21051 10591
rect 21836 10588 21864 10687
rect 30745 10659 30803 10665
rect 30745 10625 30757 10659
rect 30791 10656 30803 10659
rect 32600 10656 32628 10755
rect 32950 10752 32956 10764
rect 33008 10752 33014 10804
rect 30791 10628 32628 10656
rect 30791 10625 30803 10628
rect 30745 10619 30803 10625
rect 22002 10588 22008 10600
rect 21039 10560 21864 10588
rect 21963 10560 22008 10588
rect 21039 10557 21051 10560
rect 20993 10551 21051 10557
rect 22002 10548 22008 10560
rect 22060 10548 22066 10600
rect 22554 10548 22560 10600
rect 22612 10588 22618 10600
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22612 10560 23029 10588
rect 22612 10548 22618 10560
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 23934 10548 23940 10600
rect 23992 10588 23998 10600
rect 24765 10591 24823 10597
rect 24765 10588 24777 10591
rect 23992 10560 24777 10588
rect 23992 10548 23998 10560
rect 24765 10557 24777 10560
rect 24811 10557 24823 10591
rect 25590 10588 25596 10600
rect 25551 10560 25596 10588
rect 24765 10551 24823 10557
rect 25590 10548 25596 10560
rect 25648 10548 25654 10600
rect 27433 10591 27491 10597
rect 27433 10557 27445 10591
rect 27479 10588 27491 10591
rect 29270 10588 29276 10600
rect 27479 10560 29276 10588
rect 27479 10557 27491 10560
rect 27433 10551 27491 10557
rect 29270 10548 29276 10560
rect 29328 10548 29334 10600
rect 29362 10548 29368 10600
rect 29420 10588 29426 10600
rect 30193 10591 30251 10597
rect 30193 10588 30205 10591
rect 29420 10560 30205 10588
rect 29420 10548 29426 10560
rect 30193 10557 30205 10560
rect 30239 10557 30251 10591
rect 30193 10551 30251 10557
rect 31021 10591 31079 10597
rect 31021 10557 31033 10591
rect 31067 10588 31079 10591
rect 31110 10588 31116 10600
rect 31067 10560 31116 10588
rect 31067 10557 31079 10560
rect 31021 10551 31079 10557
rect 31110 10548 31116 10560
rect 31168 10548 31174 10600
rect 34514 10548 34520 10600
rect 34572 10588 34578 10600
rect 35805 10591 35863 10597
rect 35805 10588 35817 10591
rect 34572 10560 35817 10588
rect 34572 10548 34578 10560
rect 35805 10557 35817 10560
rect 35851 10557 35863 10591
rect 35805 10551 35863 10557
rect 3160 10492 7788 10520
rect 3160 10461 3188 10492
rect 3145 10455 3203 10461
rect 3145 10421 3157 10455
rect 3191 10421 3203 10455
rect 3145 10415 3203 10421
rect 3234 10412 3240 10464
rect 3292 10452 3298 10464
rect 4157 10455 4215 10461
rect 4157 10452 4169 10455
rect 3292 10424 4169 10452
rect 3292 10412 3298 10424
rect 4157 10421 4169 10424
rect 4203 10421 4215 10455
rect 5166 10452 5172 10464
rect 5127 10424 5172 10452
rect 4157 10415 4215 10421
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 7561 10455 7619 10461
rect 7561 10452 7573 10455
rect 5592 10424 7573 10452
rect 5592 10412 5598 10424
rect 7561 10421 7573 10424
rect 7607 10421 7619 10455
rect 7561 10415 7619 10421
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 10413 10455 10471 10461
rect 10413 10452 10425 10455
rect 9548 10424 10425 10452
rect 9548 10412 9554 10424
rect 10413 10421 10425 10424
rect 10459 10421 10471 10455
rect 10413 10415 10471 10421
rect 15197 10455 15255 10461
rect 15197 10421 15209 10455
rect 15243 10452 15255 10455
rect 16114 10452 16120 10464
rect 15243 10424 16120 10452
rect 15243 10421 15255 10424
rect 15197 10415 15255 10421
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16209 10455 16267 10461
rect 16209 10421 16221 10455
rect 16255 10452 16267 10455
rect 17402 10452 17408 10464
rect 16255 10424 17408 10452
rect 16255 10421 16267 10424
rect 16209 10415 16267 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19797 10455 19855 10461
rect 19797 10452 19809 10455
rect 19484 10424 19809 10452
rect 19484 10412 19490 10424
rect 19797 10421 19809 10424
rect 19843 10421 19855 10455
rect 19797 10415 19855 10421
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 20312 10424 20821 10452
rect 20312 10412 20318 10424
rect 20809 10421 20821 10424
rect 20855 10421 20867 10455
rect 20809 10415 20867 10421
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22833 10455 22891 10461
rect 22833 10452 22845 10455
rect 21876 10424 22845 10452
rect 21876 10412 21882 10424
rect 22833 10421 22845 10424
rect 22879 10421 22891 10455
rect 22833 10415 22891 10421
rect 24302 10412 24308 10464
rect 24360 10452 24366 10464
rect 24581 10455 24639 10461
rect 24581 10452 24593 10455
rect 24360 10424 24593 10452
rect 24360 10412 24366 10424
rect 24581 10421 24593 10424
rect 24627 10421 24639 10455
rect 27246 10452 27252 10464
rect 27207 10424 27252 10452
rect 24581 10415 24639 10421
rect 27246 10412 27252 10424
rect 27304 10412 27310 10464
rect 28994 10412 29000 10464
rect 29052 10452 29058 10464
rect 30009 10455 30067 10461
rect 30009 10452 30021 10455
rect 29052 10424 30021 10452
rect 29052 10412 29058 10424
rect 30009 10421 30021 10424
rect 30055 10421 30067 10455
rect 30009 10415 30067 10421
rect 35621 10455 35679 10461
rect 35621 10421 35633 10455
rect 35667 10452 35679 10455
rect 37182 10452 37188 10464
rect 35667 10424 37188 10452
rect 35667 10421 35679 10424
rect 35621 10415 35679 10421
rect 37182 10412 37188 10424
rect 37240 10412 37246 10464
rect 1104 10362 54832 10384
rect 1104 10310 18912 10362
rect 18964 10310 18976 10362
rect 19028 10310 19040 10362
rect 19092 10310 19104 10362
rect 19156 10310 36843 10362
rect 36895 10310 36907 10362
rect 36959 10310 36971 10362
rect 37023 10310 37035 10362
rect 37087 10310 54832 10362
rect 1104 10288 54832 10310
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 3326 10248 3332 10260
rect 2271 10220 3332 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7282 10248 7288 10260
rect 7055 10220 7288 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10217 8079 10251
rect 11514 10248 11520 10260
rect 11475 10220 11520 10248
rect 8021 10211 8079 10217
rect 2409 10115 2467 10121
rect 2409 10081 2421 10115
rect 2455 10112 2467 10115
rect 3234 10112 3240 10124
rect 2455 10084 3240 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 4798 10112 4804 10124
rect 3467 10084 4804 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 5994 10112 6000 10124
rect 5031 10084 5856 10112
rect 5955 10084 6000 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 5828 9985 5856 10084
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 8036 10112 8064 10211
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 12526 10248 12532 10260
rect 12487 10220 12532 10248
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 13538 10248 13544 10260
rect 13499 10220 13544 10248
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 16022 10248 16028 10260
rect 15983 10220 16028 10248
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 17034 10248 17040 10260
rect 16995 10220 17040 10248
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 18046 10248 18052 10260
rect 18007 10220 18052 10248
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 20070 10248 20076 10260
rect 20031 10220 20076 10248
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 21637 10251 21695 10257
rect 21637 10217 21649 10251
rect 21683 10248 21695 10251
rect 22002 10248 22008 10260
rect 21683 10220 22008 10248
rect 21683 10217 21695 10220
rect 21637 10211 21695 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 22649 10251 22707 10257
rect 22649 10248 22661 10251
rect 22152 10220 22661 10248
rect 22152 10208 22158 10220
rect 22649 10217 22661 10220
rect 22695 10217 22707 10251
rect 22649 10211 22707 10217
rect 25409 10251 25467 10257
rect 25409 10217 25421 10251
rect 25455 10248 25467 10251
rect 27430 10248 27436 10260
rect 25455 10220 27436 10248
rect 25455 10217 25467 10220
rect 25409 10211 25467 10217
rect 27430 10208 27436 10220
rect 27488 10208 27494 10260
rect 29270 10248 29276 10260
rect 29231 10220 29276 10248
rect 29270 10208 29276 10220
rect 29328 10208 29334 10260
rect 8202 10112 8208 10124
rect 7239 10084 8064 10112
rect 8163 10084 8208 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 9490 10112 9496 10124
rect 9451 10084 9496 10112
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10081 10747 10115
rect 10689 10075 10747 10081
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10112 11759 10115
rect 12618 10112 12624 10124
rect 11747 10084 12624 10112
rect 11747 10081 11759 10084
rect 11701 10075 11759 10081
rect 10704 10044 10732 10075
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10081 12771 10115
rect 13722 10112 13728 10124
rect 13683 10084 13728 10112
rect 12713 10075 12771 10081
rect 9324 10016 10732 10044
rect 12728 10044 12756 10075
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 16209 10115 16267 10121
rect 16209 10081 16221 10115
rect 16255 10112 16267 10115
rect 17126 10112 17132 10124
rect 16255 10084 17132 10112
rect 16255 10081 16267 10084
rect 16209 10075 16267 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 17276 10084 17321 10112
rect 17276 10072 17282 10084
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18104 10084 18245 10112
rect 18104 10072 18110 10084
rect 18233 10081 18245 10084
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 19245 10115 19303 10121
rect 19245 10081 19257 10115
rect 19291 10112 19303 10115
rect 20070 10112 20076 10124
rect 19291 10084 20076 10112
rect 19291 10081 19303 10084
rect 19245 10075 19303 10081
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 20254 10112 20260 10124
rect 20215 10084 20260 10112
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 21818 10112 21824 10124
rect 21779 10084 21824 10112
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 22830 10112 22836 10124
rect 22791 10084 22836 10112
rect 22830 10072 22836 10084
rect 22888 10072 22894 10124
rect 24210 10072 24216 10124
rect 24268 10112 24274 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 24268 10084 24593 10112
rect 24268 10072 24274 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 25590 10112 25596 10124
rect 25551 10084 25596 10112
rect 24581 10075 24639 10081
rect 25590 10072 25596 10084
rect 25648 10072 25654 10124
rect 27430 10112 27436 10124
rect 27391 10084 27436 10112
rect 27430 10072 27436 10084
rect 27488 10072 27494 10124
rect 27522 10072 27528 10124
rect 27580 10112 27586 10124
rect 28445 10115 28503 10121
rect 28445 10112 28457 10115
rect 27580 10084 28457 10112
rect 27580 10072 27586 10084
rect 28445 10081 28457 10084
rect 28491 10081 28503 10115
rect 29454 10112 29460 10124
rect 29415 10084 29460 10112
rect 28445 10075 28503 10081
rect 29454 10072 29460 10084
rect 29512 10072 29518 10124
rect 29546 10072 29552 10124
rect 29604 10112 29610 10124
rect 30469 10115 30527 10121
rect 30469 10112 30481 10115
rect 29604 10084 30481 10112
rect 29604 10072 29610 10084
rect 30469 10081 30481 10084
rect 30515 10081 30527 10115
rect 30469 10075 30527 10081
rect 32858 10072 32864 10124
rect 32916 10112 32922 10124
rect 33229 10115 33287 10121
rect 33229 10112 33241 10115
rect 32916 10084 33241 10112
rect 32916 10072 32922 10084
rect 33229 10081 33241 10084
rect 33275 10081 33287 10115
rect 34238 10112 34244 10124
rect 34199 10084 34244 10112
rect 33229 10075 33287 10081
rect 34238 10072 34244 10084
rect 34296 10072 34302 10124
rect 35253 10115 35311 10121
rect 35253 10081 35265 10115
rect 35299 10112 35311 10115
rect 36170 10112 36176 10124
rect 35299 10084 36176 10112
rect 35299 10081 35311 10084
rect 35253 10075 35311 10081
rect 36170 10072 36176 10084
rect 36228 10072 36234 10124
rect 36265 10115 36323 10121
rect 36265 10081 36277 10115
rect 36311 10112 36323 10115
rect 37642 10112 37648 10124
rect 36311 10084 37648 10112
rect 36311 10081 36323 10084
rect 36265 10075 36323 10081
rect 37642 10072 37648 10084
rect 37700 10072 37706 10124
rect 14182 10044 14188 10056
rect 12728 10016 14188 10044
rect 9324 9985 9352 10016
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 5813 9979 5871 9985
rect 5813 9945 5825 9979
rect 5859 9945 5871 9979
rect 5813 9939 5871 9945
rect 9309 9979 9367 9985
rect 9309 9945 9321 9979
rect 9355 9945 9367 9979
rect 9309 9939 9367 9945
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4801 9911 4859 9917
rect 4801 9908 4813 9911
rect 4212 9880 4813 9908
rect 4212 9868 4218 9880
rect 4801 9877 4813 9880
rect 4847 9877 4859 9911
rect 4801 9871 4859 9877
rect 10505 9911 10563 9917
rect 10505 9877 10517 9911
rect 10551 9908 10563 9911
rect 11422 9908 11428 9920
rect 10551 9880 11428 9908
rect 10551 9877 10563 9880
rect 10505 9871 10563 9877
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 19061 9911 19119 9917
rect 19061 9877 19073 9911
rect 19107 9908 19119 9911
rect 20622 9908 20628 9920
rect 19107 9880 20628 9908
rect 19107 9877 19119 9880
rect 19061 9871 19119 9877
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 24397 9911 24455 9917
rect 24397 9877 24409 9911
rect 24443 9908 24455 9911
rect 24578 9908 24584 9920
rect 24443 9880 24584 9908
rect 24443 9877 24455 9880
rect 24397 9871 24455 9877
rect 24578 9868 24584 9880
rect 24636 9868 24642 9920
rect 26234 9868 26240 9920
rect 26292 9908 26298 9920
rect 27249 9911 27307 9917
rect 27249 9908 27261 9911
rect 26292 9880 27261 9908
rect 26292 9868 26298 9880
rect 27249 9877 27261 9880
rect 27295 9877 27307 9911
rect 27249 9871 27307 9877
rect 27614 9868 27620 9920
rect 27672 9908 27678 9920
rect 28261 9911 28319 9917
rect 28261 9908 28273 9911
rect 27672 9880 28273 9908
rect 27672 9868 27678 9880
rect 28261 9877 28273 9880
rect 28307 9877 28319 9911
rect 28261 9871 28319 9877
rect 30285 9911 30343 9917
rect 30285 9877 30297 9911
rect 30331 9908 30343 9911
rect 30742 9908 30748 9920
rect 30331 9880 30748 9908
rect 30331 9877 30343 9880
rect 30285 9871 30343 9877
rect 30742 9868 30748 9880
rect 30800 9868 30806 9920
rect 32950 9868 32956 9920
rect 33008 9908 33014 9920
rect 33045 9911 33103 9917
rect 33045 9908 33057 9911
rect 33008 9880 33057 9908
rect 33008 9868 33014 9880
rect 33045 9877 33057 9880
rect 33091 9877 33103 9911
rect 33045 9871 33103 9877
rect 33318 9868 33324 9920
rect 33376 9908 33382 9920
rect 34057 9911 34115 9917
rect 34057 9908 34069 9911
rect 33376 9880 34069 9908
rect 33376 9868 33382 9880
rect 34057 9877 34069 9880
rect 34103 9877 34115 9911
rect 34057 9871 34115 9877
rect 35069 9911 35127 9917
rect 35069 9877 35081 9911
rect 35115 9908 35127 9911
rect 35986 9908 35992 9920
rect 35115 9880 35992 9908
rect 35115 9877 35127 9880
rect 35069 9871 35127 9877
rect 35986 9868 35992 9880
rect 36044 9868 36050 9920
rect 36081 9911 36139 9917
rect 36081 9877 36093 9911
rect 36127 9908 36139 9911
rect 36814 9908 36820 9920
rect 36127 9880 36820 9908
rect 36127 9877 36139 9880
rect 36081 9871 36139 9877
rect 36814 9868 36820 9880
rect 36872 9868 36878 9920
rect 1104 9818 54832 9840
rect 1104 9766 9947 9818
rect 9999 9766 10011 9818
rect 10063 9766 10075 9818
rect 10127 9766 10139 9818
rect 10191 9766 27878 9818
rect 27930 9766 27942 9818
rect 27994 9766 28006 9818
rect 28058 9766 28070 9818
rect 28122 9766 45808 9818
rect 45860 9766 45872 9818
rect 45924 9766 45936 9818
rect 45988 9766 46000 9818
rect 46052 9766 54832 9818
rect 1104 9744 54832 9766
rect 5350 9704 5356 9716
rect 4356 9676 5356 9704
rect 3421 9639 3479 9645
rect 3421 9605 3433 9639
rect 3467 9636 3479 9639
rect 4356 9636 4384 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 7561 9707 7619 9713
rect 7561 9673 7573 9707
rect 7607 9704 7619 9707
rect 8202 9704 8208 9716
rect 7607 9676 8208 9704
rect 7607 9673 7619 9676
rect 7561 9667 7619 9673
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 12676 9676 13185 9704
rect 12676 9664 12682 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 27430 9704 27436 9716
rect 27391 9676 27436 9704
rect 13173 9667 13231 9673
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 3467 9608 4384 9636
rect 4433 9639 4491 9645
rect 3467 9605 3479 9608
rect 3421 9599 3479 9605
rect 4433 9605 4445 9639
rect 4479 9636 4491 9639
rect 5994 9636 6000 9648
rect 4479 9608 6000 9636
rect 4479 9605 4491 9608
rect 4433 9599 4491 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 14182 9636 14188 9648
rect 14143 9608 14188 9636
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 17126 9596 17132 9648
rect 17184 9636 17190 9648
rect 17221 9639 17279 9645
rect 17221 9636 17233 9639
rect 17184 9608 17233 9636
rect 17184 9596 17190 9608
rect 17221 9605 17233 9608
rect 17267 9605 17279 9639
rect 17221 9599 17279 9605
rect 21821 9639 21879 9645
rect 21821 9605 21833 9639
rect 21867 9636 21879 9639
rect 22830 9636 22836 9648
rect 21867 9608 22836 9636
rect 21867 9605 21879 9608
rect 21821 9599 21879 9605
rect 22830 9596 22836 9608
rect 22888 9596 22894 9648
rect 24397 9639 24455 9645
rect 24397 9605 24409 9639
rect 24443 9636 24455 9639
rect 25590 9636 25596 9648
rect 24443 9608 25596 9636
rect 24443 9605 24455 9608
rect 24397 9599 24455 9605
rect 25590 9596 25596 9608
rect 25648 9596 25654 9648
rect 28905 9639 28963 9645
rect 28905 9605 28917 9639
rect 28951 9636 28963 9639
rect 29546 9636 29552 9648
rect 28951 9608 29552 9636
rect 28951 9605 28963 9608
rect 28905 9599 28963 9605
rect 29546 9596 29552 9608
rect 29604 9596 29610 9648
rect 32769 9639 32827 9645
rect 32769 9605 32781 9639
rect 32815 9636 32827 9639
rect 34238 9636 34244 9648
rect 32815 9608 34244 9636
rect 32815 9605 32827 9608
rect 32769 9599 32827 9605
rect 34238 9596 34244 9608
rect 34296 9596 34302 9648
rect 36170 9596 36176 9648
rect 36228 9636 36234 9648
rect 36633 9639 36691 9645
rect 36633 9636 36645 9639
rect 36228 9608 36645 9636
rect 36228 9596 36234 9608
rect 36633 9605 36645 9608
rect 36679 9605 36691 9639
rect 37642 9636 37648 9648
rect 37603 9608 37648 9636
rect 36633 9599 36691 9605
rect 37642 9596 37648 9608
rect 37700 9596 37706 9648
rect 5166 9568 5172 9580
rect 2608 9540 5172 9568
rect 2608 9509 2636 9540
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9469 2651 9503
rect 2593 9463 2651 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 4154 9500 4160 9512
rect 3651 9472 4160 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4614 9500 4620 9512
rect 4575 9472 4620 9500
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5905 9503 5963 9509
rect 5905 9500 5917 9503
rect 5500 9472 5917 9500
rect 5500 9460 5506 9472
rect 5905 9469 5917 9472
rect 5951 9469 5963 9503
rect 5905 9463 5963 9469
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7524 9472 7757 9500
rect 7524 9460 7530 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 8754 9500 8760 9512
rect 8715 9472 8760 9500
rect 7745 9463 7803 9469
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9500 10747 9503
rect 12434 9500 12440 9512
rect 10735 9472 12440 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 13446 9500 13452 9512
rect 13403 9472 13452 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 13964 9472 14381 9500
rect 13964 9460 13970 9472
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9500 15439 9503
rect 16022 9500 16028 9512
rect 15427 9472 16028 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 16114 9460 16120 9512
rect 16172 9500 16178 9512
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 16172 9472 16405 9500
rect 16172 9460 16178 9472
rect 16393 9469 16405 9472
rect 16439 9469 16451 9503
rect 17402 9500 17408 9512
rect 17363 9472 17408 9500
rect 16393 9463 16451 9469
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9469 19027 9503
rect 19978 9500 19984 9512
rect 19939 9472 19984 9500
rect 18969 9463 19027 9469
rect 10778 9432 10784 9444
rect 5736 9404 10784 9432
rect 2409 9367 2467 9373
rect 2409 9333 2421 9367
rect 2455 9364 2467 9367
rect 4338 9364 4344 9376
rect 2455 9336 4344 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 5736 9373 5764 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 18984 9432 19012 9463
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 20806 9460 20812 9512
rect 20864 9500 20870 9512
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 20864 9472 21005 9500
rect 20864 9460 20870 9472
rect 20993 9469 21005 9472
rect 21039 9469 21051 9503
rect 20993 9463 21051 9469
rect 21726 9460 21732 9512
rect 21784 9500 21790 9512
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 21784 9472 22017 9500
rect 21784 9460 21790 9472
rect 22005 9469 22017 9472
rect 22051 9469 22063 9503
rect 23014 9500 23020 9512
rect 22975 9472 23020 9500
rect 22005 9463 22063 9469
rect 23014 9460 23020 9472
rect 23072 9460 23078 9512
rect 24578 9500 24584 9512
rect 24539 9472 24584 9500
rect 24578 9460 24584 9472
rect 24636 9460 24642 9512
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 25682 9500 25688 9512
rect 25639 9472 25688 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 26602 9500 26608 9512
rect 26563 9472 26608 9500
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 27614 9500 27620 9512
rect 27575 9472 27620 9500
rect 27614 9460 27620 9472
rect 27672 9460 27678 9512
rect 28718 9460 28724 9512
rect 28776 9500 28782 9512
rect 29089 9503 29147 9509
rect 29089 9500 29101 9503
rect 28776 9472 29101 9500
rect 28776 9460 28782 9472
rect 29089 9469 29101 9472
rect 29135 9469 29147 9503
rect 29089 9463 29147 9469
rect 29730 9460 29736 9512
rect 29788 9500 29794 9512
rect 30929 9503 30987 9509
rect 30929 9500 30941 9503
rect 29788 9472 30941 9500
rect 29788 9460 29794 9472
rect 30929 9469 30941 9472
rect 30975 9469 30987 9503
rect 30929 9463 30987 9469
rect 31754 9460 31760 9512
rect 31812 9500 31818 9512
rect 31941 9503 31999 9509
rect 31941 9500 31953 9503
rect 31812 9472 31953 9500
rect 31812 9460 31818 9472
rect 31941 9469 31953 9472
rect 31987 9469 31999 9503
rect 31941 9463 31999 9469
rect 32122 9460 32128 9512
rect 32180 9500 32186 9512
rect 32953 9503 33011 9509
rect 32953 9500 32965 9503
rect 32180 9472 32965 9500
rect 32180 9460 32186 9472
rect 32953 9469 32965 9472
rect 32999 9469 33011 9503
rect 32953 9463 33011 9469
rect 33134 9460 33140 9512
rect 33192 9500 33198 9512
rect 33965 9503 34023 9509
rect 33965 9500 33977 9503
rect 33192 9472 33977 9500
rect 33192 9460 33198 9472
rect 33965 9469 33977 9472
rect 34011 9469 34023 9503
rect 35802 9500 35808 9512
rect 35763 9472 35808 9500
rect 33965 9463 34023 9469
rect 35802 9460 35808 9472
rect 35860 9460 35866 9512
rect 36814 9500 36820 9512
rect 36775 9472 36820 9500
rect 36814 9460 36820 9472
rect 36872 9460 36878 9512
rect 37829 9503 37887 9509
rect 37829 9469 37841 9503
rect 37875 9500 37887 9503
rect 38470 9500 38476 9512
rect 37875 9472 38476 9500
rect 37875 9469 37887 9472
rect 37829 9463 37887 9469
rect 38470 9460 38476 9472
rect 38528 9460 38534 9512
rect 20714 9432 20720 9444
rect 18984 9404 20720 9432
rect 20714 9392 20720 9404
rect 20772 9392 20778 9444
rect 29454 9432 29460 9444
rect 25424 9404 29460 9432
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9333 5779 9367
rect 5721 9327 5779 9333
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 7708 9336 8585 9364
rect 7708 9324 7714 9336
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 8573 9327 8631 9333
rect 10505 9367 10563 9373
rect 10505 9333 10517 9367
rect 10551 9364 10563 9367
rect 11606 9364 11612 9376
rect 10551 9336 11612 9364
rect 10551 9333 10563 9336
rect 10505 9327 10563 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 15197 9367 15255 9373
rect 15197 9364 15209 9367
rect 13872 9336 15209 9364
rect 13872 9324 13878 9336
rect 15197 9333 15209 9336
rect 15243 9333 15255 9367
rect 16206 9364 16212 9376
rect 16167 9336 16212 9364
rect 15197 9327 15255 9333
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 18785 9367 18843 9373
rect 18785 9333 18797 9367
rect 18831 9364 18843 9367
rect 19242 9364 19248 9376
rect 18831 9336 19248 9364
rect 18831 9333 18843 9336
rect 18785 9327 18843 9333
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 19797 9367 19855 9373
rect 19797 9333 19809 9367
rect 19843 9364 19855 9367
rect 20254 9364 20260 9376
rect 19843 9336 20260 9364
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 20809 9367 20867 9373
rect 20809 9333 20821 9367
rect 20855 9364 20867 9367
rect 22002 9364 22008 9376
rect 20855 9336 22008 9364
rect 20855 9333 20867 9336
rect 20809 9327 20867 9333
rect 22002 9324 22008 9336
rect 22060 9324 22066 9376
rect 22830 9364 22836 9376
rect 22791 9336 22836 9364
rect 22830 9324 22836 9336
rect 22888 9324 22894 9376
rect 25424 9373 25452 9404
rect 29454 9392 29460 9404
rect 29512 9392 29518 9444
rect 25409 9367 25467 9373
rect 25409 9333 25421 9367
rect 25455 9333 25467 9367
rect 25409 9327 25467 9333
rect 26326 9324 26332 9376
rect 26384 9364 26390 9376
rect 26421 9367 26479 9373
rect 26421 9364 26433 9367
rect 26384 9336 26433 9364
rect 26384 9324 26390 9336
rect 26421 9333 26433 9336
rect 26467 9333 26479 9367
rect 26421 9327 26479 9333
rect 30745 9367 30803 9373
rect 30745 9333 30757 9367
rect 30791 9364 30803 9367
rect 30926 9364 30932 9376
rect 30791 9336 30932 9364
rect 30791 9333 30803 9336
rect 30745 9327 30803 9333
rect 30926 9324 30932 9336
rect 30984 9324 30990 9376
rect 31757 9367 31815 9373
rect 31757 9333 31769 9367
rect 31803 9364 31815 9367
rect 32306 9364 32312 9376
rect 31803 9336 32312 9364
rect 31803 9333 31815 9336
rect 31757 9327 31815 9333
rect 32306 9324 32312 9336
rect 32364 9324 32370 9376
rect 33781 9367 33839 9373
rect 33781 9333 33793 9367
rect 33827 9364 33839 9367
rect 34514 9364 34520 9376
rect 33827 9336 34520 9364
rect 33827 9333 33839 9336
rect 33781 9327 33839 9333
rect 34514 9324 34520 9336
rect 34572 9324 34578 9376
rect 35621 9367 35679 9373
rect 35621 9333 35633 9367
rect 35667 9364 35679 9367
rect 36722 9364 36728 9376
rect 35667 9336 36728 9364
rect 35667 9333 35679 9336
rect 35621 9327 35679 9333
rect 36722 9324 36728 9336
rect 36780 9324 36786 9376
rect 1104 9274 54832 9296
rect 1104 9222 18912 9274
rect 18964 9222 18976 9274
rect 19028 9222 19040 9274
rect 19092 9222 19104 9274
rect 19156 9222 36843 9274
rect 36895 9222 36907 9274
rect 36959 9222 36971 9274
rect 37023 9222 37035 9274
rect 37087 9222 54832 9274
rect 1104 9200 54832 9222
rect 4798 9160 4804 9172
rect 4759 9132 4804 9160
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 7466 9160 7472 9172
rect 7427 9132 7472 9160
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 13446 9160 13452 9172
rect 12492 9132 12537 9160
rect 13407 9132 13452 9160
rect 12492 9120 12498 9132
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 16022 9160 16028 9172
rect 15983 9132 16028 9160
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 20070 9160 20076 9172
rect 20031 9132 20076 9160
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 21637 9163 21695 9169
rect 21637 9129 21649 9163
rect 21683 9160 21695 9163
rect 21910 9160 21916 9172
rect 21683 9132 21916 9160
rect 21683 9129 21695 9132
rect 21637 9123 21695 9129
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 24121 9163 24179 9169
rect 24121 9129 24133 9163
rect 24167 9160 24179 9163
rect 24210 9160 24216 9172
rect 24167 9132 24216 9160
rect 24167 9129 24179 9132
rect 24121 9123 24179 9129
rect 24210 9120 24216 9132
rect 24268 9120 24274 9172
rect 25133 9163 25191 9169
rect 25133 9129 25145 9163
rect 25179 9160 25191 9163
rect 27522 9160 27528 9172
rect 25179 9132 27528 9160
rect 25179 9129 25191 9132
rect 25133 9123 25191 9129
rect 27522 9120 27528 9132
rect 27580 9120 27586 9172
rect 28718 9160 28724 9172
rect 28679 9132 28724 9160
rect 28718 9120 28724 9132
rect 28776 9120 28782 9172
rect 29730 9160 29736 9172
rect 29691 9132 29736 9160
rect 29730 9120 29736 9132
rect 29788 9120 29794 9172
rect 31757 9163 31815 9169
rect 31757 9129 31769 9163
rect 31803 9160 31815 9163
rect 32122 9160 32128 9172
rect 31803 9132 32128 9160
rect 31803 9129 31815 9132
rect 31757 9123 31815 9129
rect 32122 9120 32128 9132
rect 32180 9120 32186 9172
rect 33134 9160 33140 9172
rect 33095 9132 33140 9160
rect 33134 9120 33140 9132
rect 33192 9120 33198 9172
rect 38470 9160 38476 9172
rect 38431 9132 38476 9160
rect 38470 9120 38476 9132
rect 38528 9120 38534 9172
rect 2130 9052 2136 9104
rect 2188 9092 2194 9104
rect 10502 9092 10508 9104
rect 2188 9064 10508 9092
rect 2188 9052 2194 9064
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 16853 9095 16911 9101
rect 16853 9092 16865 9095
rect 10744 9064 12296 9092
rect 10744 9052 10750 9064
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 2924 8996 3157 9024
rect 2924 8984 2930 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5534 9024 5540 9036
rect 5031 8996 5540 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 7466 9024 7472 9036
rect 6687 8996 7472 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 7650 9024 7656 9036
rect 7611 8996 7656 9024
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8662 9024 8668 9036
rect 8623 8996 8668 9024
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 11606 9024 11612 9036
rect 10643 8996 11468 9024
rect 11567 8996 11612 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 2961 8891 3019 8897
rect 2961 8857 2973 8891
rect 3007 8888 3019 8891
rect 8018 8888 8024 8900
rect 3007 8860 8024 8888
rect 3007 8857 3019 8860
rect 2961 8851 3019 8857
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 11238 8888 11244 8900
rect 8260 8860 11244 8888
rect 8260 8848 8266 8860
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 11440 8897 11468 8996
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 12268 9024 12296 9064
rect 12544 9064 16865 9092
rect 12544 9024 12572 9064
rect 16853 9061 16865 9064
rect 16899 9061 16911 9095
rect 27246 9092 27252 9104
rect 16853 9055 16911 9061
rect 25332 9064 27252 9092
rect 12268 8996 12572 9024
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 13170 9024 13176 9036
rect 12667 8996 13176 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13630 9024 13636 9036
rect 13591 8996 13636 9024
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 16206 9024 16212 9036
rect 16167 8996 16212 9024
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 16868 9024 16896 9055
rect 17221 9027 17279 9033
rect 17221 9024 17233 9027
rect 16868 8996 17233 9024
rect 17221 8993 17233 8996
rect 17267 8993 17279 9027
rect 18230 9024 18236 9036
rect 18191 8996 18236 9024
rect 17221 8987 17279 8993
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 19242 9024 19248 9036
rect 19203 8996 19248 9024
rect 19242 8984 19248 8996
rect 19300 8984 19306 9036
rect 20254 9024 20260 9036
rect 20215 8996 20260 9024
rect 20254 8984 20260 8996
rect 20312 8984 20318 9036
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 9024 21879 9027
rect 22830 9024 22836 9036
rect 21867 8996 22836 9024
rect 21867 8993 21879 8996
rect 21821 8987 21879 8993
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 23106 8984 23112 9036
rect 23164 9024 23170 9036
rect 23293 9027 23351 9033
rect 23293 9024 23305 9027
rect 23164 8996 23305 9024
rect 23164 8984 23170 8996
rect 23293 8993 23305 8996
rect 23339 8993 23351 9027
rect 24302 9024 24308 9036
rect 24263 8996 24308 9024
rect 23293 8987 23351 8993
rect 24302 8984 24308 8996
rect 24360 8984 24366 9036
rect 25332 9033 25360 9064
rect 27246 9052 27252 9064
rect 27304 9052 27310 9104
rect 37182 9052 37188 9104
rect 37240 9092 37246 9104
rect 37240 9064 38700 9092
rect 37240 9052 37246 9064
rect 25317 9027 25375 9033
rect 25317 8993 25329 9027
rect 25363 8993 25375 9027
rect 26326 9024 26332 9036
rect 26287 8996 26332 9024
rect 25317 8987 25375 8993
rect 26326 8984 26332 8996
rect 26384 8984 26390 9036
rect 27154 8984 27160 9036
rect 27212 9024 27218 9036
rect 27893 9027 27951 9033
rect 27893 9024 27905 9027
rect 27212 8996 27905 9024
rect 27212 8984 27218 8996
rect 27893 8993 27905 8996
rect 27939 8993 27951 9027
rect 27893 8987 27951 8993
rect 28905 9027 28963 9033
rect 28905 8993 28917 9027
rect 28951 9024 28963 9027
rect 29546 9024 29552 9036
rect 28951 8996 29552 9024
rect 28951 8993 28963 8996
rect 28905 8987 28963 8993
rect 29546 8984 29552 8996
rect 29604 8984 29610 9036
rect 29917 9027 29975 9033
rect 29917 8993 29929 9027
rect 29963 9024 29975 9027
rect 30558 9024 30564 9036
rect 29963 8996 30564 9024
rect 29963 8993 29975 8996
rect 29917 8987 29975 8993
rect 30558 8984 30564 8996
rect 30616 8984 30622 9036
rect 30926 9024 30932 9036
rect 30887 8996 30932 9024
rect 30926 8984 30932 8996
rect 30984 8984 30990 9036
rect 31941 9027 31999 9033
rect 31941 8993 31953 9027
rect 31987 9024 31999 9027
rect 32766 9024 32772 9036
rect 31987 8996 32772 9024
rect 31987 8993 31999 8996
rect 31941 8987 31999 8993
rect 32766 8984 32772 8996
rect 32824 8984 32830 9036
rect 33318 9024 33324 9036
rect 33279 8996 33324 9024
rect 33318 8984 33324 8996
rect 33376 8984 33382 9036
rect 34333 9027 34391 9033
rect 34333 8993 34345 9027
rect 34379 8993 34391 9027
rect 35342 9024 35348 9036
rect 35303 8996 35348 9024
rect 34333 8987 34391 8993
rect 34348 8956 34376 8987
rect 35342 8984 35348 8996
rect 35400 8984 35406 9036
rect 36357 9027 36415 9033
rect 36357 8993 36369 9027
rect 36403 9024 36415 9027
rect 37642 9024 37648 9036
rect 36403 8996 37648 9024
rect 36403 8993 36415 8996
rect 36357 8987 36415 8993
rect 37642 8984 37648 8996
rect 37700 8984 37706 9036
rect 38672 9033 38700 9064
rect 38657 9027 38715 9033
rect 38657 8993 38669 9027
rect 38703 8993 38715 9027
rect 38657 8987 38715 8993
rect 34348 8928 36216 8956
rect 11425 8891 11483 8897
rect 11425 8857 11437 8891
rect 11471 8857 11483 8891
rect 17034 8888 17040 8900
rect 16995 8860 17040 8888
rect 11425 8851 11483 8857
rect 17034 8848 17040 8860
rect 17092 8848 17098 8900
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 36188 8897 36216 8928
rect 19061 8891 19119 8897
rect 19061 8888 19073 8891
rect 18012 8860 19073 8888
rect 18012 8848 18018 8860
rect 19061 8857 19073 8860
rect 19107 8857 19119 8891
rect 19061 8851 19119 8857
rect 36173 8891 36231 8897
rect 36173 8857 36185 8891
rect 36219 8857 36231 8891
rect 36173 8851 36231 8857
rect 6457 8823 6515 8829
rect 6457 8789 6469 8823
rect 6503 8820 6515 8823
rect 7650 8820 7656 8832
rect 6503 8792 7656 8820
rect 6503 8789 6515 8792
rect 6457 8783 6515 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 7800 8792 8493 8820
rect 7800 8780 7806 8792
rect 8481 8789 8493 8792
rect 8527 8789 8539 8823
rect 8481 8783 8539 8789
rect 10413 8823 10471 8829
rect 10413 8789 10425 8823
rect 10459 8820 10471 8823
rect 11698 8820 11704 8832
rect 10459 8792 11704 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 18049 8823 18107 8829
rect 18049 8789 18061 8823
rect 18095 8820 18107 8823
rect 18966 8820 18972 8832
rect 18095 8792 18972 8820
rect 18095 8789 18107 8792
rect 18049 8783 18107 8789
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 23109 8823 23167 8829
rect 23109 8789 23121 8823
rect 23155 8820 23167 8823
rect 24026 8820 24032 8832
rect 23155 8792 24032 8820
rect 23155 8789 23167 8792
rect 23109 8783 23167 8789
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 26142 8820 26148 8832
rect 26103 8792 26148 8820
rect 26142 8780 26148 8792
rect 26200 8780 26206 8832
rect 27709 8823 27767 8829
rect 27709 8789 27721 8823
rect 27755 8820 27767 8823
rect 28718 8820 28724 8832
rect 27755 8792 28724 8820
rect 27755 8789 27767 8792
rect 27709 8783 27767 8789
rect 28718 8780 28724 8792
rect 28776 8780 28782 8832
rect 30745 8823 30803 8829
rect 30745 8789 30757 8823
rect 30791 8820 30803 8823
rect 31202 8820 31208 8832
rect 30791 8792 31208 8820
rect 30791 8789 30803 8792
rect 30745 8783 30803 8789
rect 31202 8780 31208 8792
rect 31260 8780 31266 8832
rect 33962 8780 33968 8832
rect 34020 8820 34026 8832
rect 34149 8823 34207 8829
rect 34149 8820 34161 8823
rect 34020 8792 34161 8820
rect 34020 8780 34026 8792
rect 34149 8789 34161 8792
rect 34195 8789 34207 8823
rect 35158 8820 35164 8832
rect 35119 8792 35164 8820
rect 34149 8783 34207 8789
rect 35158 8780 35164 8792
rect 35216 8780 35222 8832
rect 1104 8730 54832 8752
rect 1104 8678 9947 8730
rect 9999 8678 10011 8730
rect 10063 8678 10075 8730
rect 10127 8678 10139 8730
rect 10191 8678 27878 8730
rect 27930 8678 27942 8730
rect 27994 8678 28006 8730
rect 28058 8678 28070 8730
rect 28122 8678 45808 8730
rect 45860 8678 45872 8730
rect 45924 8678 45936 8730
rect 45988 8678 46000 8730
rect 46052 8678 54832 8730
rect 1104 8656 54832 8678
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 5442 8616 5448 8628
rect 5403 8588 5448 8616
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 7524 8588 8585 8616
rect 7524 8576 7530 8588
rect 8573 8585 8585 8588
rect 8619 8585 8631 8619
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 8573 8579 8631 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 16945 8619 17003 8625
rect 16945 8585 16957 8619
rect 16991 8616 17003 8619
rect 18230 8616 18236 8628
rect 16991 8588 18236 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 20036 8588 21833 8616
rect 20036 8576 20042 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 25133 8619 25191 8625
rect 25133 8585 25145 8619
rect 25179 8616 25191 8619
rect 26602 8616 26608 8628
rect 25179 8588 26608 8616
rect 25179 8585 25191 8588
rect 25133 8579 25191 8585
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 27154 8616 27160 8628
rect 27115 8588 27160 8616
rect 27154 8576 27160 8588
rect 27212 8576 27218 8628
rect 30558 8616 30564 8628
rect 30519 8588 30564 8616
rect 30558 8576 30564 8588
rect 30616 8576 30622 8628
rect 31754 8576 31760 8628
rect 31812 8616 31818 8628
rect 32766 8616 32772 8628
rect 31812 8588 31857 8616
rect 32727 8588 32772 8616
rect 31812 8576 31818 8588
rect 32766 8576 32772 8588
rect 32824 8576 32830 8628
rect 33781 8619 33839 8625
rect 33781 8585 33793 8619
rect 33827 8616 33839 8619
rect 35802 8616 35808 8628
rect 33827 8588 35808 8616
rect 33827 8585 33839 8588
rect 33781 8579 33839 8585
rect 35802 8576 35808 8588
rect 35860 8576 35866 8628
rect 37642 8616 37648 8628
rect 37603 8588 37648 8616
rect 37642 8576 37648 8588
rect 37700 8576 37706 8628
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 6270 8548 6276 8560
rect 4479 8520 6276 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 6457 8551 6515 8557
rect 6457 8517 6469 8551
rect 6503 8517 6515 8551
rect 6457 8511 6515 8517
rect 7561 8551 7619 8557
rect 7561 8517 7573 8551
rect 7607 8548 7619 8551
rect 8754 8548 8760 8560
rect 7607 8520 8760 8548
rect 7607 8517 7619 8520
rect 7561 8511 7619 8517
rect 3050 8412 3056 8424
rect 3011 8384 3056 8412
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8412 4675 8415
rect 5534 8412 5540 8424
rect 4663 8384 5540 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8412 5687 8415
rect 6472 8412 6500 8511
rect 8754 8508 8760 8520
rect 8812 8508 8818 8560
rect 10597 8551 10655 8557
rect 10597 8517 10609 8551
rect 10643 8548 10655 8551
rect 11514 8548 11520 8560
rect 10643 8520 11520 8548
rect 10643 8517 10655 8520
rect 10597 8511 10655 8517
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 14185 8551 14243 8557
rect 14185 8548 14197 8551
rect 13780 8520 14197 8548
rect 13780 8508 13786 8520
rect 14185 8517 14197 8520
rect 14231 8517 14243 8551
rect 14185 8511 14243 8517
rect 15197 8551 15255 8557
rect 15197 8517 15209 8551
rect 15243 8548 15255 8551
rect 17218 8548 17224 8560
rect 15243 8520 17224 8548
rect 15243 8517 15255 8520
rect 15197 8511 15255 8517
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 19797 8551 19855 8557
rect 19797 8517 19809 8551
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 11422 8440 11428 8492
rect 11480 8480 11486 8492
rect 19812 8480 19840 8511
rect 20714 8508 20720 8560
rect 20772 8548 20778 8560
rect 20809 8551 20867 8557
rect 20809 8548 20821 8551
rect 20772 8520 20821 8548
rect 20772 8508 20778 8520
rect 20809 8517 20821 8520
rect 20855 8517 20867 8551
rect 20809 8511 20867 8517
rect 26145 8551 26203 8557
rect 26145 8517 26157 8551
rect 26191 8548 26203 8551
rect 26326 8548 26332 8560
rect 26191 8520 26332 8548
rect 26191 8517 26203 8520
rect 26145 8511 26203 8517
rect 26326 8508 26332 8520
rect 26384 8508 26390 8560
rect 28169 8551 28227 8557
rect 28169 8517 28181 8551
rect 28215 8548 28227 8551
rect 29730 8548 29736 8560
rect 28215 8520 29736 8548
rect 28215 8517 28227 8520
rect 28169 8511 28227 8517
rect 29730 8508 29736 8520
rect 29788 8508 29794 8560
rect 34514 8508 34520 8560
rect 34572 8548 34578 8560
rect 36633 8551 36691 8557
rect 36633 8548 36645 8551
rect 34572 8520 36645 8548
rect 34572 8508 34578 8520
rect 36633 8517 36645 8520
rect 36679 8517 36691 8551
rect 36633 8511 36691 8517
rect 26234 8480 26240 8492
rect 11480 8452 13400 8480
rect 11480 8440 11486 8452
rect 6638 8412 6644 8424
rect 5675 8384 6500 8412
rect 6599 8384 6644 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 6638 8372 6644 8384
rect 6696 8372 6702 8424
rect 7742 8412 7748 8424
rect 7703 8384 7748 8412
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8352 8384 8769 8412
rect 8352 8372 8358 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11606 8412 11612 8424
rect 10827 8384 11612 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 9784 8344 9812 8375
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 13372 8421 13400 8452
rect 17144 8452 19840 8480
rect 25332 8452 26240 8480
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 14366 8412 14372 8424
rect 14327 8384 14372 8412
rect 13357 8375 13415 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 15378 8412 15384 8424
rect 15339 8384 15384 8412
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 17144 8421 17172 8452
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8381 17187 8415
rect 18966 8412 18972 8424
rect 18927 8384 18972 8412
rect 17129 8375 17187 8381
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19978 8412 19984 8424
rect 19939 8384 19984 8412
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20680 8384 21005 8412
rect 20680 8372 20686 8384
rect 20993 8381 21005 8384
rect 21039 8381 21051 8415
rect 22002 8412 22008 8424
rect 21963 8384 22008 8412
rect 20993 8375 21051 8381
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 23014 8412 23020 8424
rect 22975 8384 23020 8412
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 25332 8421 25360 8452
rect 26234 8440 26240 8452
rect 26292 8440 26298 8492
rect 35986 8440 35992 8492
rect 36044 8480 36050 8492
rect 36044 8452 37872 8480
rect 36044 8440 36050 8452
rect 25317 8415 25375 8421
rect 25317 8381 25329 8415
rect 25363 8381 25375 8415
rect 25317 8375 25375 8381
rect 26142 8372 26148 8424
rect 26200 8412 26206 8424
rect 26329 8415 26387 8421
rect 26329 8412 26341 8415
rect 26200 8384 26341 8412
rect 26200 8372 26206 8384
rect 26329 8381 26341 8384
rect 26375 8381 26387 8415
rect 27338 8412 27344 8424
rect 27299 8384 27344 8412
rect 26329 8375 26387 8381
rect 27338 8372 27344 8384
rect 27396 8372 27402 8424
rect 28350 8412 28356 8424
rect 28311 8384 28356 8412
rect 28350 8372 28356 8384
rect 28408 8372 28414 8424
rect 30742 8412 30748 8424
rect 30703 8384 30748 8412
rect 30742 8372 30748 8384
rect 30800 8372 30806 8424
rect 31202 8372 31208 8424
rect 31260 8412 31266 8424
rect 31941 8415 31999 8421
rect 31941 8412 31953 8415
rect 31260 8384 31953 8412
rect 31260 8372 31266 8384
rect 31941 8381 31953 8384
rect 31987 8381 31999 8415
rect 32950 8412 32956 8424
rect 32911 8384 32956 8412
rect 31941 8375 31999 8381
rect 32950 8372 32956 8384
rect 33008 8372 33014 8424
rect 33962 8412 33968 8424
rect 33923 8384 33968 8412
rect 33962 8372 33968 8384
rect 34020 8372 34026 8424
rect 34606 8372 34612 8424
rect 34664 8412 34670 8424
rect 35805 8415 35863 8421
rect 35805 8412 35817 8415
rect 34664 8384 35817 8412
rect 34664 8372 34670 8384
rect 35805 8381 35817 8384
rect 35851 8381 35863 8415
rect 35805 8375 35863 8381
rect 36722 8372 36728 8424
rect 36780 8412 36786 8424
rect 37844 8421 37872 8452
rect 36817 8415 36875 8421
rect 36817 8412 36829 8415
rect 36780 8384 36829 8412
rect 36780 8372 36786 8384
rect 36817 8381 36829 8384
rect 36863 8381 36875 8415
rect 36817 8375 36875 8381
rect 37829 8415 37887 8421
rect 37829 8381 37841 8415
rect 37875 8381 37887 8415
rect 37829 8375 37887 8381
rect 11422 8344 11428 8356
rect 9784 8316 11428 8344
rect 11422 8304 11428 8316
rect 11480 8304 11486 8356
rect 9585 8279 9643 8285
rect 9585 8245 9597 8279
rect 9631 8276 9643 8279
rect 10778 8276 10784 8288
rect 9631 8248 10784 8276
rect 9631 8245 9643 8248
rect 9585 8239 9643 8245
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 18782 8276 18788 8288
rect 18743 8248 18788 8276
rect 18782 8236 18788 8248
rect 18840 8236 18846 8288
rect 22833 8279 22891 8285
rect 22833 8245 22845 8279
rect 22879 8276 22891 8279
rect 23290 8276 23296 8288
rect 22879 8248 23296 8276
rect 22879 8245 22891 8248
rect 22833 8239 22891 8245
rect 23290 8236 23296 8248
rect 23348 8236 23354 8288
rect 34974 8236 34980 8288
rect 35032 8276 35038 8288
rect 35621 8279 35679 8285
rect 35621 8276 35633 8279
rect 35032 8248 35633 8276
rect 35032 8236 35038 8248
rect 35621 8245 35633 8248
rect 35667 8245 35679 8279
rect 35621 8239 35679 8245
rect 1104 8186 54832 8208
rect 1104 8134 18912 8186
rect 18964 8134 18976 8186
rect 19028 8134 19040 8186
rect 19092 8134 19104 8186
rect 19156 8134 36843 8186
rect 36895 8134 36907 8186
rect 36959 8134 36971 8186
rect 37023 8134 37035 8186
rect 37087 8134 54832 8186
rect 1104 8112 54832 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 3050 8072 3056 8084
rect 2179 8044 3056 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 8662 8072 8668 8084
rect 7607 8044 8668 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 11422 8072 11428 8084
rect 11383 8044 11428 8072
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11606 8032 11612 8084
rect 11664 8072 11670 8084
rect 12437 8075 12495 8081
rect 12437 8072 12449 8075
rect 11664 8044 12449 8072
rect 11664 8032 11670 8044
rect 12437 8041 12449 8044
rect 12483 8041 12495 8075
rect 12437 8035 12495 8041
rect 13449 8075 13507 8081
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 14366 8072 14372 8084
rect 13495 8044 14372 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14921 8075 14979 8081
rect 14921 8041 14933 8075
rect 14967 8041 14979 8075
rect 14921 8035 14979 8041
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 19978 8072 19984 8084
rect 19659 8044 19984 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 14936 8004 14964 8035
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 21637 8075 21695 8081
rect 21637 8041 21649 8075
rect 21683 8072 21695 8075
rect 22370 8072 22376 8084
rect 21683 8044 22376 8072
rect 21683 8041 21695 8044
rect 21637 8035 21695 8041
rect 22370 8032 22376 8044
rect 22428 8032 22434 8084
rect 23106 8072 23112 8084
rect 23067 8044 23112 8072
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 24118 8072 24124 8084
rect 24079 8044 24124 8072
rect 24118 8032 24124 8044
rect 24176 8032 24182 8084
rect 25133 8075 25191 8081
rect 25133 8041 25145 8075
rect 25179 8072 25191 8075
rect 25222 8072 25228 8084
rect 25179 8044 25228 8072
rect 25179 8041 25191 8044
rect 25133 8035 25191 8041
rect 25222 8032 25228 8044
rect 25280 8032 25286 8084
rect 27338 8032 27344 8084
rect 27396 8072 27402 8084
rect 27525 8075 27583 8081
rect 27525 8072 27537 8075
rect 27396 8044 27537 8072
rect 27396 8032 27402 8044
rect 27525 8041 27537 8044
rect 27571 8041 27583 8075
rect 27525 8035 27583 8041
rect 28350 8032 28356 8084
rect 28408 8072 28414 8084
rect 28537 8075 28595 8081
rect 28537 8072 28549 8075
rect 28408 8044 28549 8072
rect 28408 8032 28414 8044
rect 28537 8041 28549 8044
rect 28583 8041 28595 8075
rect 29546 8072 29552 8084
rect 29507 8044 29552 8072
rect 28537 8035 28595 8041
rect 29546 8032 29552 8044
rect 29604 8032 29610 8084
rect 33781 8075 33839 8081
rect 33781 8041 33793 8075
rect 33827 8072 33839 8075
rect 35342 8072 35348 8084
rect 33827 8044 35348 8072
rect 33827 8041 33839 8044
rect 33781 8035 33839 8041
rect 35342 8032 35348 8044
rect 35400 8032 35406 8084
rect 28994 8004 29000 8016
rect 14936 7976 19840 8004
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 3234 7936 3240 7948
rect 2363 7908 3240 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3510 7936 3516 7948
rect 3375 7908 3516 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 5718 7936 5724 7948
rect 5679 7908 5724 7936
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 6748 7868 6776 7899
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7708 7908 7757 7936
rect 7708 7896 7714 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8757 7939 8815 7945
rect 8757 7936 8769 7939
rect 8444 7908 8769 7936
rect 8444 7896 8450 7908
rect 8757 7905 8769 7908
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 10597 7939 10655 7945
rect 10597 7936 10609 7939
rect 9732 7908 10609 7936
rect 9732 7896 9738 7908
rect 10597 7905 10609 7908
rect 10643 7905 10655 7939
rect 10597 7899 10655 7905
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11572 7908 11621 7936
rect 11572 7896 11578 7908
rect 11609 7905 11621 7908
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 11756 7908 12633 7936
rect 11756 7896 11762 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 13814 7936 13820 7948
rect 13679 7908 13820 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7905 15163 7939
rect 16206 7936 16212 7948
rect 16167 7908 16212 7936
rect 15105 7899 15163 7905
rect 15120 7868 15148 7899
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 17218 7936 17224 7948
rect 17179 7908 17224 7936
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 18785 7939 18843 7945
rect 18785 7905 18797 7939
rect 18831 7936 18843 7939
rect 19702 7936 19708 7948
rect 18831 7908 19708 7936
rect 18831 7905 18843 7908
rect 18785 7899 18843 7905
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 19812 7945 19840 7976
rect 25332 7976 29000 8004
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7905 19855 7939
rect 21818 7936 21824 7948
rect 21779 7908 21824 7936
rect 19797 7899 19855 7905
rect 21818 7896 21824 7908
rect 21876 7896 21882 7948
rect 23290 7936 23296 7948
rect 23251 7908 23296 7936
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 24026 7896 24032 7948
rect 24084 7936 24090 7948
rect 25332 7945 25360 7976
rect 28994 7964 29000 7976
rect 29052 7964 29058 8016
rect 24305 7939 24363 7945
rect 24305 7936 24317 7939
rect 24084 7908 24317 7936
rect 24084 7896 24090 7908
rect 24305 7905 24317 7908
rect 24351 7905 24363 7939
rect 24305 7899 24363 7905
rect 25317 7939 25375 7945
rect 25317 7905 25329 7939
rect 25363 7905 25375 7939
rect 26326 7936 26332 7948
rect 26287 7908 26332 7936
rect 25317 7899 25375 7905
rect 26326 7896 26332 7908
rect 26384 7896 26390 7948
rect 27338 7896 27344 7948
rect 27396 7936 27402 7948
rect 27709 7939 27767 7945
rect 27709 7936 27721 7939
rect 27396 7908 27721 7936
rect 27396 7896 27402 7908
rect 27709 7905 27721 7908
rect 27755 7905 27767 7939
rect 28718 7936 28724 7948
rect 28679 7908 28724 7936
rect 27709 7899 27767 7905
rect 28718 7896 28724 7908
rect 28776 7896 28782 7948
rect 29733 7939 29791 7945
rect 29733 7905 29745 7939
rect 29779 7936 29791 7939
rect 30006 7936 30012 7948
rect 29779 7908 30012 7936
rect 29779 7905 29791 7908
rect 29733 7899 29791 7905
rect 30006 7896 30012 7908
rect 30064 7896 30070 7948
rect 33965 7939 34023 7945
rect 33965 7905 33977 7939
rect 34011 7936 34023 7939
rect 34514 7936 34520 7948
rect 34011 7908 34520 7936
rect 34011 7905 34023 7908
rect 33965 7899 34023 7905
rect 34514 7896 34520 7908
rect 34572 7896 34578 7948
rect 34974 7936 34980 7948
rect 34935 7908 34980 7936
rect 34974 7896 34980 7908
rect 35032 7896 35038 7948
rect 35066 7896 35072 7948
rect 35124 7936 35130 7948
rect 35989 7939 36047 7945
rect 35989 7936 36001 7939
rect 35124 7908 36001 7936
rect 35124 7896 35130 7908
rect 35989 7905 36001 7908
rect 36035 7905 36047 7939
rect 35989 7899 36047 7905
rect 36078 7896 36084 7948
rect 36136 7936 36142 7948
rect 37001 7939 37059 7945
rect 37001 7936 37013 7939
rect 36136 7908 37013 7936
rect 36136 7896 36142 7908
rect 37001 7905 37013 7908
rect 37047 7905 37059 7939
rect 37001 7899 37059 7905
rect 17954 7868 17960 7880
rect 6748 7840 8616 7868
rect 15120 7840 17960 7868
rect 8588 7809 8616 7840
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 8573 7803 8631 7809
rect 8573 7769 8585 7803
rect 8619 7769 8631 7803
rect 8573 7763 8631 7769
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 5534 7732 5540 7744
rect 3191 7704 5540 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 6546 7732 6552 7744
rect 6507 7704 6552 7732
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 10413 7735 10471 7741
rect 10413 7732 10425 7735
rect 8812 7704 10425 7732
rect 8812 7692 8818 7704
rect 10413 7701 10425 7704
rect 10459 7701 10471 7735
rect 10413 7695 10471 7701
rect 16025 7735 16083 7741
rect 16025 7701 16037 7735
rect 16071 7732 16083 7735
rect 16390 7732 16396 7744
rect 16071 7704 16396 7732
rect 16071 7701 16083 7704
rect 16025 7695 16083 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 17037 7735 17095 7741
rect 17037 7701 17049 7735
rect 17083 7732 17095 7735
rect 18230 7732 18236 7744
rect 17083 7704 18236 7732
rect 17083 7701 17095 7704
rect 17037 7695 17095 7701
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7732 18659 7735
rect 19978 7732 19984 7744
rect 18647 7704 19984 7732
rect 18647 7701 18659 7704
rect 18601 7695 18659 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 26145 7735 26203 7741
rect 26145 7701 26157 7735
rect 26191 7732 26203 7735
rect 27522 7732 27528 7744
rect 26191 7704 27528 7732
rect 26191 7701 26203 7704
rect 26145 7695 26203 7701
rect 27522 7692 27528 7704
rect 27580 7692 27586 7744
rect 34514 7692 34520 7744
rect 34572 7732 34578 7744
rect 34793 7735 34851 7741
rect 34793 7732 34805 7735
rect 34572 7704 34805 7732
rect 34572 7692 34578 7704
rect 34793 7701 34805 7704
rect 34839 7701 34851 7735
rect 35802 7732 35808 7744
rect 35763 7704 35808 7732
rect 34793 7695 34851 7701
rect 35802 7692 35808 7704
rect 35860 7692 35866 7744
rect 35894 7692 35900 7744
rect 35952 7732 35958 7744
rect 36817 7735 36875 7741
rect 36817 7732 36829 7735
rect 35952 7704 36829 7732
rect 35952 7692 35958 7704
rect 36817 7701 36829 7704
rect 36863 7701 36875 7735
rect 36817 7695 36875 7701
rect 1104 7642 54832 7664
rect 1104 7590 9947 7642
rect 9999 7590 10011 7642
rect 10063 7590 10075 7642
rect 10127 7590 10139 7642
rect 10191 7590 27878 7642
rect 27930 7590 27942 7642
rect 27994 7590 28006 7642
rect 28058 7590 28070 7642
rect 28122 7590 45808 7642
rect 45860 7590 45872 7642
rect 45924 7590 45936 7642
rect 45988 7590 46000 7642
rect 46052 7590 54832 7642
rect 1104 7568 54832 7590
rect 3510 7528 3516 7540
rect 3471 7500 3516 7528
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 8294 7528 8300 7540
rect 7607 7500 8300 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 13173 7531 13231 7537
rect 13173 7497 13185 7531
rect 13219 7528 13231 7531
rect 18046 7528 18052 7540
rect 13219 7500 18052 7528
rect 13219 7497 13231 7500
rect 13173 7491 13231 7497
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 19702 7488 19708 7540
rect 19760 7528 19766 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 19760 7500 20821 7528
rect 19760 7488 19766 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 22557 7531 22615 7537
rect 22557 7497 22569 7531
rect 22603 7528 22615 7531
rect 23014 7528 23020 7540
rect 22603 7500 23020 7528
rect 22603 7497 22615 7500
rect 22557 7491 22615 7497
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 27338 7528 27344 7540
rect 27299 7500 27344 7528
rect 27338 7488 27344 7500
rect 27396 7488 27402 7540
rect 30006 7528 30012 7540
rect 29967 7500 30012 7528
rect 30006 7488 30012 7500
rect 30064 7488 30070 7540
rect 32769 7531 32827 7537
rect 32769 7497 32781 7531
rect 32815 7528 32827 7531
rect 32858 7528 32864 7540
rect 32815 7500 32864 7528
rect 32815 7497 32827 7500
rect 32769 7491 32827 7497
rect 32858 7488 32864 7500
rect 32916 7488 32922 7540
rect 33781 7531 33839 7537
rect 33781 7497 33793 7531
rect 33827 7528 33839 7531
rect 34606 7528 34612 7540
rect 33827 7500 34612 7528
rect 33827 7497 33839 7500
rect 33781 7491 33839 7497
rect 34606 7488 34612 7500
rect 34664 7488 34670 7540
rect 2133 7463 2191 7469
rect 2133 7429 2145 7463
rect 2179 7429 2191 7463
rect 2133 7423 2191 7429
rect 2148 7392 2176 7423
rect 23842 7420 23848 7472
rect 23900 7460 23906 7472
rect 25409 7463 25467 7469
rect 25409 7460 25421 7463
rect 23900 7432 25421 7460
rect 23900 7420 23906 7432
rect 25409 7429 25421 7432
rect 25455 7429 25467 7463
rect 25409 7423 25467 7429
rect 14642 7392 14648 7404
rect 2148 7364 3740 7392
rect 3712 7333 3740 7364
rect 13372 7364 14648 7392
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 3705 7327 3763 7333
rect 3705 7293 3717 7327
rect 3751 7293 3763 7327
rect 4706 7324 4712 7336
rect 4667 7296 4712 7324
rect 3705 7287 3763 7293
rect 2332 7256 2360 7287
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5902 7324 5908 7336
rect 5863 7296 5908 7324
rect 5902 7284 5908 7296
rect 5960 7284 5966 7336
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 6604 7296 7757 7324
rect 6604 7284 6610 7296
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 8754 7324 8760 7336
rect 8715 7296 8760 7324
rect 7745 7287 7803 7293
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 8996 7296 9781 7324
rect 8996 7284 9002 7296
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 10778 7324 10784 7336
rect 10739 7296 10784 7324
rect 9769 7287 9827 7293
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 13372 7333 13400 7364
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 13538 7284 13544 7336
rect 13596 7324 13602 7336
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 13596 7296 14381 7324
rect 13596 7284 13602 7296
rect 14369 7293 14381 7296
rect 14415 7293 14427 7327
rect 15378 7324 15384 7336
rect 15339 7296 15384 7324
rect 14369 7287 14427 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 16390 7324 16396 7336
rect 16351 7296 16396 7324
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 17773 7327 17831 7333
rect 17773 7293 17785 7327
rect 17819 7324 17831 7327
rect 18782 7324 18788 7336
rect 17819 7296 18788 7324
rect 17819 7293 17831 7296
rect 17773 7287 17831 7293
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18932 7296 18981 7324
rect 18932 7284 18938 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 19978 7324 19984 7336
rect 19939 7296 19984 7324
rect 18969 7287 19027 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20990 7324 20996 7336
rect 20951 7296 20996 7324
rect 20990 7284 20996 7296
rect 21048 7284 21054 7336
rect 22738 7324 22744 7336
rect 22699 7296 22744 7324
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 24578 7324 24584 7336
rect 24539 7296 24584 7324
rect 24578 7284 24584 7296
rect 24636 7284 24642 7336
rect 25038 7284 25044 7336
rect 25096 7324 25102 7336
rect 25593 7327 25651 7333
rect 25593 7324 25605 7327
rect 25096 7296 25605 7324
rect 25096 7284 25102 7296
rect 25593 7293 25605 7296
rect 25639 7293 25651 7327
rect 27522 7324 27528 7336
rect 27483 7296 27528 7324
rect 25593 7287 25651 7293
rect 27522 7284 27528 7296
rect 27580 7284 27586 7336
rect 30190 7324 30196 7336
rect 30151 7296 30196 7324
rect 30190 7284 30196 7296
rect 30248 7284 30254 7336
rect 32306 7284 32312 7336
rect 32364 7324 32370 7336
rect 32953 7327 33011 7333
rect 32953 7324 32965 7327
rect 32364 7296 32965 7324
rect 32364 7284 32370 7296
rect 32953 7293 32965 7296
rect 32999 7293 33011 7327
rect 32953 7287 33011 7293
rect 33965 7327 34023 7333
rect 33965 7293 33977 7327
rect 34011 7324 34023 7327
rect 35158 7324 35164 7336
rect 34011 7296 35164 7324
rect 34011 7293 34023 7296
rect 33965 7287 34023 7293
rect 35158 7284 35164 7296
rect 35216 7284 35222 7336
rect 35802 7324 35808 7336
rect 35763 7296 35808 7324
rect 35802 7284 35808 7296
rect 35860 7284 35866 7336
rect 36170 7284 36176 7336
rect 36228 7324 36234 7336
rect 36817 7327 36875 7333
rect 36817 7324 36829 7327
rect 36228 7296 36829 7324
rect 36228 7284 36234 7296
rect 36817 7293 36829 7296
rect 36863 7293 36875 7327
rect 38010 7324 38016 7336
rect 37971 7296 38016 7324
rect 36817 7287 36875 7293
rect 38010 7284 38016 7296
rect 38068 7284 38074 7336
rect 4798 7256 4804 7268
rect 2332 7228 4804 7256
rect 4798 7216 4804 7228
rect 4856 7216 4862 7268
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 5810 7188 5816 7200
rect 4571 7160 5816 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8352 7160 8585 7188
rect 8352 7148 8358 7160
rect 8573 7157 8585 7160
rect 8619 7157 8631 7191
rect 8573 7151 8631 7157
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 8720 7160 9597 7188
rect 8720 7148 8726 7160
rect 9585 7157 9597 7160
rect 9631 7157 9643 7191
rect 10594 7188 10600 7200
rect 10555 7160 10600 7188
rect 9585 7151 9643 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 14185 7191 14243 7197
rect 14185 7157 14197 7191
rect 14231 7188 14243 7191
rect 14366 7188 14372 7200
rect 14231 7160 14372 7188
rect 14231 7157 14243 7160
rect 14185 7151 14243 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 15194 7188 15200 7200
rect 15155 7160 15200 7188
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 15344 7160 16221 7188
rect 15344 7148 15350 7160
rect 16209 7157 16221 7160
rect 16255 7157 16267 7191
rect 16209 7151 16267 7157
rect 17589 7191 17647 7197
rect 17589 7157 17601 7191
rect 17635 7188 17647 7191
rect 18690 7188 18696 7200
rect 17635 7160 18696 7188
rect 17635 7157 17647 7160
rect 17589 7151 17647 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 18785 7191 18843 7197
rect 18785 7157 18797 7191
rect 18831 7188 18843 7191
rect 19334 7188 19340 7200
rect 18831 7160 19340 7188
rect 18831 7157 18843 7160
rect 18785 7151 18843 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 19797 7191 19855 7197
rect 19797 7157 19809 7191
rect 19843 7188 19855 7191
rect 20254 7188 20260 7200
rect 19843 7160 20260 7188
rect 19843 7157 19855 7160
rect 19797 7151 19855 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 22646 7148 22652 7200
rect 22704 7188 22710 7200
rect 24397 7191 24455 7197
rect 24397 7188 24409 7191
rect 22704 7160 24409 7188
rect 22704 7148 22710 7160
rect 24397 7157 24409 7160
rect 24443 7157 24455 7191
rect 24397 7151 24455 7157
rect 35621 7191 35679 7197
rect 35621 7157 35633 7191
rect 35667 7188 35679 7191
rect 35802 7188 35808 7200
rect 35667 7160 35808 7188
rect 35667 7157 35679 7160
rect 35621 7151 35679 7157
rect 35802 7148 35808 7160
rect 35860 7148 35866 7200
rect 35986 7148 35992 7200
rect 36044 7188 36050 7200
rect 36633 7191 36691 7197
rect 36633 7188 36645 7191
rect 36044 7160 36645 7188
rect 36044 7148 36050 7160
rect 36633 7157 36645 7160
rect 36679 7157 36691 7191
rect 36633 7151 36691 7157
rect 37829 7191 37887 7197
rect 37829 7157 37841 7191
rect 37875 7188 37887 7191
rect 39850 7188 39856 7200
rect 37875 7160 39856 7188
rect 37875 7157 37887 7160
rect 37829 7151 37887 7157
rect 39850 7148 39856 7160
rect 39908 7148 39914 7200
rect 1104 7098 54832 7120
rect 1104 7046 18912 7098
rect 18964 7046 18976 7098
rect 19028 7046 19040 7098
rect 19092 7046 19104 7098
rect 19156 7046 36843 7098
rect 36895 7046 36907 7098
rect 36959 7046 36971 7098
rect 37023 7046 37035 7098
rect 37087 7046 54832 7098
rect 1104 7024 54832 7046
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5902 6984 5908 6996
rect 5675 6956 5908 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 16025 6987 16083 6993
rect 16025 6953 16037 6987
rect 16071 6984 16083 6987
rect 16206 6984 16212 6996
rect 16071 6956 16212 6984
rect 16071 6953 16083 6956
rect 16025 6947 16083 6953
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 20990 6944 20996 6996
rect 21048 6984 21054 6996
rect 21637 6987 21695 6993
rect 21637 6984 21649 6987
rect 21048 6956 21649 6984
rect 21048 6944 21054 6956
rect 21637 6953 21649 6956
rect 21683 6953 21695 6987
rect 22738 6984 22744 6996
rect 22699 6956 22744 6984
rect 21637 6947 21695 6953
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 24578 6944 24584 6996
rect 24636 6984 24642 6996
rect 24765 6987 24823 6993
rect 24765 6984 24777 6987
rect 24636 6956 24777 6984
rect 24636 6944 24642 6956
rect 24765 6953 24777 6956
rect 24811 6953 24823 6987
rect 24765 6947 24823 6953
rect 29549 6987 29607 6993
rect 29549 6953 29561 6987
rect 29595 6984 29607 6987
rect 30190 6984 30196 6996
rect 29595 6956 30196 6984
rect 29595 6953 29607 6956
rect 29549 6947 29607 6953
rect 30190 6944 30196 6956
rect 30248 6944 30254 6996
rect 33597 6987 33655 6993
rect 33597 6953 33609 6987
rect 33643 6984 33655 6987
rect 33643 6956 34836 6984
rect 33643 6953 33655 6956
rect 33597 6947 33655 6953
rect 34514 6916 34520 6928
rect 34440 6888 34520 6916
rect 2869 6851 2927 6857
rect 2869 6817 2881 6851
rect 2915 6848 2927 6851
rect 3786 6848 3792 6860
rect 2915 6820 3792 6848
rect 2915 6817 2927 6820
rect 2869 6811 2927 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 5626 6848 5632 6860
rect 3927 6820 5632 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5810 6848 5816 6860
rect 5771 6820 5816 6848
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 8294 6848 8300 6860
rect 7699 6820 8300 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 8662 6848 8668 6860
rect 8623 6820 8668 6848
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 10594 6848 10600 6860
rect 10555 6820 10600 6848
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11204 6820 11621 6848
rect 11204 6808 11210 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6848 12771 6851
rect 12759 6820 13400 6848
rect 12759 6817 12771 6820
rect 12713 6811 12771 6817
rect 7469 6715 7527 6721
rect 7469 6681 7481 6715
rect 7515 6712 7527 6715
rect 8386 6712 8392 6724
rect 7515 6684 8392 6712
rect 7515 6681 7527 6684
rect 7469 6675 7527 6681
rect 8386 6672 8392 6684
rect 8444 6672 8450 6724
rect 8481 6715 8539 6721
rect 8481 6681 8493 6715
rect 8527 6712 8539 6715
rect 9674 6712 9680 6724
rect 8527 6684 9680 6712
rect 8527 6681 8539 6684
rect 8481 6675 8539 6681
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 12529 6715 12587 6721
rect 12529 6681 12541 6715
rect 12575 6712 12587 6715
rect 12710 6712 12716 6724
rect 12575 6684 12716 6712
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 13372 6712 13400 6820
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13504 6820 13737 6848
rect 13504 6808 13510 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 16206 6848 16212 6860
rect 16167 6820 16212 6848
rect 13725 6811 13783 6817
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 16356 6820 17233 6848
rect 16356 6808 16362 6820
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 18230 6848 18236 6860
rect 18191 6820 18236 6848
rect 17221 6811 17279 6817
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 18340 6820 19257 6848
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 18340 6780 18368 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 20128 6820 20269 6848
rect 20128 6808 20134 6820
rect 20257 6817 20269 6820
rect 20303 6817 20315 6851
rect 20257 6811 20315 6817
rect 21821 6851 21879 6857
rect 21821 6817 21833 6851
rect 21867 6817 21879 6851
rect 21821 6811 21879 6817
rect 16632 6752 18368 6780
rect 16632 6740 16638 6752
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 21836 6780 21864 6811
rect 22554 6808 22560 6860
rect 22612 6848 22618 6860
rect 22925 6851 22983 6857
rect 22925 6848 22937 6851
rect 22612 6820 22937 6848
rect 22612 6808 22618 6820
rect 22925 6817 22937 6820
rect 22971 6817 22983 6851
rect 22925 6811 22983 6817
rect 23750 6808 23756 6860
rect 23808 6848 23814 6860
rect 23937 6851 23995 6857
rect 23937 6848 23949 6851
rect 23808 6820 23949 6848
rect 23808 6808 23814 6820
rect 23937 6817 23949 6820
rect 23983 6817 23995 6851
rect 23937 6811 23995 6817
rect 24854 6808 24860 6860
rect 24912 6848 24918 6860
rect 24949 6851 25007 6857
rect 24949 6848 24961 6851
rect 24912 6820 24961 6848
rect 24912 6808 24918 6820
rect 24949 6817 24961 6820
rect 24995 6817 25007 6851
rect 24949 6811 25007 6817
rect 25961 6851 26019 6857
rect 25961 6817 25973 6851
rect 26007 6817 26019 6851
rect 25961 6811 26019 6817
rect 18748 6752 21864 6780
rect 18748 6740 18754 6752
rect 23474 6740 23480 6792
rect 23532 6780 23538 6792
rect 25976 6780 26004 6811
rect 26418 6808 26424 6860
rect 26476 6848 26482 6860
rect 27433 6851 27491 6857
rect 27433 6848 27445 6851
rect 26476 6820 27445 6848
rect 26476 6808 26482 6820
rect 27433 6817 27445 6820
rect 27479 6817 27491 6851
rect 29730 6848 29736 6860
rect 29691 6820 29736 6848
rect 27433 6811 27491 6817
rect 29730 6808 29736 6820
rect 29788 6808 29794 6860
rect 33781 6851 33839 6857
rect 33781 6817 33793 6851
rect 33827 6848 33839 6851
rect 34440 6848 34468 6888
rect 34514 6876 34520 6888
rect 34572 6876 34578 6928
rect 34808 6857 34836 6956
rect 33827 6820 34468 6848
rect 34793 6851 34851 6857
rect 33827 6817 33839 6820
rect 33781 6811 33839 6817
rect 34793 6817 34805 6851
rect 34839 6817 34851 6851
rect 35802 6848 35808 6860
rect 35763 6820 35808 6848
rect 34793 6811 34851 6817
rect 35802 6808 35808 6820
rect 35860 6808 35866 6860
rect 36262 6808 36268 6860
rect 36320 6848 36326 6860
rect 36909 6851 36967 6857
rect 36909 6848 36921 6851
rect 36320 6820 36921 6848
rect 36320 6808 36326 6820
rect 36909 6817 36921 6820
rect 36955 6817 36967 6851
rect 38654 6848 38660 6860
rect 38615 6820 38660 6848
rect 36909 6811 36967 6817
rect 38654 6808 38660 6820
rect 38712 6808 38718 6860
rect 39669 6851 39727 6857
rect 39669 6817 39681 6851
rect 39715 6848 39727 6851
rect 40494 6848 40500 6860
rect 39715 6820 40500 6848
rect 39715 6817 39727 6820
rect 39669 6811 39727 6817
rect 40494 6808 40500 6820
rect 40552 6808 40558 6860
rect 23532 6752 26004 6780
rect 23532 6740 23538 6752
rect 26970 6740 26976 6792
rect 27028 6780 27034 6792
rect 34422 6780 34428 6792
rect 27028 6752 34428 6780
rect 27028 6740 27034 6752
rect 34422 6740 34428 6752
rect 34480 6740 34486 6792
rect 34606 6740 34612 6792
rect 34664 6780 34670 6792
rect 51074 6780 51080 6792
rect 34664 6752 51080 6780
rect 34664 6740 34670 6752
rect 51074 6740 51080 6752
rect 51132 6740 51138 6792
rect 18414 6712 18420 6724
rect 13372 6684 18420 6712
rect 18414 6672 18420 6684
rect 18472 6672 18478 6724
rect 35621 6715 35679 6721
rect 35621 6681 35633 6715
rect 35667 6712 35679 6715
rect 36078 6712 36084 6724
rect 35667 6684 36084 6712
rect 35667 6681 35679 6684
rect 35621 6675 35679 6681
rect 36078 6672 36084 6684
rect 36136 6672 36142 6724
rect 36725 6715 36783 6721
rect 36725 6681 36737 6715
rect 36771 6712 36783 6715
rect 38010 6712 38016 6724
rect 36771 6684 38016 6712
rect 36771 6681 36783 6684
rect 36725 6675 36783 6681
rect 38010 6672 38016 6684
rect 38068 6672 38074 6724
rect 2685 6647 2743 6653
rect 2685 6613 2697 6647
rect 2731 6644 2743 6647
rect 3326 6644 3332 6656
rect 2731 6616 3332 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 3697 6647 3755 6653
rect 3697 6613 3709 6647
rect 3743 6644 3755 6647
rect 4890 6644 4896 6656
rect 3743 6616 4896 6644
rect 3743 6613 3755 6616
rect 3697 6607 3755 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 10413 6647 10471 6653
rect 10413 6644 10425 6647
rect 8628 6616 10425 6644
rect 8628 6604 8634 6616
rect 10413 6613 10425 6616
rect 10459 6613 10471 6647
rect 10413 6607 10471 6613
rect 10502 6604 10508 6656
rect 10560 6644 10566 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10560 6616 11437 6644
rect 10560 6604 10566 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 13541 6647 13599 6653
rect 13541 6644 13553 6647
rect 12676 6616 13553 6644
rect 12676 6604 12682 6616
rect 13541 6613 13553 6616
rect 13587 6613 13599 6647
rect 13541 6607 13599 6613
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16448 6616 17049 6644
rect 16448 6604 16454 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 17402 6604 17408 6656
rect 17460 6644 17466 6656
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 17460 6616 18061 6644
rect 17460 6604 17466 6616
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 19061 6647 19119 6653
rect 19061 6644 19073 6647
rect 18196 6616 19073 6644
rect 18196 6604 18202 6616
rect 19061 6613 19073 6616
rect 19107 6613 19119 6647
rect 19061 6607 19119 6613
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6644 20131 6647
rect 20990 6644 20996 6656
rect 20119 6616 20996 6644
rect 20119 6613 20131 6616
rect 20073 6607 20131 6613
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 22738 6604 22744 6656
rect 22796 6644 22802 6656
rect 23753 6647 23811 6653
rect 23753 6644 23765 6647
rect 22796 6616 23765 6644
rect 22796 6604 22802 6616
rect 23753 6613 23765 6616
rect 23799 6613 23811 6647
rect 23753 6607 23811 6613
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25777 6647 25835 6653
rect 25777 6644 25789 6647
rect 24912 6616 25789 6644
rect 24912 6604 24918 6616
rect 25777 6613 25789 6616
rect 25823 6613 25835 6647
rect 25777 6607 25835 6613
rect 27249 6647 27307 6653
rect 27249 6613 27261 6647
rect 27295 6644 27307 6647
rect 27614 6644 27620 6656
rect 27295 6616 27620 6644
rect 27295 6613 27307 6616
rect 27249 6607 27307 6613
rect 27614 6604 27620 6616
rect 27672 6604 27678 6656
rect 33962 6604 33968 6656
rect 34020 6644 34026 6656
rect 34609 6647 34667 6653
rect 34609 6644 34621 6647
rect 34020 6616 34621 6644
rect 34020 6604 34026 6616
rect 34609 6613 34621 6616
rect 34655 6613 34667 6647
rect 34609 6607 34667 6613
rect 38473 6647 38531 6653
rect 38473 6613 38485 6647
rect 38519 6644 38531 6647
rect 38838 6644 38844 6656
rect 38519 6616 38844 6644
rect 38519 6613 38531 6616
rect 38473 6607 38531 6613
rect 38838 6604 38844 6616
rect 38896 6604 38902 6656
rect 38930 6604 38936 6656
rect 38988 6644 38994 6656
rect 39485 6647 39543 6653
rect 39485 6644 39497 6647
rect 38988 6616 39497 6644
rect 38988 6604 38994 6616
rect 39485 6613 39497 6616
rect 39531 6613 39543 6647
rect 39485 6607 39543 6613
rect 1104 6554 54832 6576
rect 1104 6502 9947 6554
rect 9999 6502 10011 6554
rect 10063 6502 10075 6554
rect 10127 6502 10139 6554
rect 10191 6502 27878 6554
rect 27930 6502 27942 6554
rect 27994 6502 28006 6554
rect 28058 6502 28070 6554
rect 28122 6502 45808 6554
rect 45860 6502 45872 6554
rect 45924 6502 45936 6554
rect 45988 6502 46000 6554
rect 46052 6502 54832 6554
rect 1104 6480 54832 6502
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 5684 6412 5733 6440
rect 5684 6400 5690 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 5721 6403 5779 6409
rect 8205 6443 8263 6449
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8938 6440 8944 6452
rect 8251 6412 8944 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9217 6443 9275 6449
rect 9217 6409 9229 6443
rect 9263 6440 9275 6443
rect 11330 6440 11336 6452
rect 9263 6412 11336 6440
rect 9263 6409 9275 6412
rect 9217 6403 9275 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 15378 6440 15384 6452
rect 15243 6412 15384 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 16206 6440 16212 6452
rect 16167 6412 16212 6440
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 22554 6440 22560 6452
rect 22515 6412 22560 6440
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 22830 6400 22836 6452
rect 22888 6440 22894 6452
rect 29362 6440 29368 6452
rect 22888 6412 29368 6440
rect 22888 6400 22894 6412
rect 29362 6400 29368 6412
rect 29420 6400 29426 6452
rect 33781 6443 33839 6449
rect 33781 6409 33793 6443
rect 33827 6440 33839 6443
rect 35066 6440 35072 6452
rect 33827 6412 35072 6440
rect 33827 6409 33839 6412
rect 33781 6403 33839 6409
rect 35066 6400 35072 6412
rect 35124 6400 35130 6452
rect 35621 6443 35679 6449
rect 35621 6409 35633 6443
rect 35667 6440 35679 6443
rect 36170 6440 36176 6452
rect 35667 6412 36176 6440
rect 35667 6409 35679 6412
rect 35621 6403 35679 6409
rect 36170 6400 36176 6412
rect 36228 6400 36234 6452
rect 36633 6443 36691 6449
rect 36633 6409 36645 6443
rect 36679 6440 36691 6443
rect 38654 6440 38660 6452
rect 36679 6412 38660 6440
rect 36679 6409 36691 6412
rect 36633 6403 36691 6409
rect 38654 6400 38660 6412
rect 38712 6400 38718 6452
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6372 2743 6375
rect 5350 6372 5356 6384
rect 2731 6344 5356 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 10410 6372 10416 6384
rect 9416 6344 10416 6372
rect 2866 6236 2872 6248
rect 2827 6208 2872 6236
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 3384 6208 3893 6236
rect 3384 6196 3390 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 4890 6236 4896 6248
rect 4851 6208 4896 6236
rect 3881 6199 3939 6205
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5905 6239 5963 6245
rect 5905 6236 5917 6239
rect 5592 6208 5917 6236
rect 5592 6196 5598 6208
rect 5905 6205 5917 6208
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8570 6236 8576 6248
rect 8435 6208 8576 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9416 6245 9444 6344
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 25409 6375 25467 6381
rect 25409 6341 25421 6375
rect 25455 6341 25467 6375
rect 25409 6335 25467 6341
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6205 9459 6239
rect 10410 6236 10416 6248
rect 10371 6208 10416 6236
rect 9401 6199 9459 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11425 6239 11483 6245
rect 11425 6236 11437 6239
rect 11112 6208 11437 6236
rect 11112 6196 11118 6208
rect 11425 6205 11437 6208
rect 11471 6205 11483 6239
rect 13354 6236 13360 6248
rect 13315 6208 13360 6236
rect 11425 6199 11483 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 14366 6236 14372 6248
rect 14327 6208 14372 6236
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 14516 6208 15393 6236
rect 14516 6196 14522 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 16390 6236 16396 6248
rect 16351 6208 16396 6236
rect 15381 6199 15439 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 17402 6236 17408 6248
rect 17363 6208 17408 6236
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 18046 6196 18052 6248
rect 18104 6236 18110 6248
rect 18969 6239 19027 6245
rect 18969 6236 18981 6239
rect 18104 6208 18981 6236
rect 18104 6196 18110 6208
rect 18969 6205 18981 6208
rect 19015 6205 19027 6239
rect 18969 6199 19027 6205
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19392 6208 19993 6236
rect 19392 6196 19398 6208
rect 19981 6205 19993 6208
rect 20027 6205 20039 6239
rect 20990 6236 20996 6248
rect 20951 6208 20996 6236
rect 19981 6199 20039 6205
rect 20990 6196 20996 6208
rect 21048 6196 21054 6248
rect 22738 6236 22744 6248
rect 22699 6208 22744 6236
rect 22738 6196 22744 6208
rect 22796 6196 22802 6248
rect 24581 6239 24639 6245
rect 24581 6205 24593 6239
rect 24627 6236 24639 6239
rect 25424 6236 25452 6335
rect 25590 6236 25596 6248
rect 24627 6208 25452 6236
rect 25551 6208 25596 6236
rect 24627 6205 24639 6208
rect 24581 6199 24639 6205
rect 25590 6196 25596 6208
rect 25648 6196 25654 6248
rect 25682 6196 25688 6248
rect 25740 6236 25746 6248
rect 26605 6239 26663 6245
rect 26605 6236 26617 6239
rect 25740 6208 26617 6236
rect 25740 6196 25746 6208
rect 26605 6205 26617 6208
rect 26651 6205 26663 6239
rect 27614 6236 27620 6248
rect 27575 6208 27620 6236
rect 26605 6199 26663 6205
rect 27614 6196 27620 6208
rect 27672 6196 27678 6248
rect 28629 6239 28687 6245
rect 28629 6205 28641 6239
rect 28675 6205 28687 6239
rect 30190 6236 30196 6248
rect 30151 6208 30196 6236
rect 28629 6199 28687 6205
rect 28644 6168 28672 6199
rect 30190 6196 30196 6208
rect 30248 6196 30254 6248
rect 33962 6236 33968 6248
rect 33923 6208 33968 6236
rect 33962 6196 33968 6208
rect 34020 6196 34026 6248
rect 35805 6239 35863 6245
rect 35805 6205 35817 6239
rect 35851 6236 35863 6239
rect 35894 6236 35900 6248
rect 35851 6208 35900 6236
rect 35851 6205 35863 6208
rect 35805 6199 35863 6205
rect 35894 6196 35900 6208
rect 35952 6196 35958 6248
rect 36817 6239 36875 6245
rect 36817 6205 36829 6239
rect 36863 6205 36875 6239
rect 36817 6199 36875 6205
rect 34330 6168 34336 6180
rect 28644 6140 34336 6168
rect 34330 6128 34336 6140
rect 34388 6128 34394 6180
rect 36832 6168 36860 6199
rect 37182 6196 37188 6248
rect 37240 6236 37246 6248
rect 37921 6239 37979 6245
rect 37921 6236 37933 6239
rect 37240 6208 37933 6236
rect 37240 6196 37246 6208
rect 37921 6205 37933 6208
rect 37967 6205 37979 6239
rect 38930 6236 38936 6248
rect 38891 6208 38936 6236
rect 37921 6199 37979 6205
rect 38930 6196 38936 6208
rect 38988 6196 38994 6248
rect 38562 6168 38568 6180
rect 36832 6140 38568 6168
rect 38562 6128 38568 6140
rect 38620 6128 38626 6180
rect 3697 6103 3755 6109
rect 3697 6069 3709 6103
rect 3743 6100 3755 6103
rect 4982 6100 4988 6112
rect 3743 6072 4988 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 9824 6072 10241 6100
rect 9824 6060 9830 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10229 6063 10287 6069
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 11241 6103 11299 6109
rect 11241 6100 11253 6103
rect 10376 6072 11253 6100
rect 10376 6060 10382 6072
rect 11241 6069 11253 6072
rect 11287 6069 11299 6103
rect 11241 6063 11299 6069
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 13173 6103 13231 6109
rect 13173 6100 13185 6103
rect 11664 6072 13185 6100
rect 11664 6060 11670 6072
rect 13173 6069 13185 6072
rect 13219 6069 13231 6103
rect 13173 6063 13231 6069
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 13688 6072 14197 6100
rect 13688 6060 13694 6072
rect 14185 6069 14197 6072
rect 14231 6069 14243 6103
rect 14185 6063 14243 6069
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 17221 6103 17279 6109
rect 17221 6100 17233 6103
rect 16264 6072 17233 6100
rect 16264 6060 16270 6072
rect 17221 6069 17233 6072
rect 17267 6069 17279 6103
rect 17221 6063 17279 6069
rect 17402 6060 17408 6112
rect 17460 6100 17466 6112
rect 18785 6103 18843 6109
rect 18785 6100 18797 6103
rect 17460 6072 18797 6100
rect 17460 6060 17466 6072
rect 18785 6069 18797 6072
rect 18831 6069 18843 6103
rect 18785 6063 18843 6069
rect 19242 6060 19248 6112
rect 19300 6100 19306 6112
rect 19797 6103 19855 6109
rect 19797 6100 19809 6103
rect 19300 6072 19809 6100
rect 19300 6060 19306 6072
rect 19797 6069 19809 6072
rect 19843 6069 19855 6103
rect 19797 6063 19855 6069
rect 19886 6060 19892 6112
rect 19944 6100 19950 6112
rect 20809 6103 20867 6109
rect 20809 6100 20821 6103
rect 19944 6072 20821 6100
rect 19944 6060 19950 6072
rect 20809 6069 20821 6072
rect 20855 6069 20867 6103
rect 20809 6063 20867 6069
rect 20990 6060 20996 6112
rect 21048 6100 21054 6112
rect 24397 6103 24455 6109
rect 24397 6100 24409 6103
rect 21048 6072 24409 6100
rect 21048 6060 21054 6072
rect 24397 6069 24409 6072
rect 24443 6069 24455 6103
rect 24397 6063 24455 6069
rect 25866 6060 25872 6112
rect 25924 6100 25930 6112
rect 26421 6103 26479 6109
rect 26421 6100 26433 6103
rect 25924 6072 26433 6100
rect 25924 6060 25930 6072
rect 26421 6069 26433 6072
rect 26467 6069 26479 6103
rect 26421 6063 26479 6069
rect 26510 6060 26516 6112
rect 26568 6100 26574 6112
rect 27433 6103 27491 6109
rect 27433 6100 27445 6103
rect 26568 6072 27445 6100
rect 26568 6060 26574 6072
rect 27433 6069 27445 6072
rect 27479 6069 27491 6103
rect 27433 6063 27491 6069
rect 28445 6103 28503 6109
rect 28445 6069 28457 6103
rect 28491 6100 28503 6103
rect 29822 6100 29828 6112
rect 28491 6072 29828 6100
rect 28491 6069 28503 6072
rect 28445 6063 28503 6069
rect 29822 6060 29828 6072
rect 29880 6060 29886 6112
rect 30009 6103 30067 6109
rect 30009 6069 30021 6103
rect 30055 6100 30067 6103
rect 31478 6100 31484 6112
rect 30055 6072 31484 6100
rect 30055 6069 30067 6072
rect 30009 6063 30067 6069
rect 31478 6060 31484 6072
rect 31536 6060 31542 6112
rect 37274 6060 37280 6112
rect 37332 6100 37338 6112
rect 37737 6103 37795 6109
rect 37737 6100 37749 6103
rect 37332 6072 37749 6100
rect 37332 6060 37338 6072
rect 37737 6069 37749 6072
rect 37783 6069 37795 6103
rect 37737 6063 37795 6069
rect 38749 6103 38807 6109
rect 38749 6069 38761 6103
rect 38795 6100 38807 6103
rect 40034 6100 40040 6112
rect 38795 6072 40040 6100
rect 38795 6069 38807 6072
rect 38749 6063 38807 6069
rect 40034 6060 40040 6072
rect 40092 6060 40098 6112
rect 1104 6010 54832 6032
rect 1104 5958 18912 6010
rect 18964 5958 18976 6010
rect 19028 5958 19040 6010
rect 19092 5958 19104 6010
rect 19156 5958 36843 6010
rect 36895 5958 36907 6010
rect 36959 5958 36971 6010
rect 37023 5958 37035 6010
rect 37087 5958 54832 6010
rect 1104 5936 54832 5958
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 2314 5896 2320 5908
rect 2179 5868 2320 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 2924 5868 7849 5896
rect 2924 5856 2930 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 10410 5896 10416 5908
rect 10371 5868 10416 5896
rect 7837 5859 7895 5865
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 13446 5896 13452 5908
rect 13407 5868 13452 5896
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 14458 5896 14464 5908
rect 14419 5868 14464 5896
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 16025 5899 16083 5905
rect 16025 5865 16037 5899
rect 16071 5896 16083 5899
rect 16298 5896 16304 5908
rect 16071 5868 16304 5896
rect 16071 5865 16083 5868
rect 16025 5859 16083 5865
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 17037 5899 17095 5905
rect 17037 5865 17049 5899
rect 17083 5896 17095 5899
rect 17218 5896 17224 5908
rect 17083 5868 17224 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 18046 5896 18052 5908
rect 18007 5868 18052 5896
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 20070 5896 20076 5908
rect 20031 5868 20076 5896
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 21637 5899 21695 5905
rect 21637 5865 21649 5899
rect 21683 5896 21695 5899
rect 22462 5896 22468 5908
rect 21683 5868 22468 5896
rect 21683 5865 21695 5868
rect 21637 5859 21695 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 22649 5899 22707 5905
rect 22649 5865 22661 5899
rect 22695 5896 22707 5899
rect 22738 5896 22744 5908
rect 22695 5868 22744 5896
rect 22695 5865 22707 5868
rect 22649 5859 22707 5865
rect 22738 5856 22744 5868
rect 22796 5856 22802 5908
rect 24394 5896 24400 5908
rect 22848 5868 24400 5896
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 5592 5800 7052 5828
rect 5592 5788 5598 5800
rect 2314 5760 2320 5772
rect 2275 5732 2320 5760
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 4982 5760 4988 5772
rect 4943 5732 4988 5760
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 6043 5732 6592 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3844 5664 5856 5692
rect 3844 5652 3850 5664
rect 4798 5624 4804 5636
rect 4759 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 5828 5633 5856 5664
rect 5813 5627 5871 5633
rect 5813 5593 5825 5627
rect 5859 5593 5871 5627
rect 6564 5624 6592 5732
rect 6914 5720 6920 5772
rect 6972 5720 6978 5772
rect 7024 5769 7052 5800
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 9030 5760 9036 5772
rect 8991 5732 9036 5760
rect 8021 5723 8079 5729
rect 6932 5692 6960 5720
rect 8036 5692 8064 5723
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 10594 5760 10600 5772
rect 10555 5732 10600 5760
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 11606 5760 11612 5772
rect 11567 5732 11612 5760
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 12618 5760 12624 5772
rect 12579 5732 12624 5760
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 13630 5760 13636 5772
rect 13591 5732 13636 5760
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15286 5760 15292 5772
rect 14691 5732 15292 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 16206 5760 16212 5772
rect 16167 5732 16212 5760
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 17221 5763 17279 5769
rect 17221 5729 17233 5763
rect 17267 5760 17279 5763
rect 18138 5760 18144 5772
rect 17267 5732 18144 5760
rect 17267 5729 17279 5732
rect 17221 5723 17279 5729
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 18233 5763 18291 5769
rect 18233 5729 18245 5763
rect 18279 5760 18291 5763
rect 19242 5760 19248 5772
rect 18279 5732 19104 5760
rect 19203 5732 19248 5760
rect 18279 5729 18291 5732
rect 18233 5723 18291 5729
rect 6932 5664 8064 5692
rect 6825 5627 6883 5633
rect 6825 5624 6837 5627
rect 6564 5596 6837 5624
rect 5813 5587 5871 5593
rect 6825 5593 6837 5596
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 6914 5584 6920 5636
rect 6972 5624 6978 5636
rect 19076 5633 19104 5732
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 21821 5763 21879 5769
rect 21821 5729 21833 5763
rect 21867 5760 21879 5763
rect 22646 5760 22652 5772
rect 21867 5732 22652 5760
rect 21867 5729 21879 5732
rect 21821 5723 21879 5729
rect 22646 5720 22652 5732
rect 22704 5720 22710 5772
rect 22848 5769 22876 5868
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 24673 5899 24731 5905
rect 24673 5865 24685 5899
rect 24719 5896 24731 5899
rect 25590 5896 25596 5908
rect 24719 5868 25596 5896
rect 24719 5865 24731 5868
rect 24673 5859 24731 5865
rect 25590 5856 25596 5868
rect 25648 5856 25654 5908
rect 35345 5899 35403 5905
rect 35345 5865 35357 5899
rect 35391 5896 35403 5899
rect 36262 5896 36268 5908
rect 35391 5868 36268 5896
rect 35391 5865 35403 5868
rect 35345 5859 35403 5865
rect 36262 5856 36268 5868
rect 36320 5856 36326 5908
rect 36357 5899 36415 5905
rect 36357 5865 36369 5899
rect 36403 5896 36415 5899
rect 37182 5896 37188 5908
rect 36403 5868 37188 5896
rect 36403 5865 36415 5868
rect 36357 5859 36415 5865
rect 37182 5856 37188 5868
rect 37240 5856 37246 5908
rect 37369 5899 37427 5905
rect 37369 5865 37381 5899
rect 37415 5865 37427 5899
rect 40494 5896 40500 5908
rect 40455 5868 40500 5896
rect 37369 5859 37427 5865
rect 37384 5828 37412 5859
rect 40494 5856 40500 5868
rect 40552 5856 40558 5908
rect 37384 5800 38700 5828
rect 22833 5763 22891 5769
rect 22833 5729 22845 5763
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 23842 5720 23848 5772
rect 23900 5769 23906 5772
rect 23900 5760 23911 5769
rect 24854 5760 24860 5772
rect 23900 5732 23945 5760
rect 24815 5732 24860 5760
rect 23900 5723 23911 5732
rect 23900 5720 23906 5723
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 25866 5760 25872 5772
rect 25827 5732 25872 5760
rect 25866 5720 25872 5732
rect 25924 5720 25930 5772
rect 26329 5763 26387 5769
rect 26329 5729 26341 5763
rect 26375 5760 26387 5763
rect 27433 5763 27491 5769
rect 27433 5760 27445 5763
rect 26375 5732 27445 5760
rect 26375 5729 26387 5732
rect 26329 5723 26387 5729
rect 27433 5729 27445 5732
rect 27479 5729 27491 5763
rect 27433 5723 27491 5729
rect 28445 5763 28503 5769
rect 28445 5729 28457 5763
rect 28491 5729 28503 5763
rect 28445 5723 28503 5729
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 28460 5692 28488 5723
rect 29086 5720 29092 5772
rect 29144 5760 29150 5772
rect 29457 5763 29515 5769
rect 29457 5760 29469 5763
rect 29144 5732 29469 5760
rect 29144 5720 29150 5732
rect 29457 5729 29469 5732
rect 29503 5729 29515 5763
rect 30466 5760 30472 5772
rect 30427 5732 30472 5760
rect 29457 5723 29515 5729
rect 30466 5720 30472 5732
rect 30524 5720 30530 5772
rect 35529 5763 35587 5769
rect 35529 5729 35541 5763
rect 35575 5760 35587 5763
rect 35986 5760 35992 5772
rect 35575 5732 35992 5760
rect 35575 5729 35587 5732
rect 35529 5723 35587 5729
rect 35986 5720 35992 5732
rect 36044 5720 36050 5772
rect 36541 5763 36599 5769
rect 36541 5729 36553 5763
rect 36587 5729 36599 5763
rect 36541 5723 36599 5729
rect 24820 5664 28488 5692
rect 36556 5692 36584 5723
rect 37366 5720 37372 5772
rect 37424 5760 37430 5772
rect 38672 5769 38700 5800
rect 39850 5788 39856 5840
rect 39908 5828 39914 5840
rect 39908 5800 40724 5828
rect 39908 5788 39914 5800
rect 37553 5763 37611 5769
rect 37553 5760 37565 5763
rect 37424 5732 37565 5760
rect 37424 5720 37430 5732
rect 37553 5729 37565 5732
rect 37599 5729 37611 5763
rect 37553 5723 37611 5729
rect 38657 5763 38715 5769
rect 38657 5729 38669 5763
rect 38703 5729 38715 5763
rect 38657 5723 38715 5729
rect 39669 5763 39727 5769
rect 39669 5729 39681 5763
rect 39715 5760 39727 5763
rect 40586 5760 40592 5772
rect 39715 5732 40592 5760
rect 39715 5729 39727 5732
rect 39669 5723 39727 5729
rect 40586 5720 40592 5732
rect 40644 5720 40650 5772
rect 40696 5769 40724 5800
rect 40681 5763 40739 5769
rect 40681 5729 40693 5763
rect 40727 5729 40739 5763
rect 40681 5723 40739 5729
rect 36556 5664 39528 5692
rect 24820 5652 24826 5664
rect 8849 5627 8907 5633
rect 8849 5624 8861 5627
rect 6972 5596 8861 5624
rect 6972 5584 6978 5596
rect 8849 5593 8861 5596
rect 8895 5593 8907 5627
rect 8849 5587 8907 5593
rect 19061 5627 19119 5633
rect 19061 5593 19073 5627
rect 19107 5593 19119 5627
rect 19061 5587 19119 5593
rect 22922 5584 22928 5636
rect 22980 5624 22986 5636
rect 22980 5596 23796 5624
rect 22980 5584 22986 5596
rect 11422 5556 11428 5568
rect 11383 5528 11428 5556
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 23658 5556 23664 5568
rect 12492 5528 12537 5556
rect 23619 5528 23664 5556
rect 12492 5516 12498 5528
rect 23658 5516 23664 5528
rect 23716 5516 23722 5568
rect 23768 5556 23796 5596
rect 23842 5584 23848 5636
rect 23900 5624 23906 5636
rect 39500 5633 39528 5664
rect 25685 5627 25743 5633
rect 25685 5624 25697 5627
rect 23900 5596 25697 5624
rect 23900 5584 23906 5596
rect 25685 5593 25697 5596
rect 25731 5593 25743 5627
rect 25685 5587 25743 5593
rect 39485 5627 39543 5633
rect 39485 5593 39497 5627
rect 39531 5593 39543 5627
rect 39485 5587 39543 5593
rect 26329 5559 26387 5565
rect 26329 5556 26341 5559
rect 23768 5528 26341 5556
rect 26329 5525 26341 5528
rect 26375 5525 26387 5559
rect 26329 5519 26387 5525
rect 26602 5516 26608 5568
rect 26660 5556 26666 5568
rect 27249 5559 27307 5565
rect 27249 5556 27261 5559
rect 26660 5528 27261 5556
rect 26660 5516 26666 5528
rect 27249 5525 27261 5528
rect 27295 5525 27307 5559
rect 27249 5519 27307 5525
rect 27338 5516 27344 5568
rect 27396 5556 27402 5568
rect 28261 5559 28319 5565
rect 28261 5556 28273 5559
rect 27396 5528 28273 5556
rect 27396 5516 27402 5528
rect 28261 5525 28273 5528
rect 28307 5525 28319 5559
rect 29270 5556 29276 5568
rect 29231 5528 29276 5556
rect 28261 5519 28319 5525
rect 29270 5516 29276 5528
rect 29328 5516 29334 5568
rect 30285 5559 30343 5565
rect 30285 5525 30297 5559
rect 30331 5556 30343 5559
rect 34514 5556 34520 5568
rect 30331 5528 34520 5556
rect 30331 5525 30343 5528
rect 30285 5519 30343 5525
rect 34514 5516 34520 5528
rect 34572 5516 34578 5568
rect 37550 5516 37556 5568
rect 37608 5556 37614 5568
rect 38473 5559 38531 5565
rect 38473 5556 38485 5559
rect 37608 5528 38485 5556
rect 37608 5516 37614 5528
rect 38473 5525 38485 5528
rect 38519 5525 38531 5559
rect 38473 5519 38531 5525
rect 1104 5466 54832 5488
rect 1104 5414 9947 5466
rect 9999 5414 10011 5466
rect 10063 5414 10075 5466
rect 10127 5414 10139 5466
rect 10191 5414 27878 5466
rect 27930 5414 27942 5466
rect 27994 5414 28006 5466
rect 28058 5414 28070 5466
rect 28122 5414 45808 5466
rect 45860 5414 45872 5466
rect 45924 5414 45936 5466
rect 45988 5414 46000 5466
rect 46052 5414 54832 5466
rect 1104 5392 54832 5414
rect 2130 5352 2136 5364
rect 2091 5324 2136 5352
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5534 5352 5540 5364
rect 5215 5324 5540 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 9030 5352 9036 5364
rect 8619 5324 9036 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 11054 5352 11060 5364
rect 10643 5324 11060 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11609 5355 11667 5361
rect 11609 5321 11621 5355
rect 11655 5352 11667 5355
rect 13354 5352 13360 5364
rect 11655 5324 13360 5352
rect 11655 5321 11667 5324
rect 11609 5315 11667 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 16117 5355 16175 5361
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 16574 5352 16580 5364
rect 16163 5324 16580 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 18782 5352 18788 5364
rect 18743 5324 18788 5352
rect 18782 5312 18788 5324
rect 18840 5312 18846 5364
rect 21085 5355 21143 5361
rect 21085 5321 21097 5355
rect 21131 5352 21143 5355
rect 21818 5352 21824 5364
rect 21131 5324 21824 5352
rect 21131 5321 21143 5324
rect 21085 5315 21143 5321
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 24397 5355 24455 5361
rect 24397 5321 24409 5355
rect 24443 5352 24455 5355
rect 25682 5352 25688 5364
rect 24443 5324 25688 5352
rect 24443 5321 24455 5324
rect 24397 5315 24455 5321
rect 25682 5312 25688 5324
rect 25740 5312 25746 5364
rect 36357 5355 36415 5361
rect 36357 5321 36369 5355
rect 36403 5352 36415 5355
rect 37366 5352 37372 5364
rect 36403 5324 37372 5352
rect 36403 5321 36415 5324
rect 36357 5315 36415 5321
rect 37366 5312 37372 5324
rect 37424 5312 37430 5364
rect 38562 5312 38568 5364
rect 38620 5352 38626 5364
rect 41233 5355 41291 5361
rect 41233 5352 41245 5355
rect 38620 5324 41245 5352
rect 38620 5312 38626 5324
rect 41233 5321 41245 5324
rect 41279 5321 41291 5355
rect 41233 5315 41291 5321
rect 13173 5287 13231 5293
rect 13173 5253 13185 5287
rect 13219 5284 13231 5287
rect 13538 5284 13544 5296
rect 13219 5256 13544 5284
rect 13219 5253 13231 5256
rect 13173 5247 13231 5253
rect 13538 5244 13544 5256
rect 13596 5244 13602 5296
rect 15105 5287 15163 5293
rect 15105 5253 15117 5287
rect 15151 5284 15163 5287
rect 20806 5284 20812 5296
rect 15151 5256 20812 5284
rect 15151 5253 15163 5256
rect 15105 5247 15163 5253
rect 20806 5244 20812 5256
rect 20864 5244 20870 5296
rect 22097 5287 22155 5293
rect 22097 5253 22109 5287
rect 22143 5253 22155 5287
rect 22097 5247 22155 5253
rect 30009 5287 30067 5293
rect 30009 5253 30021 5287
rect 30055 5284 30067 5287
rect 33502 5284 33508 5296
rect 30055 5256 33508 5284
rect 30055 5253 30067 5256
rect 30009 5247 30067 5253
rect 10502 5216 10508 5228
rect 8772 5188 10508 5216
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5117 2375 5151
rect 5350 5148 5356 5160
rect 5311 5120 5356 5148
rect 2317 5111 2375 5117
rect 2332 5080 2360 5111
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 8772 5157 8800 5188
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 15194 5216 15200 5228
rect 13372 5188 15200 5216
rect 7745 5151 7803 5157
rect 7745 5148 7757 5151
rect 6420 5120 7757 5148
rect 6420 5108 6426 5120
rect 7745 5117 7757 5120
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5117 8815 5151
rect 9766 5148 9772 5160
rect 9727 5120 9772 5148
rect 8757 5111 8815 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5148 10839 5151
rect 11422 5148 11428 5160
rect 10827 5120 11428 5148
rect 10827 5117 10839 5120
rect 10781 5111 10839 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5148 11851 5151
rect 12434 5148 12440 5160
rect 11839 5120 12440 5148
rect 11839 5117 11851 5120
rect 11793 5111 11851 5117
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 13372 5157 13400 5188
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 22112 5216 22140 5247
rect 33502 5244 33508 5256
rect 33560 5244 33566 5296
rect 29270 5216 29276 5228
rect 19996 5188 22140 5216
rect 27632 5188 29276 5216
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5117 13415 5151
rect 13357 5111 13415 5117
rect 14090 5108 14096 5160
rect 14148 5148 14154 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 14148 5120 15301 5148
rect 14148 5108 14154 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 16301 5151 16359 5157
rect 16301 5117 16313 5151
rect 16347 5148 16359 5151
rect 17402 5148 17408 5160
rect 16347 5120 17408 5148
rect 16347 5117 16359 5120
rect 16301 5111 16359 5117
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 18969 5151 19027 5157
rect 18969 5117 18981 5151
rect 19015 5148 19027 5151
rect 19886 5148 19892 5160
rect 19015 5120 19892 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 19996 5157 20024 5188
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5117 21327 5151
rect 22278 5148 22284 5160
rect 22239 5120 22284 5148
rect 21269 5111 21327 5117
rect 6454 5080 6460 5092
rect 2332 5052 6460 5080
rect 6454 5040 6460 5052
rect 6512 5040 6518 5092
rect 21284 5080 21312 5111
rect 22278 5108 22284 5120
rect 22336 5108 22342 5160
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5117 23351 5151
rect 23293 5111 23351 5117
rect 19812 5052 21312 5080
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 5592 4984 7573 5012
rect 5592 4972 5598 4984
rect 7561 4981 7573 4984
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 19812 5021 19840 5052
rect 22186 5040 22192 5092
rect 22244 5080 22250 5092
rect 23308 5080 23336 5111
rect 23382 5108 23388 5160
rect 23440 5148 23446 5160
rect 24581 5151 24639 5157
rect 24581 5148 24593 5151
rect 23440 5120 24593 5148
rect 23440 5108 23446 5120
rect 24581 5117 24593 5120
rect 24627 5117 24639 5151
rect 24581 5111 24639 5117
rect 24946 5108 24952 5160
rect 25004 5148 25010 5160
rect 25593 5151 25651 5157
rect 25593 5148 25605 5151
rect 25004 5120 25605 5148
rect 25004 5108 25010 5120
rect 25593 5117 25605 5120
rect 25639 5117 25651 5151
rect 26602 5148 26608 5160
rect 26563 5120 26608 5148
rect 25593 5111 25651 5117
rect 26602 5108 26608 5120
rect 26660 5108 26666 5160
rect 27632 5157 27660 5188
rect 29270 5176 29276 5188
rect 29328 5176 29334 5228
rect 29822 5176 29828 5228
rect 29880 5216 29886 5228
rect 29880 5188 31248 5216
rect 29880 5176 29886 5188
rect 27617 5151 27675 5157
rect 27617 5117 27629 5151
rect 27663 5117 27675 5151
rect 27617 5111 27675 5117
rect 27706 5108 27712 5160
rect 27764 5148 27770 5160
rect 28629 5151 28687 5157
rect 28629 5148 28641 5151
rect 27764 5120 28641 5148
rect 27764 5108 27770 5120
rect 28629 5117 28641 5120
rect 28675 5117 28687 5151
rect 28629 5111 28687 5117
rect 29178 5108 29184 5160
rect 29236 5148 29242 5160
rect 31220 5157 31248 5188
rect 30193 5151 30251 5157
rect 30193 5148 30205 5151
rect 29236 5120 30205 5148
rect 29236 5108 29242 5120
rect 30193 5117 30205 5120
rect 30239 5117 30251 5151
rect 30193 5111 30251 5117
rect 31205 5151 31263 5157
rect 31205 5117 31217 5151
rect 31251 5117 31263 5151
rect 31205 5111 31263 5117
rect 36541 5151 36599 5157
rect 36541 5117 36553 5151
rect 36587 5148 36599 5151
rect 37274 5148 37280 5160
rect 36587 5120 37280 5148
rect 36587 5117 36599 5120
rect 36541 5111 36599 5117
rect 37274 5108 37280 5120
rect 37332 5108 37338 5160
rect 37550 5148 37556 5160
rect 37511 5120 37556 5148
rect 37550 5108 37556 5120
rect 37608 5108 37614 5160
rect 38565 5151 38623 5157
rect 38565 5117 38577 5151
rect 38611 5117 38623 5151
rect 38565 5111 38623 5117
rect 38580 5080 38608 5111
rect 38746 5108 38752 5160
rect 38804 5148 38810 5160
rect 39577 5151 39635 5157
rect 39577 5148 39589 5151
rect 38804 5120 39589 5148
rect 38804 5108 38810 5120
rect 39577 5117 39589 5120
rect 39623 5117 39635 5151
rect 39577 5111 39635 5117
rect 40034 5108 40040 5160
rect 40092 5148 40098 5160
rect 41417 5151 41475 5157
rect 41417 5148 41429 5151
rect 40092 5120 41429 5148
rect 40092 5108 40098 5120
rect 41417 5117 41429 5120
rect 41463 5117 41475 5151
rect 41417 5111 41475 5117
rect 22244 5052 23336 5080
rect 37384 5052 38608 5080
rect 22244 5040 22250 5052
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 7708 4984 9597 5012
rect 7708 4972 7714 4984
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 19797 5015 19855 5021
rect 19797 4981 19809 5015
rect 19843 4981 19855 5015
rect 19797 4975 19855 4981
rect 21818 4972 21824 5024
rect 21876 5012 21882 5024
rect 23109 5015 23167 5021
rect 23109 5012 23121 5015
rect 21876 4984 23121 5012
rect 21876 4972 21882 4984
rect 23109 4981 23121 4984
rect 23155 4981 23167 5015
rect 23109 4975 23167 4981
rect 24486 4972 24492 5024
rect 24544 5012 24550 5024
rect 25409 5015 25467 5021
rect 25409 5012 25421 5015
rect 24544 4984 25421 5012
rect 24544 4972 24550 4984
rect 25409 4981 25421 4984
rect 25455 4981 25467 5015
rect 25409 4975 25467 4981
rect 25498 4972 25504 5024
rect 25556 5012 25562 5024
rect 26421 5015 26479 5021
rect 26421 5012 26433 5015
rect 25556 4984 26433 5012
rect 25556 4972 25562 4984
rect 26421 4981 26433 4984
rect 26467 4981 26479 5015
rect 26421 4975 26479 4981
rect 26602 4972 26608 5024
rect 26660 5012 26666 5024
rect 27433 5015 27491 5021
rect 27433 5012 27445 5015
rect 26660 4984 27445 5012
rect 26660 4972 26666 4984
rect 27433 4981 27445 4984
rect 27479 4981 27491 5015
rect 27433 4975 27491 4981
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 28445 5015 28503 5021
rect 28445 5012 28457 5015
rect 27580 4984 28457 5012
rect 27580 4972 27586 4984
rect 28445 4981 28457 4984
rect 28491 4981 28503 5015
rect 28445 4975 28503 4981
rect 30374 4972 30380 5024
rect 30432 5012 30438 5024
rect 37384 5021 37412 5052
rect 31021 5015 31079 5021
rect 31021 5012 31033 5015
rect 30432 4984 31033 5012
rect 30432 4972 30438 4984
rect 31021 4981 31033 4984
rect 31067 4981 31079 5015
rect 31021 4975 31079 4981
rect 37369 5015 37427 5021
rect 37369 4981 37381 5015
rect 37415 4981 37427 5015
rect 37369 4975 37427 4981
rect 37550 4972 37556 5024
rect 37608 5012 37614 5024
rect 38381 5015 38439 5021
rect 38381 5012 38393 5015
rect 37608 4984 38393 5012
rect 37608 4972 37614 4984
rect 38381 4981 38393 4984
rect 38427 4981 38439 5015
rect 39390 5012 39396 5024
rect 39351 4984 39396 5012
rect 38381 4975 38439 4981
rect 39390 4972 39396 4984
rect 39448 4972 39454 5024
rect 1104 4922 54832 4944
rect 1104 4870 18912 4922
rect 18964 4870 18976 4922
rect 19028 4870 19040 4922
rect 19092 4870 19104 4922
rect 19156 4870 36843 4922
rect 36895 4870 36907 4922
rect 36959 4870 36971 4922
rect 37023 4870 37035 4922
rect 37087 4870 54832 4922
rect 1104 4848 54832 4870
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 10594 4808 10600 4820
rect 8435 4780 10600 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 15930 4808 15936 4820
rect 15891 4780 15936 4808
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 17865 4811 17923 4817
rect 17865 4777 17877 4811
rect 17911 4808 17923 4811
rect 18322 4808 18328 4820
rect 17911 4780 18328 4808
rect 17911 4777 17923 4780
rect 17865 4771 17923 4777
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 18877 4811 18935 4817
rect 18877 4777 18889 4811
rect 18923 4808 18935 4811
rect 22278 4808 22284 4820
rect 18923 4780 22284 4808
rect 18923 4777 18935 4780
rect 18877 4771 18935 4777
rect 22278 4768 22284 4780
rect 22336 4768 22342 4820
rect 22649 4811 22707 4817
rect 22649 4777 22661 4811
rect 22695 4808 22707 4811
rect 23474 4808 23480 4820
rect 22695 4780 23480 4808
rect 22695 4777 22707 4780
rect 22649 4771 22707 4777
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 24946 4808 24952 4820
rect 24907 4780 24952 4808
rect 24946 4768 24952 4780
rect 25004 4768 25010 4820
rect 30466 4768 30472 4820
rect 30524 4808 30530 4820
rect 31297 4811 31355 4817
rect 31297 4808 31309 4811
rect 30524 4780 31309 4808
rect 30524 4768 30530 4780
rect 31297 4777 31309 4780
rect 31343 4777 31355 4811
rect 38746 4808 38752 4820
rect 38707 4780 38752 4808
rect 31297 4771 31355 4777
rect 38746 4768 38752 4780
rect 38804 4768 38810 4820
rect 40586 4768 40592 4820
rect 40644 4808 40650 4820
rect 40773 4811 40831 4817
rect 40773 4808 40785 4811
rect 40644 4780 40785 4808
rect 40644 4768 40650 4780
rect 40773 4777 40785 4780
rect 40819 4777 40831 4811
rect 40773 4771 40831 4777
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 6914 4672 6920 4684
rect 6595 4644 6920 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4672 7619 4675
rect 7650 4672 7656 4684
rect 7607 4644 7656 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 10318 4672 10324 4684
rect 8619 4644 10324 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 14274 4672 14280 4684
rect 14235 4644 14280 4672
rect 14274 4632 14280 4644
rect 14332 4632 14338 4684
rect 15948 4672 15976 4768
rect 23658 4740 23664 4752
rect 20640 4712 23664 4740
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 15948 4644 16221 4672
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16209 4635 16267 4641
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4641 18107 4675
rect 19058 4672 19064 4684
rect 19019 4644 19064 4672
rect 18049 4635 18107 4641
rect 18064 4604 18092 4635
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 20640 4681 20668 4712
rect 23658 4700 23664 4712
rect 23716 4700 23722 4752
rect 26510 4740 26516 4752
rect 25148 4712 26516 4740
rect 20625 4675 20683 4681
rect 20625 4641 20637 4675
rect 20671 4641 20683 4675
rect 21818 4672 21824 4684
rect 21779 4644 21824 4672
rect 20625 4635 20683 4641
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 22830 4672 22836 4684
rect 22791 4644 22836 4672
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 23845 4675 23903 4681
rect 23845 4641 23857 4675
rect 23891 4672 23903 4675
rect 24486 4672 24492 4684
rect 23891 4644 24492 4672
rect 23891 4641 23903 4644
rect 23845 4635 23903 4641
rect 24486 4632 24492 4644
rect 24544 4632 24550 4684
rect 25148 4681 25176 4712
rect 26510 4700 26516 4712
rect 26568 4700 26574 4752
rect 38838 4700 38844 4752
rect 38896 4740 38902 4752
rect 38896 4712 41000 4740
rect 38896 4700 38902 4712
rect 25133 4675 25191 4681
rect 25133 4641 25145 4675
rect 25179 4641 25191 4675
rect 25133 4635 25191 4641
rect 26145 4675 26203 4681
rect 26145 4641 26157 4675
rect 26191 4672 26203 4675
rect 27338 4672 27344 4684
rect 26191 4644 27344 4672
rect 26191 4641 26203 4644
rect 26145 4635 26203 4641
rect 27338 4632 27344 4644
rect 27396 4632 27402 4684
rect 27433 4675 27491 4681
rect 27433 4641 27445 4675
rect 27479 4672 27491 4675
rect 27522 4672 27528 4684
rect 27479 4644 27528 4672
rect 27479 4641 27491 4644
rect 27433 4635 27491 4641
rect 27522 4632 27528 4644
rect 27580 4632 27586 4684
rect 28445 4675 28503 4681
rect 28445 4641 28457 4675
rect 28491 4641 28503 4675
rect 28445 4635 28503 4641
rect 18064 4576 20484 4604
rect 5353 4539 5411 4545
rect 5353 4505 5365 4539
rect 5399 4536 5411 4539
rect 6822 4536 6828 4548
rect 5399 4508 6828 4536
rect 5399 4505 5411 4508
rect 5353 4499 5411 4505
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 7377 4539 7435 4545
rect 7377 4505 7389 4539
rect 7423 4536 7435 4539
rect 11146 4536 11152 4548
rect 7423 4508 11152 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 16025 4539 16083 4545
rect 16025 4505 16037 4539
rect 16071 4536 16083 4539
rect 18598 4536 18604 4548
rect 16071 4508 18604 4536
rect 16071 4505 16083 4508
rect 16025 4499 16083 4505
rect 18598 4496 18604 4508
rect 18656 4496 18662 4548
rect 20456 4545 20484 4576
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 28460 4604 28488 4635
rect 28994 4632 29000 4684
rect 29052 4672 29058 4684
rect 29457 4675 29515 4681
rect 29457 4672 29469 4675
rect 29052 4644 29469 4672
rect 29052 4632 29058 4644
rect 29457 4641 29469 4644
rect 29503 4641 29515 4675
rect 30466 4672 30472 4684
rect 30427 4644 30472 4672
rect 29457 4635 29515 4641
rect 30466 4632 30472 4644
rect 30524 4632 30530 4684
rect 31478 4672 31484 4684
rect 31439 4644 31484 4672
rect 31478 4632 31484 4644
rect 31536 4632 31542 4684
rect 33042 4672 33048 4684
rect 33003 4644 33048 4672
rect 33042 4632 33048 4644
rect 33100 4632 33106 4684
rect 35805 4675 35863 4681
rect 35805 4641 35817 4675
rect 35851 4672 35863 4675
rect 36170 4672 36176 4684
rect 35851 4644 36176 4672
rect 35851 4641 35863 4644
rect 35805 4635 35863 4641
rect 36170 4632 36176 4644
rect 36228 4632 36234 4684
rect 37550 4672 37556 4684
rect 37511 4644 37556 4672
rect 37550 4632 37556 4644
rect 37608 4632 37614 4684
rect 38933 4675 38991 4681
rect 38933 4641 38945 4675
rect 38979 4641 38991 4675
rect 38933 4635 38991 4641
rect 39945 4675 40003 4681
rect 39945 4641 39957 4675
rect 39991 4672 40003 4675
rect 40678 4672 40684 4684
rect 39991 4644 40684 4672
rect 39991 4641 40003 4644
rect 39945 4635 40003 4641
rect 38948 4604 38976 4635
rect 40678 4632 40684 4644
rect 40736 4632 40742 4684
rect 40972 4681 41000 4712
rect 40957 4675 41015 4681
rect 40957 4641 40969 4675
rect 41003 4641 41015 4675
rect 40957 4635 41015 4641
rect 26384 4576 28488 4604
rect 37384 4576 38976 4604
rect 26384 4564 26390 4576
rect 37384 4545 37412 4576
rect 20441 4539 20499 4545
rect 20441 4505 20453 4539
rect 20487 4505 20499 4539
rect 20441 4499 20499 4505
rect 37369 4539 37427 4545
rect 37369 4505 37381 4539
rect 37415 4505 37427 4539
rect 37369 4499 37427 4505
rect 13081 4471 13139 4477
rect 13081 4437 13093 4471
rect 13127 4468 13139 4471
rect 14182 4468 14188 4480
rect 13127 4440 14188 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 21637 4471 21695 4477
rect 21637 4468 21649 4471
rect 20864 4440 21649 4468
rect 20864 4428 20870 4440
rect 21637 4437 21649 4440
rect 21683 4437 21695 4471
rect 21637 4431 21695 4437
rect 22738 4428 22744 4480
rect 22796 4468 22802 4480
rect 23661 4471 23719 4477
rect 23661 4468 23673 4471
rect 22796 4440 23673 4468
rect 22796 4428 22802 4440
rect 23661 4437 23673 4440
rect 23707 4437 23719 4471
rect 23661 4431 23719 4437
rect 25590 4428 25596 4480
rect 25648 4468 25654 4480
rect 25961 4471 26019 4477
rect 25961 4468 25973 4471
rect 25648 4440 25973 4468
rect 25648 4428 25654 4440
rect 25961 4437 25973 4440
rect 26007 4437 26019 4471
rect 25961 4431 26019 4437
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 27249 4471 27307 4477
rect 27249 4468 27261 4471
rect 26292 4440 27261 4468
rect 26292 4428 26298 4440
rect 27249 4437 27261 4440
rect 27295 4437 27307 4471
rect 27249 4431 27307 4437
rect 27614 4428 27620 4480
rect 27672 4468 27678 4480
rect 28261 4471 28319 4477
rect 28261 4468 28273 4471
rect 27672 4440 28273 4468
rect 27672 4428 27678 4440
rect 28261 4437 28273 4440
rect 28307 4437 28319 4471
rect 28261 4431 28319 4437
rect 28350 4428 28356 4480
rect 28408 4468 28414 4480
rect 29273 4471 29331 4477
rect 29273 4468 29285 4471
rect 28408 4440 29285 4468
rect 28408 4428 28414 4440
rect 29273 4437 29285 4440
rect 29319 4437 29331 4471
rect 29273 4431 29331 4437
rect 29454 4428 29460 4480
rect 29512 4468 29518 4480
rect 30285 4471 30343 4477
rect 30285 4468 30297 4471
rect 29512 4440 30297 4468
rect 29512 4428 29518 4440
rect 30285 4437 30297 4440
rect 30331 4437 30343 4471
rect 30285 4431 30343 4437
rect 32861 4471 32919 4477
rect 32861 4437 32873 4471
rect 32907 4468 32919 4471
rect 34054 4468 34060 4480
rect 32907 4440 34060 4468
rect 32907 4437 32919 4440
rect 32861 4431 32919 4437
rect 34054 4428 34060 4440
rect 34112 4428 34118 4480
rect 35621 4471 35679 4477
rect 35621 4437 35633 4471
rect 35667 4468 35679 4471
rect 36538 4468 36544 4480
rect 35667 4440 36544 4468
rect 35667 4437 35679 4440
rect 35621 4431 35679 4437
rect 36538 4428 36544 4440
rect 36596 4428 36602 4480
rect 39761 4471 39819 4477
rect 39761 4437 39773 4471
rect 39807 4468 39819 4471
rect 40586 4468 40592 4480
rect 39807 4440 40592 4468
rect 39807 4437 39819 4440
rect 39761 4431 39819 4437
rect 40586 4428 40592 4440
rect 40644 4428 40650 4480
rect 1104 4378 54832 4400
rect 1104 4326 9947 4378
rect 9999 4326 10011 4378
rect 10063 4326 10075 4378
rect 10127 4326 10139 4378
rect 10191 4326 27878 4378
rect 27930 4326 27942 4378
rect 27994 4326 28006 4378
rect 28058 4326 28070 4378
rect 28122 4326 45808 4378
rect 45860 4326 45872 4378
rect 45924 4326 45936 4378
rect 45988 4326 46000 4378
rect 46052 4326 54832 4378
rect 1104 4304 54832 4326
rect 6454 4264 6460 4276
rect 6415 4236 6460 4264
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 13173 4267 13231 4273
rect 13173 4233 13185 4267
rect 13219 4264 13231 4267
rect 13262 4264 13268 4276
rect 13219 4236 13268 4264
rect 13219 4233 13231 4236
rect 13173 4227 13231 4233
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 14185 4267 14243 4273
rect 14185 4233 14197 4267
rect 14231 4264 14243 4267
rect 14274 4264 14280 4276
rect 14231 4236 14280 4264
rect 14231 4233 14243 4236
rect 14185 4227 14243 4233
rect 14274 4224 14280 4236
rect 14332 4224 14338 4276
rect 18785 4267 18843 4273
rect 18785 4233 18797 4267
rect 18831 4264 18843 4267
rect 19058 4264 19064 4276
rect 18831 4236 19064 4264
rect 18831 4233 18843 4236
rect 18785 4227 18843 4233
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 22465 4267 22523 4273
rect 22465 4233 22477 4267
rect 22511 4264 22523 4267
rect 22830 4264 22836 4276
rect 22511 4236 22836 4264
rect 22511 4233 22523 4236
rect 22465 4227 22523 4233
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 32677 4267 32735 4273
rect 32677 4233 32689 4267
rect 32723 4264 32735 4267
rect 33042 4264 33048 4276
rect 32723 4236 33048 4264
rect 32723 4233 32735 4236
rect 32677 4227 32735 4233
rect 33042 4224 33048 4236
rect 33100 4224 33106 4276
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 7837 4199 7895 4205
rect 7837 4196 7849 4199
rect 2372 4168 7849 4196
rect 2372 4156 2378 4168
rect 7837 4165 7849 4168
rect 7883 4165 7895 4199
rect 7837 4159 7895 4165
rect 25498 4128 25504 4140
rect 24596 4100 25504 4128
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6641 4063 6699 4069
rect 6641 4060 6653 4063
rect 6328 4032 6653 4060
rect 6328 4020 6334 4032
rect 6641 4029 6653 4032
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8202 4060 8208 4072
rect 8067 4032 8208 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 13722 4060 13728 4072
rect 13403 4032 13728 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 14056 4032 14381 4060
rect 14056 4020 14062 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16574 4060 16580 4072
rect 15611 4032 16436 4060
rect 16535 4032 16580 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 16408 3933 16436 4032
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 18506 4020 18512 4072
rect 18564 4060 18570 4072
rect 18969 4063 19027 4069
rect 18969 4060 18981 4063
rect 18564 4032 18981 4060
rect 18564 4020 18570 4032
rect 18969 4029 18981 4032
rect 19015 4029 19027 4063
rect 18969 4023 19027 4029
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20806 4060 20812 4072
rect 20027 4032 20812 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 20990 4060 20996 4072
rect 20951 4032 20996 4060
rect 20990 4020 20996 4032
rect 21048 4020 21054 4072
rect 22649 4063 22707 4069
rect 22649 4029 22661 4063
rect 22695 4060 22707 4063
rect 23842 4060 23848 4072
rect 22695 4032 23848 4060
rect 22695 4029 22707 4032
rect 22649 4023 22707 4029
rect 23842 4020 23848 4032
rect 23900 4020 23906 4072
rect 24596 4069 24624 4100
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 24581 4063 24639 4069
rect 24581 4029 24593 4063
rect 24627 4029 24639 4063
rect 25590 4060 25596 4072
rect 25551 4032 25596 4060
rect 24581 4023 24639 4029
rect 25590 4020 25596 4032
rect 25648 4020 25654 4072
rect 26602 4060 26608 4072
rect 26563 4032 26608 4060
rect 26602 4020 26608 4032
rect 26660 4020 26666 4072
rect 27614 4060 27620 4072
rect 27575 4032 27620 4060
rect 27614 4020 27620 4032
rect 27672 4020 27678 4072
rect 28258 4020 28264 4072
rect 28316 4060 28322 4072
rect 28629 4063 28687 4069
rect 28629 4060 28641 4063
rect 28316 4032 28641 4060
rect 28316 4020 28322 4032
rect 28629 4029 28641 4032
rect 28675 4029 28687 4063
rect 28629 4023 28687 4029
rect 30837 4063 30895 4069
rect 30837 4029 30849 4063
rect 30883 4029 30895 4063
rect 31846 4060 31852 4072
rect 31807 4032 31852 4060
rect 30837 4023 30895 4029
rect 22186 3992 22192 4004
rect 20824 3964 22192 3992
rect 15381 3927 15439 3933
rect 15381 3924 15393 3927
rect 14792 3896 15393 3924
rect 14792 3884 14798 3896
rect 15381 3893 15393 3896
rect 15427 3893 15439 3927
rect 15381 3887 15439 3893
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3893 16451 3927
rect 19794 3924 19800 3936
rect 19755 3896 19800 3924
rect 16393 3887 16451 3893
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 20824 3933 20852 3964
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 30852 3992 30880 4023
rect 31846 4020 31852 4032
rect 31904 4020 31910 4072
rect 32861 4063 32919 4069
rect 32861 4029 32873 4063
rect 32907 4060 32919 4063
rect 33686 4060 33692 4072
rect 32907 4032 33692 4060
rect 32907 4029 32919 4032
rect 32861 4023 32919 4029
rect 33686 4020 33692 4032
rect 33744 4020 33750 4072
rect 33870 4060 33876 4072
rect 33831 4032 33876 4060
rect 33870 4020 33876 4032
rect 33928 4020 33934 4072
rect 35618 4020 35624 4072
rect 35676 4060 35682 4072
rect 35805 4063 35863 4069
rect 35805 4060 35817 4063
rect 35676 4032 35817 4060
rect 35676 4020 35682 4032
rect 35805 4029 35817 4032
rect 35851 4029 35863 4063
rect 35805 4023 35863 4029
rect 36722 4020 36728 4072
rect 36780 4060 36786 4072
rect 36817 4063 36875 4069
rect 36817 4060 36829 4063
rect 36780 4032 36829 4060
rect 36780 4020 36786 4032
rect 36817 4029 36829 4032
rect 36863 4029 36875 4063
rect 36817 4023 36875 4029
rect 38565 4063 38623 4069
rect 38565 4029 38577 4063
rect 38611 4060 38623 4063
rect 39390 4060 39396 4072
rect 38611 4032 39396 4060
rect 38611 4029 38623 4032
rect 38565 4023 38623 4029
rect 39390 4020 39396 4032
rect 39448 4020 39454 4072
rect 39577 4063 39635 4069
rect 39577 4029 39589 4063
rect 39623 4060 39635 4063
rect 40402 4060 40408 4072
rect 39623 4032 40408 4060
rect 39623 4029 39635 4032
rect 39577 4023 39635 4029
rect 40402 4020 40408 4032
rect 40460 4020 40466 4072
rect 40586 4020 40592 4072
rect 40644 4060 40650 4072
rect 41417 4063 41475 4069
rect 41417 4060 41429 4063
rect 40644 4032 41429 4060
rect 40644 4020 40650 4032
rect 41417 4029 41429 4032
rect 41463 4029 41475 4063
rect 41417 4023 41475 4029
rect 33042 3992 33048 4004
rect 22388 3964 24440 3992
rect 30852 3964 33048 3992
rect 20809 3927 20867 3933
rect 20809 3893 20821 3927
rect 20855 3893 20867 3927
rect 20809 3887 20867 3893
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22388 3924 22416 3964
rect 24412 3933 24440 3964
rect 33042 3952 33048 3964
rect 33100 3952 33106 4004
rect 21968 3896 22416 3924
rect 24397 3927 24455 3933
rect 21968 3884 21974 3896
rect 24397 3893 24409 3927
rect 24443 3893 24455 3927
rect 24397 3887 24455 3893
rect 24486 3884 24492 3936
rect 24544 3924 24550 3936
rect 25409 3927 25467 3933
rect 25409 3924 25421 3927
rect 24544 3896 25421 3924
rect 24544 3884 24550 3896
rect 25409 3893 25421 3896
rect 25455 3893 25467 3927
rect 25409 3887 25467 3893
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 26421 3927 26479 3933
rect 26421 3924 26433 3927
rect 25556 3896 26433 3924
rect 25556 3884 25562 3896
rect 26421 3893 26433 3896
rect 26467 3893 26479 3927
rect 26421 3887 26479 3893
rect 27433 3927 27491 3933
rect 27433 3893 27445 3927
rect 27479 3924 27491 3927
rect 27706 3924 27712 3936
rect 27479 3896 27712 3924
rect 27479 3893 27491 3896
rect 27433 3887 27491 3893
rect 27706 3884 27712 3896
rect 27764 3884 27770 3936
rect 28445 3927 28503 3933
rect 28445 3893 28457 3927
rect 28491 3924 28503 3927
rect 28994 3924 29000 3936
rect 28491 3896 29000 3924
rect 28491 3893 28503 3896
rect 28445 3887 28503 3893
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 30653 3927 30711 3933
rect 30653 3893 30665 3927
rect 30699 3924 30711 3927
rect 31294 3924 31300 3936
rect 30699 3896 31300 3924
rect 30699 3893 30711 3896
rect 30653 3887 30711 3893
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 31662 3924 31668 3936
rect 31623 3896 31668 3924
rect 31662 3884 31668 3896
rect 31720 3884 31726 3936
rect 33689 3927 33747 3933
rect 33689 3893 33701 3927
rect 33735 3924 33747 3927
rect 34238 3924 34244 3936
rect 33735 3896 34244 3924
rect 33735 3893 33747 3896
rect 33689 3887 33747 3893
rect 34238 3884 34244 3896
rect 34296 3884 34302 3936
rect 35621 3927 35679 3933
rect 35621 3893 35633 3927
rect 35667 3924 35679 3927
rect 36078 3924 36084 3936
rect 35667 3896 36084 3924
rect 35667 3893 35679 3896
rect 35621 3887 35679 3893
rect 36078 3884 36084 3896
rect 36136 3884 36142 3936
rect 36630 3924 36636 3936
rect 36591 3896 36636 3924
rect 36630 3884 36636 3896
rect 36688 3884 36694 3936
rect 38378 3924 38384 3936
rect 38339 3896 38384 3924
rect 38378 3884 38384 3896
rect 38436 3884 38442 3936
rect 39393 3927 39451 3933
rect 39393 3893 39405 3927
rect 39439 3924 39451 3927
rect 40310 3924 40316 3936
rect 39439 3896 40316 3924
rect 39439 3893 39451 3896
rect 39393 3887 39451 3893
rect 40310 3884 40316 3896
rect 40368 3884 40374 3936
rect 41233 3927 41291 3933
rect 41233 3893 41245 3927
rect 41279 3924 41291 3927
rect 42426 3924 42432 3936
rect 41279 3896 42432 3924
rect 41279 3893 41291 3896
rect 41233 3887 41291 3893
rect 42426 3884 42432 3896
rect 42484 3884 42490 3936
rect 1104 3834 54832 3856
rect 1104 3782 18912 3834
rect 18964 3782 18976 3834
rect 19028 3782 19040 3834
rect 19092 3782 19104 3834
rect 19156 3782 36843 3834
rect 36895 3782 36907 3834
rect 36959 3782 36971 3834
rect 37023 3782 37035 3834
rect 37087 3782 54832 3834
rect 1104 3760 54832 3782
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 16393 3723 16451 3729
rect 16393 3689 16405 3723
rect 16439 3720 16451 3723
rect 16574 3720 16580 3732
rect 16439 3692 16580 3720
rect 16439 3689 16451 3692
rect 16393 3683 16451 3689
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 21637 3723 21695 3729
rect 21637 3689 21649 3723
rect 21683 3720 21695 3723
rect 23382 3720 23388 3732
rect 21683 3692 23388 3720
rect 21683 3689 21695 3692
rect 21637 3683 21695 3689
rect 23382 3680 23388 3692
rect 23440 3680 23446 3732
rect 24762 3720 24768 3732
rect 24723 3692 24768 3720
rect 24762 3680 24768 3692
rect 24820 3680 24826 3732
rect 28258 3720 28264 3732
rect 28219 3692 28264 3720
rect 28258 3680 28264 3692
rect 28316 3680 28322 3732
rect 33870 3680 33876 3732
rect 33928 3720 33934 3732
rect 35897 3723 35955 3729
rect 35897 3720 35909 3723
rect 33928 3692 35909 3720
rect 33928 3680 33934 3692
rect 35897 3689 35909 3692
rect 35943 3689 35955 3723
rect 35897 3683 35955 3689
rect 40678 3680 40684 3732
rect 40736 3720 40742 3732
rect 42521 3723 42579 3729
rect 42521 3720 42533 3723
rect 40736 3692 42533 3720
rect 40736 3680 40742 3692
rect 42521 3689 42533 3692
rect 42567 3689 42579 3723
rect 42521 3683 42579 3689
rect 19426 3652 19432 3664
rect 16592 3624 19432 3652
rect 14182 3584 14188 3596
rect 14143 3556 14188 3584
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 16592 3593 16620 3624
rect 19426 3612 19432 3624
rect 19484 3612 19490 3664
rect 25038 3652 25044 3664
rect 22848 3624 25044 3652
rect 16577 3587 16635 3593
rect 16577 3553 16589 3587
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 18877 3587 18935 3593
rect 18877 3553 18889 3587
rect 18923 3584 18935 3587
rect 19794 3584 19800 3596
rect 18923 3556 19800 3584
rect 18923 3553 18935 3556
rect 18877 3547 18935 3553
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 21821 3587 21879 3593
rect 21821 3553 21833 3587
rect 21867 3584 21879 3587
rect 22738 3584 22744 3596
rect 21867 3556 22744 3584
rect 21867 3553 21879 3556
rect 21821 3547 21879 3553
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 22848 3516 22876 3624
rect 25038 3612 25044 3624
rect 25096 3612 25102 3664
rect 38378 3612 38384 3664
rect 38436 3652 38442 3664
rect 38436 3624 42748 3652
rect 38436 3612 38442 3624
rect 22925 3587 22983 3593
rect 22925 3553 22937 3587
rect 22971 3584 22983 3587
rect 23937 3587 23995 3593
rect 22971 3556 23796 3584
rect 22971 3553 22983 3556
rect 22925 3547 22983 3553
rect 18616 3488 22876 3516
rect 18616 3380 18644 3488
rect 22741 3451 22799 3457
rect 22741 3417 22753 3451
rect 22787 3448 22799 3451
rect 22922 3448 22928 3460
rect 22787 3420 22928 3448
rect 22787 3417 22799 3420
rect 22741 3411 22799 3417
rect 22922 3408 22928 3420
rect 22980 3408 22986 3460
rect 23768 3457 23796 3556
rect 23937 3553 23949 3587
rect 23983 3584 23995 3587
rect 24486 3584 24492 3596
rect 23983 3556 24492 3584
rect 23983 3553 23995 3556
rect 23937 3547 23995 3553
rect 24486 3544 24492 3556
rect 24544 3544 24550 3596
rect 24949 3587 25007 3593
rect 24949 3553 24961 3587
rect 24995 3584 25007 3587
rect 25498 3584 25504 3596
rect 24995 3556 25504 3584
rect 24995 3553 25007 3556
rect 24949 3547 25007 3553
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 25961 3587 26019 3593
rect 25961 3553 25973 3587
rect 26007 3584 26019 3587
rect 26234 3584 26240 3596
rect 26007 3556 26240 3584
rect 26007 3553 26019 3556
rect 25961 3547 26019 3553
rect 26234 3544 26240 3556
rect 26292 3544 26298 3596
rect 26786 3544 26792 3596
rect 26844 3584 26850 3596
rect 27433 3587 27491 3593
rect 27433 3584 27445 3587
rect 26844 3556 27445 3584
rect 26844 3544 26850 3556
rect 27433 3553 27445 3556
rect 27479 3553 27491 3587
rect 28442 3584 28448 3596
rect 28403 3556 28448 3584
rect 27433 3547 27491 3553
rect 28442 3544 28448 3556
rect 28500 3544 28506 3596
rect 29454 3584 29460 3596
rect 29415 3556 29460 3584
rect 29454 3544 29460 3556
rect 29512 3544 29518 3596
rect 30558 3584 30564 3596
rect 30519 3556 30564 3584
rect 30558 3544 30564 3556
rect 30616 3544 30622 3596
rect 31662 3544 31668 3596
rect 31720 3584 31726 3596
rect 33045 3587 33103 3593
rect 33045 3584 33057 3587
rect 31720 3556 33057 3584
rect 31720 3544 31726 3556
rect 33045 3553 33057 3556
rect 33091 3553 33103 3587
rect 34054 3584 34060 3596
rect 34015 3556 34060 3584
rect 33045 3547 33103 3553
rect 34054 3544 34060 3556
rect 34112 3544 34118 3596
rect 35066 3584 35072 3596
rect 35027 3556 35072 3584
rect 35066 3544 35072 3556
rect 35124 3544 35130 3596
rect 36078 3584 36084 3596
rect 36039 3556 36084 3584
rect 36078 3544 36084 3556
rect 36136 3544 36142 3596
rect 36630 3544 36636 3596
rect 36688 3584 36694 3596
rect 37093 3587 37151 3593
rect 37093 3584 37105 3587
rect 36688 3556 37105 3584
rect 36688 3544 36694 3556
rect 37093 3553 37105 3556
rect 37139 3553 37151 3587
rect 38654 3584 38660 3596
rect 38615 3556 38660 3584
rect 37093 3547 37151 3553
rect 38654 3544 38660 3556
rect 38712 3544 38718 3596
rect 39669 3587 39727 3593
rect 39669 3553 39681 3587
rect 39715 3584 39727 3587
rect 40586 3584 40592 3596
rect 39715 3556 40592 3584
rect 39715 3553 39727 3556
rect 39669 3547 39727 3553
rect 40586 3544 40592 3556
rect 40644 3544 40650 3596
rect 40681 3587 40739 3593
rect 40681 3553 40693 3587
rect 40727 3584 40739 3587
rect 41230 3584 41236 3596
rect 40727 3556 41236 3584
rect 40727 3553 40739 3556
rect 40681 3547 40739 3553
rect 41230 3544 41236 3556
rect 41288 3544 41294 3596
rect 41693 3587 41751 3593
rect 41693 3553 41705 3587
rect 41739 3584 41751 3587
rect 42242 3584 42248 3596
rect 41739 3556 42248 3584
rect 41739 3553 41751 3556
rect 41693 3547 41751 3553
rect 42242 3544 42248 3556
rect 42300 3544 42306 3596
rect 42720 3593 42748 3624
rect 42705 3587 42763 3593
rect 42705 3553 42717 3587
rect 42751 3553 42763 3587
rect 42705 3547 42763 3553
rect 23753 3451 23811 3457
rect 23753 3417 23765 3451
rect 23799 3417 23811 3451
rect 23753 3411 23811 3417
rect 31846 3408 31852 3460
rect 31904 3448 31910 3460
rect 31904 3420 33364 3448
rect 31904 3408 31910 3420
rect 18693 3383 18751 3389
rect 18693 3380 18705 3383
rect 18616 3352 18705 3380
rect 18693 3349 18705 3352
rect 18739 3349 18751 3383
rect 18693 3343 18751 3349
rect 24946 3340 24952 3392
rect 25004 3380 25010 3392
rect 25777 3383 25835 3389
rect 25777 3380 25789 3383
rect 25004 3352 25789 3380
rect 25004 3340 25010 3352
rect 25777 3349 25789 3352
rect 25823 3349 25835 3383
rect 25777 3343 25835 3349
rect 25958 3340 25964 3392
rect 26016 3380 26022 3392
rect 27249 3383 27307 3389
rect 27249 3380 27261 3383
rect 26016 3352 27261 3380
rect 26016 3340 26022 3352
rect 27249 3349 27261 3352
rect 27295 3349 27307 3383
rect 29270 3380 29276 3392
rect 29231 3352 29276 3380
rect 27249 3343 27307 3349
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 30377 3383 30435 3389
rect 30377 3349 30389 3383
rect 30423 3380 30435 3383
rect 31202 3380 31208 3392
rect 30423 3352 31208 3380
rect 30423 3349 30435 3352
rect 30377 3343 30435 3349
rect 31202 3340 31208 3352
rect 31260 3340 31266 3392
rect 32861 3383 32919 3389
rect 32861 3349 32873 3383
rect 32907 3380 32919 3383
rect 33226 3380 33232 3392
rect 32907 3352 33232 3380
rect 32907 3349 32919 3352
rect 32861 3343 32919 3349
rect 33226 3340 33232 3352
rect 33284 3340 33290 3392
rect 33336 3380 33364 3420
rect 33686 3408 33692 3460
rect 33744 3448 33750 3460
rect 34885 3451 34943 3457
rect 34885 3448 34897 3451
rect 33744 3420 34897 3448
rect 33744 3408 33750 3420
rect 34885 3417 34897 3420
rect 34931 3417 34943 3451
rect 34885 3411 34943 3417
rect 41509 3451 41567 3457
rect 41509 3417 41521 3451
rect 41555 3448 41567 3451
rect 43070 3448 43076 3460
rect 41555 3420 43076 3448
rect 41555 3417 41567 3420
rect 41509 3411 41567 3417
rect 43070 3408 43076 3420
rect 43128 3408 43134 3460
rect 33873 3383 33931 3389
rect 33873 3380 33885 3383
rect 33336 3352 33885 3380
rect 33873 3349 33885 3352
rect 33919 3349 33931 3383
rect 33873 3343 33931 3349
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 36909 3383 36967 3389
rect 36909 3380 36921 3383
rect 36044 3352 36921 3380
rect 36044 3340 36050 3352
rect 36909 3349 36921 3352
rect 36955 3349 36967 3383
rect 36909 3343 36967 3349
rect 38473 3383 38531 3389
rect 38473 3349 38485 3383
rect 38519 3380 38531 3383
rect 39206 3380 39212 3392
rect 38519 3352 39212 3380
rect 38519 3349 38531 3352
rect 38473 3343 38531 3349
rect 39206 3340 39212 3352
rect 39264 3340 39270 3392
rect 39485 3383 39543 3389
rect 39485 3349 39497 3383
rect 39531 3380 39543 3383
rect 40218 3380 40224 3392
rect 39531 3352 40224 3380
rect 39531 3349 39543 3352
rect 39485 3343 39543 3349
rect 40218 3340 40224 3352
rect 40276 3340 40282 3392
rect 40497 3383 40555 3389
rect 40497 3349 40509 3383
rect 40543 3380 40555 3383
rect 41414 3380 41420 3392
rect 40543 3352 41420 3380
rect 40543 3349 40555 3352
rect 40497 3343 40555 3349
rect 41414 3340 41420 3352
rect 41472 3340 41478 3392
rect 1104 3290 54832 3312
rect 1104 3238 9947 3290
rect 9999 3238 10011 3290
rect 10063 3238 10075 3290
rect 10127 3238 10139 3290
rect 10191 3238 27878 3290
rect 27930 3238 27942 3290
rect 27994 3238 28006 3290
rect 28058 3238 28070 3290
rect 28122 3238 45808 3290
rect 45860 3238 45872 3290
rect 45924 3238 45936 3290
rect 45988 3238 46000 3290
rect 46052 3238 54832 3290
rect 1104 3216 54832 3238
rect 21729 3179 21787 3185
rect 21729 3145 21741 3179
rect 21775 3176 21787 3179
rect 25777 3179 25835 3185
rect 21775 3148 24716 3176
rect 21775 3145 21787 3148
rect 21729 3139 21787 3145
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3108 20775 3111
rect 22830 3108 22836 3120
rect 20763 3080 22836 3108
rect 20763 3077 20775 3080
rect 20717 3071 20775 3077
rect 22830 3068 22836 3080
rect 22888 3068 22894 3120
rect 24688 3040 24716 3148
rect 25777 3145 25789 3179
rect 25823 3176 25835 3179
rect 26326 3176 26332 3188
rect 25823 3148 26332 3176
rect 25823 3145 25835 3148
rect 25777 3139 25835 3145
rect 26326 3136 26332 3148
rect 26384 3136 26390 3188
rect 26786 3176 26792 3188
rect 26747 3148 26792 3176
rect 26786 3136 26792 3148
rect 26844 3136 26850 3188
rect 30558 3136 30564 3188
rect 30616 3176 30622 3188
rect 32033 3179 32091 3185
rect 32033 3176 32045 3179
rect 30616 3148 32045 3176
rect 30616 3136 30622 3148
rect 32033 3145 32045 3148
rect 32079 3145 32091 3179
rect 33042 3176 33048 3188
rect 33003 3148 33048 3176
rect 32033 3139 32091 3145
rect 33042 3136 33048 3148
rect 33100 3136 33106 3188
rect 34057 3179 34115 3185
rect 34057 3145 34069 3179
rect 34103 3176 34115 3179
rect 35066 3176 35072 3188
rect 34103 3148 35072 3176
rect 34103 3145 34115 3148
rect 34057 3139 34115 3145
rect 35066 3136 35072 3148
rect 35124 3136 35130 3188
rect 35618 3176 35624 3188
rect 35579 3148 35624 3176
rect 35618 3136 35624 3148
rect 35676 3136 35682 3188
rect 36633 3179 36691 3185
rect 36633 3145 36645 3179
rect 36679 3176 36691 3179
rect 36722 3176 36728 3188
rect 36679 3148 36728 3176
rect 36679 3145 36691 3148
rect 36633 3139 36691 3145
rect 36722 3136 36728 3148
rect 36780 3136 36786 3188
rect 38654 3136 38660 3188
rect 38712 3176 38718 3188
rect 39669 3179 39727 3185
rect 39669 3176 39681 3179
rect 38712 3148 39681 3176
rect 38712 3136 38718 3148
rect 39669 3145 39681 3148
rect 39715 3145 39727 3179
rect 41230 3176 41236 3188
rect 41191 3148 41236 3176
rect 39669 3139 39727 3145
rect 41230 3136 41236 3148
rect 41288 3136 41294 3188
rect 42242 3176 42248 3188
rect 42203 3148 42248 3176
rect 42242 3136 42248 3148
rect 42300 3136 42306 3188
rect 24765 3111 24823 3117
rect 24765 3077 24777 3111
rect 24811 3108 24823 3111
rect 29086 3108 29092 3120
rect 24811 3080 29092 3108
rect 24811 3077 24823 3080
rect 24765 3071 24823 3077
rect 29086 3068 29092 3080
rect 29144 3068 29150 3120
rect 26418 3040 26424 3052
rect 24688 3012 26424 3040
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 28350 3040 28356 3052
rect 26988 3012 28356 3040
rect 20898 2972 20904 2984
rect 20859 2944 20904 2972
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 21910 2972 21916 2984
rect 21871 2944 21916 2972
rect 21910 2932 21916 2944
rect 21968 2932 21974 2984
rect 22922 2972 22928 2984
rect 22883 2944 22928 2972
rect 22922 2932 22928 2944
rect 22980 2932 22986 2984
rect 24946 2972 24952 2984
rect 24907 2944 24952 2972
rect 24946 2932 24952 2944
rect 25004 2932 25010 2984
rect 25958 2972 25964 2984
rect 25919 2944 25964 2972
rect 25958 2932 25964 2944
rect 26016 2932 26022 2984
rect 26988 2981 27016 3012
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 26973 2975 27031 2981
rect 26973 2941 26985 2975
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 27985 2975 28043 2981
rect 27985 2941 27997 2975
rect 28031 2972 28043 2975
rect 29270 2972 29276 2984
rect 28031 2944 29276 2972
rect 28031 2941 28043 2944
rect 27985 2935 28043 2941
rect 29270 2932 29276 2944
rect 29328 2932 29334 2984
rect 30193 2975 30251 2981
rect 30193 2941 30205 2975
rect 30239 2972 30251 2975
rect 31018 2972 31024 2984
rect 30239 2944 31024 2972
rect 30239 2941 30251 2944
rect 30193 2935 30251 2941
rect 31018 2932 31024 2944
rect 31076 2932 31082 2984
rect 31202 2972 31208 2984
rect 31163 2944 31208 2972
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 31294 2932 31300 2984
rect 31352 2972 31358 2984
rect 32217 2975 32275 2981
rect 32217 2972 32229 2975
rect 31352 2944 32229 2972
rect 31352 2932 31358 2944
rect 32217 2941 32229 2944
rect 32263 2941 32275 2975
rect 33226 2972 33232 2984
rect 33187 2944 33232 2972
rect 32217 2935 32275 2941
rect 33226 2932 33232 2944
rect 33284 2932 33290 2984
rect 34238 2972 34244 2984
rect 34199 2944 34244 2972
rect 34238 2932 34244 2944
rect 34296 2932 34302 2984
rect 35805 2975 35863 2981
rect 35805 2941 35817 2975
rect 35851 2972 35863 2975
rect 35986 2972 35992 2984
rect 35851 2944 35992 2972
rect 35851 2941 35863 2944
rect 35805 2935 35863 2941
rect 35986 2932 35992 2944
rect 36044 2932 36050 2984
rect 36538 2932 36544 2984
rect 36596 2972 36602 2984
rect 36817 2975 36875 2981
rect 36817 2972 36829 2975
rect 36596 2944 36829 2972
rect 36596 2932 36602 2944
rect 36817 2941 36829 2944
rect 36863 2941 36875 2975
rect 37826 2972 37832 2984
rect 37787 2944 37832 2972
rect 36817 2935 36875 2941
rect 37826 2932 37832 2944
rect 37884 2932 37890 2984
rect 38838 2972 38844 2984
rect 38799 2944 38844 2972
rect 38838 2932 38844 2944
rect 38896 2932 38902 2984
rect 39853 2975 39911 2981
rect 39853 2941 39865 2975
rect 39899 2972 39911 2975
rect 40034 2972 40040 2984
rect 39899 2944 40040 2972
rect 39899 2941 39911 2944
rect 39853 2935 39911 2941
rect 40034 2932 40040 2944
rect 40092 2932 40098 2984
rect 40310 2932 40316 2984
rect 40368 2972 40374 2984
rect 41417 2975 41475 2981
rect 41417 2972 41429 2975
rect 40368 2944 41429 2972
rect 40368 2932 40374 2944
rect 41417 2941 41429 2944
rect 41463 2941 41475 2975
rect 42426 2972 42432 2984
rect 42387 2944 42432 2972
rect 41417 2935 41475 2941
rect 42426 2932 42432 2944
rect 42484 2932 42490 2984
rect 22741 2839 22799 2845
rect 22741 2805 22753 2839
rect 22787 2836 22799 2839
rect 23842 2836 23848 2848
rect 22787 2808 23848 2836
rect 22787 2805 22799 2808
rect 22741 2799 22799 2805
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 27798 2836 27804 2848
rect 27759 2808 27804 2836
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 30009 2839 30067 2845
rect 30009 2805 30021 2839
rect 30055 2836 30067 2839
rect 30650 2836 30656 2848
rect 30055 2808 30656 2836
rect 30055 2805 30067 2808
rect 30009 2799 30067 2805
rect 30650 2796 30656 2808
rect 30708 2796 30714 2848
rect 31021 2839 31079 2845
rect 31021 2805 31033 2839
rect 31067 2836 31079 2839
rect 31662 2836 31668 2848
rect 31067 2808 31668 2836
rect 31067 2805 31079 2808
rect 31021 2799 31079 2805
rect 31662 2796 31668 2808
rect 31720 2796 31726 2848
rect 37274 2796 37280 2848
rect 37332 2836 37338 2848
rect 37645 2839 37703 2845
rect 37645 2836 37657 2839
rect 37332 2808 37657 2836
rect 37332 2796 37338 2808
rect 37645 2805 37657 2808
rect 37691 2805 37703 2839
rect 38654 2836 38660 2848
rect 38615 2808 38660 2836
rect 37645 2799 37703 2805
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 1104 2746 54832 2768
rect 1104 2694 18912 2746
rect 18964 2694 18976 2746
rect 19028 2694 19040 2746
rect 19092 2694 19104 2746
rect 19156 2694 36843 2746
rect 36895 2694 36907 2746
rect 36959 2694 36971 2746
rect 37023 2694 37035 2746
rect 37087 2694 54832 2746
rect 1104 2672 54832 2694
rect 20809 2635 20867 2641
rect 20809 2601 20821 2635
rect 20855 2632 20867 2635
rect 20898 2632 20904 2644
rect 20855 2604 20904 2632
rect 20855 2601 20867 2604
rect 20809 2595 20867 2601
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 22649 2635 22707 2641
rect 22649 2601 22661 2635
rect 22695 2632 22707 2635
rect 22922 2632 22928 2644
rect 22695 2604 22928 2632
rect 22695 2601 22707 2604
rect 22649 2595 22707 2601
rect 22922 2592 22928 2604
rect 22980 2592 22986 2644
rect 27617 2635 27675 2641
rect 27617 2601 27629 2635
rect 27663 2632 27675 2635
rect 28442 2632 28448 2644
rect 27663 2604 28448 2632
rect 27663 2601 27675 2604
rect 27617 2595 27675 2601
rect 28442 2592 28448 2604
rect 28500 2592 28506 2644
rect 28629 2635 28687 2641
rect 28629 2601 28641 2635
rect 28675 2632 28687 2635
rect 30190 2632 30196 2644
rect 28675 2604 30196 2632
rect 28675 2601 28687 2604
rect 28629 2595 28687 2601
rect 30190 2592 30196 2604
rect 30248 2592 30254 2644
rect 30469 2635 30527 2641
rect 30469 2601 30481 2635
rect 30515 2601 30527 2635
rect 30469 2595 30527 2601
rect 23474 2564 23480 2576
rect 21008 2536 23480 2564
rect 21008 2505 21036 2536
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 30374 2564 30380 2576
rect 23584 2536 30380 2564
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2465 21051 2499
rect 22830 2496 22836 2508
rect 22791 2468 22836 2496
rect 20993 2459 21051 2465
rect 19794 2292 19800 2304
rect 19755 2264 19800 2292
rect 19794 2252 19800 2264
rect 19852 2252 19858 2304
rect 19996 2292 20024 2459
rect 22830 2456 22836 2468
rect 22888 2456 22894 2508
rect 23584 2496 23612 2536
rect 30374 2524 30380 2536
rect 30432 2524 30438 2576
rect 23842 2496 23848 2508
rect 23400 2468 23612 2496
rect 23803 2468 23848 2496
rect 23400 2292 23428 2468
rect 23842 2456 23848 2468
rect 23900 2456 23906 2508
rect 24949 2499 25007 2505
rect 24949 2496 24961 2499
rect 24688 2468 24961 2496
rect 23661 2363 23719 2369
rect 23661 2329 23673 2363
rect 23707 2360 23719 2363
rect 24688 2360 24716 2468
rect 24949 2465 24961 2468
rect 24995 2465 25007 2499
rect 24949 2459 25007 2465
rect 25961 2499 26019 2505
rect 25961 2465 25973 2499
rect 26007 2465 26019 2499
rect 27798 2496 27804 2508
rect 27759 2468 27804 2496
rect 25961 2459 26019 2465
rect 25976 2428 26004 2459
rect 27798 2456 27804 2468
rect 27856 2456 27862 2508
rect 28813 2499 28871 2505
rect 28813 2465 28825 2499
rect 28859 2496 28871 2499
rect 30484 2496 30512 2595
rect 31018 2592 31024 2644
rect 31076 2632 31082 2644
rect 31481 2635 31539 2641
rect 31481 2632 31493 2635
rect 31076 2604 31493 2632
rect 31076 2592 31082 2604
rect 31481 2601 31493 2604
rect 31527 2601 31539 2635
rect 34330 2632 34336 2644
rect 34291 2604 34336 2632
rect 31481 2595 31539 2601
rect 34330 2592 34336 2604
rect 34388 2592 34394 2644
rect 36170 2632 36176 2644
rect 36131 2604 36176 2632
rect 36170 2592 36176 2604
rect 36228 2592 36234 2644
rect 37185 2635 37243 2641
rect 37185 2601 37197 2635
rect 37231 2632 37243 2635
rect 37826 2632 37832 2644
rect 37231 2604 37832 2632
rect 37231 2601 37243 2604
rect 37185 2595 37243 2601
rect 37826 2592 37832 2604
rect 37884 2592 37890 2644
rect 38838 2592 38844 2644
rect 38896 2632 38902 2644
rect 39025 2635 39083 2641
rect 39025 2632 39037 2635
rect 38896 2604 39037 2632
rect 38896 2592 38902 2604
rect 39025 2601 39037 2604
rect 39071 2601 39083 2635
rect 40034 2632 40040 2644
rect 39995 2604 40040 2632
rect 39025 2595 39083 2601
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 40586 2592 40592 2644
rect 40644 2632 40650 2644
rect 41877 2635 41935 2641
rect 41877 2632 41889 2635
rect 40644 2604 41889 2632
rect 40644 2592 40650 2604
rect 41877 2601 41889 2604
rect 41923 2601 41935 2635
rect 41877 2595 41935 2601
rect 30650 2496 30656 2508
rect 28859 2468 30512 2496
rect 30611 2468 30656 2496
rect 28859 2465 28871 2468
rect 28813 2459 28871 2465
rect 30650 2456 30656 2468
rect 30708 2456 30714 2508
rect 31662 2496 31668 2508
rect 31623 2468 31668 2496
rect 31662 2456 31668 2468
rect 31720 2456 31726 2508
rect 33502 2496 33508 2508
rect 33463 2468 33508 2496
rect 33502 2456 33508 2468
rect 33560 2456 33566 2508
rect 34514 2496 34520 2508
rect 34475 2468 34520 2496
rect 34514 2456 34520 2468
rect 34572 2456 34578 2508
rect 36357 2499 36415 2505
rect 36357 2465 36369 2499
rect 36403 2496 36415 2499
rect 37274 2496 37280 2508
rect 36403 2468 37280 2496
rect 36403 2465 36415 2468
rect 36357 2459 36415 2465
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 37369 2499 37427 2505
rect 37369 2465 37381 2499
rect 37415 2496 37427 2499
rect 38654 2496 38660 2508
rect 37415 2468 38660 2496
rect 37415 2465 37427 2468
rect 37369 2459 37427 2465
rect 38654 2456 38660 2468
rect 38712 2456 38718 2508
rect 39206 2496 39212 2508
rect 39167 2468 39212 2496
rect 39206 2456 39212 2468
rect 39264 2456 39270 2508
rect 40218 2496 40224 2508
rect 40179 2468 40224 2496
rect 40218 2456 40224 2468
rect 40276 2456 40282 2508
rect 41414 2456 41420 2508
rect 41472 2496 41478 2508
rect 42061 2499 42119 2505
rect 42061 2496 42073 2499
rect 41472 2468 42073 2496
rect 41472 2456 41478 2468
rect 42061 2465 42073 2468
rect 42107 2465 42119 2499
rect 43070 2496 43076 2508
rect 43031 2468 43076 2496
rect 42061 2459 42119 2465
rect 43070 2456 43076 2468
rect 43128 2456 43134 2508
rect 24780 2400 26004 2428
rect 24780 2369 24808 2400
rect 23707 2332 24716 2360
rect 24765 2363 24823 2369
rect 23707 2329 23719 2332
rect 23661 2323 23719 2329
rect 24765 2329 24777 2363
rect 24811 2329 24823 2363
rect 24765 2323 24823 2329
rect 25777 2363 25835 2369
rect 25777 2329 25789 2363
rect 25823 2360 25835 2363
rect 30466 2360 30472 2372
rect 25823 2332 30472 2360
rect 25823 2329 25835 2332
rect 25777 2323 25835 2329
rect 30466 2320 30472 2332
rect 30524 2320 30530 2372
rect 40402 2320 40408 2372
rect 40460 2360 40466 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 40460 2332 42901 2360
rect 40460 2320 40466 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 42889 2323 42947 2329
rect 19996 2264 23428 2292
rect 23474 2252 23480 2304
rect 23532 2292 23538 2304
rect 33321 2295 33379 2301
rect 33321 2292 33333 2295
rect 23532 2264 33333 2292
rect 23532 2252 23538 2264
rect 33321 2261 33333 2264
rect 33367 2261 33379 2295
rect 33321 2255 33379 2261
rect 1104 2202 54832 2224
rect 1104 2150 9947 2202
rect 9999 2150 10011 2202
rect 10063 2150 10075 2202
rect 10127 2150 10139 2202
rect 10191 2150 27878 2202
rect 27930 2150 27942 2202
rect 27994 2150 28006 2202
rect 28058 2150 28070 2202
rect 28122 2150 45808 2202
rect 45860 2150 45872 2202
rect 45924 2150 45936 2202
rect 45988 2150 46000 2202
rect 46052 2150 54832 2202
rect 1104 2128 54832 2150
rect 19794 2048 19800 2100
rect 19852 2088 19858 2100
rect 29178 2088 29184 2100
rect 19852 2060 29184 2088
rect 19852 2048 19858 2060
rect 29178 2048 29184 2060
rect 29236 2048 29242 2100
<< via1 >>
rect 9947 24998 9999 25050
rect 10011 24998 10063 25050
rect 10075 24998 10127 25050
rect 10139 24998 10191 25050
rect 27878 24998 27930 25050
rect 27942 24998 27994 25050
rect 28006 24998 28058 25050
rect 28070 24998 28122 25050
rect 45808 24998 45860 25050
rect 45872 24998 45924 25050
rect 45936 24998 45988 25050
rect 46000 24998 46052 25050
rect 8852 24760 8904 24812
rect 21824 24760 21876 24812
rect 34980 24760 35032 24812
rect 7196 24735 7248 24744
rect 6552 24556 6604 24608
rect 7196 24701 7205 24735
rect 7205 24701 7239 24735
rect 7239 24701 7248 24735
rect 7196 24692 7248 24701
rect 8668 24599 8720 24608
rect 8668 24565 8677 24599
rect 8677 24565 8711 24599
rect 8711 24565 8720 24599
rect 8668 24556 8720 24565
rect 22468 24692 22520 24744
rect 40500 24760 40552 24812
rect 43352 24760 43404 24812
rect 47492 24760 47544 24812
rect 48504 24760 48556 24812
rect 40408 24692 40460 24744
rect 41236 24735 41288 24744
rect 41236 24701 41245 24735
rect 41245 24701 41279 24735
rect 41279 24701 41288 24735
rect 41236 24692 41288 24701
rect 41972 24692 42024 24744
rect 21548 24556 21600 24608
rect 24400 24556 24452 24608
rect 39948 24599 40000 24608
rect 39948 24565 39957 24599
rect 39957 24565 39991 24599
rect 39991 24565 40000 24599
rect 39948 24556 40000 24565
rect 42892 24556 42944 24608
rect 42984 24599 43036 24608
rect 42984 24565 42993 24599
rect 42993 24565 43027 24599
rect 43027 24565 43036 24599
rect 44272 24735 44324 24744
rect 44272 24701 44281 24735
rect 44281 24701 44315 24735
rect 44315 24701 44324 24735
rect 44272 24692 44324 24701
rect 42984 24556 43036 24565
rect 44548 24556 44600 24608
rect 45560 24599 45612 24608
rect 45560 24565 45569 24599
rect 45569 24565 45603 24599
rect 45603 24565 45612 24599
rect 45560 24556 45612 24565
rect 48596 24556 48648 24608
rect 50620 24692 50672 24744
rect 51080 24599 51132 24608
rect 51080 24565 51089 24599
rect 51089 24565 51123 24599
rect 51123 24565 51132 24599
rect 51080 24556 51132 24565
rect 18912 24454 18964 24506
rect 18976 24454 19028 24506
rect 19040 24454 19092 24506
rect 19104 24454 19156 24506
rect 36843 24454 36895 24506
rect 36907 24454 36959 24506
rect 36971 24454 37023 24506
rect 37035 24454 37087 24506
rect 1676 24352 1728 24404
rect 7472 24352 7524 24404
rect 13176 24352 13228 24404
rect 16028 24352 16080 24404
rect 17500 24352 17552 24404
rect 20352 24352 20404 24404
rect 23480 24352 23532 24404
rect 27620 24352 27672 24404
rect 30380 24395 30432 24404
rect 30380 24361 30389 24395
rect 30389 24361 30423 24395
rect 30423 24361 30432 24395
rect 30380 24352 30432 24361
rect 33324 24352 33376 24404
rect 34704 24352 34756 24404
rect 39028 24352 39080 24404
rect 50528 24352 50580 24404
rect 6000 24284 6052 24336
rect 11704 24284 11756 24336
rect 42892 24284 42944 24336
rect 50620 24327 50672 24336
rect 4252 24148 4304 24200
rect 5908 24259 5960 24268
rect 5908 24225 5917 24259
rect 5917 24225 5951 24259
rect 5951 24225 5960 24259
rect 6552 24259 6604 24268
rect 5908 24216 5960 24225
rect 6552 24225 6561 24259
rect 6561 24225 6595 24259
rect 6595 24225 6604 24259
rect 6552 24216 6604 24225
rect 8668 24216 8720 24268
rect 9772 24216 9824 24268
rect 13636 24216 13688 24268
rect 15384 24216 15436 24268
rect 19432 24216 19484 24268
rect 21548 24216 21600 24268
rect 25228 24216 25280 24268
rect 31484 24216 31536 24268
rect 35900 24216 35952 24268
rect 41236 24216 41288 24268
rect 42984 24216 43036 24268
rect 50620 24293 50629 24327
rect 50629 24293 50663 24327
rect 50663 24293 50672 24327
rect 50620 24284 50672 24293
rect 6828 24191 6880 24200
rect 4068 24012 4120 24064
rect 5816 24012 5868 24064
rect 6828 24157 6837 24191
rect 6837 24157 6871 24191
rect 6871 24157 6880 24191
rect 6828 24148 6880 24157
rect 10416 24148 10468 24200
rect 12624 24148 12676 24200
rect 17776 24191 17828 24200
rect 17776 24157 17785 24191
rect 17785 24157 17819 24191
rect 17819 24157 17828 24191
rect 17776 24148 17828 24157
rect 20812 24148 20864 24200
rect 21180 24191 21232 24200
rect 21180 24157 21189 24191
rect 21189 24157 21223 24191
rect 21223 24157 21232 24191
rect 21180 24148 21232 24157
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 9680 24080 9732 24132
rect 32220 24148 32272 24200
rect 32312 24191 32364 24200
rect 32312 24157 32321 24191
rect 32321 24157 32355 24191
rect 32355 24157 32364 24191
rect 32312 24148 32364 24157
rect 33692 24148 33744 24200
rect 35072 24191 35124 24200
rect 35072 24157 35081 24191
rect 35081 24157 35115 24191
rect 35115 24157 35124 24191
rect 35072 24148 35124 24157
rect 38752 24191 38804 24200
rect 38752 24157 38761 24191
rect 38761 24157 38795 24191
rect 38795 24157 38804 24191
rect 38752 24148 38804 24157
rect 29368 24012 29420 24064
rect 30748 24055 30800 24064
rect 30748 24021 30757 24055
rect 30757 24021 30791 24055
rect 30791 24021 30800 24055
rect 30748 24012 30800 24021
rect 44548 24012 44600 24064
rect 45376 24012 45428 24064
rect 46572 24148 46624 24200
rect 54852 24216 54904 24268
rect 46664 24012 46716 24064
rect 9947 23910 9999 23962
rect 10011 23910 10063 23962
rect 10075 23910 10127 23962
rect 10139 23910 10191 23962
rect 27878 23910 27930 23962
rect 27942 23910 27994 23962
rect 28006 23910 28058 23962
rect 28070 23910 28122 23962
rect 45808 23910 45860 23962
rect 45872 23910 45924 23962
rect 45936 23910 45988 23962
rect 46000 23910 46052 23962
rect 10324 23808 10376 23860
rect 14648 23808 14700 23860
rect 15108 23808 15160 23860
rect 15384 23851 15436 23860
rect 15384 23817 15393 23851
rect 15393 23817 15427 23851
rect 15427 23817 15436 23851
rect 15384 23808 15436 23817
rect 19340 23808 19392 23860
rect 22468 23851 22520 23860
rect 22468 23817 22477 23851
rect 22477 23817 22511 23851
rect 22511 23817 22520 23851
rect 22468 23808 22520 23817
rect 25228 23851 25280 23860
rect 25228 23817 25237 23851
rect 25237 23817 25271 23851
rect 25271 23817 25280 23851
rect 25228 23808 25280 23817
rect 26148 23808 26200 23860
rect 31852 23808 31904 23860
rect 32220 23808 32272 23860
rect 35900 23851 35952 23860
rect 35900 23817 35909 23851
rect 35909 23817 35943 23851
rect 35943 23817 35952 23851
rect 35900 23808 35952 23817
rect 36268 23808 36320 23860
rect 38752 23808 38804 23860
rect 41972 23851 42024 23860
rect 41972 23817 41981 23851
rect 41981 23817 42015 23851
rect 42015 23817 42024 23851
rect 41972 23808 42024 23817
rect 44272 23851 44324 23860
rect 44272 23817 44281 23851
rect 44281 23817 44315 23851
rect 44315 23817 44324 23851
rect 44272 23808 44324 23817
rect 46572 23851 46624 23860
rect 46572 23817 46581 23851
rect 46581 23817 46615 23851
rect 46615 23817 46624 23851
rect 46572 23808 46624 23817
rect 49056 23808 49108 23860
rect 7196 23672 7248 23724
rect 9772 23672 9824 23724
rect 13636 23715 13688 23724
rect 13636 23681 13645 23715
rect 13645 23681 13679 23715
rect 13679 23681 13688 23715
rect 13636 23672 13688 23681
rect 21364 23740 21416 23792
rect 7104 23604 7156 23656
rect 7656 23604 7708 23656
rect 8760 23647 8812 23656
rect 8760 23613 8769 23647
rect 8769 23613 8803 23647
rect 8803 23613 8812 23647
rect 8760 23604 8812 23613
rect 7196 23536 7248 23588
rect 6828 23468 6880 23520
rect 12716 23511 12768 23520
rect 12716 23477 12725 23511
rect 12725 23477 12759 23511
rect 12759 23477 12768 23511
rect 12716 23468 12768 23477
rect 13268 23468 13320 23520
rect 24400 23672 24452 23724
rect 29368 23672 29420 23724
rect 30748 23672 30800 23724
rect 34244 23672 34296 23724
rect 45376 23740 45428 23792
rect 39948 23672 40000 23724
rect 17776 23604 17828 23656
rect 18604 23604 18656 23656
rect 21548 23536 21600 23588
rect 19524 23468 19576 23520
rect 21732 23468 21784 23520
rect 22192 23579 22244 23588
rect 22192 23545 22201 23579
rect 22201 23545 22235 23579
rect 22235 23545 22244 23579
rect 22192 23536 22244 23545
rect 22100 23468 22152 23520
rect 29552 23604 29604 23656
rect 48596 23672 48648 23724
rect 32312 23647 32364 23656
rect 32312 23613 32321 23647
rect 32321 23613 32355 23647
rect 32355 23613 32364 23647
rect 32312 23604 32364 23613
rect 33324 23647 33376 23656
rect 33324 23613 33333 23647
rect 33333 23613 33367 23647
rect 33367 23613 33376 23647
rect 33324 23604 33376 23613
rect 33784 23604 33836 23656
rect 34980 23647 35032 23656
rect 34980 23613 34989 23647
rect 34989 23613 35023 23647
rect 35023 23613 35032 23647
rect 34980 23604 35032 23613
rect 36360 23647 36412 23656
rect 36360 23613 36369 23647
rect 36369 23613 36403 23647
rect 36403 23613 36412 23647
rect 36360 23604 36412 23613
rect 40040 23604 40092 23656
rect 40132 23604 40184 23656
rect 41788 23647 41840 23656
rect 41788 23613 41797 23647
rect 41797 23613 41831 23647
rect 41831 23613 41840 23647
rect 41788 23604 41840 23613
rect 44180 23604 44232 23656
rect 46204 23647 46256 23656
rect 46204 23613 46213 23647
rect 46213 23613 46247 23647
rect 46247 23613 46256 23647
rect 46204 23604 46256 23613
rect 46388 23647 46440 23656
rect 46388 23613 46397 23647
rect 46397 23613 46431 23647
rect 46431 23613 46440 23647
rect 46388 23604 46440 23613
rect 33416 23579 33468 23588
rect 33416 23545 33425 23579
rect 33425 23545 33459 23579
rect 33459 23545 33468 23579
rect 33416 23536 33468 23545
rect 28632 23468 28684 23520
rect 31576 23468 31628 23520
rect 37372 23536 37424 23588
rect 34520 23468 34572 23520
rect 35164 23511 35216 23520
rect 35164 23477 35173 23511
rect 35173 23477 35207 23511
rect 35207 23477 35216 23511
rect 35164 23468 35216 23477
rect 38844 23468 38896 23520
rect 41052 23468 41104 23520
rect 51816 23468 51868 23520
rect 52368 23647 52420 23656
rect 52368 23613 52377 23647
rect 52377 23613 52411 23647
rect 52411 23613 52420 23647
rect 52368 23604 52420 23613
rect 53472 23511 53524 23520
rect 53472 23477 53481 23511
rect 53481 23477 53515 23511
rect 53515 23477 53524 23511
rect 53472 23468 53524 23477
rect 18912 23366 18964 23418
rect 18976 23366 19028 23418
rect 19040 23366 19092 23418
rect 19104 23366 19156 23418
rect 36843 23366 36895 23418
rect 36907 23366 36959 23418
rect 36971 23366 37023 23418
rect 37035 23366 37087 23418
rect 3884 23264 3936 23316
rect 7012 23264 7064 23316
rect 13268 23307 13320 23316
rect 13268 23273 13277 23307
rect 13277 23273 13311 23307
rect 13311 23273 13320 23307
rect 13268 23264 13320 23273
rect 5908 23239 5960 23248
rect 5908 23205 5917 23239
rect 5917 23205 5951 23239
rect 5951 23205 5960 23239
rect 5908 23196 5960 23205
rect 8760 23239 8812 23248
rect 8760 23205 8769 23239
rect 8769 23205 8803 23239
rect 8803 23205 8812 23239
rect 8760 23196 8812 23205
rect 12624 23196 12676 23248
rect 940 23128 992 23180
rect 6920 23128 6972 23180
rect 7104 23128 7156 23180
rect 8024 23171 8076 23180
rect 8024 23137 8033 23171
rect 8033 23137 8067 23171
rect 8067 23137 8076 23171
rect 8024 23128 8076 23137
rect 11060 23171 11112 23180
rect 11060 23137 11069 23171
rect 11069 23137 11103 23171
rect 11103 23137 11112 23171
rect 11060 23128 11112 23137
rect 11428 23171 11480 23180
rect 11428 23137 11437 23171
rect 11437 23137 11471 23171
rect 11471 23137 11480 23171
rect 11428 23128 11480 23137
rect 4068 23103 4120 23112
rect 4068 23069 4077 23103
rect 4077 23069 4111 23103
rect 4111 23069 4120 23103
rect 4068 23060 4120 23069
rect 4344 23103 4396 23112
rect 4344 23069 4353 23103
rect 4353 23069 4387 23103
rect 4387 23069 4396 23103
rect 4344 23060 4396 23069
rect 4528 23060 4580 23112
rect 8760 23060 8812 23112
rect 11520 22992 11572 23044
rect 19524 23264 19576 23316
rect 19708 23264 19760 23316
rect 21088 23264 21140 23316
rect 21640 23264 21692 23316
rect 32496 23264 32548 23316
rect 32588 23264 32640 23316
rect 33232 23264 33284 23316
rect 19432 23196 19484 23248
rect 2412 22924 2464 22976
rect 5724 22924 5776 22976
rect 14832 22924 14884 22976
rect 15844 23171 15896 23180
rect 15844 23137 15853 23171
rect 15853 23137 15887 23171
rect 15887 23137 15896 23171
rect 15844 23128 15896 23137
rect 18512 23171 18564 23180
rect 18512 23137 18521 23171
rect 18521 23137 18555 23171
rect 18555 23137 18564 23171
rect 18512 23128 18564 23137
rect 16120 23103 16172 23112
rect 16120 23069 16129 23103
rect 16129 23069 16163 23103
rect 16163 23069 16172 23103
rect 16120 23060 16172 23069
rect 21088 23128 21140 23180
rect 19340 23060 19392 23112
rect 20904 23060 20956 23112
rect 21272 23171 21324 23180
rect 21272 23137 21281 23171
rect 21281 23137 21315 23171
rect 21315 23137 21324 23171
rect 21272 23128 21324 23137
rect 23480 23196 23532 23248
rect 23664 23196 23716 23248
rect 23940 23196 23992 23248
rect 25320 23196 25372 23248
rect 23296 23171 23348 23180
rect 23296 23137 23305 23171
rect 23305 23137 23339 23171
rect 23339 23137 23348 23171
rect 23296 23128 23348 23137
rect 15384 23035 15436 23044
rect 15384 23001 15393 23035
rect 15393 23001 15427 23035
rect 15427 23001 15436 23035
rect 15384 22992 15436 23001
rect 16672 22992 16724 23044
rect 21732 22992 21784 23044
rect 22100 22992 22152 23044
rect 25596 23128 25648 23180
rect 27620 23196 27672 23248
rect 27804 23128 27856 23180
rect 28080 23128 28132 23180
rect 30748 23171 30800 23180
rect 30748 23137 30757 23171
rect 30757 23137 30791 23171
rect 30791 23137 30800 23171
rect 30748 23128 30800 23137
rect 37372 23196 37424 23248
rect 32128 23171 32180 23180
rect 32128 23137 32137 23171
rect 32137 23137 32171 23171
rect 32171 23137 32180 23171
rect 32128 23128 32180 23137
rect 33416 23128 33468 23180
rect 23848 23060 23900 23112
rect 27620 23060 27672 23112
rect 29276 23060 29328 23112
rect 31576 23060 31628 23112
rect 33324 22992 33376 23044
rect 34520 22992 34572 23044
rect 35164 23128 35216 23180
rect 41604 23264 41656 23316
rect 41880 23264 41932 23316
rect 45560 23264 45612 23316
rect 46112 23264 46164 23316
rect 53472 23264 53524 23316
rect 37648 23196 37700 23248
rect 44548 23239 44600 23248
rect 39764 23128 39816 23180
rect 41144 23128 41196 23180
rect 41880 23128 41932 23180
rect 42340 23128 42392 23180
rect 44548 23205 44557 23239
rect 44557 23205 44591 23239
rect 44591 23205 44600 23239
rect 44548 23196 44600 23205
rect 46388 23196 46440 23248
rect 48504 23196 48556 23248
rect 52368 23239 52420 23248
rect 52368 23205 52377 23239
rect 52377 23205 52411 23239
rect 52411 23205 52420 23239
rect 52368 23196 52420 23205
rect 46664 23128 46716 23180
rect 47400 23128 47452 23180
rect 35440 23060 35492 23112
rect 38108 23060 38160 23112
rect 37280 22992 37332 23044
rect 18604 22924 18656 22976
rect 20720 22924 20772 22976
rect 21640 22924 21692 22976
rect 21916 22924 21968 22976
rect 22560 22924 22612 22976
rect 23940 22924 23992 22976
rect 25596 22924 25648 22976
rect 26700 22967 26752 22976
rect 26700 22933 26709 22967
rect 26709 22933 26743 22967
rect 26743 22933 26752 22967
rect 26700 22924 26752 22933
rect 28172 22924 28224 22976
rect 29368 22924 29420 22976
rect 29552 22924 29604 22976
rect 32220 22924 32272 22976
rect 34244 22967 34296 22976
rect 34244 22933 34253 22967
rect 34253 22933 34287 22967
rect 34287 22933 34296 22967
rect 34244 22924 34296 22933
rect 36360 22924 36412 22976
rect 38200 22924 38252 22976
rect 38752 23060 38804 23112
rect 44548 23060 44600 23112
rect 44916 23103 44968 23112
rect 44916 23069 44925 23103
rect 44925 23069 44959 23103
rect 44959 23069 44968 23103
rect 44916 23060 44968 23069
rect 46204 23060 46256 23112
rect 47860 23128 47912 23180
rect 51724 23128 51776 23180
rect 52000 23128 52052 23180
rect 40592 22992 40644 23044
rect 40132 22967 40184 22976
rect 40132 22933 40141 22967
rect 40141 22933 40175 22967
rect 40175 22933 40184 22967
rect 40132 22924 40184 22933
rect 44364 22924 44416 22976
rect 47492 22992 47544 23044
rect 51080 22992 51132 23044
rect 47400 22924 47452 22976
rect 47860 22924 47912 22976
rect 51448 22967 51500 22976
rect 51448 22933 51457 22967
rect 51457 22933 51491 22967
rect 51491 22933 51500 22967
rect 51448 22924 51500 22933
rect 9947 22822 9999 22874
rect 10011 22822 10063 22874
rect 10075 22822 10127 22874
rect 10139 22822 10191 22874
rect 27878 22822 27930 22874
rect 27942 22822 27994 22874
rect 28006 22822 28058 22874
rect 28070 22822 28122 22874
rect 45808 22822 45860 22874
rect 45872 22822 45924 22874
rect 45936 22822 45988 22874
rect 46000 22822 46052 22874
rect 296 22720 348 22772
rect 6920 22695 6972 22704
rect 6920 22661 6929 22695
rect 6929 22661 6963 22695
rect 6963 22661 6972 22695
rect 6920 22652 6972 22661
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 2044 22516 2096 22568
rect 4068 22584 4120 22636
rect 4344 22584 4396 22636
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 7104 22584 7156 22636
rect 4896 22448 4948 22500
rect 3332 22380 3384 22432
rect 7012 22516 7064 22568
rect 8024 22516 8076 22568
rect 11060 22652 11112 22704
rect 11244 22652 11296 22704
rect 10416 22584 10468 22636
rect 9772 22516 9824 22568
rect 11152 22516 11204 22568
rect 12716 22516 12768 22568
rect 15108 22652 15160 22704
rect 16672 22695 16724 22704
rect 16672 22661 16681 22695
rect 16681 22661 16715 22695
rect 16715 22661 16724 22695
rect 16672 22652 16724 22661
rect 15384 22627 15436 22636
rect 15384 22593 15393 22627
rect 15393 22593 15427 22627
rect 15427 22593 15436 22627
rect 15384 22584 15436 22593
rect 5724 22448 5776 22500
rect 7380 22448 7432 22500
rect 9588 22448 9640 22500
rect 10508 22380 10560 22432
rect 11060 22380 11112 22432
rect 13084 22423 13136 22432
rect 13084 22389 13093 22423
rect 13093 22389 13127 22423
rect 13127 22389 13136 22423
rect 13084 22380 13136 22389
rect 18512 22720 18564 22772
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 23204 22720 23256 22772
rect 23480 22720 23532 22772
rect 24676 22720 24728 22772
rect 31484 22720 31536 22772
rect 33324 22720 33376 22772
rect 33692 22763 33744 22772
rect 33692 22729 33701 22763
rect 33701 22729 33735 22763
rect 33735 22729 33744 22763
rect 33692 22720 33744 22729
rect 34520 22720 34572 22772
rect 35072 22720 35124 22772
rect 37372 22720 37424 22772
rect 37740 22720 37792 22772
rect 38384 22720 38436 22772
rect 38752 22763 38804 22772
rect 38752 22729 38761 22763
rect 38761 22729 38795 22763
rect 38795 22729 38804 22763
rect 38752 22720 38804 22729
rect 41880 22720 41932 22772
rect 42800 22720 42852 22772
rect 43076 22720 43128 22772
rect 20720 22695 20772 22704
rect 20720 22661 20729 22695
rect 20729 22661 20763 22695
rect 20763 22661 20772 22695
rect 20720 22652 20772 22661
rect 20812 22652 20864 22704
rect 21640 22695 21692 22704
rect 21180 22584 21232 22636
rect 21640 22661 21649 22695
rect 21649 22661 21683 22695
rect 21683 22661 21692 22695
rect 21640 22652 21692 22661
rect 23296 22652 23348 22704
rect 21916 22584 21968 22636
rect 26700 22584 26752 22636
rect 28264 22652 28316 22704
rect 31576 22652 31628 22704
rect 28172 22584 28224 22636
rect 40592 22652 40644 22704
rect 51448 22720 51500 22772
rect 32128 22584 32180 22636
rect 20996 22559 21048 22568
rect 20996 22525 21005 22559
rect 21005 22525 21039 22559
rect 21039 22525 21048 22559
rect 20996 22516 21048 22525
rect 21088 22516 21140 22568
rect 24032 22559 24084 22568
rect 22192 22448 22244 22500
rect 23296 22448 23348 22500
rect 24032 22525 24041 22559
rect 24041 22525 24075 22559
rect 24075 22525 24084 22559
rect 24032 22516 24084 22525
rect 24216 22559 24268 22568
rect 24216 22525 24225 22559
rect 24225 22525 24259 22559
rect 24259 22525 24268 22559
rect 24216 22516 24268 22525
rect 24308 22559 24360 22568
rect 24308 22525 24317 22559
rect 24317 22525 24351 22559
rect 24351 22525 24360 22559
rect 25596 22559 25648 22568
rect 24308 22516 24360 22525
rect 25596 22525 25605 22559
rect 25605 22525 25639 22559
rect 25639 22525 25648 22559
rect 25596 22516 25648 22525
rect 27160 22516 27212 22568
rect 29276 22559 29328 22568
rect 22376 22380 22428 22432
rect 24216 22380 24268 22432
rect 25228 22448 25280 22500
rect 25504 22380 25556 22432
rect 26516 22380 26568 22432
rect 29276 22525 29285 22559
rect 29285 22525 29319 22559
rect 29319 22525 29328 22559
rect 29276 22516 29328 22525
rect 33508 22559 33560 22568
rect 28172 22491 28224 22500
rect 28172 22457 28181 22491
rect 28181 22457 28215 22491
rect 28215 22457 28224 22491
rect 28172 22448 28224 22457
rect 28264 22448 28316 22500
rect 29460 22448 29512 22500
rect 33508 22525 33517 22559
rect 33517 22525 33551 22559
rect 33551 22525 33560 22559
rect 33508 22516 33560 22525
rect 37188 22584 37240 22636
rect 38752 22584 38804 22636
rect 41604 22584 41656 22636
rect 42248 22584 42300 22636
rect 44364 22584 44416 22636
rect 48964 22584 49016 22636
rect 37740 22559 37792 22568
rect 28356 22423 28408 22432
rect 28356 22389 28365 22423
rect 28365 22389 28399 22423
rect 28399 22389 28408 22423
rect 28356 22380 28408 22389
rect 28816 22380 28868 22432
rect 32312 22448 32364 22500
rect 33416 22491 33468 22500
rect 33416 22457 33425 22491
rect 33425 22457 33459 22491
rect 33459 22457 33468 22491
rect 33416 22448 33468 22457
rect 37740 22525 37749 22559
rect 37749 22525 37783 22559
rect 37783 22525 37792 22559
rect 37740 22516 37792 22525
rect 38844 22516 38896 22568
rect 39488 22516 39540 22568
rect 40408 22516 40460 22568
rect 41880 22516 41932 22568
rect 42616 22516 42668 22568
rect 32220 22380 32272 22432
rect 37280 22448 37332 22500
rect 40224 22448 40276 22500
rect 41972 22448 42024 22500
rect 43076 22516 43128 22568
rect 46388 22516 46440 22568
rect 48596 22559 48648 22568
rect 48596 22525 48605 22559
rect 48605 22525 48639 22559
rect 48639 22525 48648 22559
rect 48596 22516 48648 22525
rect 43536 22491 43588 22500
rect 43536 22457 43545 22491
rect 43545 22457 43579 22491
rect 43579 22457 43588 22491
rect 43536 22448 43588 22457
rect 41236 22380 41288 22432
rect 44824 22380 44876 22432
rect 46296 22380 46348 22432
rect 49976 22423 50028 22432
rect 49976 22389 49985 22423
rect 49985 22389 50019 22423
rect 50019 22389 50028 22423
rect 49976 22380 50028 22389
rect 51816 22448 51868 22500
rect 52460 22516 52512 22568
rect 54116 22380 54168 22432
rect 18912 22278 18964 22330
rect 18976 22278 19028 22330
rect 19040 22278 19092 22330
rect 19104 22278 19156 22330
rect 36843 22278 36895 22330
rect 36907 22278 36959 22330
rect 36971 22278 37023 22330
rect 37035 22278 37087 22330
rect 2044 22219 2096 22228
rect 2044 22185 2053 22219
rect 2053 22185 2087 22219
rect 2087 22185 2096 22219
rect 2044 22176 2096 22185
rect 4252 22176 4304 22228
rect 4896 22219 4948 22228
rect 4896 22185 4905 22219
rect 4905 22185 4939 22219
rect 4939 22185 4948 22219
rect 4896 22176 4948 22185
rect 6644 22176 6696 22228
rect 6920 22176 6972 22228
rect 7104 22176 7156 22228
rect 13084 22176 13136 22228
rect 14832 22176 14884 22228
rect 20904 22176 20956 22228
rect 21916 22219 21968 22228
rect 2504 22083 2556 22092
rect 2504 22049 2513 22083
rect 2513 22049 2547 22083
rect 2547 22049 2556 22083
rect 2504 22040 2556 22049
rect 5724 22108 5776 22160
rect 4620 22083 4672 22092
rect 4620 22049 4629 22083
rect 4629 22049 4663 22083
rect 4663 22049 4672 22083
rect 4620 22040 4672 22049
rect 6184 22040 6236 22092
rect 6736 22040 6788 22092
rect 7012 22040 7064 22092
rect 8576 22083 8628 22092
rect 5816 21972 5868 22024
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 9680 22040 9732 22092
rect 10600 22083 10652 22092
rect 10600 22049 10609 22083
rect 10609 22049 10643 22083
rect 10643 22049 10652 22083
rect 10600 22040 10652 22049
rect 10876 22040 10928 22092
rect 11060 22040 11112 22092
rect 11612 22040 11664 22092
rect 12716 22040 12768 22092
rect 21916 22185 21925 22219
rect 21925 22185 21959 22219
rect 21959 22185 21968 22219
rect 21916 22176 21968 22185
rect 23204 22176 23256 22228
rect 29092 22176 29144 22228
rect 29460 22176 29512 22228
rect 42156 22176 42208 22228
rect 42340 22219 42392 22228
rect 42340 22185 42349 22219
rect 42349 22185 42383 22219
rect 42383 22185 42392 22219
rect 42340 22176 42392 22185
rect 45008 22176 45060 22228
rect 48964 22176 49016 22228
rect 51448 22176 51500 22228
rect 21640 22108 21692 22160
rect 33508 22108 33560 22160
rect 21456 22040 21508 22092
rect 22560 22083 22612 22092
rect 22560 22049 22569 22083
rect 22569 22049 22603 22083
rect 22603 22049 22612 22083
rect 22560 22040 22612 22049
rect 23756 22083 23808 22092
rect 23756 22049 23765 22083
rect 23765 22049 23799 22083
rect 23799 22049 23808 22083
rect 23756 22040 23808 22049
rect 24308 22083 24360 22092
rect 24308 22049 24317 22083
rect 24317 22049 24351 22083
rect 24351 22049 24360 22083
rect 24308 22040 24360 22049
rect 26700 22040 26752 22092
rect 28172 22040 28224 22092
rect 33968 22083 34020 22092
rect 33968 22049 33977 22083
rect 33977 22049 34011 22083
rect 34011 22049 34020 22083
rect 33968 22040 34020 22049
rect 34152 22083 34204 22092
rect 34152 22049 34161 22083
rect 34161 22049 34195 22083
rect 34195 22049 34204 22083
rect 34152 22040 34204 22049
rect 34888 22083 34940 22092
rect 34888 22049 34897 22083
rect 34897 22049 34931 22083
rect 34931 22049 34940 22083
rect 34888 22040 34940 22049
rect 41328 22108 41380 22160
rect 40132 22040 40184 22092
rect 17132 22015 17184 22024
rect 7104 21904 7156 21956
rect 7288 21904 7340 21956
rect 9404 21836 9456 21888
rect 9588 21904 9640 21956
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 11244 21904 11296 21956
rect 21640 21904 21692 21956
rect 22284 21904 22336 21956
rect 23480 21904 23532 21956
rect 23664 21947 23716 21956
rect 23664 21913 23673 21947
rect 23673 21913 23707 21947
rect 23707 21913 23716 21947
rect 23664 21904 23716 21913
rect 23848 21972 23900 22024
rect 24768 21972 24820 22024
rect 28264 21972 28316 22024
rect 9680 21836 9732 21888
rect 11520 21879 11572 21888
rect 11520 21845 11529 21879
rect 11529 21845 11563 21879
rect 11563 21845 11572 21879
rect 11520 21836 11572 21845
rect 15568 21836 15620 21888
rect 15844 21836 15896 21888
rect 21364 21879 21416 21888
rect 21364 21845 21373 21879
rect 21373 21845 21407 21879
rect 21407 21845 21416 21879
rect 21364 21836 21416 21845
rect 22744 21836 22796 21888
rect 26700 21836 26752 21888
rect 27160 21879 27212 21888
rect 27160 21845 27169 21879
rect 27169 21845 27203 21879
rect 27203 21845 27212 21879
rect 27160 21836 27212 21845
rect 27620 21904 27672 21956
rect 29000 21972 29052 22024
rect 29368 21972 29420 22024
rect 31024 21972 31076 22024
rect 32772 21972 32824 22024
rect 29092 21836 29144 21888
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 35624 21836 35676 21888
rect 38200 21836 38252 21888
rect 39856 22015 39908 22024
rect 39856 21981 39865 22015
rect 39865 21981 39899 22015
rect 39899 21981 39908 22015
rect 39856 21972 39908 21981
rect 44916 22108 44968 22160
rect 51724 22151 51776 22160
rect 51724 22117 51733 22151
rect 51733 22117 51767 22151
rect 51767 22117 51776 22151
rect 51724 22108 51776 22117
rect 42248 22083 42300 22092
rect 42248 22049 42257 22083
rect 42257 22049 42291 22083
rect 42291 22049 42300 22083
rect 42248 22040 42300 22049
rect 42616 22040 42668 22092
rect 42800 22040 42852 22092
rect 44272 22083 44324 22092
rect 44272 22049 44281 22083
rect 44281 22049 44315 22083
rect 44315 22049 44324 22083
rect 44824 22083 44876 22092
rect 44272 22040 44324 22049
rect 44824 22049 44833 22083
rect 44833 22049 44867 22083
rect 44867 22049 44876 22083
rect 44824 22040 44876 22049
rect 46112 22040 46164 22092
rect 49792 22040 49844 22092
rect 50068 22083 50120 22092
rect 50068 22049 50077 22083
rect 50077 22049 50111 22083
rect 50111 22049 50120 22083
rect 50068 22040 50120 22049
rect 50712 22040 50764 22092
rect 46296 22015 46348 22024
rect 41328 21836 41380 21888
rect 42616 21879 42668 21888
rect 42616 21845 42625 21879
rect 42625 21845 42659 21879
rect 42659 21845 42668 21879
rect 42616 21836 42668 21845
rect 45376 21836 45428 21888
rect 46296 21981 46305 22015
rect 46305 21981 46339 22015
rect 46339 21981 46348 22015
rect 46296 21972 46348 21981
rect 47676 22015 47728 22024
rect 47676 21981 47685 22015
rect 47685 21981 47719 22015
rect 47719 21981 47728 22015
rect 47676 21972 47728 21981
rect 52276 21904 52328 21956
rect 46112 21879 46164 21888
rect 46112 21845 46121 21879
rect 46121 21845 46155 21879
rect 46155 21845 46164 21879
rect 46112 21836 46164 21845
rect 52000 21836 52052 21888
rect 52460 21836 52512 21888
rect 9947 21734 9999 21786
rect 10011 21734 10063 21786
rect 10075 21734 10127 21786
rect 10139 21734 10191 21786
rect 27878 21734 27930 21786
rect 27942 21734 27994 21786
rect 28006 21734 28058 21786
rect 28070 21734 28122 21786
rect 45808 21734 45860 21786
rect 45872 21734 45924 21786
rect 45936 21734 45988 21786
rect 46000 21734 46052 21786
rect 5816 21675 5868 21684
rect 5816 21641 5825 21675
rect 5825 21641 5859 21675
rect 5859 21641 5868 21675
rect 5816 21632 5868 21641
rect 6828 21632 6880 21684
rect 10600 21632 10652 21684
rect 14832 21675 14884 21684
rect 14832 21641 14841 21675
rect 14841 21641 14875 21675
rect 14875 21641 14884 21675
rect 14832 21632 14884 21641
rect 7104 21607 7156 21616
rect 7104 21573 7113 21607
rect 7113 21573 7147 21607
rect 7147 21573 7156 21607
rect 7104 21564 7156 21573
rect 3332 21496 3384 21548
rect 5632 21428 5684 21480
rect 6920 21496 6972 21548
rect 10968 21564 11020 21616
rect 7012 21471 7064 21480
rect 7012 21437 7021 21471
rect 7021 21437 7055 21471
rect 7055 21437 7064 21471
rect 7012 21428 7064 21437
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 9588 21496 9640 21548
rect 12256 21496 12308 21548
rect 7472 21428 7524 21480
rect 4620 21360 4672 21412
rect 10324 21360 10376 21412
rect 5724 21292 5776 21344
rect 10968 21428 11020 21480
rect 12348 21428 12400 21480
rect 17040 21632 17092 21684
rect 17132 21632 17184 21684
rect 20996 21675 21048 21684
rect 20996 21641 21005 21675
rect 21005 21641 21039 21675
rect 21039 21641 21048 21675
rect 20996 21632 21048 21641
rect 22376 21675 22428 21684
rect 22376 21641 22385 21675
rect 22385 21641 22419 21675
rect 22419 21641 22428 21675
rect 22376 21632 22428 21641
rect 28264 21632 28316 21684
rect 46112 21632 46164 21684
rect 46296 21632 46348 21684
rect 48596 21632 48648 21684
rect 17408 21564 17460 21616
rect 22560 21564 22612 21616
rect 12716 21496 12768 21548
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 14832 21428 14884 21480
rect 15568 21471 15620 21480
rect 15568 21437 15577 21471
rect 15577 21437 15611 21471
rect 15611 21437 15620 21471
rect 15568 21428 15620 21437
rect 16028 21471 16080 21480
rect 16028 21437 16037 21471
rect 16037 21437 16071 21471
rect 16071 21437 16080 21471
rect 16028 21428 16080 21437
rect 17132 21428 17184 21480
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 19800 21428 19852 21480
rect 22376 21428 22428 21480
rect 23848 21496 23900 21548
rect 26792 21564 26844 21616
rect 27712 21607 27764 21616
rect 27712 21573 27721 21607
rect 27721 21573 27755 21607
rect 27755 21573 27764 21607
rect 27712 21564 27764 21573
rect 32772 21607 32824 21616
rect 32772 21573 32781 21607
rect 32781 21573 32815 21607
rect 32815 21573 32824 21607
rect 32772 21564 32824 21573
rect 34888 21564 34940 21616
rect 27804 21496 27856 21548
rect 41052 21564 41104 21616
rect 38292 21539 38344 21548
rect 38292 21505 38301 21539
rect 38301 21505 38335 21539
rect 38335 21505 38344 21539
rect 38292 21496 38344 21505
rect 39856 21496 39908 21548
rect 43536 21539 43588 21548
rect 43536 21505 43545 21539
rect 43545 21505 43579 21539
rect 43579 21505 43588 21539
rect 43536 21496 43588 21505
rect 51724 21539 51776 21548
rect 51724 21505 51733 21539
rect 51733 21505 51767 21539
rect 51767 21505 51776 21539
rect 51724 21496 51776 21505
rect 52000 21539 52052 21548
rect 52000 21505 52009 21539
rect 52009 21505 52043 21539
rect 52043 21505 52052 21539
rect 52000 21496 52052 21505
rect 52092 21496 52144 21548
rect 23572 21428 23624 21480
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 25228 21471 25280 21480
rect 12716 21360 12768 21412
rect 18604 21360 18656 21412
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 26424 21428 26476 21480
rect 27160 21428 27212 21480
rect 28816 21428 28868 21480
rect 29736 21471 29788 21480
rect 29736 21437 29745 21471
rect 29745 21437 29779 21471
rect 29779 21437 29788 21471
rect 29736 21428 29788 21437
rect 31024 21471 31076 21480
rect 31024 21437 31033 21471
rect 31033 21437 31067 21471
rect 31067 21437 31076 21471
rect 31024 21428 31076 21437
rect 31116 21428 31168 21480
rect 33784 21471 33836 21480
rect 33784 21437 33793 21471
rect 33793 21437 33827 21471
rect 33827 21437 33836 21471
rect 33784 21428 33836 21437
rect 35348 21471 35400 21480
rect 35348 21437 35357 21471
rect 35357 21437 35391 21471
rect 35391 21437 35400 21471
rect 35348 21428 35400 21437
rect 35624 21471 35676 21480
rect 35624 21437 35633 21471
rect 35633 21437 35667 21471
rect 35667 21437 35676 21471
rect 35624 21428 35676 21437
rect 35992 21428 36044 21480
rect 38200 21428 38252 21480
rect 38384 21471 38436 21480
rect 38384 21437 38393 21471
rect 38393 21437 38427 21471
rect 38427 21437 38436 21471
rect 38384 21428 38436 21437
rect 38752 21428 38804 21480
rect 24124 21360 24176 21412
rect 28908 21360 28960 21412
rect 16948 21292 17000 21344
rect 17040 21292 17092 21344
rect 22284 21292 22336 21344
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 23848 21292 23900 21344
rect 25228 21292 25280 21344
rect 27804 21292 27856 21344
rect 30748 21292 30800 21344
rect 30932 21292 30984 21344
rect 37188 21360 37240 21412
rect 41052 21428 41104 21480
rect 41144 21292 41196 21344
rect 42984 21292 43036 21344
rect 47032 21471 47084 21480
rect 47032 21437 47041 21471
rect 47041 21437 47075 21471
rect 47075 21437 47084 21471
rect 47032 21428 47084 21437
rect 43168 21292 43220 21344
rect 47860 21292 47912 21344
rect 18912 21190 18964 21242
rect 18976 21190 19028 21242
rect 19040 21190 19092 21242
rect 19104 21190 19156 21242
rect 36843 21190 36895 21242
rect 36907 21190 36959 21242
rect 36971 21190 37023 21242
rect 37035 21190 37087 21242
rect 5632 21131 5684 21140
rect 5632 21097 5641 21131
rect 5641 21097 5675 21131
rect 5675 21097 5684 21131
rect 5632 21088 5684 21097
rect 6644 21020 6696 21072
rect 7012 21020 7064 21072
rect 5816 20952 5868 21004
rect 7380 20995 7432 21004
rect 7380 20961 7386 20995
rect 7386 20961 7432 20995
rect 7380 20952 7432 20961
rect 4804 20884 4856 20936
rect 9588 21088 9640 21140
rect 12348 21088 12400 21140
rect 13820 21088 13872 21140
rect 10876 21020 10928 21072
rect 9404 20952 9456 21004
rect 10968 20952 11020 21004
rect 13268 20952 13320 21004
rect 15108 21088 15160 21140
rect 16028 21088 16080 21140
rect 17040 21131 17092 21140
rect 17040 21097 17049 21131
rect 17049 21097 17083 21131
rect 17083 21097 17092 21131
rect 17040 21088 17092 21097
rect 19800 21131 19852 21140
rect 19800 21097 19809 21131
rect 19809 21097 19843 21131
rect 19843 21097 19852 21131
rect 19800 21088 19852 21097
rect 17132 21020 17184 21072
rect 15844 20995 15896 21004
rect 15844 20961 15853 20995
rect 15853 20961 15887 20995
rect 15887 20961 15896 20995
rect 15844 20952 15896 20961
rect 12624 20927 12676 20936
rect 7472 20859 7524 20868
rect 7472 20825 7481 20859
rect 7481 20825 7515 20859
rect 7515 20825 7524 20859
rect 7472 20816 7524 20825
rect 7932 20816 7984 20868
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 16948 20952 17000 21004
rect 18052 20952 18104 21004
rect 18512 20952 18564 21004
rect 19708 21020 19760 21072
rect 17040 20884 17092 20936
rect 25688 21088 25740 21140
rect 21548 21020 21600 21072
rect 20996 20952 21048 21004
rect 23756 21020 23808 21072
rect 24768 21063 24820 21072
rect 24768 21029 24777 21063
rect 24777 21029 24811 21063
rect 24811 21029 24820 21063
rect 24768 21020 24820 21029
rect 22744 20995 22796 21004
rect 22744 20961 22753 20995
rect 22753 20961 22787 20995
rect 22787 20961 22796 20995
rect 22744 20952 22796 20961
rect 26792 21020 26844 21072
rect 26884 20952 26936 21004
rect 17776 20816 17828 20868
rect 17960 20816 18012 20868
rect 28724 21020 28776 21072
rect 29000 21020 29052 21072
rect 31116 21063 31168 21072
rect 29828 20995 29880 21004
rect 29828 20961 29837 20995
rect 29837 20961 29871 20995
rect 29871 20961 29880 20995
rect 29828 20952 29880 20961
rect 30196 20952 30248 21004
rect 30748 20995 30800 21004
rect 30748 20961 30757 20995
rect 30757 20961 30791 20995
rect 30791 20961 30800 20995
rect 30748 20952 30800 20961
rect 31116 21029 31125 21063
rect 31125 21029 31159 21063
rect 31159 21029 31168 21063
rect 31116 21020 31168 21029
rect 35348 21088 35400 21140
rect 35992 21131 36044 21140
rect 35992 21097 36001 21131
rect 36001 21097 36035 21131
rect 36035 21097 36044 21131
rect 35992 21088 36044 21097
rect 33232 20995 33284 21004
rect 33232 20961 33241 20995
rect 33241 20961 33275 20995
rect 33275 20961 33284 20995
rect 33232 20952 33284 20961
rect 34796 21020 34848 21072
rect 32036 20884 32088 20936
rect 34152 20952 34204 21004
rect 36452 21088 36504 21140
rect 40224 21131 40276 21140
rect 40224 21097 40233 21131
rect 40233 21097 40267 21131
rect 40267 21097 40276 21131
rect 40224 21088 40276 21097
rect 41696 21088 41748 21140
rect 42800 21088 42852 21140
rect 42984 21088 43036 21140
rect 45376 21088 45428 21140
rect 45652 21088 45704 21140
rect 40040 21020 40092 21072
rect 40776 21020 40828 21072
rect 43168 21020 43220 21072
rect 34796 20927 34848 20936
rect 34796 20893 34805 20927
rect 34805 20893 34839 20927
rect 34839 20893 34848 20927
rect 34796 20884 34848 20893
rect 44456 20952 44508 21004
rect 45928 20995 45980 21004
rect 45928 20961 45937 20995
rect 45937 20961 45971 20995
rect 45971 20961 45980 20995
rect 45928 20952 45980 20961
rect 46940 21088 46992 21140
rect 51724 21088 51776 21140
rect 47032 21063 47084 21072
rect 23572 20816 23624 20868
rect 24952 20816 25004 20868
rect 11152 20748 11204 20800
rect 11336 20748 11388 20800
rect 17500 20791 17552 20800
rect 17500 20757 17509 20791
rect 17509 20757 17543 20791
rect 17543 20757 17552 20791
rect 17500 20748 17552 20757
rect 18052 20748 18104 20800
rect 25228 20748 25280 20800
rect 26700 20748 26752 20800
rect 28632 20791 28684 20800
rect 28632 20757 28641 20791
rect 28641 20757 28675 20791
rect 28675 20757 28684 20791
rect 28632 20748 28684 20757
rect 35808 20748 35860 20800
rect 36176 20816 36228 20868
rect 38936 20927 38988 20936
rect 36452 20791 36504 20800
rect 36452 20757 36461 20791
rect 36461 20757 36495 20791
rect 36495 20757 36504 20791
rect 36452 20748 36504 20757
rect 38292 20748 38344 20800
rect 38936 20893 38945 20927
rect 38945 20893 38979 20927
rect 38979 20893 38988 20927
rect 38936 20884 38988 20893
rect 40224 20884 40276 20936
rect 44272 20884 44324 20936
rect 46664 20995 46716 21004
rect 46664 20961 46673 20995
rect 46673 20961 46707 20995
rect 46707 20961 46716 20995
rect 46664 20952 46716 20961
rect 47032 21029 47041 21063
rect 47041 21029 47075 21063
rect 47075 21029 47084 21063
rect 47032 21020 47084 21029
rect 48412 20952 48464 21004
rect 50068 21020 50120 21072
rect 50160 20995 50212 21004
rect 50160 20961 50169 20995
rect 50169 20961 50203 20995
rect 50203 20961 50212 20995
rect 50160 20952 50212 20961
rect 39120 20748 39172 20800
rect 44456 20791 44508 20800
rect 44456 20757 44465 20791
rect 44465 20757 44499 20791
rect 44499 20757 44508 20791
rect 44456 20748 44508 20757
rect 46664 20748 46716 20800
rect 52276 20748 52328 20800
rect 9947 20646 9999 20698
rect 10011 20646 10063 20698
rect 10075 20646 10127 20698
rect 10139 20646 10191 20698
rect 27878 20646 27930 20698
rect 27942 20646 27994 20698
rect 28006 20646 28058 20698
rect 28070 20646 28122 20698
rect 45808 20646 45860 20698
rect 45872 20646 45924 20698
rect 45936 20646 45988 20698
rect 46000 20646 46052 20698
rect 5816 20587 5868 20596
rect 5816 20553 5825 20587
rect 5825 20553 5859 20587
rect 5859 20553 5868 20587
rect 5816 20544 5868 20553
rect 12624 20544 12676 20596
rect 15108 20587 15160 20596
rect 15108 20553 15117 20587
rect 15117 20553 15151 20587
rect 15151 20553 15160 20587
rect 15108 20544 15160 20553
rect 16120 20544 16172 20596
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 24952 20587 25004 20596
rect 24952 20553 24961 20587
rect 24961 20553 24995 20587
rect 24995 20553 25004 20587
rect 24952 20544 25004 20553
rect 26976 20544 27028 20596
rect 44456 20544 44508 20596
rect 50160 20544 50212 20596
rect 4804 20476 4856 20528
rect 5264 20476 5316 20528
rect 3516 20383 3568 20392
rect 3516 20349 3525 20383
rect 3525 20349 3559 20383
rect 3559 20349 3568 20383
rect 3516 20340 3568 20349
rect 3700 20383 3752 20392
rect 3700 20349 3709 20383
rect 3709 20349 3743 20383
rect 3743 20349 3752 20383
rect 3700 20340 3752 20349
rect 4252 20383 4304 20392
rect 4252 20349 4261 20383
rect 4261 20349 4295 20383
rect 4295 20349 4304 20383
rect 5724 20383 5776 20392
rect 4252 20340 4304 20349
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 6920 20340 6972 20392
rect 7932 20383 7984 20392
rect 7932 20349 7941 20383
rect 7941 20349 7975 20383
rect 7975 20349 7984 20383
rect 7932 20340 7984 20349
rect 8392 20340 8444 20392
rect 12716 20476 12768 20528
rect 16488 20476 16540 20528
rect 24032 20476 24084 20528
rect 24308 20519 24360 20528
rect 24308 20485 24332 20519
rect 24332 20485 24360 20519
rect 24308 20476 24360 20485
rect 26792 20519 26844 20528
rect 26792 20485 26801 20519
rect 26801 20485 26835 20519
rect 26835 20485 26844 20519
rect 26792 20476 26844 20485
rect 30196 20519 30248 20528
rect 30196 20485 30205 20519
rect 30205 20485 30239 20519
rect 30239 20485 30248 20519
rect 30196 20476 30248 20485
rect 11336 20408 11388 20460
rect 13268 20383 13320 20392
rect 5908 20272 5960 20324
rect 13268 20349 13277 20383
rect 13277 20349 13311 20383
rect 13311 20349 13320 20383
rect 13268 20340 13320 20349
rect 13544 20383 13596 20392
rect 13544 20349 13553 20383
rect 13553 20349 13587 20383
rect 13587 20349 13596 20383
rect 13544 20340 13596 20349
rect 15844 20408 15896 20460
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 17960 20340 18012 20392
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 18512 20340 18564 20392
rect 10416 20204 10468 20256
rect 20536 20272 20588 20324
rect 21272 20340 21324 20392
rect 23020 20408 23072 20460
rect 24124 20408 24176 20460
rect 24952 20408 25004 20460
rect 25412 20408 25464 20460
rect 27712 20408 27764 20460
rect 28632 20408 28684 20460
rect 31208 20408 31260 20460
rect 38936 20476 38988 20528
rect 25872 20383 25924 20392
rect 25872 20349 25881 20383
rect 25881 20349 25915 20383
rect 25915 20349 25924 20383
rect 25872 20340 25924 20349
rect 26332 20383 26384 20392
rect 26332 20349 26341 20383
rect 26341 20349 26375 20383
rect 26375 20349 26384 20383
rect 26332 20340 26384 20349
rect 26424 20383 26476 20392
rect 26424 20349 26433 20383
rect 26433 20349 26467 20383
rect 26467 20349 26476 20383
rect 26424 20340 26476 20349
rect 24124 20315 24176 20324
rect 24124 20281 24133 20315
rect 24133 20281 24167 20315
rect 24167 20281 24176 20315
rect 24124 20272 24176 20281
rect 25412 20272 25464 20324
rect 25688 20272 25740 20324
rect 28908 20272 28960 20324
rect 12164 20204 12216 20256
rect 14188 20204 14240 20256
rect 18328 20204 18380 20256
rect 20352 20247 20404 20256
rect 20352 20213 20361 20247
rect 20361 20213 20395 20247
rect 20395 20213 20404 20247
rect 20352 20204 20404 20213
rect 23388 20204 23440 20256
rect 32036 20340 32088 20392
rect 32404 20383 32456 20392
rect 32404 20349 32413 20383
rect 32413 20349 32447 20383
rect 32447 20349 32456 20383
rect 32404 20340 32456 20349
rect 35808 20408 35860 20460
rect 38108 20451 38160 20460
rect 38108 20417 38117 20451
rect 38117 20417 38151 20451
rect 38151 20417 38160 20451
rect 38108 20408 38160 20417
rect 33232 20272 33284 20324
rect 38016 20340 38068 20392
rect 38292 20383 38344 20392
rect 38292 20349 38301 20383
rect 38301 20349 38335 20383
rect 38335 20349 38344 20383
rect 38292 20340 38344 20349
rect 40040 20340 40092 20392
rect 41788 20408 41840 20460
rect 45560 20408 45612 20460
rect 50712 20519 50764 20528
rect 50712 20485 50721 20519
rect 50721 20485 50755 20519
rect 50755 20485 50764 20519
rect 50712 20476 50764 20485
rect 37280 20315 37332 20324
rect 31116 20204 31168 20256
rect 37280 20281 37289 20315
rect 37289 20281 37323 20315
rect 37323 20281 37332 20315
rect 37280 20272 37332 20281
rect 38476 20272 38528 20324
rect 35900 20204 35952 20256
rect 42892 20340 42944 20392
rect 46756 20383 46808 20392
rect 46112 20272 46164 20324
rect 46756 20349 46765 20383
rect 46765 20349 46799 20383
rect 46799 20349 46808 20383
rect 46756 20340 46808 20349
rect 48412 20383 48464 20392
rect 48412 20349 48421 20383
rect 48421 20349 48455 20383
rect 48455 20349 48464 20383
rect 48412 20340 48464 20349
rect 46940 20272 46992 20324
rect 50712 20340 50764 20392
rect 52092 20340 52144 20392
rect 53380 20340 53432 20392
rect 42984 20204 43036 20256
rect 46296 20204 46348 20256
rect 49240 20204 49292 20256
rect 51356 20272 51408 20324
rect 52000 20272 52052 20324
rect 52276 20204 52328 20256
rect 52920 20247 52972 20256
rect 52920 20213 52929 20247
rect 52929 20213 52963 20247
rect 52963 20213 52972 20247
rect 52920 20204 52972 20213
rect 18912 20102 18964 20154
rect 18976 20102 19028 20154
rect 19040 20102 19092 20154
rect 19104 20102 19156 20154
rect 36843 20102 36895 20154
rect 36907 20102 36959 20154
rect 36971 20102 37023 20154
rect 37035 20102 37087 20154
rect 3516 20000 3568 20052
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 9680 20000 9732 20052
rect 16304 20000 16356 20052
rect 18052 20000 18104 20052
rect 21272 20000 21324 20052
rect 23388 20043 23440 20052
rect 23388 20009 23397 20043
rect 23397 20009 23431 20043
rect 23431 20009 23440 20043
rect 23388 20000 23440 20009
rect 24124 20000 24176 20052
rect 30472 20000 30524 20052
rect 30748 20000 30800 20052
rect 31116 20000 31168 20052
rect 32220 20000 32272 20052
rect 32312 20000 32364 20052
rect 36176 20000 36228 20052
rect 38476 20043 38528 20052
rect 38476 20009 38485 20043
rect 38485 20009 38519 20043
rect 38519 20009 38528 20043
rect 38476 20000 38528 20009
rect 3332 19907 3384 19916
rect 3332 19873 3341 19907
rect 3341 19873 3375 19907
rect 3375 19873 3384 19907
rect 3332 19864 3384 19873
rect 6644 19864 6696 19916
rect 6736 19864 6788 19916
rect 11336 19932 11388 19984
rect 12164 19907 12216 19916
rect 1768 19839 1820 19848
rect 1768 19805 1771 19839
rect 1771 19805 1805 19839
rect 1805 19805 1820 19839
rect 1768 19796 1820 19805
rect 6184 19839 6236 19848
rect 6184 19805 6193 19839
rect 6193 19805 6227 19839
rect 6227 19805 6236 19839
rect 6184 19796 6236 19805
rect 1768 19660 1820 19712
rect 5908 19660 5960 19712
rect 8576 19796 8628 19848
rect 9588 19796 9640 19848
rect 12164 19873 12173 19907
rect 12173 19873 12207 19907
rect 12207 19873 12216 19907
rect 12164 19864 12216 19873
rect 12900 19907 12952 19916
rect 12900 19873 12909 19907
rect 12909 19873 12943 19907
rect 12943 19873 12952 19907
rect 12900 19864 12952 19873
rect 13544 19932 13596 19984
rect 14188 19907 14240 19916
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 16304 19864 16356 19916
rect 17500 19864 17552 19916
rect 16488 19796 16540 19848
rect 17224 19796 17276 19848
rect 18236 19864 18288 19916
rect 18512 19864 18564 19916
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 20352 19864 20404 19916
rect 27712 19932 27764 19984
rect 29000 19932 29052 19984
rect 34796 19932 34848 19984
rect 38384 19932 38436 19984
rect 19708 19796 19760 19848
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 21548 19796 21600 19848
rect 12900 19728 12952 19780
rect 17868 19728 17920 19780
rect 15752 19703 15804 19712
rect 15752 19669 15761 19703
rect 15761 19669 15795 19703
rect 15795 19669 15804 19703
rect 15752 19660 15804 19669
rect 18052 19660 18104 19712
rect 18328 19660 18380 19712
rect 30932 19907 30984 19916
rect 30932 19873 30941 19907
rect 30941 19873 30975 19907
rect 30975 19873 30984 19907
rect 30932 19864 30984 19873
rect 31300 19864 31352 19916
rect 32772 19864 32824 19916
rect 33232 19907 33284 19916
rect 26332 19796 26384 19848
rect 27712 19796 27764 19848
rect 29000 19796 29052 19848
rect 29184 19839 29236 19848
rect 29184 19805 29193 19839
rect 29193 19805 29227 19839
rect 29227 19805 29236 19839
rect 29184 19796 29236 19805
rect 33232 19873 33241 19907
rect 33241 19873 33275 19907
rect 33275 19873 33284 19907
rect 33232 19864 33284 19873
rect 37372 19864 37424 19916
rect 45560 20000 45612 20052
rect 45652 20000 45704 20052
rect 46020 20000 46072 20052
rect 46388 20000 46440 20052
rect 52920 20000 52972 20052
rect 53380 20043 53432 20052
rect 53380 20009 53389 20043
rect 53389 20009 53423 20043
rect 53423 20009 53432 20043
rect 53380 20000 53432 20009
rect 35348 19796 35400 19848
rect 38292 19796 38344 19848
rect 39764 19907 39816 19916
rect 39764 19873 39773 19907
rect 39773 19873 39807 19907
rect 39807 19873 39816 19907
rect 39764 19864 39816 19873
rect 50712 19932 50764 19984
rect 51724 19932 51776 19984
rect 41052 19864 41104 19916
rect 45744 19864 45796 19916
rect 46296 19907 46348 19916
rect 46020 19839 46072 19848
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 24308 19660 24360 19712
rect 32588 19728 32640 19780
rect 40132 19771 40184 19780
rect 40132 19737 40141 19771
rect 40141 19737 40175 19771
rect 40175 19737 40184 19771
rect 40132 19728 40184 19737
rect 46020 19805 46029 19839
rect 46029 19805 46063 19839
rect 46063 19805 46072 19839
rect 46020 19796 46072 19805
rect 46296 19873 46305 19907
rect 46305 19873 46339 19907
rect 46339 19873 46348 19907
rect 46296 19864 46348 19873
rect 48596 19864 48648 19916
rect 49240 19907 49292 19916
rect 49240 19873 49249 19907
rect 49249 19873 49283 19907
rect 49283 19873 49292 19907
rect 49240 19864 49292 19873
rect 48504 19796 48556 19848
rect 52736 19796 52788 19848
rect 41052 19703 41104 19712
rect 41052 19669 41061 19703
rect 41061 19669 41095 19703
rect 41095 19669 41104 19703
rect 41052 19660 41104 19669
rect 41420 19703 41472 19712
rect 41420 19669 41429 19703
rect 41429 19669 41463 19703
rect 41463 19669 41472 19703
rect 41420 19660 41472 19669
rect 46940 19660 46992 19712
rect 47400 19703 47452 19712
rect 47400 19669 47409 19703
rect 47409 19669 47443 19703
rect 47443 19669 47452 19703
rect 47400 19660 47452 19669
rect 9947 19558 9999 19610
rect 10011 19558 10063 19610
rect 10075 19558 10127 19610
rect 10139 19558 10191 19610
rect 27878 19558 27930 19610
rect 27942 19558 27994 19610
rect 28006 19558 28058 19610
rect 28070 19558 28122 19610
rect 45808 19558 45860 19610
rect 45872 19558 45924 19610
rect 45936 19558 45988 19610
rect 46000 19558 46052 19610
rect 3700 19456 3752 19508
rect 10508 19499 10560 19508
rect 10508 19465 10517 19499
rect 10517 19465 10551 19499
rect 10551 19465 10560 19499
rect 10508 19456 10560 19465
rect 16488 19499 16540 19508
rect 16488 19465 16497 19499
rect 16497 19465 16531 19499
rect 16531 19465 16540 19499
rect 16488 19456 16540 19465
rect 18512 19499 18564 19508
rect 18512 19465 18521 19499
rect 18521 19465 18555 19499
rect 18555 19465 18564 19499
rect 18512 19456 18564 19465
rect 18604 19456 18656 19508
rect 27344 19456 27396 19508
rect 30472 19499 30524 19508
rect 30472 19465 30481 19499
rect 30481 19465 30515 19499
rect 30515 19465 30524 19499
rect 30472 19456 30524 19465
rect 32220 19456 32272 19508
rect 41052 19456 41104 19508
rect 42892 19499 42944 19508
rect 42892 19465 42901 19499
rect 42901 19465 42935 19499
rect 42935 19465 42944 19499
rect 42892 19456 42944 19465
rect 44824 19456 44876 19508
rect 47400 19456 47452 19508
rect 6184 19388 6236 19440
rect 11980 19388 12032 19440
rect 17960 19388 18012 19440
rect 18236 19388 18288 19440
rect 20536 19388 20588 19440
rect 26516 19388 26568 19440
rect 27804 19388 27856 19440
rect 52368 19388 52420 19440
rect 10416 19320 10468 19372
rect 22008 19320 22060 19372
rect 27620 19320 27672 19372
rect 34520 19320 34572 19372
rect 2964 19252 3016 19304
rect 4160 19252 4212 19304
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 6644 19252 6696 19304
rect 6736 19184 6788 19236
rect 8300 19252 8352 19304
rect 10140 19252 10192 19304
rect 3148 19116 3200 19168
rect 6920 19116 6972 19168
rect 8852 19184 8904 19236
rect 8668 19116 8720 19168
rect 9588 19116 9640 19168
rect 11336 19252 11388 19304
rect 13084 19252 13136 19304
rect 16304 19295 16356 19304
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 19432 19295 19484 19304
rect 19432 19261 19441 19295
rect 19441 19261 19475 19295
rect 19475 19261 19484 19295
rect 19432 19252 19484 19261
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 21456 19252 21508 19304
rect 23664 19252 23716 19304
rect 13452 19116 13504 19168
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 18328 19116 18380 19168
rect 23940 19295 23992 19304
rect 23940 19261 23949 19295
rect 23949 19261 23983 19295
rect 23983 19261 23992 19295
rect 23940 19252 23992 19261
rect 25228 19252 25280 19304
rect 25320 19252 25372 19304
rect 25872 19184 25924 19236
rect 30012 19252 30064 19304
rect 30748 19252 30800 19304
rect 27712 19227 27764 19236
rect 27712 19193 27721 19227
rect 27721 19193 27755 19227
rect 27755 19193 27764 19227
rect 27712 19184 27764 19193
rect 31116 19252 31168 19304
rect 31300 19295 31352 19304
rect 31300 19261 31309 19295
rect 31309 19261 31343 19295
rect 31343 19261 31352 19295
rect 31300 19252 31352 19261
rect 31392 19252 31444 19304
rect 31944 19184 31996 19236
rect 32312 19295 32364 19304
rect 32312 19261 32321 19295
rect 32321 19261 32355 19295
rect 32355 19261 32364 19295
rect 36268 19295 36320 19304
rect 32312 19252 32364 19261
rect 36268 19261 36277 19295
rect 36277 19261 36311 19295
rect 36311 19261 36320 19295
rect 36268 19252 36320 19261
rect 39396 19320 39448 19372
rect 39672 19320 39724 19372
rect 36176 19184 36228 19236
rect 36820 19295 36872 19304
rect 36820 19261 36829 19295
rect 36829 19261 36863 19295
rect 36863 19261 36872 19295
rect 36820 19252 36872 19261
rect 37280 19252 37332 19304
rect 38292 19295 38344 19304
rect 38292 19261 38301 19295
rect 38301 19261 38335 19295
rect 38335 19261 38344 19295
rect 38292 19252 38344 19261
rect 38384 19295 38436 19304
rect 38384 19261 38393 19295
rect 38393 19261 38427 19295
rect 38427 19261 38436 19295
rect 38384 19252 38436 19261
rect 39764 19252 39816 19304
rect 41420 19252 41472 19304
rect 42340 19295 42392 19304
rect 41604 19184 41656 19236
rect 20720 19116 20772 19168
rect 24216 19116 24268 19168
rect 32404 19159 32456 19168
rect 32404 19125 32413 19159
rect 32413 19125 32447 19159
rect 32447 19125 32456 19159
rect 32404 19116 32456 19125
rect 32772 19116 32824 19168
rect 37280 19159 37332 19168
rect 37280 19125 37289 19159
rect 37289 19125 37323 19159
rect 37323 19125 37332 19159
rect 37280 19116 37332 19125
rect 37648 19159 37700 19168
rect 37648 19125 37657 19159
rect 37657 19125 37691 19159
rect 37691 19125 37700 19159
rect 37648 19116 37700 19125
rect 38752 19116 38804 19168
rect 39764 19116 39816 19168
rect 41328 19116 41380 19168
rect 42340 19261 42349 19295
rect 42349 19261 42383 19295
rect 42383 19261 42392 19295
rect 42340 19252 42392 19261
rect 42432 19295 42484 19304
rect 42432 19261 42441 19295
rect 42441 19261 42475 19295
rect 42475 19261 42484 19295
rect 46020 19320 46072 19372
rect 48504 19320 48556 19372
rect 42432 19252 42484 19261
rect 44180 19252 44232 19304
rect 44824 19252 44876 19304
rect 46112 19295 46164 19304
rect 46112 19261 46121 19295
rect 46121 19261 46155 19295
rect 46155 19261 46164 19295
rect 46112 19252 46164 19261
rect 47860 19252 47912 19304
rect 48412 19252 48464 19304
rect 48596 19295 48648 19304
rect 48596 19261 48605 19295
rect 48605 19261 48639 19295
rect 48639 19261 48648 19295
rect 48596 19252 48648 19261
rect 49240 19320 49292 19372
rect 44088 19184 44140 19236
rect 46756 19184 46808 19236
rect 47124 19184 47176 19236
rect 49056 19295 49108 19304
rect 49056 19261 49065 19295
rect 49065 19261 49099 19295
rect 49099 19261 49108 19295
rect 49056 19252 49108 19261
rect 50712 19252 50764 19304
rect 52460 19320 52512 19372
rect 49608 19184 49660 19236
rect 52644 19184 52696 19236
rect 42432 19116 42484 19168
rect 42524 19116 42576 19168
rect 46112 19116 46164 19168
rect 46204 19159 46256 19168
rect 46204 19125 46213 19159
rect 46213 19125 46247 19159
rect 46247 19125 46256 19159
rect 46204 19116 46256 19125
rect 46664 19116 46716 19168
rect 49240 19116 49292 19168
rect 53380 19159 53432 19168
rect 53380 19125 53389 19159
rect 53389 19125 53423 19159
rect 53423 19125 53432 19159
rect 53380 19116 53432 19125
rect 18912 19014 18964 19066
rect 18976 19014 19028 19066
rect 19040 19014 19092 19066
rect 19104 19014 19156 19066
rect 36843 19014 36895 19066
rect 36907 19014 36959 19066
rect 36971 19014 37023 19066
rect 37035 19014 37087 19066
rect 2964 18955 3016 18964
rect 2964 18921 2973 18955
rect 2973 18921 3007 18955
rect 3007 18921 3016 18955
rect 2964 18912 3016 18921
rect 10324 18912 10376 18964
rect 16580 18912 16632 18964
rect 17224 18955 17276 18964
rect 17224 18921 17233 18955
rect 17233 18921 17267 18955
rect 17267 18921 17276 18955
rect 17224 18912 17276 18921
rect 5080 18844 5132 18896
rect 3148 18819 3200 18828
rect 3148 18785 3157 18819
rect 3157 18785 3191 18819
rect 3191 18785 3200 18819
rect 3148 18776 3200 18785
rect 4252 18819 4304 18828
rect 4252 18785 4261 18819
rect 4261 18785 4295 18819
rect 4295 18785 4304 18819
rect 4252 18776 4304 18785
rect 6736 18776 6788 18828
rect 9588 18844 9640 18896
rect 8852 18776 8904 18828
rect 10140 18819 10192 18828
rect 10140 18785 10149 18819
rect 10149 18785 10183 18819
rect 10183 18785 10192 18819
rect 10140 18776 10192 18785
rect 13268 18776 13320 18828
rect 13452 18819 13504 18828
rect 13452 18785 13461 18819
rect 13461 18785 13495 18819
rect 13495 18785 13504 18819
rect 13452 18776 13504 18785
rect 13820 18776 13872 18828
rect 15752 18776 15804 18828
rect 18052 18912 18104 18964
rect 25504 18955 25556 18964
rect 25504 18921 25513 18955
rect 25513 18921 25547 18955
rect 25547 18921 25556 18955
rect 25504 18912 25556 18921
rect 29184 18912 29236 18964
rect 29920 18912 29972 18964
rect 24216 18819 24268 18828
rect 11336 18708 11388 18760
rect 6920 18640 6972 18692
rect 7380 18615 7432 18624
rect 7380 18581 7389 18615
rect 7389 18581 7423 18615
rect 7423 18581 7432 18615
rect 7380 18572 7432 18581
rect 9680 18572 9732 18624
rect 12624 18640 12676 18692
rect 15016 18572 15068 18624
rect 20996 18708 21048 18760
rect 24216 18785 24225 18819
rect 24225 18785 24259 18819
rect 24259 18785 24268 18819
rect 24216 18776 24268 18785
rect 25504 18776 25556 18828
rect 28356 18819 28408 18828
rect 28356 18785 28365 18819
rect 28365 18785 28399 18819
rect 28399 18785 28408 18819
rect 28356 18776 28408 18785
rect 25964 18708 26016 18760
rect 29920 18819 29972 18828
rect 29920 18785 29929 18819
rect 29929 18785 29963 18819
rect 29963 18785 29972 18819
rect 29920 18776 29972 18785
rect 30012 18819 30064 18828
rect 30012 18785 30021 18819
rect 30021 18785 30055 18819
rect 30055 18785 30064 18819
rect 32312 18819 32364 18828
rect 30012 18776 30064 18785
rect 32312 18785 32321 18819
rect 32321 18785 32355 18819
rect 32355 18785 32364 18819
rect 32312 18776 32364 18785
rect 32404 18819 32456 18828
rect 32404 18785 32413 18819
rect 32413 18785 32447 18819
rect 32447 18785 32456 18819
rect 33508 18844 33560 18896
rect 33692 18955 33744 18964
rect 33692 18921 33701 18955
rect 33701 18921 33735 18955
rect 33735 18921 33744 18955
rect 36176 18955 36228 18964
rect 33692 18912 33744 18921
rect 36176 18921 36185 18955
rect 36185 18921 36219 18955
rect 36219 18921 36228 18955
rect 36176 18912 36228 18921
rect 36268 18912 36320 18964
rect 37648 18912 37700 18964
rect 41512 18912 41564 18964
rect 41696 18955 41748 18964
rect 41696 18921 41705 18955
rect 41705 18921 41739 18955
rect 41739 18921 41748 18955
rect 41696 18912 41748 18921
rect 48596 18912 48648 18964
rect 32404 18776 32456 18785
rect 36176 18776 36228 18828
rect 36728 18776 36780 18828
rect 33600 18708 33652 18760
rect 33692 18708 33744 18760
rect 34336 18708 34388 18760
rect 38844 18776 38896 18828
rect 39304 18819 39356 18828
rect 39304 18785 39313 18819
rect 39313 18785 39347 18819
rect 39347 18785 39356 18819
rect 39304 18776 39356 18785
rect 39488 18819 39540 18828
rect 39488 18785 39497 18819
rect 39497 18785 39531 18819
rect 39531 18785 39540 18819
rect 39488 18776 39540 18785
rect 39856 18887 39908 18896
rect 39856 18853 39865 18887
rect 39865 18853 39899 18887
rect 39899 18853 39908 18887
rect 39856 18844 39908 18853
rect 40040 18844 40092 18896
rect 49608 18887 49660 18896
rect 41696 18776 41748 18828
rect 44456 18776 44508 18828
rect 49608 18853 49617 18887
rect 49617 18853 49651 18887
rect 49651 18853 49660 18887
rect 49608 18844 49660 18853
rect 44640 18819 44692 18828
rect 44640 18785 44649 18819
rect 44649 18785 44683 18819
rect 44683 18785 44692 18819
rect 47860 18819 47912 18828
rect 44640 18776 44692 18785
rect 47860 18785 47869 18819
rect 47869 18785 47903 18819
rect 47903 18785 47912 18819
rect 47860 18776 47912 18785
rect 48872 18776 48924 18828
rect 49056 18819 49108 18828
rect 49056 18785 49065 18819
rect 49065 18785 49099 18819
rect 49099 18785 49108 18819
rect 49056 18776 49108 18785
rect 49240 18819 49292 18828
rect 49240 18785 49249 18819
rect 49249 18785 49283 18819
rect 49283 18785 49292 18819
rect 49240 18776 49292 18785
rect 49976 18776 50028 18828
rect 51356 18819 51408 18828
rect 18328 18640 18380 18692
rect 21364 18572 21416 18624
rect 25228 18640 25280 18692
rect 36452 18640 36504 18692
rect 26700 18572 26752 18624
rect 27344 18572 27396 18624
rect 29000 18615 29052 18624
rect 29000 18581 29009 18615
rect 29009 18581 29043 18615
rect 29043 18581 29052 18615
rect 29000 18572 29052 18581
rect 29276 18572 29328 18624
rect 33692 18572 33744 18624
rect 33876 18615 33928 18624
rect 33876 18581 33885 18615
rect 33885 18581 33919 18615
rect 33919 18581 33928 18615
rect 33876 18572 33928 18581
rect 37372 18572 37424 18624
rect 38292 18640 38344 18692
rect 44180 18708 44232 18760
rect 46940 18708 46992 18760
rect 51356 18785 51365 18819
rect 51365 18785 51399 18819
rect 51399 18785 51408 18819
rect 51356 18776 51408 18785
rect 52460 18776 52512 18828
rect 53380 18912 53432 18964
rect 53288 18776 53340 18828
rect 38844 18572 38896 18624
rect 39120 18572 39172 18624
rect 39580 18572 39632 18624
rect 44456 18640 44508 18692
rect 45008 18683 45060 18692
rect 45008 18649 45017 18683
rect 45017 18649 45051 18683
rect 45051 18649 45060 18683
rect 45008 18640 45060 18649
rect 45652 18640 45704 18692
rect 40224 18572 40276 18624
rect 41512 18572 41564 18624
rect 47952 18615 48004 18624
rect 47952 18581 47961 18615
rect 47961 18581 47995 18615
rect 47995 18581 48004 18615
rect 47952 18572 48004 18581
rect 52552 18572 52604 18624
rect 9947 18470 9999 18522
rect 10011 18470 10063 18522
rect 10075 18470 10127 18522
rect 10139 18470 10191 18522
rect 27878 18470 27930 18522
rect 27942 18470 27994 18522
rect 28006 18470 28058 18522
rect 28070 18470 28122 18522
rect 45808 18470 45860 18522
rect 45872 18470 45924 18522
rect 45936 18470 45988 18522
rect 46000 18470 46052 18522
rect 6920 18368 6972 18420
rect 8116 18368 8168 18420
rect 4160 18343 4212 18352
rect 4160 18309 4169 18343
rect 4169 18309 4203 18343
rect 4203 18309 4212 18343
rect 4160 18300 4212 18309
rect 10324 18368 10376 18420
rect 13084 18368 13136 18420
rect 17776 18368 17828 18420
rect 7380 18232 7432 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 18052 18300 18104 18352
rect 20996 18343 21048 18352
rect 15016 18275 15068 18284
rect 2872 18164 2924 18216
rect 4344 18207 4396 18216
rect 4344 18173 4353 18207
rect 4353 18173 4387 18207
rect 4387 18173 4396 18207
rect 4344 18164 4396 18173
rect 5080 18207 5132 18216
rect 4252 18096 4304 18148
rect 5080 18173 5089 18207
rect 5089 18173 5123 18207
rect 5123 18173 5132 18207
rect 5080 18164 5132 18173
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 9680 18164 9732 18216
rect 13084 18207 13136 18216
rect 11980 18096 12032 18148
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 13268 18164 13320 18216
rect 6368 18028 6420 18080
rect 14372 18028 14424 18080
rect 15016 18241 15025 18275
rect 15025 18241 15059 18275
rect 15059 18241 15068 18275
rect 15016 18232 15068 18241
rect 18788 18164 18840 18216
rect 20996 18309 21005 18343
rect 21005 18309 21039 18343
rect 21039 18309 21048 18343
rect 23020 18368 23072 18420
rect 29368 18368 29420 18420
rect 20996 18300 21048 18309
rect 31392 18368 31444 18420
rect 32404 18368 32456 18420
rect 32128 18300 32180 18352
rect 34980 18368 35032 18420
rect 32956 18343 33008 18352
rect 32956 18309 32965 18343
rect 32965 18309 32999 18343
rect 32999 18309 33008 18343
rect 32956 18300 33008 18309
rect 21364 18275 21416 18284
rect 21364 18241 21373 18275
rect 21373 18241 21407 18275
rect 21407 18241 21416 18275
rect 21364 18232 21416 18241
rect 25228 18275 25280 18284
rect 25228 18241 25237 18275
rect 25237 18241 25271 18275
rect 25271 18241 25280 18275
rect 25228 18232 25280 18241
rect 25504 18232 25556 18284
rect 29000 18232 29052 18284
rect 29644 18275 29696 18284
rect 29644 18241 29653 18275
rect 29653 18241 29687 18275
rect 29687 18241 29696 18275
rect 29644 18232 29696 18241
rect 16488 18096 16540 18148
rect 19708 18139 19760 18148
rect 19708 18105 19717 18139
rect 19717 18105 19751 18139
rect 19751 18105 19760 18139
rect 19708 18096 19760 18105
rect 23480 18096 23532 18148
rect 23940 18096 23992 18148
rect 22008 18028 22060 18080
rect 23020 18028 23072 18080
rect 25228 18028 25280 18080
rect 25964 18164 26016 18216
rect 31208 18207 31260 18216
rect 26608 18096 26660 18148
rect 26976 18096 27028 18148
rect 28264 18096 28316 18148
rect 28908 18096 28960 18148
rect 29000 18096 29052 18148
rect 27436 18028 27488 18080
rect 28816 18028 28868 18080
rect 31208 18173 31217 18207
rect 31217 18173 31251 18207
rect 31251 18173 31260 18207
rect 31208 18164 31260 18173
rect 31760 18207 31812 18216
rect 31760 18173 31769 18207
rect 31769 18173 31803 18207
rect 31803 18173 31812 18207
rect 31760 18164 31812 18173
rect 32404 18232 32456 18284
rect 33600 18275 33652 18284
rect 33600 18241 33609 18275
rect 33609 18241 33643 18275
rect 33643 18241 33652 18275
rect 33600 18232 33652 18241
rect 32312 18164 32364 18216
rect 34980 18207 35032 18216
rect 34980 18173 34989 18207
rect 34989 18173 35023 18207
rect 35023 18173 35032 18207
rect 34980 18164 35032 18173
rect 35164 18207 35216 18216
rect 35164 18173 35173 18207
rect 35173 18173 35207 18207
rect 35207 18173 35216 18207
rect 35164 18164 35216 18173
rect 35624 18207 35676 18216
rect 35624 18173 35633 18207
rect 35633 18173 35667 18207
rect 35667 18173 35676 18207
rect 35624 18164 35676 18173
rect 35716 18207 35768 18216
rect 35716 18173 35725 18207
rect 35725 18173 35759 18207
rect 35759 18173 35768 18207
rect 37280 18300 37332 18352
rect 39672 18368 39724 18420
rect 39764 18411 39816 18420
rect 39764 18377 39773 18411
rect 39773 18377 39807 18411
rect 39807 18377 39816 18411
rect 39764 18368 39816 18377
rect 39948 18368 40000 18420
rect 41604 18368 41656 18420
rect 45008 18368 45060 18420
rect 47952 18368 48004 18420
rect 39120 18343 39172 18352
rect 39120 18309 39129 18343
rect 39129 18309 39163 18343
rect 39163 18309 39172 18343
rect 39120 18300 39172 18309
rect 39304 18300 39356 18352
rect 39028 18232 39080 18284
rect 40132 18232 40184 18284
rect 35716 18164 35768 18173
rect 38936 18164 38988 18216
rect 39948 18164 40000 18216
rect 40776 18207 40828 18216
rect 40776 18173 40785 18207
rect 40785 18173 40819 18207
rect 40819 18173 40828 18207
rect 40776 18164 40828 18173
rect 42524 18207 42576 18216
rect 38844 18139 38896 18148
rect 33048 18028 33100 18080
rect 35164 18028 35216 18080
rect 38844 18105 38853 18139
rect 38853 18105 38887 18139
rect 38887 18105 38896 18139
rect 38844 18096 38896 18105
rect 42524 18173 42533 18207
rect 42533 18173 42567 18207
rect 42567 18173 42576 18207
rect 42524 18164 42576 18173
rect 42616 18164 42668 18216
rect 52736 18368 52788 18420
rect 44456 18275 44508 18284
rect 44456 18241 44465 18275
rect 44465 18241 44499 18275
rect 44499 18241 44508 18275
rect 46112 18275 46164 18284
rect 44456 18232 44508 18241
rect 46112 18241 46121 18275
rect 46121 18241 46155 18275
rect 46155 18241 46164 18275
rect 46112 18232 46164 18241
rect 49056 18275 49108 18284
rect 44272 18164 44324 18216
rect 44732 18164 44784 18216
rect 46296 18207 46348 18216
rect 42984 18096 43036 18148
rect 45652 18096 45704 18148
rect 46296 18173 46305 18207
rect 46305 18173 46339 18207
rect 46339 18173 46348 18207
rect 46296 18164 46348 18173
rect 48320 18207 48372 18216
rect 48320 18173 48329 18207
rect 48329 18173 48363 18207
rect 48363 18173 48372 18207
rect 48320 18164 48372 18173
rect 48596 18207 48648 18216
rect 48596 18173 48605 18207
rect 48605 18173 48639 18207
rect 48639 18173 48648 18207
rect 48596 18164 48648 18173
rect 49056 18241 49065 18275
rect 49065 18241 49099 18275
rect 49099 18241 49108 18275
rect 49056 18232 49108 18241
rect 49056 18096 49108 18148
rect 36452 18028 36504 18080
rect 40040 18028 40092 18080
rect 41972 18028 42024 18080
rect 47308 18071 47360 18080
rect 47308 18037 47317 18071
rect 47317 18037 47351 18071
rect 47351 18037 47360 18071
rect 47308 18028 47360 18037
rect 51356 18164 51408 18216
rect 52644 18207 52696 18216
rect 52644 18173 52653 18207
rect 52653 18173 52687 18207
rect 52687 18173 52696 18207
rect 52644 18164 52696 18173
rect 49884 18139 49936 18148
rect 49884 18105 49893 18139
rect 49893 18105 49927 18139
rect 49927 18105 49936 18139
rect 49884 18096 49936 18105
rect 51632 18096 51684 18148
rect 52552 18139 52604 18148
rect 52552 18105 52561 18139
rect 52561 18105 52595 18139
rect 52595 18105 52604 18139
rect 52552 18096 52604 18105
rect 49976 18028 50028 18080
rect 18912 17926 18964 17978
rect 18976 17926 19028 17978
rect 19040 17926 19092 17978
rect 19104 17926 19156 17978
rect 36843 17926 36895 17978
rect 36907 17926 36959 17978
rect 36971 17926 37023 17978
rect 37035 17926 37087 17978
rect 4344 17824 4396 17876
rect 11244 17824 11296 17876
rect 11796 17824 11848 17876
rect 2136 17688 2188 17740
rect 8300 17756 8352 17808
rect 12348 17756 12400 17808
rect 6828 17688 6880 17740
rect 8576 17688 8628 17740
rect 10968 17688 11020 17740
rect 11796 17731 11848 17740
rect 11796 17697 11805 17731
rect 11805 17697 11839 17731
rect 11839 17697 11848 17731
rect 11796 17688 11848 17697
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 12624 17824 12676 17876
rect 15936 17824 15988 17876
rect 18052 17824 18104 17876
rect 19248 17867 19300 17876
rect 19248 17833 19257 17867
rect 19257 17833 19291 17867
rect 19291 17833 19300 17867
rect 19248 17824 19300 17833
rect 19340 17824 19392 17876
rect 13820 17756 13872 17808
rect 6736 17484 6788 17536
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 10692 17527 10744 17536
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 12992 17527 13044 17536
rect 12992 17493 13001 17527
rect 13001 17493 13035 17527
rect 13035 17493 13044 17527
rect 12992 17484 13044 17493
rect 16488 17688 16540 17740
rect 17224 17688 17276 17740
rect 18236 17731 18288 17740
rect 18236 17697 18245 17731
rect 18245 17697 18279 17731
rect 18279 17697 18288 17731
rect 18236 17688 18288 17697
rect 19708 17688 19760 17740
rect 21088 17731 21140 17740
rect 21088 17697 21097 17731
rect 21097 17697 21131 17731
rect 21131 17697 21140 17731
rect 21088 17688 21140 17697
rect 22008 17731 22060 17740
rect 22008 17697 22017 17731
rect 22017 17697 22051 17731
rect 22051 17697 22060 17731
rect 22008 17688 22060 17697
rect 22376 17688 22428 17740
rect 29276 17824 29328 17876
rect 30012 17824 30064 17876
rect 25780 17799 25832 17808
rect 25780 17765 25789 17799
rect 25789 17765 25823 17799
rect 25823 17765 25832 17799
rect 25780 17756 25832 17765
rect 29644 17756 29696 17808
rect 23020 17731 23072 17740
rect 23020 17697 23029 17731
rect 23029 17697 23063 17731
rect 23063 17697 23072 17731
rect 23020 17688 23072 17697
rect 28724 17731 28776 17740
rect 28724 17697 28733 17731
rect 28733 17697 28767 17731
rect 28767 17697 28776 17731
rect 28724 17688 28776 17697
rect 29460 17731 29512 17740
rect 24952 17620 25004 17672
rect 25228 17663 25280 17672
rect 25228 17629 25237 17663
rect 25237 17629 25271 17663
rect 25271 17629 25280 17663
rect 25228 17620 25280 17629
rect 29460 17697 29469 17731
rect 29469 17697 29503 17731
rect 29503 17697 29512 17731
rect 29460 17688 29512 17697
rect 31208 17756 31260 17808
rect 32312 17731 32364 17740
rect 32312 17697 32321 17731
rect 32321 17697 32355 17731
rect 32355 17697 32364 17731
rect 32772 17731 32824 17740
rect 32312 17688 32364 17697
rect 32772 17697 32781 17731
rect 32781 17697 32815 17731
rect 32815 17697 32824 17731
rect 32772 17688 32824 17697
rect 34612 17688 34664 17740
rect 35716 17688 35768 17740
rect 36636 17756 36688 17808
rect 37188 17756 37240 17808
rect 30380 17620 30432 17672
rect 33508 17620 33560 17672
rect 36360 17688 36412 17740
rect 37372 17688 37424 17740
rect 14740 17484 14792 17536
rect 17132 17527 17184 17536
rect 17132 17493 17141 17527
rect 17141 17493 17175 17527
rect 17175 17493 17184 17527
rect 17132 17484 17184 17493
rect 18052 17527 18104 17536
rect 18052 17493 18061 17527
rect 18061 17493 18095 17527
rect 18095 17493 18104 17527
rect 18052 17484 18104 17493
rect 23296 17527 23348 17536
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23296 17484 23348 17493
rect 25412 17552 25464 17604
rect 29000 17552 29052 17604
rect 35900 17595 35952 17604
rect 35900 17561 35909 17595
rect 35909 17561 35943 17595
rect 35943 17561 35952 17595
rect 35900 17552 35952 17561
rect 28632 17484 28684 17536
rect 28908 17484 28960 17536
rect 29736 17484 29788 17536
rect 33324 17527 33376 17536
rect 33324 17493 33333 17527
rect 33333 17493 33367 17527
rect 33367 17493 33376 17527
rect 33324 17484 33376 17493
rect 37924 17824 37976 17876
rect 38108 17688 38160 17740
rect 38384 17731 38436 17740
rect 38384 17697 38393 17731
rect 38393 17697 38427 17731
rect 38427 17697 38436 17731
rect 38384 17688 38436 17697
rect 38660 17756 38712 17808
rect 38844 17824 38896 17876
rect 39028 17824 39080 17876
rect 44180 17824 44232 17876
rect 44548 17824 44600 17876
rect 38568 17688 38620 17740
rect 39948 17552 40000 17604
rect 39304 17484 39356 17536
rect 40776 17688 40828 17740
rect 40868 17731 40920 17740
rect 40868 17697 40877 17731
rect 40877 17697 40911 17731
rect 40911 17697 40920 17731
rect 40868 17688 40920 17697
rect 41328 17688 41380 17740
rect 45560 17756 45612 17808
rect 46296 17756 46348 17808
rect 45652 17688 45704 17740
rect 48596 17824 48648 17876
rect 52460 17824 52512 17876
rect 40776 17552 40828 17604
rect 44088 17663 44140 17672
rect 44088 17629 44097 17663
rect 44097 17629 44131 17663
rect 44131 17629 44140 17663
rect 44088 17620 44140 17629
rect 48320 17688 48372 17740
rect 49884 17756 49936 17808
rect 50804 17688 50856 17740
rect 51632 17731 51684 17740
rect 51632 17697 51641 17731
rect 51641 17697 51675 17731
rect 51675 17697 51684 17731
rect 51632 17688 51684 17697
rect 53288 17688 53340 17740
rect 47124 17663 47176 17672
rect 47124 17629 47133 17663
rect 47133 17629 47167 17663
rect 47167 17629 47176 17663
rect 51356 17663 51408 17672
rect 47124 17620 47176 17629
rect 51356 17629 51365 17663
rect 51365 17629 51399 17663
rect 51399 17629 51408 17663
rect 51356 17620 51408 17629
rect 52368 17620 52420 17672
rect 50252 17552 50304 17604
rect 43996 17484 44048 17536
rect 45192 17484 45244 17536
rect 46480 17527 46532 17536
rect 46480 17493 46489 17527
rect 46489 17493 46523 17527
rect 46523 17493 46532 17527
rect 46480 17484 46532 17493
rect 9947 17382 9999 17434
rect 10011 17382 10063 17434
rect 10075 17382 10127 17434
rect 10139 17382 10191 17434
rect 27878 17382 27930 17434
rect 27942 17382 27994 17434
rect 28006 17382 28058 17434
rect 28070 17382 28122 17434
rect 45808 17382 45860 17434
rect 45872 17382 45924 17434
rect 45936 17382 45988 17434
rect 46000 17382 46052 17434
rect 2136 17323 2188 17332
rect 2136 17289 2145 17323
rect 2145 17289 2179 17323
rect 2179 17289 2188 17323
rect 2136 17280 2188 17289
rect 5264 17280 5316 17332
rect 8024 17212 8076 17264
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 2596 17076 2648 17128
rect 9588 17144 9640 17196
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 7564 17119 7616 17128
rect 4068 17008 4120 17060
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 8024 17076 8076 17128
rect 8300 17119 8352 17128
rect 8300 17085 8309 17119
rect 8309 17085 8343 17119
rect 8343 17085 8352 17119
rect 8300 17076 8352 17085
rect 9680 17076 9732 17128
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 10692 17076 10744 17128
rect 16028 17280 16080 17332
rect 16580 17280 16632 17332
rect 24952 17280 25004 17332
rect 14280 17255 14332 17264
rect 14280 17221 14289 17255
rect 14289 17221 14323 17255
rect 14323 17221 14332 17255
rect 14280 17212 14332 17221
rect 18696 17212 18748 17264
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 16488 17144 16540 17196
rect 8576 17008 8628 17060
rect 14372 17076 14424 17128
rect 15108 17076 15160 17128
rect 15292 17119 15344 17128
rect 15292 17085 15301 17119
rect 15301 17085 15335 17119
rect 15335 17085 15344 17119
rect 15292 17076 15344 17085
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 17132 17076 17184 17128
rect 19800 17212 19852 17264
rect 28356 17280 28408 17332
rect 28448 17280 28500 17332
rect 29828 17280 29880 17332
rect 29920 17280 29972 17332
rect 31944 17280 31996 17332
rect 33324 17280 33376 17332
rect 39028 17280 39080 17332
rect 19248 17008 19300 17060
rect 19616 17119 19668 17128
rect 19616 17085 19625 17119
rect 19625 17085 19659 17119
rect 19659 17085 19668 17119
rect 19616 17076 19668 17085
rect 22376 17076 22428 17128
rect 23296 17076 23348 17128
rect 25320 17076 25372 17128
rect 26240 17076 26292 17128
rect 36084 17212 36136 17264
rect 41696 17280 41748 17332
rect 42248 17280 42300 17332
rect 44088 17323 44140 17332
rect 44088 17289 44097 17323
rect 44097 17289 44131 17323
rect 44131 17289 44140 17323
rect 44088 17280 44140 17289
rect 44548 17280 44600 17332
rect 45192 17280 45244 17332
rect 39212 17212 39264 17264
rect 39948 17212 40000 17264
rect 43996 17212 44048 17264
rect 29276 17144 29328 17196
rect 29460 17187 29512 17196
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 28448 17076 28500 17128
rect 28540 17076 28592 17128
rect 30012 17144 30064 17196
rect 30380 17187 30432 17196
rect 30380 17153 30389 17187
rect 30389 17153 30423 17187
rect 30423 17153 30432 17187
rect 30380 17144 30432 17153
rect 34520 17144 34572 17196
rect 38016 17144 38068 17196
rect 39304 17144 39356 17196
rect 41604 17187 41656 17196
rect 29644 17076 29696 17128
rect 29920 17119 29972 17128
rect 29920 17085 29929 17119
rect 29929 17085 29963 17119
rect 29963 17085 29972 17119
rect 29920 17076 29972 17085
rect 27160 17008 27212 17060
rect 27620 17051 27672 17060
rect 27620 17017 27629 17051
rect 27629 17017 27663 17051
rect 27663 17017 27672 17051
rect 27620 17008 27672 17017
rect 29000 17008 29052 17060
rect 5632 16940 5684 16992
rect 11244 16940 11296 16992
rect 14372 16940 14424 16992
rect 15108 16983 15160 16992
rect 15108 16949 15117 16983
rect 15117 16949 15151 16983
rect 15151 16949 15160 16983
rect 15108 16940 15160 16949
rect 16488 16983 16540 16992
rect 16488 16949 16497 16983
rect 16497 16949 16531 16983
rect 16531 16949 16540 16983
rect 16488 16940 16540 16949
rect 21088 16940 21140 16992
rect 21272 16940 21324 16992
rect 24584 16940 24636 16992
rect 28264 16940 28316 16992
rect 31116 17076 31168 17128
rect 33600 17076 33652 17128
rect 35624 17119 35676 17128
rect 32220 17008 32272 17060
rect 33232 17008 33284 17060
rect 35624 17085 35633 17119
rect 35633 17085 35667 17119
rect 35667 17085 35676 17119
rect 35624 17076 35676 17085
rect 35900 17008 35952 17060
rect 36084 17076 36136 17128
rect 36452 17076 36504 17128
rect 37832 17119 37884 17128
rect 37832 17085 37841 17119
rect 37841 17085 37875 17119
rect 37875 17085 37884 17119
rect 37832 17076 37884 17085
rect 37188 17008 37240 17060
rect 39488 17076 39540 17128
rect 41604 17153 41613 17187
rect 41613 17153 41647 17187
rect 41647 17153 41656 17187
rect 41604 17144 41656 17153
rect 42248 17119 42300 17128
rect 38752 17008 38804 17060
rect 39672 17008 39724 17060
rect 35624 16940 35676 16992
rect 38108 16940 38160 16992
rect 39764 16940 39816 16992
rect 42248 17085 42257 17119
rect 42257 17085 42291 17119
rect 42291 17085 42300 17119
rect 42248 17076 42300 17085
rect 42708 17076 42760 17128
rect 46480 17144 46532 17196
rect 50896 17280 50948 17332
rect 48872 17212 48924 17264
rect 50436 17212 50488 17264
rect 50804 17187 50856 17196
rect 50804 17153 50813 17187
rect 50813 17153 50847 17187
rect 50847 17153 50856 17187
rect 50804 17144 50856 17153
rect 50988 17144 51040 17196
rect 51080 17144 51132 17196
rect 52368 17187 52420 17196
rect 45560 17076 45612 17128
rect 47492 17076 47544 17128
rect 50252 17119 50304 17128
rect 50252 17085 50261 17119
rect 50261 17085 50295 17119
rect 50295 17085 50304 17119
rect 50252 17076 50304 17085
rect 50436 17119 50488 17128
rect 50436 17085 50459 17119
rect 50459 17085 50488 17119
rect 50436 17076 50488 17085
rect 42984 17008 43036 17060
rect 44180 16940 44232 16992
rect 47952 17008 48004 17060
rect 51356 17008 51408 17060
rect 48504 16983 48556 16992
rect 48504 16949 48513 16983
rect 48513 16949 48547 16983
rect 48547 16949 48556 16983
rect 48504 16940 48556 16949
rect 51264 16940 51316 16992
rect 52368 17153 52377 17187
rect 52377 17153 52411 17187
rect 52411 17153 52420 17187
rect 52368 17144 52420 17153
rect 18912 16838 18964 16890
rect 18976 16838 19028 16890
rect 19040 16838 19092 16890
rect 19104 16838 19156 16890
rect 36843 16838 36895 16890
rect 36907 16838 36959 16890
rect 36971 16838 37023 16890
rect 37035 16838 37087 16890
rect 2596 16779 2648 16788
rect 2596 16745 2605 16779
rect 2605 16745 2639 16779
rect 2639 16745 2648 16779
rect 2596 16736 2648 16745
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 3792 16643 3844 16652
rect 2780 16600 2832 16609
rect 3792 16609 3801 16643
rect 3801 16609 3835 16643
rect 3835 16609 3844 16643
rect 3792 16600 3844 16609
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 6368 16643 6420 16652
rect 6368 16609 6377 16643
rect 6377 16609 6411 16643
rect 6411 16609 6420 16643
rect 6368 16600 6420 16609
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 7564 16600 7616 16652
rect 11428 16736 11480 16788
rect 12348 16736 12400 16788
rect 10692 16668 10744 16720
rect 10416 16600 10468 16652
rect 13176 16600 13228 16652
rect 14280 16600 14332 16652
rect 14924 16600 14976 16652
rect 16488 16643 16540 16652
rect 16488 16609 16497 16643
rect 16497 16609 16531 16643
rect 16531 16609 16540 16643
rect 16488 16600 16540 16609
rect 17224 16736 17276 16788
rect 21272 16736 21324 16788
rect 17868 16668 17920 16720
rect 18052 16600 18104 16652
rect 19340 16643 19392 16652
rect 19340 16609 19349 16643
rect 19349 16609 19383 16643
rect 19383 16609 19392 16643
rect 19340 16600 19392 16609
rect 22560 16600 22612 16652
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 23388 16600 23440 16652
rect 24400 16643 24452 16652
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 28540 16736 28592 16788
rect 28632 16736 28684 16788
rect 24676 16668 24728 16720
rect 24584 16600 24636 16652
rect 26516 16643 26568 16652
rect 26516 16609 26525 16643
rect 26525 16609 26559 16643
rect 26559 16609 26568 16643
rect 29000 16668 29052 16720
rect 26516 16600 26568 16609
rect 12348 16532 12400 16584
rect 15108 16532 15160 16584
rect 11704 16464 11756 16516
rect 18512 16464 18564 16516
rect 18788 16464 18840 16516
rect 25320 16507 25372 16516
rect 25320 16473 25329 16507
rect 25329 16473 25363 16507
rect 25363 16473 25372 16507
rect 25320 16464 25372 16473
rect 3148 16396 3200 16448
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 6920 16396 6972 16448
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 26240 16464 26292 16516
rect 27160 16643 27212 16652
rect 27160 16609 27169 16643
rect 27169 16609 27203 16643
rect 27203 16609 27212 16643
rect 27160 16600 27212 16609
rect 27712 16600 27764 16652
rect 28908 16600 28960 16652
rect 33600 16779 33652 16788
rect 33600 16745 33609 16779
rect 33609 16745 33643 16779
rect 33643 16745 33652 16779
rect 33600 16736 33652 16745
rect 29460 16600 29512 16652
rect 29552 16600 29604 16652
rect 29736 16600 29788 16652
rect 30472 16643 30524 16652
rect 30472 16609 30481 16643
rect 30481 16609 30515 16643
rect 30515 16609 30524 16643
rect 30472 16600 30524 16609
rect 32956 16600 33008 16652
rect 35808 16600 35860 16652
rect 32864 16532 32916 16584
rect 35900 16532 35952 16584
rect 37188 16736 37240 16788
rect 42340 16736 42392 16788
rect 47492 16779 47544 16788
rect 47492 16745 47501 16779
rect 47501 16745 47535 16779
rect 47535 16745 47544 16779
rect 47492 16736 47544 16745
rect 39948 16711 40000 16720
rect 39948 16677 39957 16711
rect 39957 16677 39991 16711
rect 39991 16677 40000 16711
rect 39948 16668 40000 16677
rect 40500 16668 40552 16720
rect 40776 16643 40828 16652
rect 38384 16575 38436 16584
rect 29276 16464 29328 16516
rect 36360 16464 36412 16516
rect 25964 16439 26016 16448
rect 25964 16405 25973 16439
rect 25973 16405 26007 16439
rect 26007 16405 26016 16439
rect 25964 16396 26016 16405
rect 26884 16396 26936 16448
rect 27068 16396 27120 16448
rect 35808 16396 35860 16448
rect 36452 16396 36504 16448
rect 38384 16541 38393 16575
rect 38393 16541 38427 16575
rect 38427 16541 38436 16575
rect 38384 16532 38436 16541
rect 38752 16532 38804 16584
rect 39120 16532 39172 16584
rect 39672 16532 39724 16584
rect 40500 16532 40552 16584
rect 40776 16609 40782 16643
rect 40782 16609 40828 16643
rect 40776 16600 40828 16609
rect 47308 16668 47360 16720
rect 49056 16668 49108 16720
rect 41052 16600 41104 16652
rect 41788 16600 41840 16652
rect 42064 16532 42116 16584
rect 44640 16600 44692 16652
rect 45468 16600 45520 16652
rect 47400 16643 47452 16652
rect 47400 16609 47409 16643
rect 47409 16609 47443 16643
rect 47443 16609 47452 16643
rect 47400 16600 47452 16609
rect 48504 16600 48556 16652
rect 50160 16600 50212 16652
rect 51448 16600 51500 16652
rect 51724 16600 51776 16652
rect 52368 16575 52420 16584
rect 52368 16541 52377 16575
rect 52377 16541 52411 16575
rect 52411 16541 52420 16575
rect 52368 16532 52420 16541
rect 42892 16464 42944 16516
rect 50896 16464 50948 16516
rect 51264 16464 51316 16516
rect 51356 16464 51408 16516
rect 53472 16507 53524 16516
rect 53472 16473 53481 16507
rect 53481 16473 53515 16507
rect 53515 16473 53524 16507
rect 53472 16464 53524 16473
rect 39948 16396 40000 16448
rect 40316 16396 40368 16448
rect 42708 16396 42760 16448
rect 48596 16396 48648 16448
rect 9947 16294 9999 16346
rect 10011 16294 10063 16346
rect 10075 16294 10127 16346
rect 10139 16294 10191 16346
rect 27878 16294 27930 16346
rect 27942 16294 27994 16346
rect 28006 16294 28058 16346
rect 28070 16294 28122 16346
rect 45808 16294 45860 16346
rect 45872 16294 45924 16346
rect 45936 16294 45988 16346
rect 46000 16294 46052 16346
rect 4160 16192 4212 16244
rect 6552 16192 6604 16244
rect 8760 16192 8812 16244
rect 11980 16192 12032 16244
rect 13912 16192 13964 16244
rect 15292 16192 15344 16244
rect 6736 16124 6788 16176
rect 6828 16056 6880 16108
rect 2872 15988 2924 16040
rect 3884 15988 3936 16040
rect 6920 15988 6972 16040
rect 8024 16124 8076 16176
rect 9036 16031 9088 16040
rect 9036 15997 9045 16031
rect 9045 15997 9079 16031
rect 9079 15997 9088 16031
rect 9036 15988 9088 15997
rect 13176 16056 13228 16108
rect 19432 16124 19484 16176
rect 3976 15963 4028 15972
rect 3976 15929 3985 15963
rect 3985 15929 4019 15963
rect 4019 15929 4028 15963
rect 3976 15920 4028 15929
rect 8576 15920 8628 15972
rect 13544 16031 13596 16040
rect 4988 15852 5040 15904
rect 7564 15852 7616 15904
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 10508 15852 10560 15904
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 14372 15852 14424 15904
rect 14924 15852 14976 15904
rect 15476 15852 15528 15904
rect 16580 15988 16632 16040
rect 19524 16056 19576 16108
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 17040 15963 17092 15972
rect 17040 15929 17049 15963
rect 17049 15929 17083 15963
rect 17083 15929 17092 15963
rect 17040 15920 17092 15929
rect 18696 15920 18748 15972
rect 19708 15988 19760 16040
rect 19892 16031 19944 16040
rect 19892 15997 19901 16031
rect 19901 15997 19935 16031
rect 19935 15997 19944 16031
rect 21548 16031 21600 16040
rect 19892 15988 19944 15997
rect 21548 15997 21557 16031
rect 21557 15997 21591 16031
rect 21591 15997 21600 16031
rect 21548 15988 21600 15997
rect 21640 15988 21692 16040
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 24676 16031 24728 16040
rect 22100 15988 22152 15997
rect 24676 15997 24685 16031
rect 24685 15997 24719 16031
rect 24719 15997 24728 16031
rect 24676 15988 24728 15997
rect 27344 16235 27396 16244
rect 27344 16201 27353 16235
rect 27353 16201 27387 16235
rect 27387 16201 27396 16235
rect 27344 16192 27396 16201
rect 28908 16192 28960 16244
rect 32864 16235 32916 16244
rect 32864 16201 32873 16235
rect 32873 16201 32907 16235
rect 32907 16201 32916 16235
rect 32864 16192 32916 16201
rect 35900 16235 35952 16244
rect 35900 16201 35909 16235
rect 35909 16201 35943 16235
rect 35943 16201 35952 16235
rect 35900 16192 35952 16201
rect 39396 16192 39448 16244
rect 47400 16192 47452 16244
rect 53472 16235 53524 16244
rect 53472 16201 53481 16235
rect 53481 16201 53515 16235
rect 53515 16201 53524 16235
rect 53472 16192 53524 16201
rect 27068 16099 27120 16108
rect 27068 16065 27077 16099
rect 27077 16065 27111 16099
rect 27111 16065 27120 16099
rect 27068 16056 27120 16065
rect 26240 15988 26292 16040
rect 26424 15988 26476 16040
rect 29552 15988 29604 16040
rect 31116 15988 31168 16040
rect 41788 16056 41840 16108
rect 42708 16056 42760 16108
rect 47032 16056 47084 16108
rect 48136 16099 48188 16108
rect 48136 16065 48145 16099
rect 48145 16065 48179 16099
rect 48179 16065 48188 16099
rect 48136 16056 48188 16065
rect 35532 16031 35584 16040
rect 35532 15997 35541 16031
rect 35541 15997 35575 16031
rect 35575 15997 35584 16031
rect 35532 15988 35584 15997
rect 35808 15988 35860 16040
rect 39120 16031 39172 16040
rect 39120 15997 39129 16031
rect 39129 15997 39163 16031
rect 39163 15997 39172 16031
rect 39120 15988 39172 15997
rect 42064 16031 42116 16040
rect 42064 15997 42073 16031
rect 42073 15997 42107 16031
rect 42107 15997 42116 16031
rect 42064 15988 42116 15997
rect 42800 15988 42852 16040
rect 43536 16031 43588 16040
rect 43536 15997 43545 16031
rect 43545 15997 43579 16031
rect 43579 15997 43588 16031
rect 43536 15988 43588 15997
rect 50620 16124 50672 16176
rect 52368 16099 52420 16108
rect 48596 16031 48648 16040
rect 48596 15997 48605 16031
rect 48605 15997 48639 16031
rect 48639 15997 48648 16031
rect 48596 15988 48648 15997
rect 52368 16065 52377 16099
rect 52377 16065 52411 16099
rect 52411 16065 52420 16099
rect 52368 16056 52420 16065
rect 16764 15852 16816 15904
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 18788 15895 18840 15904
rect 18788 15861 18797 15895
rect 18797 15861 18831 15895
rect 18831 15861 18840 15895
rect 18788 15852 18840 15861
rect 30748 15920 30800 15972
rect 33968 15920 34020 15972
rect 35624 15963 35676 15972
rect 35624 15929 35633 15963
rect 35633 15929 35667 15963
rect 35667 15929 35676 15963
rect 35624 15920 35676 15929
rect 41880 15963 41932 15972
rect 41880 15929 41889 15963
rect 41889 15929 41923 15963
rect 41923 15929 41932 15963
rect 41880 15920 41932 15929
rect 51264 15988 51316 16040
rect 48964 15920 49016 15972
rect 50160 15963 50212 15972
rect 50160 15929 50169 15963
rect 50169 15929 50203 15963
rect 50203 15929 50212 15963
rect 50160 15920 50212 15929
rect 21640 15852 21692 15904
rect 29736 15852 29788 15904
rect 42156 15895 42208 15904
rect 42156 15861 42165 15895
rect 42165 15861 42199 15895
rect 42199 15861 42208 15895
rect 42156 15852 42208 15861
rect 51816 15852 51868 15904
rect 18912 15750 18964 15802
rect 18976 15750 19028 15802
rect 19040 15750 19092 15802
rect 19104 15750 19156 15802
rect 36843 15750 36895 15802
rect 36907 15750 36959 15802
rect 36971 15750 37023 15802
rect 37035 15750 37087 15802
rect 2780 15648 2832 15700
rect 3792 15648 3844 15700
rect 7656 15691 7708 15700
rect 2504 15580 2556 15632
rect 3148 15512 3200 15564
rect 4988 15555 5040 15564
rect 4988 15521 4997 15555
rect 4997 15521 5031 15555
rect 5031 15521 5040 15555
rect 4988 15512 5040 15521
rect 6368 15580 6420 15632
rect 7656 15657 7665 15691
rect 7665 15657 7699 15691
rect 7699 15657 7708 15691
rect 7656 15648 7708 15657
rect 10416 15648 10468 15700
rect 14188 15648 14240 15700
rect 18512 15691 18564 15700
rect 8024 15580 8076 15632
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 9956 15580 10008 15632
rect 6276 15512 6328 15521
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 10324 15512 10376 15564
rect 10600 15555 10652 15564
rect 10600 15521 10609 15555
rect 10609 15521 10643 15555
rect 10643 15521 10652 15555
rect 10600 15512 10652 15521
rect 11520 15512 11572 15564
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 13544 15580 13596 15632
rect 14280 15555 14332 15564
rect 11244 15444 11296 15496
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 19892 15648 19944 15700
rect 29000 15648 29052 15700
rect 33968 15691 34020 15700
rect 20812 15580 20864 15632
rect 33968 15657 33977 15691
rect 33977 15657 34011 15691
rect 34011 15657 34020 15691
rect 33968 15648 34020 15657
rect 43996 15691 44048 15700
rect 43996 15657 44005 15691
rect 44005 15657 44039 15691
rect 44039 15657 44048 15691
rect 43996 15648 44048 15657
rect 45468 15691 45520 15700
rect 45468 15657 45477 15691
rect 45477 15657 45511 15691
rect 45511 15657 45520 15691
rect 45468 15648 45520 15657
rect 17040 15555 17092 15564
rect 17040 15521 17049 15555
rect 17049 15521 17083 15555
rect 17083 15521 17092 15555
rect 17040 15512 17092 15521
rect 19616 15512 19668 15564
rect 23940 15512 23992 15564
rect 31944 15580 31996 15632
rect 32496 15555 32548 15564
rect 32496 15521 32505 15555
rect 32505 15521 32539 15555
rect 32539 15521 32548 15555
rect 32496 15512 32548 15521
rect 32680 15512 32732 15564
rect 38384 15580 38436 15632
rect 34980 15512 35032 15564
rect 35808 15555 35860 15564
rect 35808 15521 35817 15555
rect 35817 15521 35851 15555
rect 35851 15521 35860 15555
rect 35808 15512 35860 15521
rect 36636 15512 36688 15564
rect 39028 15555 39080 15564
rect 39028 15521 39037 15555
rect 39037 15521 39071 15555
rect 39071 15521 39080 15555
rect 39028 15512 39080 15521
rect 39396 15512 39448 15564
rect 40408 15512 40460 15564
rect 41788 15580 41840 15632
rect 42156 15580 42208 15632
rect 48596 15580 48648 15632
rect 51724 15623 51776 15632
rect 46756 15555 46808 15564
rect 46756 15521 46765 15555
rect 46765 15521 46799 15555
rect 46799 15521 46808 15555
rect 46756 15512 46808 15521
rect 46940 15555 46992 15564
rect 46940 15521 46949 15555
rect 46949 15521 46983 15555
rect 46983 15521 46992 15555
rect 46940 15512 46992 15521
rect 47216 15512 47268 15564
rect 48964 15555 49016 15564
rect 48964 15521 48973 15555
rect 48973 15521 49007 15555
rect 49007 15521 49016 15555
rect 48964 15512 49016 15521
rect 49056 15555 49108 15564
rect 49056 15521 49065 15555
rect 49065 15521 49099 15555
rect 49099 15521 49108 15555
rect 51724 15589 51733 15623
rect 51733 15589 51767 15623
rect 51767 15589 51776 15623
rect 51724 15580 51776 15589
rect 49056 15512 49108 15521
rect 50620 15512 50672 15564
rect 51356 15555 51408 15564
rect 51356 15521 51365 15555
rect 51365 15521 51399 15555
rect 51399 15521 51408 15555
rect 51356 15512 51408 15521
rect 6460 15419 6512 15428
rect 6460 15385 6469 15419
rect 6469 15385 6503 15419
rect 6503 15385 6512 15419
rect 6460 15376 6512 15385
rect 12440 15376 12492 15428
rect 9772 15308 9824 15360
rect 10416 15351 10468 15360
rect 10416 15317 10425 15351
rect 10425 15317 10459 15351
rect 10459 15317 10468 15351
rect 10416 15308 10468 15317
rect 19340 15444 19392 15496
rect 21732 15444 21784 15496
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 27620 15444 27672 15496
rect 29368 15444 29420 15496
rect 19708 15308 19760 15360
rect 21732 15351 21784 15360
rect 21732 15317 21741 15351
rect 21741 15317 21775 15351
rect 21775 15317 21784 15351
rect 21732 15308 21784 15317
rect 24768 15376 24820 15428
rect 23388 15308 23440 15360
rect 23940 15308 23992 15360
rect 31208 15444 31260 15496
rect 34428 15444 34480 15496
rect 38752 15487 38804 15496
rect 38752 15453 38761 15487
rect 38761 15453 38795 15487
rect 38795 15453 38804 15487
rect 38752 15444 38804 15453
rect 43996 15444 44048 15496
rect 49608 15487 49660 15496
rect 49608 15453 49617 15487
rect 49617 15453 49651 15487
rect 49651 15453 49660 15487
rect 49608 15444 49660 15453
rect 29736 15376 29788 15428
rect 40316 15376 40368 15428
rect 30104 15308 30156 15360
rect 31116 15308 31168 15360
rect 41696 15351 41748 15360
rect 41696 15317 41705 15351
rect 41705 15317 41739 15351
rect 41739 15317 41748 15351
rect 41696 15308 41748 15317
rect 47032 15351 47084 15360
rect 47032 15317 47041 15351
rect 47041 15317 47075 15351
rect 47075 15317 47084 15351
rect 47032 15308 47084 15317
rect 9947 15206 9999 15258
rect 10011 15206 10063 15258
rect 10075 15206 10127 15258
rect 10139 15206 10191 15258
rect 27878 15206 27930 15258
rect 27942 15206 27994 15258
rect 28006 15206 28058 15258
rect 28070 15206 28122 15258
rect 45808 15206 45860 15258
rect 45872 15206 45924 15258
rect 45936 15206 45988 15258
rect 46000 15206 46052 15258
rect 2228 14900 2280 14952
rect 4068 14968 4120 15020
rect 6368 14968 6420 15020
rect 3884 14943 3936 14952
rect 3884 14909 3893 14943
rect 3893 14909 3927 14943
rect 3927 14909 3936 14943
rect 3884 14900 3936 14909
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 6552 14900 6604 14952
rect 11244 15104 11296 15156
rect 12348 15036 12400 15088
rect 12624 15036 12676 15088
rect 13176 15036 13228 15088
rect 14280 15104 14332 15156
rect 20812 15104 20864 15156
rect 24032 15104 24084 15156
rect 27528 15104 27580 15156
rect 32588 15104 32640 15156
rect 17960 15036 18012 15088
rect 18512 15036 18564 15088
rect 20720 15036 20772 15088
rect 21732 15036 21784 15088
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 13636 15011 13688 15020
rect 13636 14977 13645 15011
rect 13645 14977 13679 15011
rect 13679 14977 13688 15011
rect 13636 14968 13688 14977
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 9680 14943 9732 14952
rect 8300 14832 8352 14884
rect 9036 14832 9088 14884
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 11152 14900 11204 14952
rect 12348 14900 12400 14952
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 13084 14943 13136 14952
rect 13084 14909 13093 14943
rect 13093 14909 13127 14943
rect 13127 14909 13136 14943
rect 13084 14900 13136 14909
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 10324 14875 10376 14884
rect 10324 14841 10333 14875
rect 10333 14841 10367 14875
rect 10367 14841 10376 14875
rect 10324 14832 10376 14841
rect 12808 14832 12860 14884
rect 18236 14968 18288 15020
rect 19340 14968 19392 15020
rect 25872 15036 25924 15088
rect 33232 15036 33284 15088
rect 15844 14943 15896 14952
rect 15844 14909 15853 14943
rect 15853 14909 15887 14943
rect 15887 14909 15896 14943
rect 15844 14900 15896 14909
rect 18788 14900 18840 14952
rect 16488 14832 16540 14884
rect 18328 14832 18380 14884
rect 19892 14900 19944 14952
rect 20812 14900 20864 14952
rect 22008 14832 22060 14884
rect 23388 14900 23440 14952
rect 27436 14968 27488 15020
rect 28908 14968 28960 15020
rect 3424 14764 3476 14816
rect 7196 14764 7248 14816
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 16672 14807 16724 14816
rect 16672 14773 16681 14807
rect 16681 14773 16715 14807
rect 16715 14773 16724 14807
rect 16672 14764 16724 14773
rect 18512 14764 18564 14816
rect 19432 14764 19484 14816
rect 22928 14807 22980 14816
rect 22928 14773 22937 14807
rect 22937 14773 22971 14807
rect 22971 14773 22980 14807
rect 22928 14764 22980 14773
rect 24400 14807 24452 14816
rect 24400 14773 24409 14807
rect 24409 14773 24443 14807
rect 24443 14773 24452 14807
rect 24400 14764 24452 14773
rect 24952 14900 25004 14952
rect 25136 14943 25188 14952
rect 25136 14909 25145 14943
rect 25145 14909 25179 14943
rect 25179 14909 25188 14943
rect 25136 14900 25188 14909
rect 26608 14900 26660 14952
rect 27528 14943 27580 14952
rect 27528 14909 27537 14943
rect 27537 14909 27571 14943
rect 27571 14909 27580 14943
rect 27528 14900 27580 14909
rect 30748 14943 30800 14952
rect 30748 14909 30757 14943
rect 30757 14909 30791 14943
rect 30791 14909 30800 14943
rect 30748 14900 30800 14909
rect 31116 14943 31168 14952
rect 26516 14764 26568 14816
rect 29276 14832 29328 14884
rect 31116 14909 31125 14943
rect 31125 14909 31159 14943
rect 31159 14909 31168 14943
rect 31116 14900 31168 14909
rect 32496 14968 32548 15020
rect 32680 15011 32732 15020
rect 32680 14977 32689 15011
rect 32689 14977 32723 15011
rect 32723 14977 32732 15011
rect 32680 14968 32732 14977
rect 34428 15104 34480 15156
rect 39396 15104 39448 15156
rect 34980 14943 35032 14952
rect 34980 14909 34989 14943
rect 34989 14909 35023 14943
rect 35023 14909 35032 14943
rect 34980 14900 35032 14909
rect 35624 14968 35676 15020
rect 38752 15036 38804 15088
rect 36728 15011 36780 15020
rect 36728 14977 36737 15011
rect 36737 14977 36771 15011
rect 36771 14977 36780 15011
rect 36728 14968 36780 14977
rect 39028 14968 39080 15020
rect 41512 14968 41564 15020
rect 46940 15104 46992 15156
rect 47032 15104 47084 15156
rect 48320 15104 48372 15156
rect 50620 15147 50672 15156
rect 50620 15113 50629 15147
rect 50629 15113 50663 15147
rect 50663 15113 50672 15147
rect 50620 15104 50672 15113
rect 51448 15104 51500 15156
rect 44180 15036 44232 15088
rect 43536 14968 43588 15020
rect 45284 15011 45336 15020
rect 35716 14832 35768 14884
rect 39396 14900 39448 14952
rect 40500 14943 40552 14952
rect 40500 14909 40509 14943
rect 40509 14909 40543 14943
rect 40543 14909 40552 14943
rect 40500 14900 40552 14909
rect 41880 14900 41932 14952
rect 42524 14943 42576 14952
rect 42524 14909 42533 14943
rect 42533 14909 42567 14943
rect 42567 14909 42576 14943
rect 42524 14900 42576 14909
rect 42800 14900 42852 14952
rect 43720 14943 43772 14952
rect 43720 14909 43729 14943
rect 43729 14909 43763 14943
rect 43763 14909 43772 14943
rect 43720 14900 43772 14909
rect 44364 14900 44416 14952
rect 45284 14977 45293 15011
rect 45293 14977 45327 15011
rect 45327 14977 45336 15011
rect 45284 14968 45336 14977
rect 45652 14968 45704 15020
rect 45192 14900 45244 14952
rect 55588 14968 55640 15020
rect 47584 14900 47636 14952
rect 50160 14900 50212 14952
rect 52000 14943 52052 14952
rect 52000 14909 52009 14943
rect 52009 14909 52043 14943
rect 52043 14909 52052 14943
rect 52000 14900 52052 14909
rect 30012 14764 30064 14816
rect 31484 14807 31536 14816
rect 31484 14773 31493 14807
rect 31493 14773 31527 14807
rect 31527 14773 31536 14807
rect 31484 14764 31536 14773
rect 34060 14764 34112 14816
rect 39396 14764 39448 14816
rect 40132 14832 40184 14884
rect 45836 14832 45888 14884
rect 46940 14875 46992 14884
rect 46940 14841 46949 14875
rect 46949 14841 46983 14875
rect 46983 14841 46992 14875
rect 46940 14832 46992 14841
rect 39672 14764 39724 14816
rect 46204 14764 46256 14816
rect 52276 14832 52328 14884
rect 49700 14764 49752 14816
rect 18912 14662 18964 14714
rect 18976 14662 19028 14714
rect 19040 14662 19092 14714
rect 19104 14662 19156 14714
rect 36843 14662 36895 14714
rect 36907 14662 36959 14714
rect 36971 14662 37023 14714
rect 37035 14662 37087 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 3424 14467 3476 14476
rect 3424 14433 3433 14467
rect 3433 14433 3467 14467
rect 3467 14433 3476 14467
rect 3424 14424 3476 14433
rect 3976 14424 4028 14476
rect 6552 14603 6604 14612
rect 6552 14569 6561 14603
rect 6561 14569 6595 14603
rect 6595 14569 6604 14603
rect 6552 14560 6604 14569
rect 12808 14603 12860 14612
rect 12808 14569 12817 14603
rect 12817 14569 12851 14603
rect 12851 14569 12860 14603
rect 12808 14560 12860 14569
rect 13820 14603 13872 14612
rect 13820 14569 13829 14603
rect 13829 14569 13863 14603
rect 13863 14569 13872 14603
rect 13820 14560 13872 14569
rect 15384 14603 15436 14612
rect 15384 14569 15393 14603
rect 15393 14569 15427 14603
rect 15427 14569 15436 14603
rect 15384 14560 15436 14569
rect 15752 14560 15804 14612
rect 16948 14560 17000 14612
rect 24032 14560 24084 14612
rect 6920 14492 6972 14544
rect 8392 14492 8444 14544
rect 6460 14424 6512 14476
rect 4528 14356 4580 14408
rect 7288 14424 7340 14476
rect 10416 14424 10468 14476
rect 13728 14492 13780 14544
rect 18420 14535 18472 14544
rect 18420 14501 18429 14535
rect 18429 14501 18463 14535
rect 18463 14501 18472 14535
rect 18420 14492 18472 14501
rect 11152 14424 11204 14476
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 11704 14424 11756 14476
rect 12716 14424 12768 14476
rect 14832 14424 14884 14476
rect 20812 14492 20864 14544
rect 22008 14535 22060 14544
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 19708 14424 19760 14476
rect 22008 14501 22017 14535
rect 22017 14501 22051 14535
rect 22051 14501 22060 14535
rect 22008 14492 22060 14501
rect 23388 14535 23440 14544
rect 23388 14501 23397 14535
rect 23397 14501 23431 14535
rect 23431 14501 23440 14535
rect 23388 14492 23440 14501
rect 16028 14356 16080 14408
rect 5448 14263 5500 14272
rect 5448 14229 5457 14263
rect 5457 14229 5491 14263
rect 5491 14229 5500 14263
rect 5448 14220 5500 14229
rect 6644 14220 6696 14272
rect 12440 14220 12492 14272
rect 12992 14288 13044 14340
rect 15200 14288 15252 14340
rect 15384 14220 15436 14272
rect 19616 14288 19668 14340
rect 22928 14424 22980 14476
rect 25872 14560 25924 14612
rect 27528 14560 27580 14612
rect 30748 14560 30800 14612
rect 35716 14603 35768 14612
rect 35716 14569 35725 14603
rect 35725 14569 35759 14603
rect 35759 14569 35768 14603
rect 35716 14560 35768 14569
rect 40500 14560 40552 14612
rect 44180 14560 44232 14612
rect 48136 14560 48188 14612
rect 37740 14535 37792 14544
rect 25044 14424 25096 14476
rect 26516 14467 26568 14476
rect 26516 14433 26525 14467
rect 26525 14433 26559 14467
rect 26559 14433 26568 14467
rect 26516 14424 26568 14433
rect 27620 14424 27672 14476
rect 30104 14424 30156 14476
rect 32680 14424 32732 14476
rect 37740 14501 37749 14535
rect 37749 14501 37783 14535
rect 37783 14501 37792 14535
rect 37740 14492 37792 14501
rect 39396 14492 39448 14544
rect 42800 14492 42852 14544
rect 47584 14535 47636 14544
rect 47584 14501 47593 14535
rect 47593 14501 47627 14535
rect 47627 14501 47636 14535
rect 47584 14492 47636 14501
rect 34060 14467 34112 14476
rect 34060 14433 34069 14467
rect 34069 14433 34103 14467
rect 34103 14433 34112 14467
rect 34060 14424 34112 14433
rect 35164 14424 35216 14476
rect 28264 14356 28316 14408
rect 31484 14356 31536 14408
rect 34152 14399 34204 14408
rect 34152 14365 34161 14399
rect 34161 14365 34195 14399
rect 34195 14365 34204 14399
rect 35440 14424 35492 14476
rect 37832 14424 37884 14476
rect 38568 14424 38620 14476
rect 40132 14467 40184 14476
rect 40132 14433 40141 14467
rect 40141 14433 40175 14467
rect 40175 14433 40184 14467
rect 40132 14424 40184 14433
rect 34152 14356 34204 14365
rect 39764 14356 39816 14408
rect 42524 14424 42576 14476
rect 42892 14424 42944 14476
rect 44732 14424 44784 14476
rect 45836 14467 45888 14476
rect 45836 14433 45845 14467
rect 45845 14433 45879 14467
rect 45879 14433 45888 14467
rect 45836 14424 45888 14433
rect 46756 14424 46808 14476
rect 46940 14424 46992 14476
rect 47216 14467 47268 14476
rect 46204 14399 46256 14408
rect 46204 14365 46213 14399
rect 46213 14365 46247 14399
rect 46247 14365 46256 14399
rect 46204 14356 46256 14365
rect 47216 14433 47225 14467
rect 47225 14433 47259 14467
rect 47259 14433 47268 14467
rect 47216 14424 47268 14433
rect 49608 14492 49660 14544
rect 49700 14467 49752 14476
rect 49700 14433 49709 14467
rect 49709 14433 49743 14467
rect 49743 14433 49752 14467
rect 49700 14424 49752 14433
rect 52276 14467 52328 14476
rect 34428 14331 34480 14340
rect 34428 14297 34437 14331
rect 34437 14297 34471 14331
rect 34471 14297 34480 14331
rect 34428 14288 34480 14297
rect 35348 14331 35400 14340
rect 35348 14297 35357 14331
rect 35357 14297 35391 14331
rect 35391 14297 35400 14331
rect 35348 14288 35400 14297
rect 35532 14288 35584 14340
rect 37372 14288 37424 14340
rect 41696 14288 41748 14340
rect 42156 14288 42208 14340
rect 47216 14288 47268 14340
rect 52276 14433 52285 14467
rect 52285 14433 52319 14467
rect 52319 14433 52328 14467
rect 52276 14424 52328 14433
rect 50712 14288 50764 14340
rect 18420 14220 18472 14272
rect 22192 14220 22244 14272
rect 22744 14263 22796 14272
rect 22744 14229 22753 14263
rect 22753 14229 22787 14263
rect 22787 14229 22796 14263
rect 22744 14220 22796 14229
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 26240 14220 26292 14272
rect 30104 14220 30156 14272
rect 32036 14220 32088 14272
rect 37556 14220 37608 14272
rect 38568 14220 38620 14272
rect 40224 14263 40276 14272
rect 40224 14229 40233 14263
rect 40233 14229 40267 14263
rect 40267 14229 40276 14263
rect 40224 14220 40276 14229
rect 49608 14220 49660 14272
rect 49792 14220 49844 14272
rect 51448 14220 51500 14272
rect 51816 14263 51868 14272
rect 51816 14229 51825 14263
rect 51825 14229 51859 14263
rect 51859 14229 51868 14263
rect 51816 14220 51868 14229
rect 52460 14220 52512 14272
rect 9947 14118 9999 14170
rect 10011 14118 10063 14170
rect 10075 14118 10127 14170
rect 10139 14118 10191 14170
rect 27878 14118 27930 14170
rect 27942 14118 27994 14170
rect 28006 14118 28058 14170
rect 28070 14118 28122 14170
rect 45808 14118 45860 14170
rect 45872 14118 45924 14170
rect 45936 14118 45988 14170
rect 46000 14118 46052 14170
rect 5540 14016 5592 14068
rect 6276 14016 6328 14068
rect 8300 14016 8352 14068
rect 14280 14016 14332 14068
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 15844 14016 15896 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 25136 14016 25188 14068
rect 26424 14059 26476 14068
rect 26424 14025 26433 14059
rect 26433 14025 26467 14059
rect 26467 14025 26476 14059
rect 26424 14016 26476 14025
rect 28264 14059 28316 14068
rect 28264 14025 28273 14059
rect 28273 14025 28307 14059
rect 28307 14025 28316 14059
rect 28264 14016 28316 14025
rect 29368 14059 29420 14068
rect 29368 14025 29377 14059
rect 29377 14025 29411 14059
rect 29411 14025 29420 14059
rect 29368 14016 29420 14025
rect 2228 13812 2280 13864
rect 8760 13948 8812 14000
rect 11520 13948 11572 14000
rect 16948 13991 17000 14000
rect 16948 13957 16957 13991
rect 16957 13957 16991 13991
rect 16991 13957 17000 13991
rect 16948 13948 17000 13957
rect 4436 13855 4488 13864
rect 4436 13821 4445 13855
rect 4445 13821 4479 13855
rect 4479 13821 4488 13855
rect 4436 13812 4488 13821
rect 5448 13812 5500 13864
rect 7104 13812 7156 13864
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 2320 13676 2372 13728
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 12992 13880 13044 13932
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13636 13880 13688 13932
rect 13728 13880 13780 13932
rect 15476 13880 15528 13932
rect 15752 13923 15804 13932
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 13820 13812 13872 13864
rect 22744 13948 22796 14000
rect 41236 14016 41288 14068
rect 43720 14059 43772 14068
rect 43720 14025 43729 14059
rect 43729 14025 43763 14059
rect 43763 14025 43772 14059
rect 43720 14016 43772 14025
rect 44824 14016 44876 14068
rect 45192 14016 45244 14068
rect 49792 14016 49844 14068
rect 50712 14059 50764 14068
rect 50712 14025 50721 14059
rect 50721 14025 50755 14059
rect 50755 14025 50764 14059
rect 50712 14016 50764 14025
rect 52000 14059 52052 14068
rect 52000 14025 52009 14059
rect 52009 14025 52043 14059
rect 52043 14025 52052 14059
rect 52000 14016 52052 14025
rect 52460 14059 52512 14068
rect 52460 14025 52469 14059
rect 52469 14025 52503 14059
rect 52503 14025 52512 14059
rect 52460 14016 52512 14025
rect 32588 13991 32640 14000
rect 32588 13957 32597 13991
rect 32597 13957 32631 13991
rect 32631 13957 32640 13991
rect 32588 13948 32640 13957
rect 32956 13991 33008 14000
rect 32956 13957 32965 13991
rect 32965 13957 32999 13991
rect 32999 13957 33008 13991
rect 32956 13948 33008 13957
rect 35348 13948 35400 14000
rect 37372 13991 37424 14000
rect 37372 13957 37381 13991
rect 37381 13957 37415 13991
rect 37415 13957 37424 13991
rect 37372 13948 37424 13957
rect 16580 13812 16632 13864
rect 16672 13812 16724 13864
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 19432 13812 19484 13821
rect 19800 13855 19852 13864
rect 19800 13821 19809 13855
rect 19809 13821 19843 13855
rect 19843 13821 19852 13855
rect 19800 13812 19852 13821
rect 24860 13880 24912 13932
rect 24952 13880 25004 13932
rect 30104 13880 30156 13932
rect 22744 13855 22796 13864
rect 22744 13821 22753 13855
rect 22753 13821 22787 13855
rect 22787 13821 22796 13855
rect 22744 13812 22796 13821
rect 24216 13855 24268 13864
rect 24216 13821 24225 13855
rect 24225 13821 24259 13855
rect 24259 13821 24268 13855
rect 24216 13812 24268 13821
rect 24768 13812 24820 13864
rect 25412 13855 25464 13864
rect 20996 13787 21048 13796
rect 20996 13753 21005 13787
rect 21005 13753 21039 13787
rect 21039 13753 21048 13787
rect 20996 13744 21048 13753
rect 25412 13821 25421 13855
rect 25421 13821 25455 13855
rect 25455 13821 25464 13855
rect 25412 13812 25464 13821
rect 26516 13812 26568 13864
rect 29092 13812 29144 13864
rect 29276 13855 29328 13864
rect 29276 13821 29285 13855
rect 29285 13821 29319 13855
rect 29319 13821 29328 13855
rect 29276 13812 29328 13821
rect 31484 13855 31536 13864
rect 31484 13821 31493 13855
rect 31493 13821 31527 13855
rect 31527 13821 31536 13855
rect 31484 13812 31536 13821
rect 33048 13812 33100 13864
rect 38568 13880 38620 13932
rect 40224 13880 40276 13932
rect 42708 13880 42760 13932
rect 45284 13948 45336 14000
rect 34152 13812 34204 13864
rect 35440 13855 35492 13864
rect 35440 13821 35449 13855
rect 35449 13821 35483 13855
rect 35483 13821 35492 13855
rect 35440 13812 35492 13821
rect 35992 13812 36044 13864
rect 37556 13855 37608 13864
rect 37556 13821 37565 13855
rect 37565 13821 37599 13855
rect 37599 13821 37608 13855
rect 37556 13812 37608 13821
rect 37648 13855 37700 13864
rect 37648 13821 37657 13855
rect 37657 13821 37691 13855
rect 37691 13821 37700 13855
rect 37648 13812 37700 13821
rect 38200 13744 38252 13796
rect 40868 13812 40920 13864
rect 43076 13812 43128 13864
rect 43996 13812 44048 13864
rect 44824 13855 44876 13864
rect 44824 13821 44833 13855
rect 44833 13821 44867 13855
rect 44867 13821 44876 13855
rect 44824 13812 44876 13821
rect 49700 13880 49752 13932
rect 47308 13812 47360 13864
rect 49608 13855 49660 13864
rect 49608 13821 49617 13855
rect 49617 13821 49651 13855
rect 49651 13821 49660 13855
rect 49608 13812 49660 13821
rect 51448 13812 51500 13864
rect 41696 13744 41748 13796
rect 47124 13744 47176 13796
rect 48228 13744 48280 13796
rect 13268 13676 13320 13728
rect 14924 13676 14976 13728
rect 30932 13676 30984 13728
rect 41328 13676 41380 13728
rect 41512 13676 41564 13728
rect 49700 13719 49752 13728
rect 49700 13685 49709 13719
rect 49709 13685 49743 13719
rect 49743 13685 49752 13719
rect 49700 13676 49752 13685
rect 18912 13574 18964 13626
rect 18976 13574 19028 13626
rect 19040 13574 19092 13626
rect 19104 13574 19156 13626
rect 36843 13574 36895 13626
rect 36907 13574 36959 13626
rect 36971 13574 37023 13626
rect 37035 13574 37087 13626
rect 4436 13515 4488 13524
rect 4436 13481 4445 13515
rect 4445 13481 4479 13515
rect 4479 13481 4488 13515
rect 4436 13472 4488 13481
rect 8392 13472 8444 13524
rect 16028 13515 16080 13524
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 4896 13336 4948 13388
rect 7012 13404 7064 13456
rect 5448 13379 5500 13388
rect 5448 13345 5457 13379
rect 5457 13345 5491 13379
rect 5491 13345 5500 13379
rect 6920 13379 6972 13388
rect 5448 13336 5500 13345
rect 6920 13345 6929 13379
rect 6929 13345 6963 13379
rect 6963 13345 6972 13379
rect 6920 13336 6972 13345
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 16028 13481 16037 13515
rect 16037 13481 16071 13515
rect 16071 13481 16080 13515
rect 16028 13472 16080 13481
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 22376 13515 22428 13524
rect 22376 13481 22385 13515
rect 22385 13481 22419 13515
rect 22419 13481 22428 13515
rect 22376 13472 22428 13481
rect 24952 13472 25004 13524
rect 29552 13515 29604 13524
rect 29552 13481 29561 13515
rect 29561 13481 29595 13515
rect 29595 13481 29604 13515
rect 29552 13472 29604 13481
rect 30104 13472 30156 13524
rect 31484 13472 31536 13524
rect 42156 13515 42208 13524
rect 42156 13481 42165 13515
rect 42165 13481 42199 13515
rect 42199 13481 42208 13515
rect 42156 13472 42208 13481
rect 45652 13472 45704 13524
rect 51448 13515 51500 13524
rect 51448 13481 51457 13515
rect 51457 13481 51491 13515
rect 51491 13481 51500 13515
rect 51448 13472 51500 13481
rect 17224 13404 17276 13456
rect 24216 13404 24268 13456
rect 25688 13447 25740 13456
rect 5540 13268 5592 13320
rect 10324 13336 10376 13388
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 16672 13379 16724 13388
rect 13268 13268 13320 13320
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 21272 13379 21324 13388
rect 17684 13268 17736 13320
rect 19340 13268 19392 13320
rect 19432 13268 19484 13320
rect 21272 13345 21281 13379
rect 21281 13345 21315 13379
rect 21315 13345 21324 13379
rect 21272 13336 21324 13345
rect 25044 13379 25096 13388
rect 25044 13345 25053 13379
rect 25053 13345 25087 13379
rect 25087 13345 25096 13379
rect 25044 13336 25096 13345
rect 25228 13336 25280 13388
rect 19800 13268 19852 13320
rect 20720 13268 20772 13320
rect 25688 13413 25697 13447
rect 25697 13413 25731 13447
rect 25731 13413 25740 13447
rect 25688 13404 25740 13413
rect 26240 13336 26292 13388
rect 26884 13404 26936 13456
rect 27620 13336 27672 13388
rect 34152 13404 34204 13456
rect 35348 13404 35400 13456
rect 30932 13336 30984 13388
rect 32036 13336 32088 13388
rect 32404 13379 32456 13388
rect 28448 13311 28500 13320
rect 2320 13132 2372 13184
rect 8024 13132 8076 13184
rect 10324 13132 10376 13184
rect 10876 13132 10928 13184
rect 13544 13175 13596 13184
rect 13544 13141 13553 13175
rect 13553 13141 13587 13175
rect 13587 13141 13596 13175
rect 13544 13132 13596 13141
rect 19432 13175 19484 13184
rect 19432 13141 19456 13175
rect 19456 13141 19484 13175
rect 19432 13132 19484 13141
rect 19800 13132 19852 13184
rect 28448 13277 28457 13311
rect 28457 13277 28491 13311
rect 28491 13277 28500 13311
rect 28448 13268 28500 13277
rect 31668 13268 31720 13320
rect 32404 13345 32413 13379
rect 32413 13345 32447 13379
rect 32447 13345 32456 13379
rect 32404 13336 32456 13345
rect 33968 13336 34020 13388
rect 34520 13379 34572 13388
rect 34520 13345 34529 13379
rect 34529 13345 34563 13379
rect 34563 13345 34572 13379
rect 35992 13379 36044 13388
rect 34520 13336 34572 13345
rect 35992 13345 36001 13379
rect 36001 13345 36035 13379
rect 36035 13345 36044 13379
rect 35992 13336 36044 13345
rect 37648 13404 37700 13456
rect 41328 13404 41380 13456
rect 38200 13379 38252 13388
rect 38200 13345 38209 13379
rect 38209 13345 38243 13379
rect 38243 13345 38252 13379
rect 38200 13336 38252 13345
rect 40868 13379 40920 13388
rect 33232 13268 33284 13320
rect 33508 13268 33560 13320
rect 34980 13311 35032 13320
rect 34980 13277 34989 13311
rect 34989 13277 35023 13311
rect 35023 13277 35032 13311
rect 34980 13268 35032 13277
rect 38568 13268 38620 13320
rect 35532 13200 35584 13252
rect 40868 13345 40877 13379
rect 40877 13345 40911 13379
rect 40911 13345 40920 13379
rect 40868 13336 40920 13345
rect 41420 13336 41472 13388
rect 42708 13336 42760 13388
rect 44456 13379 44508 13388
rect 44456 13345 44465 13379
rect 44465 13345 44499 13379
rect 44499 13345 44508 13379
rect 44456 13336 44508 13345
rect 46756 13404 46808 13456
rect 43628 13311 43680 13320
rect 43628 13277 43637 13311
rect 43637 13277 43671 13311
rect 43671 13277 43680 13311
rect 43628 13268 43680 13277
rect 44088 13268 44140 13320
rect 44272 13268 44324 13320
rect 40868 13132 40920 13184
rect 41052 13175 41104 13184
rect 41052 13141 41061 13175
rect 41061 13141 41095 13175
rect 41095 13141 41104 13175
rect 41052 13132 41104 13141
rect 46204 13336 46256 13388
rect 46572 13336 46624 13388
rect 47308 13379 47360 13388
rect 47308 13345 47317 13379
rect 47317 13345 47351 13379
rect 47351 13345 47360 13379
rect 47308 13336 47360 13345
rect 49700 13336 49752 13388
rect 47860 13268 47912 13320
rect 51816 13268 51868 13320
rect 49332 13132 49384 13184
rect 9947 13030 9999 13082
rect 10011 13030 10063 13082
rect 10075 13030 10127 13082
rect 10139 13030 10191 13082
rect 27878 13030 27930 13082
rect 27942 13030 27994 13082
rect 28006 13030 28058 13082
rect 28070 13030 28122 13082
rect 45808 13030 45860 13082
rect 45872 13030 45924 13082
rect 45936 13030 45988 13082
rect 46000 13030 46052 13082
rect 2228 12971 2280 12980
rect 2228 12937 2237 12971
rect 2237 12937 2271 12971
rect 2271 12937 2280 12971
rect 2228 12928 2280 12937
rect 7104 12971 7156 12980
rect 7104 12937 7113 12971
rect 7113 12937 7147 12971
rect 7147 12937 7156 12971
rect 7104 12928 7156 12937
rect 9680 12928 9732 12980
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 11704 12928 11756 12980
rect 13360 12928 13412 12980
rect 14924 12971 14976 12980
rect 14924 12937 14933 12971
rect 14933 12937 14967 12971
rect 14967 12937 14976 12971
rect 14924 12928 14976 12937
rect 16672 12971 16724 12980
rect 16672 12937 16681 12971
rect 16681 12937 16715 12971
rect 16715 12937 16724 12971
rect 16672 12928 16724 12937
rect 19524 12928 19576 12980
rect 22744 12928 22796 12980
rect 23480 12928 23532 12980
rect 29092 12928 29144 12980
rect 8300 12860 8352 12912
rect 16488 12860 16540 12912
rect 26056 12903 26108 12912
rect 26056 12869 26065 12903
rect 26065 12869 26099 12903
rect 26099 12869 26108 12903
rect 26056 12860 26108 12869
rect 31392 12928 31444 12980
rect 34428 12928 34480 12980
rect 41696 12971 41748 12980
rect 2412 12767 2464 12776
rect 2412 12733 2413 12767
rect 2413 12733 2447 12767
rect 2447 12733 2464 12767
rect 2412 12724 2464 12733
rect 3424 12767 3476 12776
rect 3424 12733 3433 12767
rect 3433 12733 3467 12767
rect 3467 12733 3476 12767
rect 3424 12724 3476 12733
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 6184 12724 6236 12776
rect 25688 12792 25740 12844
rect 36452 12860 36504 12912
rect 33968 12835 34020 12844
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 8852 12724 8904 12776
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 13176 12724 13228 12776
rect 13544 12724 13596 12776
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 16028 12724 16080 12776
rect 17592 12724 17644 12776
rect 19616 12767 19668 12776
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 21548 12767 21600 12776
rect 21548 12733 21565 12767
rect 21565 12733 21599 12767
rect 21599 12733 21600 12767
rect 21548 12724 21600 12733
rect 22468 12724 22520 12776
rect 24032 12767 24084 12776
rect 24032 12733 24041 12767
rect 24041 12733 24075 12767
rect 24075 12733 24084 12767
rect 24032 12724 24084 12733
rect 9956 12656 10008 12708
rect 19708 12656 19760 12708
rect 24952 12724 25004 12776
rect 26424 12724 26476 12776
rect 26792 12767 26844 12776
rect 26792 12733 26801 12767
rect 26801 12733 26835 12767
rect 26835 12733 26844 12767
rect 26792 12724 26844 12733
rect 27252 12724 27304 12776
rect 28908 12724 28960 12776
rect 33968 12801 33977 12835
rect 33977 12801 34011 12835
rect 34011 12801 34020 12835
rect 33968 12792 34020 12801
rect 34980 12792 35032 12844
rect 41696 12937 41705 12971
rect 41705 12937 41739 12971
rect 41739 12937 41748 12971
rect 41696 12928 41748 12937
rect 37740 12860 37792 12912
rect 25136 12656 25188 12708
rect 27712 12656 27764 12708
rect 28172 12656 28224 12708
rect 29460 12656 29512 12708
rect 31668 12724 31720 12776
rect 32404 12724 32456 12776
rect 33416 12767 33468 12776
rect 33416 12733 33425 12767
rect 33425 12733 33459 12767
rect 33459 12733 33468 12767
rect 33416 12724 33468 12733
rect 39672 12792 39724 12844
rect 33324 12656 33376 12708
rect 2412 12588 2464 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 4988 12588 5040 12640
rect 12992 12588 13044 12640
rect 13912 12588 13964 12640
rect 23756 12588 23808 12640
rect 24032 12588 24084 12640
rect 24676 12588 24728 12640
rect 35992 12724 36044 12776
rect 39120 12767 39172 12776
rect 39120 12733 39129 12767
rect 39129 12733 39163 12767
rect 39163 12733 39172 12767
rect 39120 12724 39172 12733
rect 40040 12860 40092 12912
rect 41052 12767 41104 12776
rect 34612 12588 34664 12640
rect 41052 12733 41061 12767
rect 41061 12733 41095 12767
rect 41095 12733 41104 12767
rect 41052 12724 41104 12733
rect 44824 12928 44876 12980
rect 47860 12971 47912 12980
rect 47860 12937 47869 12971
rect 47869 12937 47903 12971
rect 47903 12937 47912 12971
rect 47860 12928 47912 12937
rect 49332 12971 49384 12980
rect 49332 12937 49341 12971
rect 49341 12937 49375 12971
rect 49375 12937 49384 12971
rect 49332 12928 49384 12937
rect 44088 12903 44140 12912
rect 44088 12869 44097 12903
rect 44097 12869 44131 12903
rect 44131 12869 44140 12903
rect 44088 12860 44140 12869
rect 44456 12792 44508 12844
rect 47124 12835 47176 12844
rect 47124 12801 47133 12835
rect 47133 12801 47167 12835
rect 47167 12801 47176 12835
rect 47124 12792 47176 12801
rect 48228 12835 48280 12844
rect 48228 12801 48237 12835
rect 48237 12801 48271 12835
rect 48271 12801 48280 12835
rect 48228 12792 48280 12801
rect 39580 12699 39632 12708
rect 39580 12665 39589 12699
rect 39589 12665 39623 12699
rect 39623 12665 39632 12699
rect 39580 12656 39632 12665
rect 39672 12656 39724 12708
rect 44272 12724 44324 12776
rect 46572 12767 46624 12776
rect 46572 12733 46581 12767
rect 46581 12733 46615 12767
rect 46615 12733 46624 12767
rect 46572 12724 46624 12733
rect 46756 12767 46808 12776
rect 46756 12733 46765 12767
rect 46765 12733 46799 12767
rect 46799 12733 46808 12767
rect 46756 12724 46808 12733
rect 40040 12588 40092 12640
rect 40316 12588 40368 12640
rect 41972 12631 42024 12640
rect 41972 12597 41981 12631
rect 41981 12597 42015 12631
rect 42015 12597 42024 12631
rect 41972 12588 42024 12597
rect 18912 12486 18964 12538
rect 18976 12486 19028 12538
rect 19040 12486 19092 12538
rect 19104 12486 19156 12538
rect 36843 12486 36895 12538
rect 36907 12486 36959 12538
rect 36971 12486 37023 12538
rect 37035 12486 37087 12538
rect 3424 12384 3476 12436
rect 4896 12384 4948 12436
rect 6184 12384 6236 12436
rect 9956 12427 10008 12436
rect 9956 12393 9965 12427
rect 9965 12393 9999 12427
rect 9999 12393 10008 12427
rect 9956 12384 10008 12393
rect 10600 12384 10652 12436
rect 3240 12248 3292 12300
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 6920 12248 6972 12300
rect 7564 12248 7616 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8576 12248 8628 12300
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 5540 12044 5592 12096
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 7932 12044 7984 12096
rect 10876 12180 10928 12232
rect 15660 12248 15712 12300
rect 16580 12248 16632 12300
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 15292 12112 15344 12164
rect 16580 12155 16632 12164
rect 16580 12121 16589 12155
rect 16589 12121 16623 12155
rect 16623 12121 16632 12155
rect 16580 12112 16632 12121
rect 13912 12044 13964 12096
rect 14648 12044 14700 12096
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 19708 12384 19760 12436
rect 26424 12384 26476 12436
rect 29092 12427 29144 12436
rect 29092 12393 29101 12427
rect 29101 12393 29135 12427
rect 29135 12393 29144 12427
rect 29092 12384 29144 12393
rect 30748 12384 30800 12436
rect 19340 12316 19392 12368
rect 20996 12316 21048 12368
rect 25044 12316 25096 12368
rect 30104 12316 30156 12368
rect 17500 12248 17552 12257
rect 19616 12291 19668 12300
rect 19616 12257 19625 12291
rect 19625 12257 19659 12291
rect 19659 12257 19668 12291
rect 19616 12248 19668 12257
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 21088 12291 21140 12300
rect 19800 12248 19852 12257
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 23480 12248 23532 12300
rect 25136 12291 25188 12300
rect 25136 12257 25145 12291
rect 25145 12257 25179 12291
rect 25179 12257 25188 12291
rect 25136 12248 25188 12257
rect 25412 12248 25464 12300
rect 26240 12248 26292 12300
rect 22008 12180 22060 12232
rect 26792 12248 26844 12300
rect 28264 12248 28316 12300
rect 30472 12291 30524 12300
rect 30472 12257 30481 12291
rect 30481 12257 30515 12291
rect 30515 12257 30524 12291
rect 30472 12248 30524 12257
rect 29460 12180 29512 12232
rect 34704 12384 34756 12436
rect 40316 12384 40368 12436
rect 40868 12384 40920 12436
rect 43076 12427 43128 12436
rect 43076 12393 43085 12427
rect 43085 12393 43119 12427
rect 43119 12393 43128 12427
rect 43076 12384 43128 12393
rect 44732 12427 44784 12436
rect 44732 12393 44741 12427
rect 44741 12393 44775 12427
rect 44775 12393 44784 12427
rect 44732 12384 44784 12393
rect 31668 12316 31720 12368
rect 32588 12248 32640 12300
rect 34336 12248 34388 12300
rect 35072 12248 35124 12300
rect 35440 12291 35492 12300
rect 35440 12257 35449 12291
rect 35449 12257 35483 12291
rect 35483 12257 35492 12291
rect 35440 12248 35492 12257
rect 43628 12291 43680 12300
rect 43628 12257 43637 12291
rect 43637 12257 43671 12291
rect 43671 12257 43680 12291
rect 43628 12248 43680 12257
rect 31116 12180 31168 12232
rect 32680 12223 32732 12232
rect 32680 12189 32689 12223
rect 32689 12189 32723 12223
rect 32723 12189 32732 12223
rect 32680 12180 32732 12189
rect 32772 12180 32824 12232
rect 39580 12180 39632 12232
rect 18880 12044 18932 12096
rect 26056 12112 26108 12164
rect 29092 12112 29144 12164
rect 23940 12044 23992 12096
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 28448 12044 28500 12096
rect 30932 12112 30984 12164
rect 32772 12044 32824 12096
rect 35624 12087 35676 12096
rect 35624 12053 35633 12087
rect 35633 12053 35667 12087
rect 35667 12053 35676 12087
rect 35624 12044 35676 12053
rect 41972 12044 42024 12096
rect 9947 11942 9999 11994
rect 10011 11942 10063 11994
rect 10075 11942 10127 11994
rect 10139 11942 10191 11994
rect 27878 11942 27930 11994
rect 27942 11942 27994 11994
rect 28006 11942 28058 11994
rect 28070 11942 28122 11994
rect 45808 11942 45860 11994
rect 45872 11942 45924 11994
rect 45936 11942 45988 11994
rect 46000 11942 46052 11994
rect 4528 11840 4580 11892
rect 7564 11883 7616 11892
rect 7564 11849 7573 11883
rect 7573 11849 7607 11883
rect 7607 11849 7616 11883
rect 7564 11840 7616 11849
rect 8576 11883 8628 11892
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 13820 11840 13872 11892
rect 15200 11883 15252 11892
rect 15200 11849 15209 11883
rect 15209 11849 15243 11883
rect 15243 11849 15252 11883
rect 15200 11840 15252 11849
rect 15292 11840 15344 11892
rect 17592 11840 17644 11892
rect 17684 11840 17736 11892
rect 18880 11840 18932 11892
rect 30012 11883 30064 11892
rect 13912 11772 13964 11824
rect 20720 11772 20772 11824
rect 22008 11772 22060 11824
rect 30012 11849 30021 11883
rect 30021 11849 30055 11883
rect 30055 11849 30064 11883
rect 30012 11840 30064 11849
rect 2136 11636 2188 11688
rect 6828 11704 6880 11756
rect 16028 11747 16080 11756
rect 16028 11713 16037 11747
rect 16037 11713 16071 11747
rect 16071 11713 16080 11747
rect 16028 11704 16080 11713
rect 16580 11747 16632 11756
rect 16580 11713 16589 11747
rect 16589 11713 16623 11747
rect 16623 11713 16632 11747
rect 16580 11704 16632 11713
rect 17132 11704 17184 11756
rect 19524 11747 19576 11756
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 7932 11636 7984 11688
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 9772 11679 9824 11688
rect 9772 11645 9781 11679
rect 9781 11645 9815 11679
rect 9815 11645 9824 11679
rect 9772 11636 9824 11645
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 11428 11636 11480 11688
rect 13452 11636 13504 11688
rect 14280 11636 14332 11688
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 17500 11636 17552 11688
rect 17960 11636 18012 11688
rect 19524 11713 19533 11747
rect 19533 11713 19567 11747
rect 19567 11713 19576 11747
rect 19524 11704 19576 11713
rect 20720 11636 20772 11688
rect 21916 11679 21968 11688
rect 21916 11645 21925 11679
rect 21925 11645 21959 11679
rect 21959 11645 21968 11679
rect 21916 11636 21968 11645
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 25136 11636 25188 11688
rect 20904 11611 20956 11620
rect 20904 11577 20913 11611
rect 20913 11577 20947 11611
rect 20947 11577 20956 11611
rect 20904 11568 20956 11577
rect 21640 11568 21692 11620
rect 26240 11636 26292 11688
rect 27252 11636 27304 11688
rect 31208 11679 31260 11688
rect 31208 11645 31217 11679
rect 31217 11645 31251 11679
rect 31251 11645 31260 11679
rect 31208 11636 31260 11645
rect 32680 11772 32732 11824
rect 33416 11840 33468 11892
rect 32772 11704 32824 11756
rect 35440 11772 35492 11824
rect 36452 11840 36504 11892
rect 36820 11883 36872 11892
rect 36820 11849 36829 11883
rect 36829 11849 36863 11883
rect 36863 11849 36872 11883
rect 36820 11840 36872 11849
rect 39120 11840 39172 11892
rect 36820 11704 36872 11756
rect 32588 11679 32640 11688
rect 32588 11645 32597 11679
rect 32597 11645 32631 11679
rect 32631 11645 32640 11679
rect 32588 11636 32640 11645
rect 33324 11636 33376 11688
rect 34612 11636 34664 11688
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 5264 11500 5316 11552
rect 7012 11500 7064 11552
rect 9036 11500 9088 11552
rect 9680 11500 9732 11552
rect 14372 11500 14424 11552
rect 21732 11543 21784 11552
rect 21732 11509 21741 11543
rect 21741 11509 21775 11543
rect 21775 11509 21784 11543
rect 21732 11500 21784 11509
rect 30472 11568 30524 11620
rect 34704 11568 34756 11620
rect 35624 11636 35676 11688
rect 25596 11500 25648 11552
rect 27252 11543 27304 11552
rect 27252 11509 27261 11543
rect 27261 11509 27295 11543
rect 27295 11509 27304 11543
rect 27252 11500 27304 11509
rect 34336 11500 34388 11552
rect 18912 11398 18964 11450
rect 18976 11398 19028 11450
rect 19040 11398 19092 11450
rect 19104 11398 19156 11450
rect 36843 11398 36895 11450
rect 36907 11398 36959 11450
rect 36971 11398 37023 11450
rect 37035 11398 37087 11450
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 4528 11296 4580 11348
rect 6920 11296 6972 11348
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 21088 11296 21140 11348
rect 3332 11228 3384 11280
rect 4252 11160 4304 11212
rect 5264 11160 5316 11212
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 14004 11228 14056 11280
rect 9036 11203 9088 11212
rect 9036 11169 9045 11203
rect 9045 11169 9079 11203
rect 9079 11169 9088 11203
rect 9036 11160 9088 11169
rect 11428 11160 11480 11212
rect 12532 11160 12584 11212
rect 6184 11092 6236 11144
rect 12992 11160 13044 11212
rect 17132 11160 17184 11212
rect 18052 11160 18104 11212
rect 18236 11203 18288 11212
rect 18236 11169 18245 11203
rect 18245 11169 18279 11203
rect 18279 11169 18288 11203
rect 18236 11160 18288 11169
rect 20076 11160 20128 11212
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 22100 11203 22152 11212
rect 22100 11169 22109 11203
rect 22109 11169 22143 11203
rect 22143 11169 22152 11203
rect 22100 11160 22152 11169
rect 22376 11160 22428 11212
rect 24124 11203 24176 11212
rect 24124 11169 24133 11203
rect 24133 11169 24167 11203
rect 24167 11169 24176 11203
rect 24124 11160 24176 11169
rect 24768 11228 24820 11280
rect 25688 11296 25740 11348
rect 32772 11296 32824 11348
rect 26056 11228 26108 11280
rect 14188 11092 14240 11144
rect 24952 11203 25004 11212
rect 24952 11169 24961 11203
rect 24961 11169 24995 11203
rect 24995 11169 25004 11203
rect 27436 11203 27488 11212
rect 24952 11160 25004 11169
rect 27436 11169 27445 11203
rect 27445 11169 27479 11203
rect 27479 11169 27488 11203
rect 27436 11160 27488 11169
rect 30104 11271 30156 11280
rect 30104 11237 30113 11271
rect 30113 11237 30147 11271
rect 30147 11237 30156 11271
rect 30104 11228 30156 11237
rect 33324 11296 33376 11348
rect 34520 11296 34572 11348
rect 35072 11271 35124 11280
rect 35072 11237 35081 11271
rect 35081 11237 35115 11271
rect 35115 11237 35124 11271
rect 35072 11228 35124 11237
rect 27252 11092 27304 11144
rect 28264 11160 28316 11212
rect 28172 11092 28224 11144
rect 32220 11160 32272 11212
rect 33232 11160 33284 11212
rect 34612 11160 34664 11212
rect 34704 11203 34756 11212
rect 34704 11169 34713 11203
rect 34713 11169 34747 11203
rect 34747 11169 34756 11203
rect 34704 11160 34756 11169
rect 4620 11024 4672 11076
rect 13636 11024 13688 11076
rect 15384 11024 15436 11076
rect 18420 11024 18472 11076
rect 22560 11024 22612 11076
rect 23020 11024 23072 11076
rect 6368 10956 6420 11008
rect 13728 10956 13780 11008
rect 17408 10956 17460 11008
rect 18972 10956 19024 11008
rect 19984 10956 20036 11008
rect 23940 10999 23992 11008
rect 23940 10965 23949 10999
rect 23949 10965 23983 10999
rect 23983 10965 23992 10999
rect 23940 10956 23992 10965
rect 9947 10854 9999 10906
rect 10011 10854 10063 10906
rect 10075 10854 10127 10906
rect 10139 10854 10191 10906
rect 27878 10854 27930 10906
rect 27942 10854 27994 10906
rect 28006 10854 28058 10906
rect 28070 10854 28122 10906
rect 45808 10854 45860 10906
rect 45872 10854 45924 10906
rect 45936 10854 45988 10906
rect 46000 10854 46052 10906
rect 4436 10752 4488 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 9772 10752 9824 10804
rect 11428 10795 11480 10804
rect 11428 10761 11437 10795
rect 11437 10761 11471 10795
rect 11471 10761 11480 10795
rect 11428 10752 11480 10761
rect 12532 10752 12584 10804
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 17132 10752 17184 10804
rect 21548 10752 21600 10804
rect 25228 10752 25280 10804
rect 26240 10752 26292 10804
rect 32220 10752 32272 10804
rect 16672 10684 16724 10736
rect 2320 10591 2372 10600
rect 2320 10557 2329 10591
rect 2329 10557 2363 10591
rect 2363 10557 2372 10591
rect 2320 10548 2372 10557
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 4344 10591 4396 10600
rect 4344 10557 4353 10591
rect 4353 10557 4387 10591
rect 4387 10557 4396 10591
rect 4344 10548 4396 10557
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 9680 10548 9732 10600
rect 11520 10548 11572 10600
rect 12532 10548 12584 10600
rect 13544 10548 13596 10600
rect 14372 10591 14424 10600
rect 14372 10557 14381 10591
rect 14381 10557 14415 10591
rect 14415 10557 14424 10591
rect 14372 10548 14424 10557
rect 16028 10548 16080 10600
rect 17040 10548 17092 10600
rect 17408 10591 17460 10600
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 17408 10548 17460 10557
rect 18972 10591 19024 10600
rect 18972 10557 18981 10591
rect 18981 10557 19015 10591
rect 19015 10557 19024 10591
rect 18972 10548 19024 10557
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 32956 10752 33008 10804
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 22560 10548 22612 10600
rect 23940 10548 23992 10600
rect 25596 10591 25648 10600
rect 25596 10557 25605 10591
rect 25605 10557 25639 10591
rect 25639 10557 25648 10591
rect 25596 10548 25648 10557
rect 29276 10548 29328 10600
rect 29368 10548 29420 10600
rect 31116 10548 31168 10600
rect 34520 10548 34572 10600
rect 3240 10412 3292 10464
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 5540 10412 5592 10464
rect 9496 10412 9548 10464
rect 16120 10412 16172 10464
rect 17408 10412 17460 10464
rect 19432 10412 19484 10464
rect 20260 10412 20312 10464
rect 21824 10412 21876 10464
rect 24308 10412 24360 10464
rect 27252 10455 27304 10464
rect 27252 10421 27261 10455
rect 27261 10421 27295 10455
rect 27295 10421 27304 10455
rect 27252 10412 27304 10421
rect 29000 10412 29052 10464
rect 37188 10412 37240 10464
rect 18912 10310 18964 10362
rect 18976 10310 19028 10362
rect 19040 10310 19092 10362
rect 19104 10310 19156 10362
rect 36843 10310 36895 10362
rect 36907 10310 36959 10362
rect 36971 10310 37023 10362
rect 37035 10310 37087 10362
rect 3332 10208 3384 10260
rect 7288 10208 7340 10260
rect 11520 10251 11572 10260
rect 3240 10072 3292 10124
rect 4804 10072 4856 10124
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 11520 10217 11529 10251
rect 11529 10217 11563 10251
rect 11563 10217 11572 10251
rect 11520 10208 11572 10217
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 13544 10251 13596 10260
rect 13544 10217 13553 10251
rect 13553 10217 13587 10251
rect 13587 10217 13596 10251
rect 13544 10208 13596 10217
rect 16028 10251 16080 10260
rect 16028 10217 16037 10251
rect 16037 10217 16071 10251
rect 16071 10217 16080 10251
rect 16028 10208 16080 10217
rect 17040 10251 17092 10260
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 18052 10251 18104 10260
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 22008 10208 22060 10260
rect 22100 10208 22152 10260
rect 27436 10208 27488 10260
rect 29276 10251 29328 10260
rect 29276 10217 29285 10251
rect 29285 10217 29319 10251
rect 29319 10217 29328 10251
rect 29276 10208 29328 10217
rect 8208 10115 8260 10124
rect 8208 10081 8217 10115
rect 8217 10081 8251 10115
rect 8251 10081 8260 10115
rect 8208 10072 8260 10081
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 12624 10072 12676 10124
rect 13728 10115 13780 10124
rect 13728 10081 13737 10115
rect 13737 10081 13771 10115
rect 13771 10081 13780 10115
rect 13728 10072 13780 10081
rect 17132 10072 17184 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 18052 10072 18104 10124
rect 20076 10072 20128 10124
rect 20260 10115 20312 10124
rect 20260 10081 20269 10115
rect 20269 10081 20303 10115
rect 20303 10081 20312 10115
rect 20260 10072 20312 10081
rect 21824 10115 21876 10124
rect 21824 10081 21833 10115
rect 21833 10081 21867 10115
rect 21867 10081 21876 10115
rect 21824 10072 21876 10081
rect 22836 10115 22888 10124
rect 22836 10081 22845 10115
rect 22845 10081 22879 10115
rect 22879 10081 22888 10115
rect 22836 10072 22888 10081
rect 24216 10072 24268 10124
rect 25596 10115 25648 10124
rect 25596 10081 25605 10115
rect 25605 10081 25639 10115
rect 25639 10081 25648 10115
rect 25596 10072 25648 10081
rect 27436 10115 27488 10124
rect 27436 10081 27445 10115
rect 27445 10081 27479 10115
rect 27479 10081 27488 10115
rect 27436 10072 27488 10081
rect 27528 10072 27580 10124
rect 29460 10115 29512 10124
rect 29460 10081 29469 10115
rect 29469 10081 29503 10115
rect 29503 10081 29512 10115
rect 29460 10072 29512 10081
rect 29552 10072 29604 10124
rect 32864 10072 32916 10124
rect 34244 10115 34296 10124
rect 34244 10081 34253 10115
rect 34253 10081 34287 10115
rect 34287 10081 34296 10115
rect 34244 10072 34296 10081
rect 36176 10072 36228 10124
rect 37648 10072 37700 10124
rect 14188 10004 14240 10056
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 4160 9868 4212 9920
rect 11428 9868 11480 9920
rect 20628 9868 20680 9920
rect 24584 9868 24636 9920
rect 26240 9868 26292 9920
rect 27620 9868 27672 9920
rect 30748 9868 30800 9920
rect 32956 9868 33008 9920
rect 33324 9868 33376 9920
rect 35992 9868 36044 9920
rect 36820 9868 36872 9920
rect 9947 9766 9999 9818
rect 10011 9766 10063 9818
rect 10075 9766 10127 9818
rect 10139 9766 10191 9818
rect 27878 9766 27930 9818
rect 27942 9766 27994 9818
rect 28006 9766 28058 9818
rect 28070 9766 28122 9818
rect 45808 9766 45860 9818
rect 45872 9766 45924 9818
rect 45936 9766 45988 9818
rect 46000 9766 46052 9818
rect 5356 9664 5408 9716
rect 8208 9664 8260 9716
rect 12624 9664 12676 9716
rect 27436 9707 27488 9716
rect 27436 9673 27445 9707
rect 27445 9673 27479 9707
rect 27479 9673 27488 9707
rect 27436 9664 27488 9673
rect 6000 9596 6052 9648
rect 14188 9639 14240 9648
rect 14188 9605 14197 9639
rect 14197 9605 14231 9639
rect 14231 9605 14240 9639
rect 14188 9596 14240 9605
rect 17132 9596 17184 9648
rect 22836 9596 22888 9648
rect 25596 9596 25648 9648
rect 29552 9596 29604 9648
rect 34244 9596 34296 9648
rect 36176 9596 36228 9648
rect 37648 9639 37700 9648
rect 37648 9605 37657 9639
rect 37657 9605 37691 9639
rect 37691 9605 37700 9639
rect 37648 9596 37700 9605
rect 5172 9528 5224 9580
rect 4160 9460 4212 9512
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 5448 9460 5500 9512
rect 7472 9460 7524 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 12440 9460 12492 9512
rect 13452 9460 13504 9512
rect 13912 9460 13964 9512
rect 16028 9460 16080 9512
rect 16120 9460 16172 9512
rect 17408 9503 17460 9512
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 19984 9503 20036 9512
rect 4344 9324 4396 9376
rect 10784 9392 10836 9444
rect 19984 9469 19993 9503
rect 19993 9469 20027 9503
rect 20027 9469 20036 9503
rect 19984 9460 20036 9469
rect 20812 9460 20864 9512
rect 21732 9460 21784 9512
rect 23020 9503 23072 9512
rect 23020 9469 23029 9503
rect 23029 9469 23063 9503
rect 23063 9469 23072 9503
rect 23020 9460 23072 9469
rect 24584 9503 24636 9512
rect 24584 9469 24593 9503
rect 24593 9469 24627 9503
rect 24627 9469 24636 9503
rect 24584 9460 24636 9469
rect 25688 9460 25740 9512
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 27620 9503 27672 9512
rect 27620 9469 27629 9503
rect 27629 9469 27663 9503
rect 27663 9469 27672 9503
rect 27620 9460 27672 9469
rect 28724 9460 28776 9512
rect 29736 9460 29788 9512
rect 31760 9460 31812 9512
rect 32128 9460 32180 9512
rect 33140 9460 33192 9512
rect 35808 9503 35860 9512
rect 35808 9469 35817 9503
rect 35817 9469 35851 9503
rect 35851 9469 35860 9503
rect 35808 9460 35860 9469
rect 36820 9503 36872 9512
rect 36820 9469 36829 9503
rect 36829 9469 36863 9503
rect 36863 9469 36872 9503
rect 36820 9460 36872 9469
rect 38476 9460 38528 9512
rect 20720 9392 20772 9444
rect 7656 9324 7708 9376
rect 11612 9324 11664 9376
rect 13820 9324 13872 9376
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 19248 9324 19300 9376
rect 20260 9324 20312 9376
rect 22008 9324 22060 9376
rect 22836 9367 22888 9376
rect 22836 9333 22845 9367
rect 22845 9333 22879 9367
rect 22879 9333 22888 9367
rect 22836 9324 22888 9333
rect 29460 9392 29512 9444
rect 26332 9324 26384 9376
rect 30932 9324 30984 9376
rect 32312 9324 32364 9376
rect 34520 9324 34572 9376
rect 36728 9324 36780 9376
rect 18912 9222 18964 9274
rect 18976 9222 19028 9274
rect 19040 9222 19092 9274
rect 19104 9222 19156 9274
rect 36843 9222 36895 9274
rect 36907 9222 36959 9274
rect 36971 9222 37023 9274
rect 37035 9222 37087 9274
rect 4804 9163 4856 9172
rect 4804 9129 4813 9163
rect 4813 9129 4847 9163
rect 4847 9129 4856 9163
rect 4804 9120 4856 9129
rect 7472 9163 7524 9172
rect 7472 9129 7481 9163
rect 7481 9129 7515 9163
rect 7515 9129 7524 9163
rect 7472 9120 7524 9129
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 13452 9163 13504 9172
rect 12440 9120 12492 9129
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 16028 9163 16080 9172
rect 16028 9129 16037 9163
rect 16037 9129 16071 9163
rect 16071 9129 16080 9163
rect 16028 9120 16080 9129
rect 20076 9163 20128 9172
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 21916 9120 21968 9172
rect 24216 9120 24268 9172
rect 27528 9120 27580 9172
rect 28724 9163 28776 9172
rect 28724 9129 28733 9163
rect 28733 9129 28767 9163
rect 28767 9129 28776 9163
rect 28724 9120 28776 9129
rect 29736 9163 29788 9172
rect 29736 9129 29745 9163
rect 29745 9129 29779 9163
rect 29779 9129 29788 9163
rect 29736 9120 29788 9129
rect 32128 9120 32180 9172
rect 33140 9163 33192 9172
rect 33140 9129 33149 9163
rect 33149 9129 33183 9163
rect 33183 9129 33192 9163
rect 33140 9120 33192 9129
rect 38476 9163 38528 9172
rect 38476 9129 38485 9163
rect 38485 9129 38519 9163
rect 38519 9129 38528 9163
rect 38476 9120 38528 9129
rect 2136 9052 2188 9104
rect 10508 9052 10560 9104
rect 10692 9052 10744 9104
rect 2872 8984 2924 9036
rect 5540 8984 5592 9036
rect 7472 8984 7524 9036
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 8668 9027 8720 9036
rect 8668 8993 8677 9027
rect 8677 8993 8711 9027
rect 8711 8993 8720 9027
rect 8668 8984 8720 8993
rect 11612 9027 11664 9036
rect 8024 8848 8076 8900
rect 8208 8848 8260 8900
rect 11244 8848 11296 8900
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 13176 8984 13228 9036
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 16212 9027 16264 9036
rect 16212 8993 16221 9027
rect 16221 8993 16255 9027
rect 16255 8993 16264 9027
rect 16212 8984 16264 8993
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 19248 9027 19300 9036
rect 19248 8993 19257 9027
rect 19257 8993 19291 9027
rect 19291 8993 19300 9027
rect 19248 8984 19300 8993
rect 20260 9027 20312 9036
rect 20260 8993 20269 9027
rect 20269 8993 20303 9027
rect 20303 8993 20312 9027
rect 20260 8984 20312 8993
rect 22836 8984 22888 9036
rect 23112 8984 23164 9036
rect 24308 9027 24360 9036
rect 24308 8993 24317 9027
rect 24317 8993 24351 9027
rect 24351 8993 24360 9027
rect 24308 8984 24360 8993
rect 27252 9052 27304 9104
rect 37188 9052 37240 9104
rect 26332 9027 26384 9036
rect 26332 8993 26341 9027
rect 26341 8993 26375 9027
rect 26375 8993 26384 9027
rect 26332 8984 26384 8993
rect 27160 8984 27212 9036
rect 29552 8984 29604 9036
rect 30564 8984 30616 9036
rect 30932 9027 30984 9036
rect 30932 8993 30941 9027
rect 30941 8993 30975 9027
rect 30975 8993 30984 9027
rect 30932 8984 30984 8993
rect 32772 8984 32824 9036
rect 33324 9027 33376 9036
rect 33324 8993 33333 9027
rect 33333 8993 33367 9027
rect 33367 8993 33376 9027
rect 33324 8984 33376 8993
rect 35348 9027 35400 9036
rect 35348 8993 35357 9027
rect 35357 8993 35391 9027
rect 35391 8993 35400 9027
rect 35348 8984 35400 8993
rect 37648 8984 37700 9036
rect 17040 8891 17092 8900
rect 17040 8857 17049 8891
rect 17049 8857 17083 8891
rect 17083 8857 17092 8891
rect 17040 8848 17092 8857
rect 17960 8848 18012 8900
rect 7656 8780 7708 8832
rect 7748 8780 7800 8832
rect 11704 8780 11756 8832
rect 18972 8780 19024 8832
rect 24032 8780 24084 8832
rect 26148 8823 26200 8832
rect 26148 8789 26157 8823
rect 26157 8789 26191 8823
rect 26191 8789 26200 8823
rect 26148 8780 26200 8789
rect 28724 8780 28776 8832
rect 31208 8780 31260 8832
rect 33968 8780 34020 8832
rect 35164 8823 35216 8832
rect 35164 8789 35173 8823
rect 35173 8789 35207 8823
rect 35207 8789 35216 8823
rect 35164 8780 35216 8789
rect 9947 8678 9999 8730
rect 10011 8678 10063 8730
rect 10075 8678 10127 8730
rect 10139 8678 10191 8730
rect 27878 8678 27930 8730
rect 27942 8678 27994 8730
rect 28006 8678 28058 8730
rect 28070 8678 28122 8730
rect 45808 8678 45860 8730
rect 45872 8678 45924 8730
rect 45936 8678 45988 8730
rect 46000 8678 46052 8730
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 7472 8576 7524 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 18236 8576 18288 8628
rect 19984 8576 20036 8628
rect 26608 8576 26660 8628
rect 27160 8619 27212 8628
rect 27160 8585 27169 8619
rect 27169 8585 27203 8619
rect 27203 8585 27212 8619
rect 27160 8576 27212 8585
rect 30564 8619 30616 8628
rect 30564 8585 30573 8619
rect 30573 8585 30607 8619
rect 30607 8585 30616 8619
rect 30564 8576 30616 8585
rect 31760 8619 31812 8628
rect 31760 8585 31769 8619
rect 31769 8585 31803 8619
rect 31803 8585 31812 8619
rect 32772 8619 32824 8628
rect 31760 8576 31812 8585
rect 32772 8585 32781 8619
rect 32781 8585 32815 8619
rect 32815 8585 32824 8619
rect 32772 8576 32824 8585
rect 35808 8576 35860 8628
rect 37648 8619 37700 8628
rect 37648 8585 37657 8619
rect 37657 8585 37691 8619
rect 37691 8585 37700 8619
rect 37648 8576 37700 8585
rect 6276 8508 6328 8560
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 5540 8372 5592 8424
rect 8760 8508 8812 8560
rect 11520 8508 11572 8560
rect 13728 8508 13780 8560
rect 17224 8508 17276 8560
rect 11428 8440 11480 8492
rect 20720 8508 20772 8560
rect 26332 8508 26384 8560
rect 29736 8508 29788 8560
rect 34520 8508 34572 8560
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 7748 8415 7800 8424
rect 7748 8381 7757 8415
rect 7757 8381 7791 8415
rect 7791 8381 7800 8415
rect 7748 8372 7800 8381
rect 8300 8372 8352 8424
rect 11612 8372 11664 8424
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 15384 8415 15436 8424
rect 15384 8381 15393 8415
rect 15393 8381 15427 8415
rect 15427 8381 15436 8415
rect 15384 8372 15436 8381
rect 18972 8415 19024 8424
rect 18972 8381 18981 8415
rect 18981 8381 19015 8415
rect 19015 8381 19024 8415
rect 18972 8372 19024 8381
rect 19984 8415 20036 8424
rect 19984 8381 19993 8415
rect 19993 8381 20027 8415
rect 20027 8381 20036 8415
rect 19984 8372 20036 8381
rect 20628 8372 20680 8424
rect 22008 8415 22060 8424
rect 22008 8381 22017 8415
rect 22017 8381 22051 8415
rect 22051 8381 22060 8415
rect 22008 8372 22060 8381
rect 23020 8415 23072 8424
rect 23020 8381 23029 8415
rect 23029 8381 23063 8415
rect 23063 8381 23072 8415
rect 23020 8372 23072 8381
rect 26240 8440 26292 8492
rect 35992 8440 36044 8492
rect 26148 8372 26200 8424
rect 27344 8415 27396 8424
rect 27344 8381 27353 8415
rect 27353 8381 27387 8415
rect 27387 8381 27396 8415
rect 27344 8372 27396 8381
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 30748 8415 30800 8424
rect 30748 8381 30757 8415
rect 30757 8381 30791 8415
rect 30791 8381 30800 8415
rect 30748 8372 30800 8381
rect 31208 8372 31260 8424
rect 32956 8415 33008 8424
rect 32956 8381 32965 8415
rect 32965 8381 32999 8415
rect 32999 8381 33008 8415
rect 32956 8372 33008 8381
rect 33968 8415 34020 8424
rect 33968 8381 33977 8415
rect 33977 8381 34011 8415
rect 34011 8381 34020 8415
rect 33968 8372 34020 8381
rect 34612 8372 34664 8424
rect 36728 8372 36780 8424
rect 11428 8304 11480 8356
rect 10784 8236 10836 8288
rect 18788 8279 18840 8288
rect 18788 8245 18797 8279
rect 18797 8245 18831 8279
rect 18831 8245 18840 8279
rect 18788 8236 18840 8245
rect 23296 8236 23348 8288
rect 34980 8236 35032 8288
rect 18912 8134 18964 8186
rect 18976 8134 19028 8186
rect 19040 8134 19092 8186
rect 19104 8134 19156 8186
rect 36843 8134 36895 8186
rect 36907 8134 36959 8186
rect 36971 8134 37023 8186
rect 37035 8134 37087 8186
rect 3056 8032 3108 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 8668 8032 8720 8084
rect 11428 8075 11480 8084
rect 11428 8041 11437 8075
rect 11437 8041 11471 8075
rect 11471 8041 11480 8075
rect 11428 8032 11480 8041
rect 11612 8032 11664 8084
rect 14372 8032 14424 8084
rect 19984 8032 20036 8084
rect 22376 8032 22428 8084
rect 23112 8075 23164 8084
rect 23112 8041 23121 8075
rect 23121 8041 23155 8075
rect 23155 8041 23164 8075
rect 23112 8032 23164 8041
rect 24124 8075 24176 8084
rect 24124 8041 24133 8075
rect 24133 8041 24167 8075
rect 24167 8041 24176 8075
rect 24124 8032 24176 8041
rect 25228 8032 25280 8084
rect 27344 8032 27396 8084
rect 28356 8032 28408 8084
rect 29552 8075 29604 8084
rect 29552 8041 29561 8075
rect 29561 8041 29595 8075
rect 29595 8041 29604 8075
rect 29552 8032 29604 8041
rect 35348 8032 35400 8084
rect 3240 7896 3292 7948
rect 3516 7896 3568 7948
rect 5724 7939 5776 7948
rect 5724 7905 5733 7939
rect 5733 7905 5767 7939
rect 5767 7905 5776 7939
rect 5724 7896 5776 7905
rect 7656 7896 7708 7948
rect 8392 7896 8444 7948
rect 9680 7896 9732 7948
rect 11520 7896 11572 7948
rect 11704 7896 11756 7948
rect 13820 7896 13872 7948
rect 16212 7939 16264 7948
rect 16212 7905 16221 7939
rect 16221 7905 16255 7939
rect 16255 7905 16264 7939
rect 16212 7896 16264 7905
rect 17224 7939 17276 7948
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 19708 7896 19760 7948
rect 21824 7939 21876 7948
rect 21824 7905 21833 7939
rect 21833 7905 21867 7939
rect 21867 7905 21876 7939
rect 21824 7896 21876 7905
rect 23296 7939 23348 7948
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 24032 7896 24084 7948
rect 29000 7964 29052 8016
rect 26332 7939 26384 7948
rect 26332 7905 26341 7939
rect 26341 7905 26375 7939
rect 26375 7905 26384 7939
rect 26332 7896 26384 7905
rect 27344 7896 27396 7948
rect 28724 7939 28776 7948
rect 28724 7905 28733 7939
rect 28733 7905 28767 7939
rect 28767 7905 28776 7939
rect 28724 7896 28776 7905
rect 30012 7896 30064 7948
rect 34520 7896 34572 7948
rect 34980 7939 35032 7948
rect 34980 7905 34989 7939
rect 34989 7905 35023 7939
rect 35023 7905 35032 7939
rect 34980 7896 35032 7905
rect 35072 7896 35124 7948
rect 36084 7896 36136 7948
rect 17960 7828 18012 7880
rect 5540 7692 5592 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 8760 7692 8812 7744
rect 16396 7692 16448 7744
rect 18236 7692 18288 7744
rect 19984 7692 20036 7744
rect 27528 7692 27580 7744
rect 34520 7692 34572 7744
rect 35808 7735 35860 7744
rect 35808 7701 35817 7735
rect 35817 7701 35851 7735
rect 35851 7701 35860 7735
rect 35808 7692 35860 7701
rect 35900 7692 35952 7744
rect 9947 7590 9999 7642
rect 10011 7590 10063 7642
rect 10075 7590 10127 7642
rect 10139 7590 10191 7642
rect 27878 7590 27930 7642
rect 27942 7590 27994 7642
rect 28006 7590 28058 7642
rect 28070 7590 28122 7642
rect 45808 7590 45860 7642
rect 45872 7590 45924 7642
rect 45936 7590 45988 7642
rect 46000 7590 46052 7642
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 8300 7488 8352 7540
rect 18052 7488 18104 7540
rect 19708 7488 19760 7540
rect 23020 7488 23072 7540
rect 27344 7531 27396 7540
rect 27344 7497 27353 7531
rect 27353 7497 27387 7531
rect 27387 7497 27396 7531
rect 27344 7488 27396 7497
rect 30012 7531 30064 7540
rect 30012 7497 30021 7531
rect 30021 7497 30055 7531
rect 30055 7497 30064 7531
rect 30012 7488 30064 7497
rect 32864 7488 32916 7540
rect 34612 7488 34664 7540
rect 23848 7420 23900 7472
rect 4712 7327 4764 7336
rect 4712 7293 4721 7327
rect 4721 7293 4755 7327
rect 4755 7293 4764 7327
rect 4712 7284 4764 7293
rect 5908 7327 5960 7336
rect 5908 7293 5917 7327
rect 5917 7293 5951 7327
rect 5951 7293 5960 7327
rect 5908 7284 5960 7293
rect 6552 7284 6604 7336
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 8944 7284 8996 7336
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 14648 7352 14700 7404
rect 13544 7284 13596 7336
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 16396 7327 16448 7336
rect 16396 7293 16405 7327
rect 16405 7293 16439 7327
rect 16439 7293 16448 7327
rect 16396 7284 16448 7293
rect 18788 7284 18840 7336
rect 18880 7284 18932 7336
rect 19984 7327 20036 7336
rect 19984 7293 19993 7327
rect 19993 7293 20027 7327
rect 20027 7293 20036 7327
rect 19984 7284 20036 7293
rect 20996 7327 21048 7336
rect 20996 7293 21005 7327
rect 21005 7293 21039 7327
rect 21039 7293 21048 7327
rect 20996 7284 21048 7293
rect 22744 7327 22796 7336
rect 22744 7293 22753 7327
rect 22753 7293 22787 7327
rect 22787 7293 22796 7327
rect 22744 7284 22796 7293
rect 24584 7327 24636 7336
rect 24584 7293 24593 7327
rect 24593 7293 24627 7327
rect 24627 7293 24636 7327
rect 24584 7284 24636 7293
rect 25044 7284 25096 7336
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 30196 7327 30248 7336
rect 30196 7293 30205 7327
rect 30205 7293 30239 7327
rect 30239 7293 30248 7327
rect 30196 7284 30248 7293
rect 32312 7284 32364 7336
rect 35164 7284 35216 7336
rect 35808 7327 35860 7336
rect 35808 7293 35817 7327
rect 35817 7293 35851 7327
rect 35851 7293 35860 7327
rect 35808 7284 35860 7293
rect 36176 7284 36228 7336
rect 38016 7327 38068 7336
rect 38016 7293 38025 7327
rect 38025 7293 38059 7327
rect 38059 7293 38068 7327
rect 38016 7284 38068 7293
rect 4804 7216 4856 7268
rect 5816 7148 5868 7200
rect 8300 7148 8352 7200
rect 8668 7148 8720 7200
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 10600 7148 10652 7157
rect 14372 7148 14424 7200
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 15292 7148 15344 7200
rect 18696 7148 18748 7200
rect 19340 7148 19392 7200
rect 20260 7148 20312 7200
rect 22652 7148 22704 7200
rect 35808 7148 35860 7200
rect 35992 7148 36044 7200
rect 39856 7148 39908 7200
rect 18912 7046 18964 7098
rect 18976 7046 19028 7098
rect 19040 7046 19092 7098
rect 19104 7046 19156 7098
rect 36843 7046 36895 7098
rect 36907 7046 36959 7098
rect 36971 7046 37023 7098
rect 37035 7046 37087 7098
rect 5908 6944 5960 6996
rect 16212 6944 16264 6996
rect 20996 6944 21048 6996
rect 22744 6987 22796 6996
rect 22744 6953 22753 6987
rect 22753 6953 22787 6987
rect 22787 6953 22796 6987
rect 22744 6944 22796 6953
rect 24584 6944 24636 6996
rect 30196 6944 30248 6996
rect 3792 6808 3844 6860
rect 5632 6808 5684 6860
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 8300 6808 8352 6860
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 11152 6808 11204 6860
rect 8392 6672 8444 6724
rect 9680 6672 9732 6724
rect 12716 6672 12768 6724
rect 13452 6808 13504 6860
rect 16212 6851 16264 6860
rect 16212 6817 16221 6851
rect 16221 6817 16255 6851
rect 16255 6817 16264 6851
rect 16212 6808 16264 6817
rect 16304 6808 16356 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 16580 6740 16632 6792
rect 20076 6808 20128 6860
rect 18696 6740 18748 6792
rect 22560 6808 22612 6860
rect 23756 6808 23808 6860
rect 24860 6808 24912 6860
rect 23480 6740 23532 6792
rect 26424 6808 26476 6860
rect 29736 6851 29788 6860
rect 29736 6817 29745 6851
rect 29745 6817 29779 6851
rect 29779 6817 29788 6851
rect 29736 6808 29788 6817
rect 34520 6876 34572 6928
rect 35808 6851 35860 6860
rect 35808 6817 35817 6851
rect 35817 6817 35851 6851
rect 35851 6817 35860 6851
rect 35808 6808 35860 6817
rect 36268 6808 36320 6860
rect 38660 6851 38712 6860
rect 38660 6817 38669 6851
rect 38669 6817 38703 6851
rect 38703 6817 38712 6851
rect 38660 6808 38712 6817
rect 40500 6808 40552 6860
rect 26976 6740 27028 6792
rect 34428 6740 34480 6792
rect 34612 6740 34664 6792
rect 51080 6740 51132 6792
rect 18420 6672 18472 6724
rect 36084 6672 36136 6724
rect 38016 6672 38068 6724
rect 3332 6604 3384 6656
rect 4896 6604 4948 6656
rect 8576 6604 8628 6656
rect 10508 6604 10560 6656
rect 12624 6604 12676 6656
rect 16396 6604 16448 6656
rect 17408 6604 17460 6656
rect 18144 6604 18196 6656
rect 20996 6604 21048 6656
rect 22744 6604 22796 6656
rect 24860 6604 24912 6656
rect 27620 6604 27672 6656
rect 33968 6604 34020 6656
rect 38844 6604 38896 6656
rect 38936 6604 38988 6656
rect 9947 6502 9999 6554
rect 10011 6502 10063 6554
rect 10075 6502 10127 6554
rect 10139 6502 10191 6554
rect 27878 6502 27930 6554
rect 27942 6502 27994 6554
rect 28006 6502 28058 6554
rect 28070 6502 28122 6554
rect 45808 6502 45860 6554
rect 45872 6502 45924 6554
rect 45936 6502 45988 6554
rect 46000 6502 46052 6554
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 5632 6400 5684 6452
rect 8944 6400 8996 6452
rect 11336 6400 11388 6452
rect 15384 6400 15436 6452
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 22560 6443 22612 6452
rect 22560 6409 22569 6443
rect 22569 6409 22603 6443
rect 22603 6409 22612 6443
rect 22560 6400 22612 6409
rect 22836 6400 22888 6452
rect 29368 6400 29420 6452
rect 35072 6400 35124 6452
rect 36176 6400 36228 6452
rect 38660 6400 38712 6452
rect 5356 6332 5408 6384
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 3332 6196 3384 6248
rect 4896 6239 4948 6248
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 5540 6196 5592 6248
rect 8576 6196 8628 6248
rect 10416 6332 10468 6384
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 11060 6196 11112 6248
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 14464 6196 14516 6248
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 18052 6196 18104 6248
rect 19340 6196 19392 6248
rect 20996 6239 21048 6248
rect 20996 6205 21005 6239
rect 21005 6205 21039 6239
rect 21039 6205 21048 6239
rect 20996 6196 21048 6205
rect 22744 6239 22796 6248
rect 22744 6205 22753 6239
rect 22753 6205 22787 6239
rect 22787 6205 22796 6239
rect 22744 6196 22796 6205
rect 25596 6239 25648 6248
rect 25596 6205 25605 6239
rect 25605 6205 25639 6239
rect 25639 6205 25648 6239
rect 25596 6196 25648 6205
rect 25688 6196 25740 6248
rect 27620 6239 27672 6248
rect 27620 6205 27629 6239
rect 27629 6205 27663 6239
rect 27663 6205 27672 6239
rect 27620 6196 27672 6205
rect 30196 6239 30248 6248
rect 30196 6205 30205 6239
rect 30205 6205 30239 6239
rect 30239 6205 30248 6239
rect 30196 6196 30248 6205
rect 33968 6239 34020 6248
rect 33968 6205 33977 6239
rect 33977 6205 34011 6239
rect 34011 6205 34020 6239
rect 33968 6196 34020 6205
rect 35900 6196 35952 6248
rect 34336 6128 34388 6180
rect 37188 6196 37240 6248
rect 38936 6239 38988 6248
rect 38936 6205 38945 6239
rect 38945 6205 38979 6239
rect 38979 6205 38988 6239
rect 38936 6196 38988 6205
rect 38568 6128 38620 6180
rect 4988 6060 5040 6112
rect 9772 6060 9824 6112
rect 10324 6060 10376 6112
rect 11612 6060 11664 6112
rect 13636 6060 13688 6112
rect 16212 6060 16264 6112
rect 17408 6060 17460 6112
rect 19248 6060 19300 6112
rect 19892 6060 19944 6112
rect 20996 6060 21048 6112
rect 25872 6060 25924 6112
rect 26516 6060 26568 6112
rect 29828 6060 29880 6112
rect 31484 6060 31536 6112
rect 37280 6060 37332 6112
rect 40040 6060 40092 6112
rect 18912 5958 18964 6010
rect 18976 5958 19028 6010
rect 19040 5958 19092 6010
rect 19104 5958 19156 6010
rect 36843 5958 36895 6010
rect 36907 5958 36959 6010
rect 36971 5958 37023 6010
rect 37035 5958 37087 6010
rect 2320 5856 2372 5908
rect 2872 5856 2924 5908
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 13452 5899 13504 5908
rect 13452 5865 13461 5899
rect 13461 5865 13495 5899
rect 13495 5865 13504 5899
rect 13452 5856 13504 5865
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 16304 5856 16356 5908
rect 17224 5856 17276 5908
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 20076 5899 20128 5908
rect 20076 5865 20085 5899
rect 20085 5865 20119 5899
rect 20119 5865 20128 5899
rect 20076 5856 20128 5865
rect 22468 5856 22520 5908
rect 22744 5856 22796 5908
rect 5540 5788 5592 5840
rect 2320 5763 2372 5772
rect 2320 5729 2329 5763
rect 2329 5729 2363 5763
rect 2363 5729 2372 5763
rect 2320 5720 2372 5729
rect 4988 5763 5040 5772
rect 4988 5729 4997 5763
rect 4997 5729 5031 5763
rect 5031 5729 5040 5763
rect 4988 5720 5040 5729
rect 3792 5652 3844 5704
rect 4804 5627 4856 5636
rect 4804 5593 4813 5627
rect 4813 5593 4847 5627
rect 4847 5593 4856 5627
rect 4804 5584 4856 5593
rect 6920 5720 6972 5772
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 12624 5763 12676 5772
rect 12624 5729 12633 5763
rect 12633 5729 12667 5763
rect 12667 5729 12676 5763
rect 12624 5720 12676 5729
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 15292 5720 15344 5772
rect 16212 5763 16264 5772
rect 16212 5729 16221 5763
rect 16221 5729 16255 5763
rect 16255 5729 16264 5763
rect 16212 5720 16264 5729
rect 18144 5720 18196 5772
rect 19248 5763 19300 5772
rect 6920 5584 6972 5636
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 22652 5720 22704 5772
rect 24400 5856 24452 5908
rect 25596 5856 25648 5908
rect 36268 5856 36320 5908
rect 37188 5856 37240 5908
rect 40500 5899 40552 5908
rect 40500 5865 40509 5899
rect 40509 5865 40543 5899
rect 40543 5865 40552 5899
rect 40500 5856 40552 5865
rect 23848 5763 23900 5772
rect 23848 5729 23865 5763
rect 23865 5729 23899 5763
rect 23899 5729 23900 5763
rect 24860 5763 24912 5772
rect 23848 5720 23900 5729
rect 24860 5729 24869 5763
rect 24869 5729 24903 5763
rect 24903 5729 24912 5763
rect 24860 5720 24912 5729
rect 25872 5763 25924 5772
rect 25872 5729 25881 5763
rect 25881 5729 25915 5763
rect 25915 5729 25924 5763
rect 25872 5720 25924 5729
rect 24768 5652 24820 5704
rect 29092 5720 29144 5772
rect 30472 5763 30524 5772
rect 30472 5729 30481 5763
rect 30481 5729 30515 5763
rect 30515 5729 30524 5763
rect 30472 5720 30524 5729
rect 35992 5720 36044 5772
rect 37372 5720 37424 5772
rect 39856 5788 39908 5840
rect 40592 5720 40644 5772
rect 22928 5584 22980 5636
rect 11428 5559 11480 5568
rect 11428 5525 11437 5559
rect 11437 5525 11471 5559
rect 11471 5525 11480 5559
rect 11428 5516 11480 5525
rect 12440 5559 12492 5568
rect 12440 5525 12449 5559
rect 12449 5525 12483 5559
rect 12483 5525 12492 5559
rect 23664 5559 23716 5568
rect 12440 5516 12492 5525
rect 23664 5525 23673 5559
rect 23673 5525 23707 5559
rect 23707 5525 23716 5559
rect 23664 5516 23716 5525
rect 23848 5584 23900 5636
rect 26608 5516 26660 5568
rect 27344 5516 27396 5568
rect 29276 5559 29328 5568
rect 29276 5525 29285 5559
rect 29285 5525 29319 5559
rect 29319 5525 29328 5559
rect 29276 5516 29328 5525
rect 34520 5516 34572 5568
rect 37556 5516 37608 5568
rect 9947 5414 9999 5466
rect 10011 5414 10063 5466
rect 10075 5414 10127 5466
rect 10139 5414 10191 5466
rect 27878 5414 27930 5466
rect 27942 5414 27994 5466
rect 28006 5414 28058 5466
rect 28070 5414 28122 5466
rect 45808 5414 45860 5466
rect 45872 5414 45924 5466
rect 45936 5414 45988 5466
rect 46000 5414 46052 5466
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 5540 5312 5592 5364
rect 9036 5312 9088 5364
rect 11060 5312 11112 5364
rect 13360 5312 13412 5364
rect 16580 5312 16632 5364
rect 18788 5355 18840 5364
rect 18788 5321 18797 5355
rect 18797 5321 18831 5355
rect 18831 5321 18840 5355
rect 18788 5312 18840 5321
rect 21824 5312 21876 5364
rect 25688 5312 25740 5364
rect 37372 5312 37424 5364
rect 38568 5312 38620 5364
rect 13544 5244 13596 5296
rect 20812 5244 20864 5296
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 6368 5108 6420 5160
rect 10508 5176 10560 5228
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 11428 5108 11480 5160
rect 12440 5108 12492 5160
rect 15200 5176 15252 5228
rect 33508 5244 33560 5296
rect 14096 5108 14148 5160
rect 17408 5108 17460 5160
rect 19892 5108 19944 5160
rect 22284 5151 22336 5160
rect 6460 5040 6512 5092
rect 22284 5117 22293 5151
rect 22293 5117 22327 5151
rect 22327 5117 22336 5151
rect 22284 5108 22336 5117
rect 5540 4972 5592 5024
rect 7656 4972 7708 5024
rect 22192 5040 22244 5092
rect 23388 5108 23440 5160
rect 24952 5108 25004 5160
rect 26608 5151 26660 5160
rect 26608 5117 26617 5151
rect 26617 5117 26651 5151
rect 26651 5117 26660 5151
rect 26608 5108 26660 5117
rect 29276 5176 29328 5228
rect 29828 5176 29880 5228
rect 27712 5108 27764 5160
rect 29184 5108 29236 5160
rect 37280 5108 37332 5160
rect 37556 5151 37608 5160
rect 37556 5117 37565 5151
rect 37565 5117 37599 5151
rect 37599 5117 37608 5151
rect 37556 5108 37608 5117
rect 38752 5108 38804 5160
rect 40040 5108 40092 5160
rect 21824 4972 21876 5024
rect 24492 4972 24544 5024
rect 25504 4972 25556 5024
rect 26608 4972 26660 5024
rect 27528 4972 27580 5024
rect 30380 4972 30432 5024
rect 37556 4972 37608 5024
rect 39396 5015 39448 5024
rect 39396 4981 39405 5015
rect 39405 4981 39439 5015
rect 39439 4981 39448 5015
rect 39396 4972 39448 4981
rect 18912 4870 18964 4922
rect 18976 4870 19028 4922
rect 19040 4870 19092 4922
rect 19104 4870 19156 4922
rect 36843 4870 36895 4922
rect 36907 4870 36959 4922
rect 36971 4870 37023 4922
rect 37035 4870 37087 4922
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 10600 4768 10652 4820
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 18328 4768 18380 4820
rect 22284 4768 22336 4820
rect 23480 4768 23532 4820
rect 24952 4811 25004 4820
rect 24952 4777 24961 4811
rect 24961 4777 24995 4811
rect 24995 4777 25004 4811
rect 24952 4768 25004 4777
rect 30472 4768 30524 4820
rect 38752 4811 38804 4820
rect 38752 4777 38761 4811
rect 38761 4777 38795 4811
rect 38795 4777 38804 4811
rect 38752 4768 38804 4777
rect 40592 4768 40644 4820
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 6920 4632 6972 4684
rect 7656 4632 7708 4684
rect 10324 4632 10376 4684
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 14280 4675 14332 4684
rect 14280 4641 14289 4675
rect 14289 4641 14323 4675
rect 14323 4641 14332 4675
rect 14280 4632 14332 4641
rect 19064 4675 19116 4684
rect 19064 4641 19073 4675
rect 19073 4641 19107 4675
rect 19107 4641 19116 4675
rect 19064 4632 19116 4641
rect 23664 4700 23716 4752
rect 21824 4675 21876 4684
rect 21824 4641 21833 4675
rect 21833 4641 21867 4675
rect 21867 4641 21876 4675
rect 21824 4632 21876 4641
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 24492 4632 24544 4684
rect 26516 4700 26568 4752
rect 38844 4700 38896 4752
rect 27344 4632 27396 4684
rect 27528 4632 27580 4684
rect 6828 4496 6880 4548
rect 11152 4496 11204 4548
rect 18604 4496 18656 4548
rect 26332 4564 26384 4616
rect 29000 4632 29052 4684
rect 30472 4675 30524 4684
rect 30472 4641 30481 4675
rect 30481 4641 30515 4675
rect 30515 4641 30524 4675
rect 30472 4632 30524 4641
rect 31484 4675 31536 4684
rect 31484 4641 31493 4675
rect 31493 4641 31527 4675
rect 31527 4641 31536 4675
rect 31484 4632 31536 4641
rect 33048 4675 33100 4684
rect 33048 4641 33057 4675
rect 33057 4641 33091 4675
rect 33091 4641 33100 4675
rect 33048 4632 33100 4641
rect 36176 4632 36228 4684
rect 37556 4675 37608 4684
rect 37556 4641 37565 4675
rect 37565 4641 37599 4675
rect 37599 4641 37608 4675
rect 37556 4632 37608 4641
rect 40684 4632 40736 4684
rect 14188 4428 14240 4480
rect 20812 4428 20864 4480
rect 22744 4428 22796 4480
rect 25596 4428 25648 4480
rect 26240 4428 26292 4480
rect 27620 4428 27672 4480
rect 28356 4428 28408 4480
rect 29460 4428 29512 4480
rect 34060 4428 34112 4480
rect 36544 4428 36596 4480
rect 40592 4428 40644 4480
rect 9947 4326 9999 4378
rect 10011 4326 10063 4378
rect 10075 4326 10127 4378
rect 10139 4326 10191 4378
rect 27878 4326 27930 4378
rect 27942 4326 27994 4378
rect 28006 4326 28058 4378
rect 28070 4326 28122 4378
rect 45808 4326 45860 4378
rect 45872 4326 45924 4378
rect 45936 4326 45988 4378
rect 46000 4326 46052 4378
rect 6460 4267 6512 4276
rect 6460 4233 6469 4267
rect 6469 4233 6503 4267
rect 6503 4233 6512 4267
rect 6460 4224 6512 4233
rect 13268 4224 13320 4276
rect 14280 4224 14332 4276
rect 19064 4224 19116 4276
rect 22836 4224 22888 4276
rect 33048 4224 33100 4276
rect 2320 4156 2372 4208
rect 6276 4020 6328 4072
rect 8208 4020 8260 4072
rect 13728 4020 13780 4072
rect 14004 4020 14056 4072
rect 16580 4063 16632 4072
rect 14740 3884 14792 3936
rect 16580 4029 16589 4063
rect 16589 4029 16623 4063
rect 16623 4029 16632 4063
rect 16580 4020 16632 4029
rect 18512 4020 18564 4072
rect 20812 4020 20864 4072
rect 20996 4063 21048 4072
rect 20996 4029 21005 4063
rect 21005 4029 21039 4063
rect 21039 4029 21048 4063
rect 20996 4020 21048 4029
rect 23848 4020 23900 4072
rect 25504 4088 25556 4140
rect 25596 4063 25648 4072
rect 25596 4029 25605 4063
rect 25605 4029 25639 4063
rect 25639 4029 25648 4063
rect 25596 4020 25648 4029
rect 26608 4063 26660 4072
rect 26608 4029 26617 4063
rect 26617 4029 26651 4063
rect 26651 4029 26660 4063
rect 26608 4020 26660 4029
rect 27620 4063 27672 4072
rect 27620 4029 27629 4063
rect 27629 4029 27663 4063
rect 27663 4029 27672 4063
rect 27620 4020 27672 4029
rect 28264 4020 28316 4072
rect 31852 4063 31904 4072
rect 19800 3927 19852 3936
rect 19800 3893 19809 3927
rect 19809 3893 19843 3927
rect 19843 3893 19852 3927
rect 19800 3884 19852 3893
rect 22192 3952 22244 4004
rect 31852 4029 31861 4063
rect 31861 4029 31895 4063
rect 31895 4029 31904 4063
rect 31852 4020 31904 4029
rect 33692 4020 33744 4072
rect 33876 4063 33928 4072
rect 33876 4029 33885 4063
rect 33885 4029 33919 4063
rect 33919 4029 33928 4063
rect 33876 4020 33928 4029
rect 35624 4020 35676 4072
rect 36728 4020 36780 4072
rect 39396 4020 39448 4072
rect 40408 4020 40460 4072
rect 40592 4020 40644 4072
rect 21916 3884 21968 3936
rect 33048 3952 33100 4004
rect 24492 3884 24544 3936
rect 25504 3884 25556 3936
rect 27712 3884 27764 3936
rect 29000 3884 29052 3936
rect 31300 3884 31352 3936
rect 31668 3927 31720 3936
rect 31668 3893 31677 3927
rect 31677 3893 31711 3927
rect 31711 3893 31720 3927
rect 31668 3884 31720 3893
rect 34244 3884 34296 3936
rect 36084 3884 36136 3936
rect 36636 3927 36688 3936
rect 36636 3893 36645 3927
rect 36645 3893 36679 3927
rect 36679 3893 36688 3927
rect 36636 3884 36688 3893
rect 38384 3927 38436 3936
rect 38384 3893 38393 3927
rect 38393 3893 38427 3927
rect 38427 3893 38436 3927
rect 38384 3884 38436 3893
rect 40316 3884 40368 3936
rect 42432 3884 42484 3936
rect 18912 3782 18964 3834
rect 18976 3782 19028 3834
rect 19040 3782 19092 3834
rect 19104 3782 19156 3834
rect 36843 3782 36895 3834
rect 36907 3782 36959 3834
rect 36971 3782 37023 3834
rect 37035 3782 37087 3834
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 16580 3680 16632 3732
rect 23388 3680 23440 3732
rect 24768 3723 24820 3732
rect 24768 3689 24777 3723
rect 24777 3689 24811 3723
rect 24811 3689 24820 3723
rect 24768 3680 24820 3689
rect 28264 3723 28316 3732
rect 28264 3689 28273 3723
rect 28273 3689 28307 3723
rect 28307 3689 28316 3723
rect 28264 3680 28316 3689
rect 33876 3680 33928 3732
rect 40684 3680 40736 3732
rect 14188 3587 14240 3596
rect 14188 3553 14197 3587
rect 14197 3553 14231 3587
rect 14231 3553 14240 3587
rect 14188 3544 14240 3553
rect 19432 3612 19484 3664
rect 19800 3544 19852 3596
rect 22744 3544 22796 3596
rect 25044 3612 25096 3664
rect 38384 3612 38436 3664
rect 22928 3408 22980 3460
rect 24492 3544 24544 3596
rect 25504 3544 25556 3596
rect 26240 3544 26292 3596
rect 26792 3544 26844 3596
rect 28448 3587 28500 3596
rect 28448 3553 28457 3587
rect 28457 3553 28491 3587
rect 28491 3553 28500 3587
rect 28448 3544 28500 3553
rect 29460 3587 29512 3596
rect 29460 3553 29469 3587
rect 29469 3553 29503 3587
rect 29503 3553 29512 3587
rect 29460 3544 29512 3553
rect 30564 3587 30616 3596
rect 30564 3553 30573 3587
rect 30573 3553 30607 3587
rect 30607 3553 30616 3587
rect 30564 3544 30616 3553
rect 31668 3544 31720 3596
rect 34060 3587 34112 3596
rect 34060 3553 34069 3587
rect 34069 3553 34103 3587
rect 34103 3553 34112 3587
rect 34060 3544 34112 3553
rect 35072 3587 35124 3596
rect 35072 3553 35081 3587
rect 35081 3553 35115 3587
rect 35115 3553 35124 3587
rect 35072 3544 35124 3553
rect 36084 3587 36136 3596
rect 36084 3553 36093 3587
rect 36093 3553 36127 3587
rect 36127 3553 36136 3587
rect 36084 3544 36136 3553
rect 36636 3544 36688 3596
rect 38660 3587 38712 3596
rect 38660 3553 38669 3587
rect 38669 3553 38703 3587
rect 38703 3553 38712 3587
rect 38660 3544 38712 3553
rect 40592 3544 40644 3596
rect 41236 3544 41288 3596
rect 42248 3544 42300 3596
rect 31852 3408 31904 3460
rect 24952 3340 25004 3392
rect 25964 3340 26016 3392
rect 29276 3383 29328 3392
rect 29276 3349 29285 3383
rect 29285 3349 29319 3383
rect 29319 3349 29328 3383
rect 29276 3340 29328 3349
rect 31208 3340 31260 3392
rect 33232 3340 33284 3392
rect 33692 3408 33744 3460
rect 43076 3408 43128 3460
rect 35992 3340 36044 3392
rect 39212 3340 39264 3392
rect 40224 3340 40276 3392
rect 41420 3340 41472 3392
rect 9947 3238 9999 3290
rect 10011 3238 10063 3290
rect 10075 3238 10127 3290
rect 10139 3238 10191 3290
rect 27878 3238 27930 3290
rect 27942 3238 27994 3290
rect 28006 3238 28058 3290
rect 28070 3238 28122 3290
rect 45808 3238 45860 3290
rect 45872 3238 45924 3290
rect 45936 3238 45988 3290
rect 46000 3238 46052 3290
rect 22836 3068 22888 3120
rect 26332 3136 26384 3188
rect 26792 3179 26844 3188
rect 26792 3145 26801 3179
rect 26801 3145 26835 3179
rect 26835 3145 26844 3179
rect 26792 3136 26844 3145
rect 30564 3136 30616 3188
rect 33048 3179 33100 3188
rect 33048 3145 33057 3179
rect 33057 3145 33091 3179
rect 33091 3145 33100 3179
rect 33048 3136 33100 3145
rect 35072 3136 35124 3188
rect 35624 3179 35676 3188
rect 35624 3145 35633 3179
rect 35633 3145 35667 3179
rect 35667 3145 35676 3179
rect 35624 3136 35676 3145
rect 36728 3136 36780 3188
rect 38660 3136 38712 3188
rect 41236 3179 41288 3188
rect 41236 3145 41245 3179
rect 41245 3145 41279 3179
rect 41279 3145 41288 3179
rect 41236 3136 41288 3145
rect 42248 3179 42300 3188
rect 42248 3145 42257 3179
rect 42257 3145 42291 3179
rect 42291 3145 42300 3179
rect 42248 3136 42300 3145
rect 29092 3068 29144 3120
rect 26424 3000 26476 3052
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 21916 2975 21968 2984
rect 21916 2941 21925 2975
rect 21925 2941 21959 2975
rect 21959 2941 21968 2975
rect 21916 2932 21968 2941
rect 22928 2975 22980 2984
rect 22928 2941 22937 2975
rect 22937 2941 22971 2975
rect 22971 2941 22980 2975
rect 22928 2932 22980 2941
rect 24952 2975 25004 2984
rect 24952 2941 24961 2975
rect 24961 2941 24995 2975
rect 24995 2941 25004 2975
rect 24952 2932 25004 2941
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 28356 3000 28408 3052
rect 29276 2932 29328 2984
rect 31024 2932 31076 2984
rect 31208 2975 31260 2984
rect 31208 2941 31217 2975
rect 31217 2941 31251 2975
rect 31251 2941 31260 2975
rect 31208 2932 31260 2941
rect 31300 2932 31352 2984
rect 33232 2975 33284 2984
rect 33232 2941 33241 2975
rect 33241 2941 33275 2975
rect 33275 2941 33284 2975
rect 33232 2932 33284 2941
rect 34244 2975 34296 2984
rect 34244 2941 34253 2975
rect 34253 2941 34287 2975
rect 34287 2941 34296 2975
rect 34244 2932 34296 2941
rect 35992 2932 36044 2984
rect 36544 2932 36596 2984
rect 37832 2975 37884 2984
rect 37832 2941 37841 2975
rect 37841 2941 37875 2975
rect 37875 2941 37884 2975
rect 37832 2932 37884 2941
rect 38844 2975 38896 2984
rect 38844 2941 38853 2975
rect 38853 2941 38887 2975
rect 38887 2941 38896 2975
rect 38844 2932 38896 2941
rect 40040 2932 40092 2984
rect 40316 2932 40368 2984
rect 42432 2975 42484 2984
rect 42432 2941 42441 2975
rect 42441 2941 42475 2975
rect 42475 2941 42484 2975
rect 42432 2932 42484 2941
rect 23848 2796 23900 2848
rect 27804 2839 27856 2848
rect 27804 2805 27813 2839
rect 27813 2805 27847 2839
rect 27847 2805 27856 2839
rect 27804 2796 27856 2805
rect 30656 2796 30708 2848
rect 31668 2796 31720 2848
rect 37280 2796 37332 2848
rect 38660 2839 38712 2848
rect 38660 2805 38669 2839
rect 38669 2805 38703 2839
rect 38703 2805 38712 2839
rect 38660 2796 38712 2805
rect 18912 2694 18964 2746
rect 18976 2694 19028 2746
rect 19040 2694 19092 2746
rect 19104 2694 19156 2746
rect 36843 2694 36895 2746
rect 36907 2694 36959 2746
rect 36971 2694 37023 2746
rect 37035 2694 37087 2746
rect 20904 2592 20956 2644
rect 22928 2592 22980 2644
rect 28448 2592 28500 2644
rect 30196 2592 30248 2644
rect 23480 2524 23532 2576
rect 22836 2499 22888 2508
rect 19800 2295 19852 2304
rect 19800 2261 19809 2295
rect 19809 2261 19843 2295
rect 19843 2261 19852 2295
rect 19800 2252 19852 2261
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 30380 2524 30432 2576
rect 23848 2499 23900 2508
rect 23848 2465 23857 2499
rect 23857 2465 23891 2499
rect 23891 2465 23900 2499
rect 23848 2456 23900 2465
rect 27804 2499 27856 2508
rect 27804 2465 27813 2499
rect 27813 2465 27847 2499
rect 27847 2465 27856 2499
rect 27804 2456 27856 2465
rect 31024 2592 31076 2644
rect 34336 2635 34388 2644
rect 34336 2601 34345 2635
rect 34345 2601 34379 2635
rect 34379 2601 34388 2635
rect 34336 2592 34388 2601
rect 36176 2635 36228 2644
rect 36176 2601 36185 2635
rect 36185 2601 36219 2635
rect 36219 2601 36228 2635
rect 36176 2592 36228 2601
rect 37832 2592 37884 2644
rect 38844 2592 38896 2644
rect 40040 2635 40092 2644
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 40592 2592 40644 2644
rect 30656 2499 30708 2508
rect 30656 2465 30665 2499
rect 30665 2465 30699 2499
rect 30699 2465 30708 2499
rect 30656 2456 30708 2465
rect 31668 2499 31720 2508
rect 31668 2465 31677 2499
rect 31677 2465 31711 2499
rect 31711 2465 31720 2499
rect 31668 2456 31720 2465
rect 33508 2499 33560 2508
rect 33508 2465 33517 2499
rect 33517 2465 33551 2499
rect 33551 2465 33560 2499
rect 33508 2456 33560 2465
rect 34520 2499 34572 2508
rect 34520 2465 34529 2499
rect 34529 2465 34563 2499
rect 34563 2465 34572 2499
rect 34520 2456 34572 2465
rect 37280 2456 37332 2508
rect 38660 2456 38712 2508
rect 39212 2499 39264 2508
rect 39212 2465 39221 2499
rect 39221 2465 39255 2499
rect 39255 2465 39264 2499
rect 39212 2456 39264 2465
rect 40224 2499 40276 2508
rect 40224 2465 40233 2499
rect 40233 2465 40267 2499
rect 40267 2465 40276 2499
rect 40224 2456 40276 2465
rect 41420 2456 41472 2508
rect 43076 2499 43128 2508
rect 43076 2465 43085 2499
rect 43085 2465 43119 2499
rect 43119 2465 43128 2499
rect 43076 2456 43128 2465
rect 30472 2320 30524 2372
rect 40408 2320 40460 2372
rect 23480 2252 23532 2304
rect 9947 2150 9999 2202
rect 10011 2150 10063 2202
rect 10075 2150 10127 2202
rect 10139 2150 10191 2202
rect 27878 2150 27930 2202
rect 27942 2150 27994 2202
rect 28006 2150 28058 2202
rect 28070 2150 28122 2202
rect 45808 2150 45860 2202
rect 45872 2150 45924 2202
rect 45936 2150 45988 2202
rect 46000 2150 46052 2202
rect 19800 2048 19852 2100
rect 29184 2048 29236 2100
<< metal2 >>
rect 294 26400 350 27200
rect 938 26400 994 27200
rect 1674 26400 1730 27200
rect 2410 26400 2466 27200
rect 3146 26400 3202 27200
rect 3882 26400 3938 27200
rect 4526 26400 4582 27200
rect 5262 26400 5318 27200
rect 5998 26400 6054 27200
rect 6734 26400 6790 27200
rect 7470 26400 7526 27200
rect 8114 26400 8170 27200
rect 8850 26400 8906 27200
rect 9586 26400 9642 27200
rect 10322 26400 10378 27200
rect 11058 26400 11114 27200
rect 11702 26400 11758 27200
rect 12438 26400 12494 27200
rect 13174 26400 13230 27200
rect 13910 26400 13966 27200
rect 14646 26400 14702 27200
rect 15290 26400 15346 27200
rect 16026 26400 16082 27200
rect 16762 26400 16818 27200
rect 17498 26400 17554 27200
rect 18234 26400 18290 27200
rect 18970 26400 19026 27200
rect 19614 26400 19670 27200
rect 20350 26400 20406 27200
rect 21086 26400 21142 27200
rect 21822 26400 21878 27200
rect 22558 26400 22614 27200
rect 23202 26400 23258 27200
rect 23938 26400 23994 27200
rect 24674 26400 24730 27200
rect 25410 26400 25466 27200
rect 26146 26400 26202 27200
rect 26790 26400 26846 27200
rect 27526 26400 27582 27200
rect 28262 26400 28318 27200
rect 28998 26400 29054 27200
rect 29734 26400 29790 27200
rect 30378 26400 30434 27200
rect 31114 26400 31170 27200
rect 31850 26400 31906 27200
rect 32586 26400 32642 27200
rect 33322 26400 33378 27200
rect 33966 26400 34022 27200
rect 34702 26400 34758 27200
rect 35438 26400 35494 27200
rect 36174 26400 36230 27200
rect 36910 26400 36966 27200
rect 37646 26400 37702 27200
rect 38290 26400 38346 27200
rect 39026 26400 39082 27200
rect 39762 26400 39818 27200
rect 40498 26400 40554 27200
rect 41234 26400 41290 27200
rect 41878 26400 41934 27200
rect 42614 26400 42670 27200
rect 43350 26400 43406 27200
rect 44086 26400 44142 27200
rect 44822 26400 44878 27200
rect 45466 26400 45522 27200
rect 46202 26400 46258 27200
rect 46938 26400 46994 27200
rect 47674 26400 47730 27200
rect 48410 26400 48466 27200
rect 49054 26400 49110 27200
rect 49790 26400 49846 27200
rect 50526 26400 50582 27200
rect 51262 26400 51318 27200
rect 51998 26400 52054 27200
rect 52642 26400 52698 27200
rect 53378 26400 53434 27200
rect 54114 26400 54170 27200
rect 54850 26400 54906 27200
rect 55586 26400 55642 27200
rect 308 22778 336 26400
rect 952 23186 980 26400
rect 1688 24410 1716 26400
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 940 23180 992 23186
rect 940 23122 992 23128
rect 2424 22982 2452 26400
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 296 22772 348 22778
rect 296 22714 348 22720
rect 3160 22642 3188 26400
rect 3896 23322 3924 26400
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 4080 23118 4108 24006
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 4080 22642 4108 23054
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 2056 22234 2084 22510
rect 3332 22432 3384 22438
rect 3332 22374 3384 22380
rect 2044 22228 2096 22234
rect 2044 22170 2096 22176
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2516 22001 2544 22034
rect 2502 21992 2558 22001
rect 2502 21927 2558 21936
rect 3344 21554 3372 22374
rect 4264 22234 4292 24142
rect 4540 23118 4568 26400
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 4356 22642 4384 23054
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4908 22506 4936 22578
rect 4896 22500 4948 22506
rect 4896 22442 4948 22448
rect 4908 22234 4936 22442
rect 4252 22228 4304 22234
rect 4252 22170 4304 22176
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3344 19922 3372 21490
rect 4632 21418 4660 22034
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4816 20534 4844 20878
rect 5276 20534 5304 26400
rect 6012 24342 6040 26400
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6000 24336 6052 24342
rect 6000 24278 6052 24284
rect 6564 24274 6592 24550
rect 5908 24268 5960 24274
rect 5908 24210 5960 24216
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 5816 24064 5868 24070
rect 5920 24018 5948 24210
rect 5868 24012 5948 24018
rect 5816 24006 5948 24012
rect 5828 23990 5948 24006
rect 5920 23254 5948 23990
rect 5908 23248 5960 23254
rect 5908 23190 5960 23196
rect 5724 22976 5776 22982
rect 5724 22918 5776 22924
rect 5736 22506 5764 22918
rect 5724 22500 5776 22506
rect 5724 22442 5776 22448
rect 5736 22166 5764 22442
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 5724 22160 5776 22166
rect 5724 22102 5776 22108
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5828 21690 5856 21966
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5644 21146 5672 21422
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5736 20398 5764 21286
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5828 20602 5856 20946
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3700 20392 3752 20398
rect 3700 20334 3752 20340
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 3528 20058 3556 20334
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19718 1808 19790
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 3712 19514 3740 20334
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 4264 19394 4292 20334
rect 5908 20324 5960 20330
rect 5908 20266 5960 20272
rect 5920 19718 5948 20266
rect 6196 19854 6224 22034
rect 6656 21978 6684 22170
rect 6748 22098 6776 26400
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 23526 6868 24142
rect 7208 23730 7236 24686
rect 7484 24410 7512 26400
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 6932 22710 6960 23122
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 6932 22234 6960 22646
rect 7024 22574 7052 23258
rect 7116 23186 7144 23598
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7024 22098 7052 22510
rect 7116 22234 7144 22578
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 6656 21950 6960 21978
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6656 19922 6684 21014
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 4172 19366 4292 19394
rect 4172 19310 4200 19366
rect 5920 19310 5948 19654
rect 6196 19446 6224 19790
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 6656 19310 6684 19858
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 2976 18970 3004 19246
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 3160 18834 3188 19110
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 4172 18358 4200 19246
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2148 17338 2176 17682
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2608 16794 2636 17070
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2792 15706 2820 16594
rect 2884 16046 2912 18158
rect 4264 18154 4292 18770
rect 5092 18222 5120 18838
rect 6656 18714 6684 19246
rect 6748 19242 6776 19858
rect 6736 19236 6788 19242
rect 6736 19178 6788 19184
rect 6748 18834 6776 19178
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6656 18686 6776 18714
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4356 17882 4384 18158
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 5276 17338 5304 18158
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4080 16658 4108 17002
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5644 16658 5672 16934
rect 6380 16658 6408 18022
rect 6748 17542 6776 18686
rect 6840 18222 6868 21626
rect 6932 21554 6960 21950
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 7024 21486 7052 22034
rect 7104 21956 7156 21962
rect 7104 21898 7156 21904
rect 7116 21622 7144 21898
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7024 21078 7052 21422
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 19174 6960 20334
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6932 18426 6960 18634
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17746 6868 18158
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2504 15632 2556 15638
rect 2504 15574 2556 15580
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2240 12986 2268 13806
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13394 2360 13670
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2148 11354 2176 11630
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2332 10606 2360 13126
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2424 12646 2452 12718
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2516 10418 2544 15574
rect 3160 15570 3188 16390
rect 3804 15706 3832 16594
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 3896 14958 3924 15982
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 14482 3464 14758
rect 3988 14482 4016 15914
rect 4080 15026 4108 16594
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4172 14958 4200 16186
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 15570 5028 15846
rect 6380 15638 6408 16594
rect 6564 16250 6592 16594
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6748 16182 6776 17478
rect 7208 17202 7236 23530
rect 7380 22500 7432 22506
rect 7380 22442 7432 22448
rect 7286 21992 7342 22001
rect 7286 21927 7288 21936
rect 7340 21927 7342 21936
rect 7288 21898 7340 21904
rect 7392 21010 7420 22442
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7484 20874 7512 21422
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18290 7420 18566
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 16658 7604 17070
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6840 16114 6868 16390
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6932 16046 6960 16390
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 4448 13870 4476 14894
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3252 12306 3280 13670
rect 4448 13530 4476 13806
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 3436 12442 3464 12718
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3344 11286 3372 11494
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 4264 11218 4292 12582
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4448 10810 4476 12718
rect 4540 11898 4568 14350
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5460 13870 5488 14214
rect 6288 14074 6316 15506
rect 6380 15026 6408 15574
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6472 14482 6500 15370
rect 7576 14958 7604 15846
rect 7668 15706 7696 23598
rect 8024 23180 8076 23186
rect 8024 23122 8076 23128
rect 8036 22574 8064 23122
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 7932 20868 7984 20874
rect 7932 20810 7984 20816
rect 7944 20398 7972 20810
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 8128 18426 8156 26400
rect 8864 24818 8892 26400
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 8680 24274 8708 24550
rect 9600 24290 9628 26400
rect 9921 25052 10217 25072
rect 9977 25050 10001 25052
rect 10057 25050 10081 25052
rect 10137 25050 10161 25052
rect 9999 24998 10001 25050
rect 10063 24998 10075 25050
rect 10137 24998 10139 25050
rect 9977 24996 10001 24998
rect 10057 24996 10081 24998
rect 10137 24996 10161 24998
rect 9921 24976 10217 24996
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 9508 24262 9628 24290
rect 9772 24268 9824 24274
rect 8760 23656 8812 23662
rect 8760 23598 8812 23604
rect 8772 23254 8800 23598
rect 8760 23248 8812 23254
rect 8760 23190 8812 23196
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8404 20058 8432 20334
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8588 19854 8616 22034
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8300 19304 8352 19310
rect 8298 19272 8300 19281
rect 8352 19272 8354 19281
rect 8298 19207 8354 19216
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8036 17270 8064 17478
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8036 17134 8064 17206
rect 8312 17134 8340 17750
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8036 16182 8064 17070
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 8036 15638 8064 16118
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 6564 14618 6592 14894
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13394 5488 13806
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 4908 12442 4936 13330
rect 5552 13326 5580 14010
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 5000 12306 5028 12582
rect 6196 12442 6224 12718
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 5552 11694 5580 12038
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 4540 11354 4568 11630
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 5276 11218 5304 11494
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 2332 10390 2544 10418
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2148 5370 2176 9046
rect 2332 5914 2360 10390
rect 3252 10130 3280 10406
rect 3344 10266 3372 10542
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2884 8634 2912 8978
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3068 8090 3096 8366
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3252 7954 3280 9862
rect 4172 9518 4200 9862
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4356 9382 4384 10542
rect 4632 9518 4660 11018
rect 6196 10810 6224 11086
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6380 10606 6408 10950
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4816 9178 4844 10066
rect 5184 9586 5212 10406
rect 5368 9722 5396 10542
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 5460 8634 5488 9454
rect 5552 9042 5580 10406
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9654 6040 10066
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5552 8090 5580 8366
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 3528 7546 3556 7890
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6254 3372 6598
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 2884 5914 2912 6190
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2332 4214 2360 5714
rect 3804 5710 3832 6802
rect 4724 6458 4752 7278
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 4816 5642 4844 7210
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6254 4936 6598
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5000 5778 5028 6054
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 5368 5166 5396 6326
rect 5552 6254 5580 7686
rect 5736 7546 5764 7890
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6866 5856 7142
rect 5920 7002 5948 7278
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5644 6458 5672 6802
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5552 5370 5580 5782
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4690 5580 4966
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 6288 4078 6316 8502
rect 6656 8430 6684 14214
rect 6932 13394 6960 14486
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13456 7064 13462
rect 7116 13410 7144 13806
rect 7064 13404 7144 13410
rect 7012 13398 7144 13404
rect 6920 13388 6972 13394
rect 7024 13382 7144 13398
rect 7208 13394 7236 14758
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 6920 13330 6972 13336
rect 7116 12986 7144 13382
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11762 6868 12038
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6932 11354 6960 12242
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7024 11218 7052 11494
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 7300 10266 7328 14418
rect 8312 14074 8340 14826
rect 8404 14550 8432 18158
rect 8588 17746 8616 19790
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8680 18290 8708 19110
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 15978 8616 17002
rect 8772 16250 8800 23054
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9416 21554 9444 21830
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9416 21010 9444 21490
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9508 19281 9536 24262
rect 9772 24210 9824 24216
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9600 21962 9628 22442
rect 9692 22098 9720 24074
rect 9784 23730 9812 24210
rect 9921 23964 10217 23984
rect 9977 23962 10001 23964
rect 10057 23962 10081 23964
rect 10137 23962 10161 23964
rect 9999 23910 10001 23962
rect 10063 23910 10075 23962
rect 10137 23910 10139 23962
rect 9977 23908 10001 23910
rect 10057 23908 10081 23910
rect 10137 23908 10161 23910
rect 9921 23888 10217 23908
rect 10336 23866 10364 26400
rect 11072 24290 11100 26400
rect 11716 24342 11744 26400
rect 11704 24336 11756 24342
rect 11072 24262 11376 24290
rect 11704 24278 11756 24284
rect 12452 24290 12480 26400
rect 13188 24410 13216 26400
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 12452 24262 12572 24290
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9921 22876 10217 22896
rect 9977 22874 10001 22876
rect 10057 22874 10081 22876
rect 10137 22874 10161 22876
rect 9999 22822 10001 22874
rect 10063 22822 10075 22874
rect 10137 22822 10139 22874
rect 9977 22820 10001 22822
rect 10057 22820 10081 22822
rect 10137 22820 10161 22822
rect 9921 22800 10217 22820
rect 10428 22642 10456 24142
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 11072 22710 11100 23122
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9600 21146 9628 21490
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9692 20058 9720 21830
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9494 19272 9550 19281
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 9416 19230 9494 19258
rect 8864 18834 8892 19178
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 9416 18612 9444 19230
rect 9494 19207 9550 19216
rect 9600 19174 9628 19790
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9600 18902 9628 19110
rect 9588 18896 9640 18902
rect 9588 18838 9640 18844
rect 9680 18624 9732 18630
rect 9416 18584 9680 18612
rect 9680 18566 9732 18572
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 17218 9720 18158
rect 9600 17202 9720 17218
rect 9784 17202 9812 22510
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 9921 21788 10217 21808
rect 9977 21786 10001 21788
rect 10057 21786 10081 21788
rect 10137 21786 10161 21788
rect 9999 21734 10001 21786
rect 10063 21734 10075 21786
rect 10137 21734 10139 21786
rect 9977 21732 10001 21734
rect 10057 21732 10081 21734
rect 10137 21732 10161 21734
rect 9921 21712 10217 21732
rect 10324 21412 10376 21418
rect 10324 21354 10376 21360
rect 9921 20700 10217 20720
rect 9977 20698 10001 20700
rect 10057 20698 10081 20700
rect 10137 20698 10161 20700
rect 9999 20646 10001 20698
rect 10063 20646 10075 20698
rect 10137 20646 10139 20698
rect 9977 20644 10001 20646
rect 10057 20644 10081 20646
rect 10137 20644 10161 20646
rect 9921 20624 10217 20644
rect 9921 19612 10217 19632
rect 9977 19610 10001 19612
rect 10057 19610 10081 19612
rect 10137 19610 10161 19612
rect 9999 19558 10001 19610
rect 10063 19558 10075 19610
rect 10137 19558 10139 19610
rect 9977 19556 10001 19558
rect 10057 19556 10081 19558
rect 10137 19556 10161 19558
rect 9921 19536 10217 19556
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10152 18834 10180 19246
rect 10336 18970 10364 21354
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10428 19378 10456 20198
rect 10520 19514 10548 22374
rect 11072 22098 11100 22374
rect 10600 22092 10652 22098
rect 10600 22034 10652 22040
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 10612 21690 10640 22034
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10888 21078 10916 22034
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 10980 21486 11008 21558
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10980 21010 11008 21422
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10152 18680 10180 18770
rect 10152 18652 10364 18680
rect 9921 18524 10217 18544
rect 9977 18522 10001 18524
rect 10057 18522 10081 18524
rect 10137 18522 10161 18524
rect 9999 18470 10001 18522
rect 10063 18470 10075 18522
rect 10137 18470 10139 18522
rect 9977 18468 10001 18470
rect 10057 18468 10081 18470
rect 10137 18468 10161 18470
rect 9921 18448 10217 18468
rect 10336 18426 10364 18652
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10980 17746 11008 20946
rect 11164 20806 11192 22510
rect 11256 21962 11284 22646
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11348 20890 11376 24262
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11256 20862 11376 20890
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11256 17882 11284 20862
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11348 20466 11376 20742
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11348 19990 11376 20402
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11348 19310 11376 19926
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11348 18766 11376 19246
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 9921 17436 10217 17456
rect 9977 17434 10001 17436
rect 10057 17434 10081 17436
rect 10137 17434 10161 17436
rect 9999 17382 10001 17434
rect 10063 17382 10075 17434
rect 10137 17382 10139 17434
rect 9977 17380 10001 17382
rect 10057 17380 10081 17382
rect 10137 17380 10161 17382
rect 9921 17360 10217 17380
rect 9588 17196 9720 17202
rect 9640 17190 9720 17196
rect 9772 17196 9824 17202
rect 9588 17138 9640 17144
rect 9772 17138 9824 17144
rect 10704 17134 10732 17478
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8576 15972 8628 15978
rect 8576 15914 8628 15920
rect 8588 15570 8616 15914
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 9048 14890 9076 15982
rect 9692 14958 9720 17070
rect 10428 16658 10456 17070
rect 10704 16726 10732 17070
rect 11256 16998 11284 17818
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11440 16794 11468 23122
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 11532 22080 11560 22986
rect 11612 22092 11664 22098
rect 11532 22052 11612 22080
rect 11532 21894 11560 22052
rect 11612 22034 11664 22040
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 12254 21584 12310 21593
rect 12254 21519 12256 21528
rect 12308 21519 12310 21528
rect 12256 21490 12308 21496
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12360 21146 12388 21422
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12176 19922 12204 20198
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11992 19446 12020 19790
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11980 18148 12032 18154
rect 11980 18090 12032 18096
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11808 17746 11836 17818
rect 11992 17746 12020 18090
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12360 16794 12388 17750
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 9921 16348 10217 16368
rect 9977 16346 10001 16348
rect 10057 16346 10081 16348
rect 10137 16346 10161 16348
rect 9999 16294 10001 16346
rect 10063 16294 10075 16346
rect 10137 16294 10139 16346
rect 9977 16292 10001 16294
rect 10057 16292 10081 16294
rect 10137 16292 10161 16294
rect 9921 16272 10217 16292
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 9968 15638 9996 15846
rect 10428 15706 10456 15846
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 9770 15464 9826 15473
rect 9770 15399 9826 15408
rect 9784 15366 9812 15399
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9921 15260 10217 15280
rect 9977 15258 10001 15260
rect 10057 15258 10081 15260
rect 10137 15258 10161 15260
rect 9999 15206 10001 15258
rect 10063 15206 10075 15258
rect 10137 15206 10139 15258
rect 9977 15204 10001 15206
rect 10057 15204 10081 15206
rect 10137 15204 10161 15206
rect 9921 15184 10217 15204
rect 10336 15065 10364 15506
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10322 15056 10378 15065
rect 10322 14991 10378 15000
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 13190 8064 13806
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12782 8064 13126
rect 8312 12918 8340 14010
rect 8404 13530 8432 14486
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 7576 11898 7604 12242
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7944 11694 7972 12038
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 9178 7512 9454
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7668 9042 7696 9318
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7484 8634 7512 8978
rect 8036 8906 8064 12242
rect 8588 11898 8616 12242
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8772 11694 8800 13942
rect 9692 12986 9720 14894
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 9921 14172 10217 14192
rect 9977 14170 10001 14172
rect 10057 14170 10081 14172
rect 10137 14170 10161 14172
rect 9999 14118 10001 14170
rect 10063 14118 10075 14170
rect 10137 14118 10139 14170
rect 9977 14116 10001 14118
rect 10057 14116 10081 14118
rect 10137 14116 10161 14118
rect 9921 14096 10217 14116
rect 10336 13394 10364 14826
rect 10428 14482 10456 15302
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 9921 13084 10217 13104
rect 9977 13082 10001 13084
rect 10057 13082 10081 13084
rect 10137 13082 10161 13084
rect 9999 13030 10001 13082
rect 10063 13030 10075 13082
rect 10137 13030 10139 13082
rect 9977 13028 10001 13030
rect 10057 13028 10081 13030
rect 10137 13028 10161 13030
rect 9921 13008 10217 13028
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 10336 12782 10364 13126
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8864 11354 8892 12718
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9968 12442 9996 12650
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 10428 12238 10456 12922
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 9921 11996 10217 12016
rect 9977 11994 10001 11996
rect 10057 11994 10081 11996
rect 10137 11994 10161 11996
rect 9999 11942 10001 11994
rect 10063 11942 10075 11994
rect 10137 11942 10139 11994
rect 9977 11940 10001 11942
rect 10057 11940 10081 11942
rect 10137 11940 10161 11942
rect 9921 11920 10217 11940
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 9048 11218 9076 11494
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9692 10606 9720 11494
rect 9784 10810 9812 11630
rect 9921 10908 10217 10928
rect 9977 10906 10001 10908
rect 10057 10906 10081 10908
rect 10137 10906 10161 10908
rect 9999 10854 10001 10906
rect 10063 10854 10075 10906
rect 10137 10854 10139 10906
rect 9977 10852 10001 10854
rect 10057 10852 10081 10854
rect 10137 10852 10161 10854
rect 9921 10832 10217 10852
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10130 9536 10406
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 8220 9722 8248 10066
rect 9921 9820 10217 9840
rect 9977 9818 10001 9820
rect 10057 9818 10081 9820
rect 10137 9818 10161 9820
rect 9999 9766 10001 9818
rect 10063 9766 10075 9818
rect 10137 9766 10139 9818
rect 9977 9764 10001 9766
rect 10057 9764 10081 9766
rect 10137 9764 10161 9766
rect 9921 9744 10217 9764
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 7668 7954 7696 8774
rect 7760 8430 7788 8774
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7342 6592 7686
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6920 5772 6972 5778
rect 6840 5732 6920 5760
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4826 6408 5102
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6472 4282 6500 5034
rect 6840 4554 6868 5732
rect 6920 5714 6972 5720
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6932 4690 6960 5578
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4690 7696 4966
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 8220 4078 8248 8842
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 7546 8340 8366
rect 8680 8090 8708 8978
rect 8772 8566 8800 9454
rect 10520 9330 10548 15846
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 10612 12442 10640 15506
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 15162 11284 15438
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11164 14482 11192 14894
rect 11152 14476 11204 14482
rect 11336 14476 11388 14482
rect 11204 14436 11336 14464
rect 11152 14418 11204 14424
rect 11336 14418 11388 14424
rect 11532 14090 11560 15506
rect 11716 14482 11744 16458
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11992 15502 12020 16186
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12360 15094 12388 16526
rect 12544 15473 12572 24262
rect 13636 24268 13688 24274
rect 13636 24210 13688 24216
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12636 23254 12664 24142
rect 13648 23730 13676 24210
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12728 22574 12756 23462
rect 13280 23322 13308 23462
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22098 12756 22510
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 13096 22234 13124 22374
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12714 21584 12770 21593
rect 12714 21519 12716 21528
rect 12768 21519 12770 21528
rect 12716 21490 12768 21496
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12636 20602 12664 20878
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12728 20534 12756 21354
rect 13832 21146 13860 21422
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 13280 20398 13308 20946
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13556 19990 13584 20334
rect 13544 19984 13596 19990
rect 13544 19926 13596 19932
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12912 19786 12940 19858
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12636 17882 12664 18634
rect 13096 18426 13124 19246
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13464 18834 13492 19110
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13096 18222 13124 18362
rect 13280 18222 13308 18770
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12636 15570 12664 17818
rect 13832 17814 13860 18770
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17202 13032 17478
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13188 16114 13216 16594
rect 13924 16250 13952 26400
rect 14660 23866 14688 26400
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14844 22234 14872 22918
rect 15120 22710 15148 23802
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14844 21690 14872 22170
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14844 21486 14872 21626
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 15120 21146 15148 22646
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15120 20602 15148 21082
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14200 19922 14228 20198
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15028 18290 15056 18566
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14292 16658 14320 17206
rect 14384 17134 14412 18022
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14384 16998 14412 17070
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14384 16454 14412 16934
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13556 15638 13584 15982
rect 14384 15910 14412 16390
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12530 15464 12586 15473
rect 12440 15428 12492 15434
rect 12530 15399 12586 15408
rect 12440 15370 12492 15376
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12348 14952 12400 14958
rect 12452 14940 12480 15370
rect 12544 15026 12572 15399
rect 12636 15094 12664 15506
rect 12624 15088 12676 15094
rect 13176 15088 13228 15094
rect 12624 15030 12676 15036
rect 13082 15056 13138 15065
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12636 14958 12664 15030
rect 13176 15030 13228 15036
rect 13082 14991 13138 15000
rect 13096 14958 13124 14991
rect 13188 14958 13216 15030
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 12400 14912 12480 14940
rect 12624 14952 12676 14958
rect 12348 14894 12400 14900
rect 12624 14894 12676 14900
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12820 14618 12848 14826
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 11348 14062 11560 14090
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10888 12238 10916 13126
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10796 9450 10824 11630
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10428 9302 10548 9330
rect 9921 8732 10217 8752
rect 9977 8730 10001 8732
rect 10057 8730 10081 8732
rect 10137 8730 10161 8732
rect 9999 8678 10001 8730
rect 10063 8678 10075 8730
rect 10137 8678 10139 8730
rect 9977 8676 10001 8678
rect 10057 8676 10081 8678
rect 10137 8676 10161 8678
rect 9921 8656 10217 8676
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 6866 8340 7142
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8404 6730 8432 7890
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7342 8800 7686
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6866 8708 7142
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6254 8616 6598
rect 8956 6458 8984 7278
rect 9692 6730 9720 7890
rect 9921 7644 10217 7664
rect 9977 7642 10001 7644
rect 10057 7642 10081 7644
rect 10137 7642 10161 7644
rect 9999 7590 10001 7642
rect 10063 7590 10075 7642
rect 10137 7590 10139 7642
rect 9977 7588 10001 7590
rect 10057 7588 10081 7590
rect 10137 7588 10161 7590
rect 9921 7568 10217 7588
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9921 6556 10217 6576
rect 9977 6554 10001 6556
rect 10057 6554 10081 6556
rect 10137 6554 10161 6556
rect 9999 6502 10001 6554
rect 10063 6502 10075 6554
rect 10137 6502 10139 6554
rect 9977 6500 10001 6502
rect 10057 6500 10081 6502
rect 10137 6500 10161 6502
rect 9921 6480 10217 6500
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 10428 6390 10456 9302
rect 10508 9104 10560 9110
rect 10692 9104 10744 9110
rect 10560 9052 10692 9058
rect 10508 9046 10744 9052
rect 10520 9030 10732 9046
rect 11242 8936 11298 8945
rect 11242 8871 11244 8880
rect 11296 8871 11298 8880
rect 11244 8842 11296 8848
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7342 10824 8230
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 6866 10640 7142
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9048 5370 9076 5714
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9784 5166 9812 6054
rect 9921 5468 10217 5488
rect 9977 5466 10001 5468
rect 10057 5466 10081 5468
rect 10137 5466 10161 5468
rect 9999 5414 10001 5466
rect 10063 5414 10075 5466
rect 10137 5414 10139 5466
rect 9977 5412 10001 5414
rect 10057 5412 10081 5414
rect 10137 5412 10161 5414
rect 9921 5392 10217 5412
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 10336 4690 10364 6054
rect 10428 5914 10456 6190
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10520 5234 10548 6598
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10612 4826 10640 5714
rect 11072 5370 11100 6190
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 11164 4554 11192 6802
rect 11348 6458 11376 14062
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11532 12782 11560 13942
rect 11716 12986 11744 14418
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 13394 12480 14214
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11440 11354 11468 11630
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 11440 10810 11468 11154
rect 12544 10810 12572 11154
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 11532 10266 11560 10542
rect 12544 10266 12572 10542
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11440 8498 11468 9862
rect 12636 9722 12664 10066
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 9042 11652 9318
rect 12452 9178 12480 9454
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11440 8090 11468 8298
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11532 7954 11560 8502
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11624 8090 11652 8366
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11716 7954 11744 8774
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 12728 6730 12756 14418
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13004 13938 13032 14282
rect 13648 13938 13676 14962
rect 13820 14612 13872 14618
rect 13872 14572 14044 14600
rect 13820 14554 13872 14560
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13740 13938 13768 14486
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13280 13734 13308 13806
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13280 13326 13308 13670
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 11218 13032 12582
rect 13188 12238 13216 12718
rect 13372 12238 13400 12922
rect 13556 12782 13584 13126
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13832 11898 13860 13806
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12102 13952 12582
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 11354 13492 11630
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13556 10266 13584 10542
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13464 9178 13492 9454
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13648 9042 13676 11018
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10130 13768 10950
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13924 9518 13952 11766
rect 14016 11286 14044 14572
rect 14200 12782 14228 15642
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14292 15162 14320 15506
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14292 11694 14320 14010
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14200 10810 14228 11086
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14384 10606 14412 11494
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9654 14228 9998
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13188 8634 13216 8978
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5778 11652 6054
rect 12636 5778 12664 6598
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 11440 5166 11468 5510
rect 12452 5166 12480 5510
rect 13372 5370 13400 6190
rect 13464 5914 13492 6802
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13556 5302 13584 7278
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5778 13676 6054
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 9921 4380 10217 4400
rect 9977 4378 10001 4380
rect 10057 4378 10081 4380
rect 10137 4378 10161 4380
rect 9999 4326 10001 4378
rect 10063 4326 10075 4378
rect 10137 4326 10139 4378
rect 9977 4324 10001 4326
rect 10057 4324 10081 4326
rect 10137 4324 10161 4326
rect 9921 4304 10217 4324
rect 13280 4282 13308 4626
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13740 4078 13768 8502
rect 13832 7954 13860 9318
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 8090 14412 8366
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 14660 7410 14688 12038
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6254 14412 7142
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14476 5914 14504 6190
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 4826 14136 5102
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14016 3738 14044 4014
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14200 3602 14228 4422
rect 14292 4282 14320 4626
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14752 3942 14780 17478
rect 15304 17134 15332 26400
rect 16040 24410 16068 26400
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 15396 23866 15424 24210
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15384 23044 15436 23050
rect 15384 22986 15436 22992
rect 15396 22642 15424 22986
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15856 21894 15884 23122
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15580 21486 15608 21830
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16040 21146 16068 21422
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15856 20466 15884 20946
rect 16132 20602 16160 23054
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16684 22710 16712 22986
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16316 19922 16344 19994
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15764 18834 15792 19654
rect 16316 19310 16344 19858
rect 16500 19854 16528 20470
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16500 19514 16528 19790
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15120 16998 15148 17070
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14936 15910 14964 16594
rect 15120 16590 15148 16934
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14844 14074 14872 14418
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14936 13734 14964 15846
rect 15304 15570 15332 16186
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15382 15056 15438 15065
rect 15382 14991 15438 15000
rect 15396 14618 15424 14991
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 12986 14964 13670
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 15212 11898 15240 14282
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15304 11898 15332 12106
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15396 11694 15424 14214
rect 15488 13938 15516 15846
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15672 12306 15700 14758
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15764 13938 15792 14554
rect 15856 14074 15884 14894
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15396 8430 15424 11018
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15212 5234 15240 7142
rect 15304 5778 15332 7142
rect 15396 6458 15424 7278
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15948 4826 15976 17818
rect 16500 17746 16528 18090
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16040 17134 16068 17274
rect 16500 17202 16528 17682
rect 16592 17338 16620 18906
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16658 16528 16934
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16592 16046 16620 17274
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16776 15910 16804 26400
rect 17512 24410 17540 26400
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17788 23662 17816 24142
rect 17776 23656 17828 23662
rect 17776 23598 17828 23604
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17144 21690 17172 21966
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17052 21350 17080 21626
rect 17420 21622 17448 21966
rect 17408 21616 17460 21622
rect 17408 21558 17460 21564
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 16960 21010 16988 21286
rect 17052 21146 17080 21286
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 17052 20942 17080 21082
rect 17144 21078 17172 21422
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 17144 20602 17172 21014
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 17788 20874 18000 20890
rect 17776 20868 18012 20874
rect 17828 20862 17960 20868
rect 17776 20810 17828 20816
rect 17960 20810 18012 20816
rect 18064 20806 18092 20946
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17512 19922 17540 20742
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17236 18970 17264 19790
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17788 18426 17816 19110
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 17134 17172 17478
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17236 16794 17264 17682
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17880 16726 17908 19722
rect 17972 19446 18000 20334
rect 18064 20058 18092 20334
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18248 19922 18276 26400
rect 18984 24698 19012 26400
rect 18984 24670 19380 24698
rect 18886 24508 19182 24528
rect 18942 24506 18966 24508
rect 19022 24506 19046 24508
rect 19102 24506 19126 24508
rect 18964 24454 18966 24506
rect 19028 24454 19040 24506
rect 19102 24454 19104 24506
rect 18942 24452 18966 24454
rect 19022 24452 19046 24454
rect 19102 24452 19126 24454
rect 18886 24432 19182 24452
rect 19352 23866 19380 24670
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18524 22778 18552 23122
rect 18616 22982 18644 23598
rect 18886 23420 19182 23440
rect 18942 23418 18966 23420
rect 19022 23418 19046 23420
rect 19102 23418 19126 23420
rect 18964 23366 18966 23418
rect 19028 23366 19040 23418
rect 19102 23366 19104 23418
rect 18942 23364 18966 23366
rect 19022 23364 19046 23366
rect 19102 23364 19126 23366
rect 18886 23344 19182 23364
rect 19444 23254 19472 24210
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19536 23322 19564 23462
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 19352 22574 19380 23054
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19628 22420 19656 26400
rect 20364 24410 20392 26400
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 19260 22392 19656 22420
rect 18886 22332 19182 22352
rect 18942 22330 18966 22332
rect 19022 22330 19046 22332
rect 19102 22330 19126 22332
rect 18964 22278 18966 22330
rect 19028 22278 19040 22330
rect 19102 22278 19104 22330
rect 18942 22276 18966 22278
rect 19022 22276 19046 22278
rect 19102 22276 19126 22278
rect 18886 22256 19182 22276
rect 18604 21412 18656 21418
rect 18604 21354 18656 21360
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18524 20398 18552 20946
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18340 19718 18368 20198
rect 18524 19922 18552 20334
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 18064 18970 18092 19654
rect 18524 19514 18552 19858
rect 18616 19514 18644 21354
rect 18886 21244 19182 21264
rect 18942 21242 18966 21244
rect 19022 21242 19046 21244
rect 19102 21242 19126 21244
rect 18964 21190 18966 21242
rect 19028 21190 19040 21242
rect 19102 21190 19104 21242
rect 18942 21188 18966 21190
rect 19022 21188 19046 21190
rect 19102 21188 19126 21190
rect 18886 21168 19182 21188
rect 19260 20466 19288 22392
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 18886 20156 19182 20176
rect 18942 20154 18966 20156
rect 19022 20154 19046 20156
rect 19102 20154 19126 20156
rect 18964 20102 18966 20154
rect 19028 20102 19040 20154
rect 19102 20102 19104 20154
rect 18942 20100 18966 20102
rect 19022 20100 19046 20102
rect 19102 20100 19126 20102
rect 18886 20080 19182 20100
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 18064 17882 18092 18294
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18248 17746 18276 19382
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18698 18368 19110
rect 18886 19068 19182 19088
rect 18942 19066 18966 19068
rect 19022 19066 19046 19068
rect 19102 19066 19126 19068
rect 18964 19014 18966 19066
rect 19028 19014 19040 19066
rect 19102 19014 19104 19066
rect 18942 19012 18966 19014
rect 19022 19012 19046 19014
rect 19102 19012 19126 19014
rect 18886 18992 19182 19012
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 18064 16658 18092 17478
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 17052 15570 17080 15914
rect 18524 15706 18552 16458
rect 18708 15978 18736 17206
rect 18800 16522 18828 18158
rect 18886 17980 19182 18000
rect 18942 17978 18966 17980
rect 19022 17978 19046 17980
rect 19102 17978 19126 17980
rect 18964 17926 18966 17978
rect 19028 17926 19040 17978
rect 19102 17926 19104 17978
rect 18942 17924 18966 17926
rect 19022 17924 19046 17926
rect 19102 17924 19126 17926
rect 18886 17904 19182 17924
rect 19352 17882 19380 19858
rect 19444 19310 19472 21422
rect 19720 21078 19748 23258
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20732 22710 20760 22918
rect 20824 22710 20852 24142
rect 21100 23322 21128 26400
rect 21836 24818 21864 26400
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21560 24274 21588 24550
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20916 22234 20944 23054
rect 21100 22574 21128 23122
rect 21192 22642 21220 24142
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 21008 21690 21036 22510
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19812 21146 19840 21422
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19708 21072 19760 21078
rect 19708 21014 19760 21020
rect 21008 21010 21036 21626
rect 20996 21004 21048 21010
rect 20996 20946 21048 20952
rect 21284 20398 21312 23122
rect 21376 21894 21404 23734
rect 21560 23594 21588 24210
rect 22480 23866 22508 24686
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 21548 23588 21600 23594
rect 21548 23530 21600 23536
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 19922 20392 20198
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19720 19310 19748 19790
rect 20548 19446 20576 20266
rect 21284 20058 21312 20334
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 20732 19174 20760 19790
rect 21468 19310 21496 22034
rect 21560 21078 21588 23530
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21652 22982 21680 23258
rect 21744 23050 21772 23462
rect 22112 23050 22140 23462
rect 21732 23044 21784 23050
rect 21732 22986 21784 22992
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21652 22710 21680 22918
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 21652 22166 21680 22646
rect 21928 22642 21956 22918
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21928 22234 21956 22578
rect 22204 22506 22232 23530
rect 22572 22982 22600 26400
rect 23216 24800 23244 26400
rect 23216 24772 23520 24800
rect 23492 24410 23520 24772
rect 23480 24404 23532 24410
rect 23480 24346 23532 24352
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23676 23254 23704 24142
rect 23952 23254 23980 26400
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24412 23730 24440 24550
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23664 23248 23716 23254
rect 23664 23190 23716 23196
rect 23940 23248 23992 23254
rect 23940 23190 23992 23196
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 21652 21962 21680 22102
rect 21640 21956 21692 21962
rect 21640 21898 21692 21904
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 21350 22324 21898
rect 22388 21690 22416 22374
rect 23216 22234 23244 22714
rect 23308 22710 23336 23122
rect 23492 22778 23520 23190
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23308 22506 23336 22646
rect 23296 22500 23348 22506
rect 23296 22442 23348 22448
rect 23204 22228 23256 22234
rect 23860 22216 23888 23054
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23204 22170 23256 22176
rect 23584 22188 23888 22216
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22388 21486 22416 21626
rect 22572 21622 22600 22034
rect 23480 21956 23532 21962
rect 23584 21944 23612 22188
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23532 21916 23612 21944
rect 23664 21956 23716 21962
rect 23480 21898 23532 21904
rect 23664 21898 23716 21904
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21560 19854 21588 21014
rect 22756 21010 22784 21830
rect 23676 21486 23704 21898
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 22006 19408 22062 19417
rect 22006 19343 22008 19352
rect 22060 19343 22062 19352
rect 22008 19314 22060 19320
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 21008 18358 21036 18702
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19260 17066 19288 17818
rect 19720 17746 19748 18090
rect 21100 17746 21128 19246
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 18290 21404 18566
rect 23032 18426 23060 20402
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23400 20058 23428 20198
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 23032 18086 23060 18362
rect 23492 18154 23520 21286
rect 23584 20874 23612 21422
rect 23768 21078 23796 22034
rect 23860 22030 23888 22188
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 21350 23888 21490
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23756 21072 23808 21078
rect 23756 21014 23808 21020
rect 23572 20868 23624 20874
rect 23572 20810 23624 20816
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23676 19310 23704 19654
rect 23952 19310 23980 22918
rect 24688 22778 24716 26400
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25240 23866 25268 24210
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25320 23248 25372 23254
rect 25320 23190 25372 23196
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24032 22568 24084 22574
rect 24030 22536 24032 22545
rect 24216 22568 24268 22574
rect 24084 22536 24086 22545
rect 24308 22568 24360 22574
rect 24216 22510 24268 22516
rect 24306 22536 24308 22545
rect 24360 22536 24362 22545
rect 24030 22471 24086 22480
rect 24228 22438 24256 22510
rect 24306 22471 24362 22480
rect 25228 22500 25280 22506
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24320 22098 24348 22471
rect 25228 22442 25280 22448
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24124 21412 24176 21418
rect 24124 21354 24176 21360
rect 24032 20528 24084 20534
rect 24030 20496 24032 20505
rect 24084 20496 24086 20505
rect 24136 20466 24164 21354
rect 24780 21078 24808 21966
rect 25240 21486 25268 22442
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24952 20868 25004 20874
rect 24952 20810 25004 20816
rect 24964 20602 24992 20810
rect 25240 20806 25268 21286
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 24308 20528 24360 20534
rect 24308 20470 24360 20476
rect 24030 20431 24086 20440
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24124 20324 24176 20330
rect 24124 20266 24176 20272
rect 24136 20058 24164 20266
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24320 19718 24348 20470
rect 24964 20466 24992 20538
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 25332 19310 25360 23190
rect 25424 20466 25452 26400
rect 26160 23866 26188 26400
rect 26148 23860 26200 23866
rect 26148 23802 26200 23808
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25608 22982 25636 23122
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 26700 22976 26752 22982
rect 26700 22918 26752 22924
rect 25608 22574 25636 22918
rect 26712 22642 26740 22918
rect 26700 22636 26752 22642
rect 26700 22578 26752 22584
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 25412 20460 25464 20466
rect 25412 20402 25464 20408
rect 25412 20324 25464 20330
rect 25412 20266 25464 20272
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 24228 18834 24256 19110
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 25240 18698 25268 19246
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25240 18290 25268 18634
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 22020 17746 22048 18022
rect 23032 17746 23060 18022
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 18886 16892 19182 16912
rect 18942 16890 18966 16892
rect 19022 16890 19046 16892
rect 19102 16890 19126 16892
rect 18964 16838 18966 16890
rect 19028 16838 19040 16890
rect 19102 16838 19104 16890
rect 18942 16836 18966 16838
rect 19022 16836 19046 16838
rect 19102 16836 19126 16838
rect 18886 16816 19182 16836
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 18524 15094 18552 15642
rect 17960 15088 18012 15094
rect 18512 15088 18564 15094
rect 17960 15030 18012 15036
rect 18432 15036 18512 15042
rect 18432 15030 18564 15036
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16040 13530 16068 14350
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16500 12918 16528 14826
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 13870 16712 14758
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16960 14006 16988 14554
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16592 13682 16620 13806
rect 16592 13654 16712 13682
rect 16684 13394 16712 13654
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16684 12986 16712 13330
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16040 11762 16068 12718
rect 17236 12322 17264 13398
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 16592 12306 16712 12322
rect 17144 12306 17264 12322
rect 16580 12300 16712 12306
rect 16632 12294 16712 12300
rect 16580 12242 16632 12248
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16592 11762 16620 12106
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16684 10742 16712 12294
rect 17132 12300 17264 12306
rect 17184 12294 17264 12300
rect 17500 12300 17552 12306
rect 17132 12242 17184 12248
rect 17500 12242 17552 12248
rect 17144 11762 17172 12242
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17512 11694 17540 12242
rect 17604 11898 17632 12718
rect 17696 11898 17724 13262
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17972 11694 18000 15030
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18432 15014 18552 15030
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 18248 11218 18276 14962
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 17144 10810 17172 11154
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 17420 10606 17448 10950
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 16040 10266 16068 10542
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16132 9518 16160 10406
rect 17052 10266 17080 10542
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17144 9654 17172 10066
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16040 9178 16068 9454
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16224 9042 16252 9318
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 17038 8936 17094 8945
rect 17038 8871 17040 8880
rect 17092 8871 17094 8880
rect 17040 8842 17092 8848
rect 17236 8566 17264 10066
rect 17420 9518 17448 10406
rect 18064 10266 18092 11154
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 16224 7002 16252 7890
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7342 16436 7686
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16224 6458 16252 6802
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5778 16252 6054
rect 16316 5914 16344 6802
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6254 16436 6598
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16592 5370 16620 6734
rect 17236 5914 17264 7890
rect 17972 7886 18000 8842
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18064 7546 18092 10066
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18248 8634 18276 8978
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18248 6866 18276 7686
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 17420 6254 17448 6598
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 17420 5166 17448 6054
rect 18064 5914 18092 6190
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18156 5778 18184 6598
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 18340 4826 18368 14826
rect 18432 14550 18460 15014
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18432 14278 18460 14486
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18432 6730 18460 11018
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18524 4078 18552 14758
rect 18616 4554 18644 15846
rect 18800 14958 18828 15846
rect 18886 15804 19182 15824
rect 18942 15802 18966 15804
rect 19022 15802 19046 15804
rect 19102 15802 19126 15804
rect 18964 15750 18966 15802
rect 19028 15750 19040 15802
rect 19102 15750 19104 15802
rect 18942 15748 18966 15750
rect 19022 15748 19046 15750
rect 19102 15748 19126 15750
rect 18886 15728 19182 15748
rect 19352 15502 19380 16594
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 16182 19472 16390
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19536 16017 19564 16050
rect 19522 16008 19578 16017
rect 19522 15943 19578 15952
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19352 15026 19380 15438
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 18886 14716 19182 14736
rect 18942 14714 18966 14716
rect 19022 14714 19046 14716
rect 19102 14714 19126 14716
rect 18964 14662 18966 14714
rect 19028 14662 19040 14714
rect 19102 14662 19104 14714
rect 18942 14660 18966 14662
rect 19022 14660 19046 14662
rect 19102 14660 19126 14662
rect 18886 14640 19182 14660
rect 19444 14482 19472 14758
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19444 13870 19472 14418
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 18886 13628 19182 13648
rect 18942 13626 18966 13628
rect 19022 13626 19046 13628
rect 19102 13626 19126 13628
rect 18964 13574 18966 13626
rect 19028 13574 19040 13626
rect 19102 13574 19104 13626
rect 18942 13572 18966 13574
rect 19022 13572 19046 13574
rect 19102 13572 19126 13574
rect 18886 13552 19182 13572
rect 19444 13326 19472 13806
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 18886 12540 19182 12560
rect 18942 12538 18966 12540
rect 19022 12538 19046 12540
rect 19102 12538 19126 12540
rect 18964 12486 18966 12538
rect 19028 12486 19040 12538
rect 19102 12486 19104 12538
rect 18942 12484 18966 12486
rect 19022 12484 19046 12486
rect 19102 12484 19126 12486
rect 18886 12464 19182 12484
rect 19352 12374 19380 13262
rect 19432 13184 19484 13190
rect 19536 13172 19564 15943
rect 19628 15570 19656 17070
rect 19720 16046 19748 17682
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19708 16040 19760 16046
rect 19708 15982 19760 15988
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19628 14346 19656 15506
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19720 14482 19748 15302
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19812 13870 19840 17206
rect 21100 16998 21128 17682
rect 22388 17134 22416 17682
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23308 17134 23336 17478
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21284 16794 21312 16934
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21640 16040 21692 16046
rect 22100 16040 22152 16046
rect 21640 15982 21692 15988
rect 22098 16008 22100 16017
rect 22152 16008 22154 16017
rect 19904 15706 19932 15982
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19904 14958 19932 15642
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20824 15162 20852 15574
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19812 13326 19840 13806
rect 20732 13530 20760 15030
rect 20824 14958 20852 15098
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20824 14074 20852 14486
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20732 13326 20760 13466
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 19484 13144 19564 13172
rect 19800 13184 19852 13190
rect 19432 13126 19484 13132
rect 19800 13126 19852 13132
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11898 18920 12038
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 19536 11762 19564 12922
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 12306 19656 12718
rect 19708 12708 19760 12714
rect 19708 12650 19760 12656
rect 19720 12442 19748 12650
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19812 12306 19840 13126
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 20732 11830 20760 13262
rect 21008 12374 21036 13738
rect 21284 13394 21312 14010
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21560 12866 21588 15982
rect 21652 15910 21680 15982
rect 22098 15943 22154 15952
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 21744 15366 21772 15438
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21744 15094 21772 15302
rect 21732 15088 21784 15094
rect 21732 15030 21784 15036
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 22020 14550 22048 14826
rect 22008 14544 22060 14550
rect 22008 14486 22060 14492
rect 22204 14278 22232 15438
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22388 13530 22416 17070
rect 22572 16658 22784 16674
rect 22560 16652 22796 16658
rect 22612 16646 22744 16652
rect 22560 16594 22612 16600
rect 22744 16594 22796 16600
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23400 15366 23428 16594
rect 23952 15570 23980 18090
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 17678 25268 18022
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 24964 17338 24992 17614
rect 25424 17610 25452 20266
rect 25516 18970 25544 22374
rect 26424 21480 26476 21486
rect 26424 21422 26476 21428
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25700 20330 25728 21082
rect 26436 20398 26464 21422
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 26332 20392 26384 20398
rect 26332 20334 26384 20340
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 25688 20324 25740 20330
rect 25688 20266 25740 20272
rect 25884 19242 25912 20334
rect 26344 19854 26372 20334
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26528 19446 26556 22374
rect 26700 22092 26752 22098
rect 26700 22034 26752 22040
rect 26712 21894 26740 22034
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 26712 20806 26740 21830
rect 26804 21622 26832 26400
rect 27540 24426 27568 26400
rect 27852 25052 28148 25072
rect 27908 25050 27932 25052
rect 27988 25050 28012 25052
rect 28068 25050 28092 25052
rect 27930 24998 27932 25050
rect 27994 24998 28006 25050
rect 28068 24998 28070 25050
rect 27908 24996 27932 24998
rect 27988 24996 28012 24998
rect 28068 24996 28092 24998
rect 27852 24976 28148 24996
rect 27540 24410 27660 24426
rect 27540 24404 27672 24410
rect 27540 24398 27620 24404
rect 27620 24346 27672 24352
rect 27852 23964 28148 23984
rect 27908 23962 27932 23964
rect 27988 23962 28012 23964
rect 28068 23962 28092 23964
rect 27930 23910 27932 23962
rect 27994 23910 28006 23962
rect 28068 23910 28070 23962
rect 27908 23908 27932 23910
rect 27988 23908 28012 23910
rect 28068 23908 28092 23910
rect 27852 23888 28148 23908
rect 27632 23310 27936 23338
rect 27632 23254 27660 23310
rect 27620 23248 27672 23254
rect 27620 23190 27672 23196
rect 27908 23202 27936 23310
rect 27908 23186 28120 23202
rect 27804 23180 27856 23186
rect 27908 23180 28132 23186
rect 27908 23174 28080 23180
rect 27804 23122 27856 23128
rect 28080 23122 28132 23128
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27160 22568 27212 22574
rect 27160 22510 27212 22516
rect 27172 21894 27200 22510
rect 27632 21962 27660 23054
rect 27816 22964 27844 23122
rect 27724 22936 27844 22964
rect 28172 22976 28224 22982
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 26792 21616 26844 21622
rect 26792 21558 26844 21564
rect 27172 21486 27200 21830
rect 27724 21622 27752 22936
rect 28172 22918 28224 22924
rect 27852 22876 28148 22896
rect 27908 22874 27932 22876
rect 27988 22874 28012 22876
rect 28068 22874 28092 22876
rect 27930 22822 27932 22874
rect 27994 22822 28006 22874
rect 28068 22822 28070 22874
rect 27908 22820 27932 22822
rect 27988 22820 28012 22822
rect 28068 22820 28092 22822
rect 27852 22800 28148 22820
rect 28184 22642 28212 22918
rect 28276 22710 28304 26400
rect 28632 23520 28684 23526
rect 28632 23462 28684 23468
rect 28264 22704 28316 22710
rect 28264 22646 28316 22652
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 28262 22536 28318 22545
rect 28172 22500 28224 22506
rect 28262 22471 28264 22480
rect 28172 22442 28224 22448
rect 28316 22471 28318 22480
rect 28264 22442 28316 22448
rect 28184 22098 28212 22442
rect 28356 22432 28408 22438
rect 28356 22374 28408 22380
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 27852 21788 28148 21808
rect 27908 21786 27932 21788
rect 27988 21786 28012 21788
rect 28068 21786 28092 21788
rect 27930 21734 27932 21786
rect 27994 21734 28006 21786
rect 28068 21734 28070 21786
rect 27908 21732 27932 21734
rect 27988 21732 28012 21734
rect 28068 21732 28092 21734
rect 27852 21712 28148 21732
rect 28276 21690 28304 21966
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 27160 21480 27212 21486
rect 27160 21422 27212 21428
rect 27816 21350 27844 21490
rect 28368 21457 28396 22374
rect 28354 21448 28410 21457
rect 28354 21383 28410 21392
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 26792 21072 26844 21078
rect 26792 21014 26844 21020
rect 26882 21040 26938 21049
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26516 19440 26568 19446
rect 26516 19382 26568 19388
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25516 18834 25544 18906
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25516 18290 25544 18770
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25976 18222 26004 18702
rect 25964 18216 26016 18222
rect 25964 18158 26016 18164
rect 25780 17808 25832 17814
rect 25778 17776 25780 17785
rect 25832 17776 25834 17785
rect 25778 17711 25834 17720
rect 25412 17604 25464 17610
rect 25412 17546 25464 17552
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24596 16658 24624 16934
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24412 16561 24440 16594
rect 24398 16552 24454 16561
rect 24398 16487 24454 16496
rect 24596 16114 24624 16594
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24688 16046 24716 16662
rect 25332 16522 25360 17070
rect 25962 16552 26018 16561
rect 25320 16516 25372 16522
rect 26252 16522 26280 17070
rect 26528 16658 26556 19382
rect 26712 18630 26740 20742
rect 26804 20534 26832 21014
rect 26882 20975 26884 20984
rect 26936 20975 26938 20984
rect 26884 20946 26936 20952
rect 28644 20806 28672 23462
rect 28816 22432 28868 22438
rect 28816 22374 28868 22380
rect 28828 21486 28856 22374
rect 29012 22114 29040 26400
rect 29748 24290 29776 26400
rect 30392 24410 30420 26400
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 31128 24290 31156 26400
rect 29748 24262 29868 24290
rect 31128 24262 31248 24290
rect 29368 24064 29420 24070
rect 29368 24006 29420 24012
rect 29380 23730 29408 24006
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29276 23112 29328 23118
rect 29276 23054 29328 23060
rect 29288 22574 29316 23054
rect 29380 22982 29408 23666
rect 29552 23656 29604 23662
rect 29552 23598 29604 23604
rect 29564 22982 29592 23598
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 29552 22976 29604 22982
rect 29552 22918 29604 22924
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 29092 22228 29144 22234
rect 29144 22188 29224 22216
rect 29092 22170 29144 22176
rect 29012 22086 29132 22114
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 29012 21706 29040 21966
rect 29104 21894 29132 22086
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 29012 21678 29132 21706
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28906 21448 28962 21457
rect 28724 21072 28776 21078
rect 28722 21040 28724 21049
rect 28776 21040 28778 21049
rect 28722 20975 28778 20984
rect 28632 20800 28684 20806
rect 28632 20742 28684 20748
rect 27852 20700 28148 20720
rect 27908 20698 27932 20700
rect 27988 20698 28012 20700
rect 28068 20698 28092 20700
rect 27930 20646 27932 20698
rect 27994 20646 28006 20698
rect 28068 20646 28070 20698
rect 27908 20644 27932 20646
rect 27988 20644 28012 20646
rect 28068 20644 28092 20646
rect 27852 20624 28148 20644
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 26792 20528 26844 20534
rect 26988 20505 27016 20538
rect 26792 20470 26844 20476
rect 26974 20496 27030 20505
rect 28644 20466 28672 20742
rect 26974 20431 27030 20440
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 27724 19990 27752 20402
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27712 19848 27764 19854
rect 27712 19790 27764 19796
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27356 19394 27384 19450
rect 27356 19378 27660 19394
rect 27356 19372 27672 19378
rect 27356 19366 27620 19372
rect 27620 19314 27672 19320
rect 27724 19242 27752 19790
rect 27852 19612 28148 19632
rect 27908 19610 27932 19612
rect 27988 19610 28012 19612
rect 28068 19610 28092 19612
rect 27930 19558 27932 19610
rect 27994 19558 28006 19610
rect 28068 19558 28070 19610
rect 27908 19556 27932 19558
rect 27988 19556 28012 19558
rect 28068 19556 28092 19558
rect 27852 19536 28148 19556
rect 27804 19440 27856 19446
rect 27802 19408 27804 19417
rect 27856 19408 27858 19417
rect 27802 19343 27858 19352
rect 27712 19236 27764 19242
rect 27712 19178 27764 19184
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 26700 18624 26752 18630
rect 26700 18566 26752 18572
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 26608 18148 26660 18154
rect 26608 18090 26660 18096
rect 26976 18148 27028 18154
rect 26976 18090 27028 18096
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 25962 16487 26018 16496
rect 26240 16516 26292 16522
rect 25320 16458 25372 16464
rect 25976 16454 26004 16487
rect 26240 16458 26292 16464
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23952 15366 23980 15506
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23400 14958 23428 15302
rect 23388 14952 23440 14958
rect 23388 14894 23440 14900
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22940 14482 22968 14758
rect 23400 14550 23428 14894
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22756 14006 22784 14214
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22756 12986 22784 13806
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 21560 12838 21680 12866
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 20732 11694 20760 11766
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20904 11620 20956 11626
rect 20904 11562 20956 11568
rect 18886 11452 19182 11472
rect 18942 11450 18966 11452
rect 19022 11450 19046 11452
rect 19102 11450 19126 11452
rect 18964 11398 18966 11450
rect 19028 11398 19040 11450
rect 19102 11398 19104 11450
rect 18942 11396 18966 11398
rect 19022 11396 19046 11398
rect 19102 11396 19126 11398
rect 18886 11376 19182 11396
rect 20916 11218 20944 11562
rect 21100 11354 21128 12242
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 18984 10606 19012 10950
rect 19996 10606 20024 10950
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 18886 10364 19182 10384
rect 18942 10362 18966 10364
rect 19022 10362 19046 10364
rect 19102 10362 19126 10364
rect 18964 10310 18966 10362
rect 19028 10310 19040 10362
rect 19102 10310 19104 10362
rect 18942 10308 18966 10310
rect 19022 10308 19046 10310
rect 19102 10308 19126 10310
rect 18886 10288 19182 10308
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 18886 9276 19182 9296
rect 18942 9274 18966 9276
rect 19022 9274 19046 9276
rect 19102 9274 19126 9276
rect 18964 9222 18966 9274
rect 19028 9222 19040 9274
rect 19102 9222 19104 9274
rect 18942 9220 18966 9222
rect 19022 9220 19046 9222
rect 19102 9220 19126 9222
rect 18886 9200 19182 9220
rect 19260 9042 19288 9318
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8430 19012 8774
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18800 7342 18828 8230
rect 18886 8188 19182 8208
rect 18942 8186 18966 8188
rect 19022 8186 19046 8188
rect 19102 8186 19126 8188
rect 18964 8134 18966 8186
rect 19028 8134 19040 8186
rect 19102 8134 19104 8186
rect 18942 8132 18966 8134
rect 19022 8132 19046 8134
rect 19102 8132 19126 8134
rect 18886 8112 19182 8132
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18696 7200 18748 7206
rect 18892 7188 18920 7278
rect 18696 7142 18748 7148
rect 18800 7160 18920 7188
rect 19340 7200 19392 7206
rect 18708 6798 18736 7142
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18800 5370 18828 7160
rect 19340 7142 19392 7148
rect 18886 7100 19182 7120
rect 18942 7098 18966 7100
rect 19022 7098 19046 7100
rect 19102 7098 19126 7100
rect 18964 7046 18966 7098
rect 19028 7046 19040 7098
rect 19102 7046 19104 7098
rect 18942 7044 18966 7046
rect 19022 7044 19046 7046
rect 19102 7044 19126 7046
rect 18886 7024 19182 7044
rect 19352 6254 19380 7142
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 18886 6012 19182 6032
rect 18942 6010 18966 6012
rect 19022 6010 19046 6012
rect 19102 6010 19126 6012
rect 18964 5958 18966 6010
rect 19028 5958 19040 6010
rect 19102 5958 19104 6010
rect 18942 5956 18966 5958
rect 19022 5956 19046 5958
rect 19102 5956 19126 5958
rect 18886 5936 19182 5956
rect 19260 5778 19288 6054
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18886 4924 19182 4944
rect 18942 4922 18966 4924
rect 19022 4922 19046 4924
rect 19102 4922 19126 4924
rect 18964 4870 18966 4922
rect 19028 4870 19040 4922
rect 19102 4870 19104 4922
rect 18942 4868 18966 4870
rect 19022 4868 19046 4870
rect 19102 4868 19126 4870
rect 18886 4848 19182 4868
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18604 4548 18656 4554
rect 18604 4490 18656 4496
rect 19076 4282 19104 4626
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 16592 3738 16620 4014
rect 18886 3836 19182 3856
rect 18942 3834 18966 3836
rect 19022 3834 19046 3836
rect 19102 3834 19126 3836
rect 18964 3782 18966 3834
rect 19028 3782 19040 3834
rect 19102 3782 19104 3834
rect 18942 3780 18966 3782
rect 19022 3780 19046 3782
rect 19102 3780 19126 3782
rect 18886 3760 19182 3780
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 19444 3670 19472 10406
rect 20088 10266 20116 11154
rect 21560 10810 21588 12718
rect 21652 11626 21680 12838
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22020 11830 22048 12174
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20272 10130 20300 10406
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19996 8634 20024 9454
rect 20088 9178 20116 10066
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20272 9042 20300 9318
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20640 8430 20668 9862
rect 21744 9518 21772 11494
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 10130 21864 10406
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20732 8566 20760 9386
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 19996 8090 20024 8366
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19720 7546 19748 7890
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19996 7342 20024 7686
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19904 5166 19932 6054
rect 20088 5914 20116 6802
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20272 5778 20300 7142
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20824 5302 20852 9454
rect 21928 9178 21956 11630
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10266 22048 10542
rect 22112 10266 22140 11154
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22020 8430 22048 9318
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22388 8090 22416 11154
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 21008 7002 21036 7278
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21008 6254 21036 6598
rect 20996 6248 21048 6254
rect 20996 6190 21048 6196
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20824 4078 20852 4422
rect 21008 4078 21036 6054
rect 21836 5370 21864 7890
rect 22480 5914 22508 12718
rect 23492 12306 23520 12922
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 23020 11076 23072 11082
rect 23020 11018 23072 11024
rect 22572 10606 22600 11018
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22848 9654 22876 10066
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 23032 9518 23060 11018
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22848 9042 22876 9318
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 23032 7546 23060 8366
rect 23124 8090 23152 8978
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23308 7954 23336 8230
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 22572 6458 22600 6802
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22664 5778 22692 7142
rect 22756 7002 22784 7278
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 23768 6866 23796 12582
rect 23952 12102 23980 15302
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 24044 14618 24072 15098
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 24228 13462 24256 13806
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 24044 12646 24072 12718
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23952 10606 23980 10950
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 7954 24072 8774
rect 24136 8090 24164 11154
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24228 9178 24256 10066
rect 24216 9172 24268 9178
rect 24216 9114 24268 9120
rect 24320 9042 24348 10406
rect 24308 9036 24360 9042
rect 24308 8978 24360 8984
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22756 6254 22784 6598
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 22848 5930 22876 6394
rect 22756 5914 22876 5930
rect 22744 5908 22876 5914
rect 22796 5902 22876 5908
rect 22744 5850 22796 5856
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21836 4690 21864 4966
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 22204 4010 22232 5034
rect 22296 4826 22324 5102
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19812 3602 19840 3878
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 9921 3292 10217 3312
rect 9977 3290 10001 3292
rect 10057 3290 10081 3292
rect 10137 3290 10161 3292
rect 9999 3238 10001 3290
rect 10063 3238 10075 3290
rect 10137 3238 10139 3290
rect 9977 3236 10001 3238
rect 10057 3236 10081 3238
rect 10137 3236 10161 3238
rect 9921 3216 10217 3236
rect 21928 2990 21956 3878
rect 22756 3602 22784 4422
rect 22848 4282 22876 4626
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22940 3466 22968 5578
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23400 3738 23428 5102
rect 23492 4826 23520 6734
rect 23860 5778 23888 7414
rect 24412 5914 24440 14758
rect 24688 12646 24716 15982
rect 24768 15428 24820 15434
rect 24768 15370 24820 15376
rect 24780 13870 24808 15370
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 24964 13938 24992 14894
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24780 11286 24808 11630
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24596 9518 24624 9862
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24596 7002 24624 7278
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 24872 6866 24900 13874
rect 25056 13818 25084 14418
rect 25148 14074 25176 14894
rect 25884 14618 25912 15030
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 26252 14278 26280 15982
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 24964 13790 25084 13818
rect 24964 13530 24992 13790
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 24964 12782 24992 13466
rect 25240 13394 25268 14214
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 25056 12374 25084 13330
rect 25136 12708 25188 12714
rect 25136 12650 25188 12656
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 25148 12306 25176 12650
rect 25424 12306 25452 13806
rect 25688 13456 25740 13462
rect 25688 13398 25740 13404
rect 25700 12850 25728 13398
rect 26252 13394 26280 14214
rect 26436 14074 26464 15982
rect 26620 14958 26648 18090
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 26528 14482 26556 14758
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26528 13870 26556 14418
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26896 13462 26924 16390
rect 26884 13456 26936 13462
rect 26884 13398 26936 13404
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26056 12912 26108 12918
rect 26056 12854 26108 12860
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11218 24992 12038
rect 25148 11694 25176 12242
rect 26068 12170 26096 12854
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26436 12442 26464 12718
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26804 12306 26832 12718
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 26056 12164 26108 12170
rect 26056 12106 26108 12112
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25240 8090 25268 10746
rect 25608 10606 25636 11494
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25608 9654 25636 10066
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25700 9518 25728 11290
rect 26068 11286 26096 12106
rect 26252 11694 26280 12242
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26056 11280 26108 11286
rect 26056 11222 26108 11228
rect 26252 10810 26280 11630
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 26160 8430 26188 8774
rect 26252 8498 26280 9862
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26344 9042 26372 9318
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26620 8634 26648 9454
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 26332 8560 26384 8566
rect 26332 8502 26384 8508
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 26148 8424 26200 8430
rect 26148 8366 26200 8372
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 26344 7954 26372 8502
rect 26332 7948 26384 7954
rect 26332 7890 26384 7896
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24872 5778 24900 6598
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23676 4758 23704 5510
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 23860 4078 23888 5578
rect 24492 5024 24544 5030
rect 24492 4966 24544 4972
rect 24504 4690 24532 4966
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 24504 3602 24532 3878
rect 24780 3738 24808 5646
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24964 4826 24992 5102
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 25056 3670 25084 7278
rect 26424 6860 26476 6866
rect 26424 6802 26476 6808
rect 25596 6248 25648 6254
rect 25596 6190 25648 6196
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25608 5914 25636 6190
rect 25596 5908 25648 5914
rect 25596 5850 25648 5856
rect 25700 5370 25728 6190
rect 25872 6112 25924 6118
rect 25872 6054 25924 6060
rect 25884 5778 25912 6054
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25688 5364 25740 5370
rect 25688 5306 25740 5312
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25516 4146 25544 4966
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 25596 4480 25648 4486
rect 25596 4422 25648 4428
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 25608 4078 25636 4422
rect 25596 4072 25648 4078
rect 25596 4014 25648 4020
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25044 3664 25096 3670
rect 25044 3606 25096 3612
rect 25516 3602 25544 3878
rect 26252 3602 26280 4422
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 25964 3392 26016 3398
rect 25964 3334 26016 3340
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 18886 2748 19182 2768
rect 18942 2746 18966 2748
rect 19022 2746 19046 2748
rect 19102 2746 19126 2748
rect 18964 2694 18966 2746
rect 19028 2694 19040 2746
rect 19102 2694 19104 2746
rect 18942 2692 18966 2694
rect 19022 2692 19046 2694
rect 19102 2692 19126 2694
rect 18886 2672 19182 2692
rect 20916 2650 20944 2926
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 22848 2514 22876 3062
rect 24964 2990 24992 3334
rect 25976 2990 26004 3334
rect 26344 3194 26372 4558
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 26436 3058 26464 6802
rect 26988 6798 27016 18090
rect 27160 17060 27212 17066
rect 27160 17002 27212 17008
rect 27172 16658 27200 17002
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27080 16114 27108 16390
rect 27356 16250 27384 18566
rect 27852 18524 28148 18544
rect 27908 18522 27932 18524
rect 27988 18522 28012 18524
rect 28068 18522 28092 18524
rect 27930 18470 27932 18522
rect 27994 18470 28006 18522
rect 28068 18470 28070 18522
rect 27908 18468 27932 18470
rect 27988 18468 28012 18470
rect 28068 18468 28092 18470
rect 27852 18448 28148 18468
rect 28264 18148 28316 18154
rect 28264 18090 28316 18096
rect 27436 18080 27488 18086
rect 27436 18022 27488 18028
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27448 15026 27476 18022
rect 27852 17436 28148 17456
rect 27908 17434 27932 17436
rect 27988 17434 28012 17436
rect 28068 17434 28092 17436
rect 27930 17382 27932 17434
rect 27994 17382 28006 17434
rect 28068 17382 28070 17434
rect 27908 17380 27932 17382
rect 27988 17380 28012 17382
rect 28068 17380 28092 17382
rect 27852 17360 28148 17380
rect 27620 17060 27672 17066
rect 27620 17002 27672 17008
rect 27632 15586 27660 17002
rect 28276 16998 28304 18090
rect 28368 17338 28396 18770
rect 28828 18086 28856 21422
rect 28906 21383 28908 21392
rect 28960 21383 28962 21392
rect 28908 21354 28960 21360
rect 29000 21072 29052 21078
rect 29104 21060 29132 21678
rect 29052 21032 29132 21060
rect 29000 21014 29052 21020
rect 28908 20324 28960 20330
rect 28908 20266 28960 20272
rect 28920 18154 28948 20266
rect 29012 19990 29040 21014
rect 29000 19984 29052 19990
rect 29000 19926 29052 19932
rect 29012 19854 29040 19926
rect 29196 19854 29224 22188
rect 29380 22030 29408 22918
rect 29460 22500 29512 22506
rect 29460 22442 29512 22448
rect 29472 22234 29500 22442
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 29368 22024 29420 22030
rect 29368 21966 29420 21972
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29748 21486 29776 21830
rect 29736 21480 29788 21486
rect 29736 21422 29788 21428
rect 29840 21010 29868 24262
rect 30748 24064 30800 24070
rect 30748 24006 30800 24012
rect 30760 23730 30788 24006
rect 30748 23724 30800 23730
rect 30748 23666 30800 23672
rect 30748 23180 30800 23186
rect 30748 23122 30800 23128
rect 30760 21350 30788 23122
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31036 21486 31064 21966
rect 31024 21480 31076 21486
rect 31024 21422 31076 21428
rect 31116 21480 31168 21486
rect 31116 21422 31168 21428
rect 30748 21344 30800 21350
rect 30748 21286 30800 21292
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 30208 20534 30236 20946
rect 30196 20528 30248 20534
rect 30196 20470 30248 20476
rect 30760 20058 30788 20946
rect 30472 20052 30524 20058
rect 30472 19994 30524 20000
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 29184 19848 29236 19854
rect 29184 19790 29236 19796
rect 29196 18970 29224 19790
rect 30484 19514 30512 19994
rect 30472 19508 30524 19514
rect 30472 19450 30524 19456
rect 30760 19310 30788 19994
rect 30944 19922 30972 21286
rect 31128 21078 31156 21422
rect 31116 21072 31168 21078
rect 31116 21014 31168 21020
rect 31220 20466 31248 24262
rect 31484 24268 31536 24274
rect 31484 24210 31536 24216
rect 31496 22778 31524 24210
rect 31864 23866 31892 26400
rect 32220 24200 32272 24206
rect 32220 24142 32272 24148
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32232 23866 32260 24142
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 32220 23860 32272 23866
rect 32220 23802 32272 23808
rect 32324 23662 32352 24142
rect 32312 23656 32364 23662
rect 32312 23598 32364 23604
rect 31576 23520 31628 23526
rect 31576 23462 31628 23468
rect 31588 23118 31616 23462
rect 32600 23322 32628 26400
rect 33336 24410 33364 26400
rect 33324 24404 33376 24410
rect 33324 24346 33376 24352
rect 33692 24200 33744 24206
rect 33692 24142 33744 24148
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 32496 23316 32548 23322
rect 32496 23258 32548 23264
rect 32588 23316 32640 23322
rect 32588 23258 32640 23264
rect 33232 23316 33284 23322
rect 33232 23258 33284 23264
rect 32128 23180 32180 23186
rect 32128 23122 32180 23128
rect 31576 23112 31628 23118
rect 31576 23054 31628 23060
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 31588 22710 31616 23054
rect 31576 22704 31628 22710
rect 31576 22646 31628 22652
rect 32140 22642 32168 23122
rect 32508 23089 32536 23258
rect 32494 23080 32550 23089
rect 32494 23015 32550 23024
rect 32220 22976 32272 22982
rect 32220 22918 32272 22924
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32232 22438 32260 22918
rect 32312 22500 32364 22506
rect 32312 22442 32364 22448
rect 32220 22432 32272 22438
rect 32220 22374 32272 22380
rect 32036 20936 32088 20942
rect 32036 20878 32088 20884
rect 31208 20460 31260 20466
rect 31208 20402 31260 20408
rect 32048 20398 32076 20878
rect 32036 20392 32088 20398
rect 32036 20334 32088 20340
rect 31116 20256 31168 20262
rect 31116 20198 31168 20204
rect 31128 20058 31156 20198
rect 32324 20058 32352 22442
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32784 21622 32812 21966
rect 32772 21616 32824 21622
rect 32772 21558 32824 21564
rect 32404 20392 32456 20398
rect 32404 20334 32456 20340
rect 31116 20052 31168 20058
rect 31116 19994 31168 20000
rect 32220 20052 32272 20058
rect 32220 19994 32272 20000
rect 32312 20052 32364 20058
rect 32312 19994 32364 20000
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 31300 19916 31352 19922
rect 31300 19858 31352 19864
rect 31312 19310 31340 19858
rect 32232 19514 32260 19994
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 32324 19310 32352 19994
rect 30012 19304 30064 19310
rect 30012 19246 30064 19252
rect 30748 19304 30800 19310
rect 30748 19246 30800 19252
rect 31116 19304 31168 19310
rect 31116 19246 31168 19252
rect 31300 19304 31352 19310
rect 31300 19246 31352 19252
rect 31392 19304 31444 19310
rect 31392 19246 31444 19252
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 29920 18964 29972 18970
rect 29920 18906 29972 18912
rect 29932 18834 29960 18906
rect 30024 18834 30052 19246
rect 29920 18828 29972 18834
rect 29920 18770 29972 18776
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 29366 18728 29422 18737
rect 29366 18663 29422 18672
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29012 18290 29040 18566
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 28908 18148 28960 18154
rect 28908 18090 28960 18096
rect 29000 18148 29052 18154
rect 29000 18090 29052 18096
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28724 17740 28776 17746
rect 28828 17728 28856 18022
rect 28776 17700 28856 17728
rect 28724 17682 28776 17688
rect 29012 17610 29040 18090
rect 29288 17882 29316 18566
rect 29380 18426 29408 18663
rect 30024 18465 30052 18770
rect 30010 18456 30066 18465
rect 29368 18420 29420 18426
rect 30010 18391 30066 18400
rect 29368 18362 29420 18368
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29656 17814 29684 18226
rect 30012 17876 30064 17882
rect 30012 17818 30064 17824
rect 29644 17808 29696 17814
rect 29644 17750 29696 17756
rect 29460 17740 29512 17746
rect 29460 17682 29512 17688
rect 29000 17604 29052 17610
rect 29000 17546 29052 17552
rect 28632 17536 28684 17542
rect 28630 17504 28632 17513
rect 28908 17536 28960 17542
rect 28684 17504 28686 17513
rect 28630 17439 28686 17448
rect 28906 17504 28908 17513
rect 28960 17504 28962 17513
rect 28906 17439 28962 17448
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28448 17332 28500 17338
rect 28448 17274 28500 17280
rect 28460 17134 28488 17274
rect 28448 17128 28500 17134
rect 28448 17070 28500 17076
rect 28540 17128 28592 17134
rect 28540 17070 28592 17076
rect 28264 16992 28316 16998
rect 28264 16934 28316 16940
rect 28552 16794 28580 17070
rect 28644 16794 28672 17439
rect 29472 17202 29500 17682
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29276 17196 29328 17202
rect 29276 17138 29328 17144
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29000 17060 29052 17066
rect 29000 17002 29052 17008
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 29012 16726 29040 17002
rect 29000 16720 29052 16726
rect 29000 16662 29052 16668
rect 27712 16652 27764 16658
rect 27712 16594 27764 16600
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 27540 15558 27660 15586
rect 27540 15162 27568 15558
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27540 14618 27568 14894
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 27632 14482 27660 15438
rect 27620 14476 27672 14482
rect 27620 14418 27672 14424
rect 27632 13394 27660 14418
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 27252 12776 27304 12782
rect 27252 12718 27304 12724
rect 27264 11694 27292 12718
rect 27724 12714 27752 16594
rect 27852 16348 28148 16368
rect 27908 16346 27932 16348
rect 27988 16346 28012 16348
rect 28068 16346 28092 16348
rect 27930 16294 27932 16346
rect 27994 16294 28006 16346
rect 28068 16294 28070 16346
rect 27908 16292 27932 16294
rect 27988 16292 28012 16294
rect 28068 16292 28092 16294
rect 27852 16272 28148 16292
rect 28920 16250 28948 16594
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 29012 15706 29040 16662
rect 29288 16522 29316 17138
rect 29644 17128 29696 17134
rect 29644 17070 29696 17076
rect 29656 16946 29684 17070
rect 29472 16918 29684 16946
rect 29472 16658 29500 16918
rect 29748 16658 29776 17478
rect 29826 17368 29882 17377
rect 29826 17303 29828 17312
rect 29880 17303 29882 17312
rect 29920 17332 29972 17338
rect 29828 17274 29880 17280
rect 29920 17274 29972 17280
rect 29932 17134 29960 17274
rect 30024 17202 30052 17818
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30392 17202 30420 17614
rect 30012 17196 30064 17202
rect 30012 17138 30064 17144
rect 30380 17196 30432 17202
rect 30380 17138 30432 17144
rect 31128 17134 31156 19246
rect 31404 18426 31432 19246
rect 31944 19236 31996 19242
rect 31944 19178 31996 19184
rect 31758 18592 31814 18601
rect 31758 18527 31814 18536
rect 31392 18420 31444 18426
rect 31392 18362 31444 18368
rect 31772 18222 31800 18527
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 31760 18216 31812 18222
rect 31760 18158 31812 18164
rect 31220 17814 31248 18158
rect 31208 17808 31260 17814
rect 31208 17750 31260 17756
rect 31956 17338 31984 19178
rect 32416 19174 32444 20334
rect 32784 19922 32812 21558
rect 33244 21010 33272 23258
rect 33336 23050 33364 23598
rect 33416 23588 33468 23594
rect 33416 23530 33468 23536
rect 33428 23186 33456 23530
rect 33416 23180 33468 23186
rect 33416 23122 33468 23128
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 33336 22778 33364 22986
rect 33324 22772 33376 22778
rect 33324 22714 33376 22720
rect 33428 22506 33456 23122
rect 33704 22778 33732 24142
rect 33784 23656 33836 23662
rect 33784 23598 33836 23604
rect 33692 22772 33744 22778
rect 33692 22714 33744 22720
rect 33508 22568 33560 22574
rect 33508 22510 33560 22516
rect 33416 22500 33468 22506
rect 33416 22442 33468 22448
rect 33520 22166 33548 22510
rect 33508 22160 33560 22166
rect 33508 22102 33560 22108
rect 33796 21486 33824 23598
rect 33980 22098 34008 26400
rect 34716 24410 34744 26400
rect 34980 24812 35032 24818
rect 34980 24754 35032 24760
rect 34704 24404 34756 24410
rect 34704 24346 34756 24352
rect 34244 23724 34296 23730
rect 34244 23666 34296 23672
rect 34256 22982 34284 23666
rect 34992 23662 35020 24754
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 34980 23656 35032 23662
rect 34980 23598 35032 23604
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34532 23050 34560 23462
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34244 22976 34296 22982
rect 34244 22918 34296 22924
rect 34532 22778 34560 22986
rect 35084 22778 35112 24142
rect 35164 23520 35216 23526
rect 35164 23462 35216 23468
rect 35176 23186 35204 23462
rect 35164 23180 35216 23186
rect 35164 23122 35216 23128
rect 35452 23118 35480 26400
rect 35900 24268 35952 24274
rect 35900 24210 35952 24216
rect 35912 23866 35940 24210
rect 36188 23882 36216 26400
rect 36924 24698 36952 26400
rect 36924 24670 37228 24698
rect 36817 24508 37113 24528
rect 36873 24506 36897 24508
rect 36953 24506 36977 24508
rect 37033 24506 37057 24508
rect 36895 24454 36897 24506
rect 36959 24454 36971 24506
rect 37033 24454 37035 24506
rect 36873 24452 36897 24454
rect 36953 24452 36977 24454
rect 37033 24452 37057 24454
rect 36817 24432 37113 24452
rect 36188 23866 36308 23882
rect 35900 23860 35952 23866
rect 36188 23860 36320 23866
rect 36188 23854 36268 23860
rect 35900 23802 35952 23808
rect 36268 23802 36320 23808
rect 36360 23656 36412 23662
rect 36360 23598 36412 23604
rect 35440 23112 35492 23118
rect 35440 23054 35492 23060
rect 36372 22982 36400 23598
rect 36817 23420 37113 23440
rect 36873 23418 36897 23420
rect 36953 23418 36977 23420
rect 37033 23418 37057 23420
rect 36895 23366 36897 23418
rect 36959 23366 36971 23418
rect 37033 23366 37035 23418
rect 36873 23364 36897 23366
rect 36953 23364 36977 23366
rect 37033 23364 37057 23366
rect 36817 23344 37113 23364
rect 36360 22976 36412 22982
rect 36360 22918 36412 22924
rect 34520 22772 34572 22778
rect 34520 22714 34572 22720
rect 35072 22772 35124 22778
rect 35072 22714 35124 22720
rect 37200 22642 37228 24670
rect 37372 23588 37424 23594
rect 37372 23530 37424 23536
rect 37384 23254 37412 23530
rect 37660 23254 37688 26400
rect 37372 23248 37424 23254
rect 37372 23190 37424 23196
rect 37648 23248 37700 23254
rect 37648 23190 37700 23196
rect 37280 23044 37332 23050
rect 37280 22986 37332 22992
rect 37188 22636 37240 22642
rect 37188 22578 37240 22584
rect 37292 22506 37320 22986
rect 37384 22778 37412 23190
rect 38108 23112 38160 23118
rect 38108 23054 38160 23060
rect 37372 22772 37424 22778
rect 37372 22714 37424 22720
rect 37740 22772 37792 22778
rect 37740 22714 37792 22720
rect 37752 22574 37780 22714
rect 37740 22568 37792 22574
rect 37740 22510 37792 22516
rect 37280 22500 37332 22506
rect 37280 22442 37332 22448
rect 36817 22332 37113 22352
rect 36873 22330 36897 22332
rect 36953 22330 36977 22332
rect 37033 22330 37057 22332
rect 36895 22278 36897 22330
rect 36959 22278 36971 22330
rect 37033 22278 37035 22330
rect 36873 22276 36897 22278
rect 36953 22276 36977 22278
rect 37033 22276 37057 22278
rect 36817 22256 37113 22276
rect 33968 22092 34020 22098
rect 33968 22034 34020 22040
rect 34152 22092 34204 22098
rect 34152 22034 34204 22040
rect 34888 22092 34940 22098
rect 34888 22034 34940 22040
rect 33784 21480 33836 21486
rect 33784 21422 33836 21428
rect 34164 21010 34192 22034
rect 34900 21622 34928 22034
rect 35624 21888 35676 21894
rect 35624 21830 35676 21836
rect 34888 21616 34940 21622
rect 34888 21558 34940 21564
rect 35636 21486 35664 21830
rect 35348 21480 35400 21486
rect 35348 21422 35400 21428
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 35992 21480 36044 21486
rect 35992 21422 36044 21428
rect 35360 21146 35388 21422
rect 36004 21146 36032 21422
rect 37188 21412 37240 21418
rect 37188 21354 37240 21360
rect 36817 21244 37113 21264
rect 36873 21242 36897 21244
rect 36953 21242 36977 21244
rect 37033 21242 37057 21244
rect 36895 21190 36897 21242
rect 36959 21190 36971 21242
rect 37033 21190 37035 21242
rect 36873 21188 36897 21190
rect 36953 21188 36977 21190
rect 37033 21188 37057 21190
rect 36817 21168 37113 21188
rect 35348 21140 35400 21146
rect 35348 21082 35400 21088
rect 35992 21140 36044 21146
rect 35992 21082 36044 21088
rect 36452 21140 36504 21146
rect 36452 21082 36504 21088
rect 34796 21072 34848 21078
rect 34796 21014 34848 21020
rect 33232 21004 33284 21010
rect 33232 20946 33284 20952
rect 34152 21004 34204 21010
rect 34152 20946 34204 20952
rect 34808 20942 34836 21014
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 33232 20324 33284 20330
rect 33232 20266 33284 20272
rect 33244 19922 33272 20266
rect 34808 19990 34836 20878
rect 34796 19984 34848 19990
rect 34796 19926 34848 19932
rect 32772 19916 32824 19922
rect 32772 19858 32824 19864
rect 33232 19916 33284 19922
rect 33232 19858 33284 19864
rect 35360 19854 35388 21082
rect 36176 20868 36228 20874
rect 36176 20810 36228 20816
rect 35808 20800 35860 20806
rect 35808 20742 35860 20748
rect 35820 20466 35848 20742
rect 35808 20460 35860 20466
rect 35808 20402 35860 20408
rect 35900 20256 35952 20262
rect 35900 20198 35952 20204
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 32588 19780 32640 19786
rect 32588 19722 32640 19728
rect 32404 19168 32456 19174
rect 32404 19110 32456 19116
rect 32402 18864 32458 18873
rect 32312 18828 32364 18834
rect 32402 18799 32404 18808
rect 32312 18770 32364 18776
rect 32456 18799 32458 18808
rect 32404 18770 32456 18776
rect 32324 18601 32352 18770
rect 32310 18592 32366 18601
rect 32310 18527 32366 18536
rect 32416 18426 32444 18770
rect 32404 18420 32456 18426
rect 32404 18362 32456 18368
rect 32128 18352 32180 18358
rect 32128 18294 32180 18300
rect 32140 18204 32168 18294
rect 32416 18290 32444 18362
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32312 18216 32364 18222
rect 32140 18176 32312 18204
rect 32312 18158 32364 18164
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 31116 17128 31168 17134
rect 31116 17070 31168 17076
rect 30470 16688 30526 16697
rect 29460 16652 29512 16658
rect 29460 16594 29512 16600
rect 29552 16652 29604 16658
rect 29552 16594 29604 16600
rect 29736 16652 29788 16658
rect 30470 16623 30472 16632
rect 29736 16594 29788 16600
rect 30524 16623 30526 16632
rect 30472 16594 30524 16600
rect 29276 16516 29328 16522
rect 29276 16458 29328 16464
rect 29564 16046 29592 16594
rect 31128 16046 31156 17070
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 31116 16040 31168 16046
rect 31116 15982 31168 15988
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 27852 15260 28148 15280
rect 27908 15258 27932 15260
rect 27988 15258 28012 15260
rect 28068 15258 28092 15260
rect 27930 15206 27932 15258
rect 27994 15206 28006 15258
rect 28068 15206 28070 15258
rect 27908 15204 27932 15206
rect 27988 15204 28012 15206
rect 28068 15204 28092 15206
rect 27852 15184 28148 15204
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 27852 14172 28148 14192
rect 27908 14170 27932 14172
rect 27988 14170 28012 14172
rect 28068 14170 28092 14172
rect 27930 14118 27932 14170
rect 27994 14118 28006 14170
rect 28068 14118 28070 14170
rect 27908 14116 27932 14118
rect 27988 14116 28012 14118
rect 28068 14116 28092 14118
rect 27852 14096 28148 14116
rect 28276 14074 28304 14350
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 27852 13084 28148 13104
rect 27908 13082 27932 13084
rect 27988 13082 28012 13084
rect 28068 13082 28092 13084
rect 27930 13030 27932 13082
rect 27994 13030 28006 13082
rect 28068 13030 28070 13082
rect 27908 13028 27932 13030
rect 27988 13028 28012 13030
rect 28068 13028 28092 13030
rect 27852 13008 28148 13028
rect 27712 12708 27764 12714
rect 27712 12650 27764 12656
rect 28172 12708 28224 12714
rect 28172 12650 28224 12656
rect 27852 11996 28148 12016
rect 27908 11994 27932 11996
rect 27988 11994 28012 11996
rect 28068 11994 28092 11996
rect 27930 11942 27932 11994
rect 27994 11942 28006 11994
rect 28068 11942 28070 11994
rect 27908 11940 27932 11942
rect 27988 11940 28012 11942
rect 28068 11940 28092 11942
rect 27852 11920 28148 11940
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27264 11150 27292 11494
rect 27436 11212 27488 11218
rect 27436 11154 27488 11160
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 27264 9110 27292 10406
rect 27448 10266 27476 11154
rect 28184 11150 28212 12650
rect 28264 12300 28316 12306
rect 28264 12242 28316 12248
rect 28276 11218 28304 12242
rect 28460 12102 28488 13262
rect 28920 12782 28948 14962
rect 29276 14884 29328 14890
rect 29276 14826 29328 14832
rect 29288 13870 29316 14826
rect 29380 14074 29408 15438
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29104 12986 29132 13806
rect 29564 13530 29592 15982
rect 30748 15972 30800 15978
rect 30748 15914 30800 15920
rect 29736 15904 29788 15910
rect 29736 15846 29788 15852
rect 29748 15434 29776 15846
rect 29736 15428 29788 15434
rect 29736 15370 29788 15376
rect 30104 15360 30156 15366
rect 30104 15302 30156 15308
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 29552 13524 29604 13530
rect 29552 13466 29604 13472
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 28908 12776 28960 12782
rect 28908 12718 28960 12724
rect 29460 12708 29512 12714
rect 29460 12650 29512 12656
rect 29092 12436 29144 12442
rect 29092 12378 29144 12384
rect 29104 12170 29132 12378
rect 29472 12238 29500 12650
rect 29460 12232 29512 12238
rect 29460 12174 29512 12180
rect 29092 12164 29144 12170
rect 29092 12106 29144 12112
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 30024 11898 30052 14758
rect 30116 14482 30144 15302
rect 30760 14958 30788 15914
rect 31956 15638 31984 17274
rect 32324 17082 32352 17682
rect 32232 17066 32352 17082
rect 32220 17060 32352 17066
rect 32272 17054 32352 17060
rect 32220 17002 32272 17008
rect 31944 15632 31996 15638
rect 31944 15574 31996 15580
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31116 15360 31168 15366
rect 31116 15302 31168 15308
rect 31128 14958 31156 15302
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 31116 14952 31168 14958
rect 31116 14894 31168 14900
rect 30760 14618 30788 14894
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30104 14476 30156 14482
rect 30104 14418 30156 14424
rect 30116 14278 30144 14418
rect 30104 14272 30156 14278
rect 30104 14214 30156 14220
rect 30116 13938 30144 14214
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 30116 13530 30144 13874
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 30944 13394 30972 13670
rect 30932 13388 30984 13394
rect 30932 13330 30984 13336
rect 30748 12436 30800 12442
rect 30800 12396 30972 12424
rect 30748 12378 30800 12384
rect 30104 12368 30156 12374
rect 30104 12310 30156 12316
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 30116 11286 30144 12310
rect 30472 12300 30524 12306
rect 30472 12242 30524 12248
rect 30484 11626 30512 12242
rect 30944 12170 30972 12396
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 30932 12164 30984 12170
rect 30932 12106 30984 12112
rect 30472 11620 30524 11626
rect 30472 11562 30524 11568
rect 30104 11280 30156 11286
rect 30104 11222 30156 11228
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 27852 10908 28148 10928
rect 27908 10906 27932 10908
rect 27988 10906 28012 10908
rect 28068 10906 28092 10908
rect 27930 10854 27932 10906
rect 27994 10854 28006 10906
rect 28068 10854 28070 10906
rect 27908 10852 27932 10854
rect 27988 10852 28012 10854
rect 28068 10852 28092 10854
rect 27852 10832 28148 10852
rect 31128 10606 31156 12174
rect 31220 11694 31248 15438
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31496 14414 31524 14758
rect 31484 14408 31536 14414
rect 31404 14368 31484 14396
rect 31404 12986 31432 14368
rect 31484 14350 31536 14356
rect 32036 14272 32088 14278
rect 32036 14214 32088 14220
rect 31484 13864 31536 13870
rect 31484 13806 31536 13812
rect 31496 13530 31524 13806
rect 31484 13524 31536 13530
rect 31484 13466 31536 13472
rect 32048 13394 32076 14214
rect 32036 13388 32088 13394
rect 32036 13330 32088 13336
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 31392 12980 31444 12986
rect 31392 12922 31444 12928
rect 31680 12782 31708 13262
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 31680 12374 31708 12718
rect 31668 12368 31720 12374
rect 31668 12310 31720 12316
rect 31208 11688 31260 11694
rect 31208 11630 31260 11636
rect 32232 11218 32260 17002
rect 32496 15564 32548 15570
rect 32496 15506 32548 15512
rect 32508 15026 32536 15506
rect 32600 15162 32628 19722
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32784 17746 32812 19110
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 33508 18896 33560 18902
rect 33704 18873 33732 18906
rect 33508 18838 33560 18844
rect 33690 18864 33746 18873
rect 32954 18592 33010 18601
rect 32954 18527 33010 18536
rect 32968 18358 32996 18527
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 33048 18080 33100 18086
rect 33048 18022 33100 18028
rect 32772 17740 32824 17746
rect 32772 17682 32824 17688
rect 32956 16652 33008 16658
rect 32956 16594 33008 16600
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32876 16250 32904 16526
rect 32864 16244 32916 16250
rect 32864 16186 32916 16192
rect 32680 15564 32732 15570
rect 32680 15506 32732 15512
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32496 15020 32548 15026
rect 32496 14962 32548 14968
rect 32600 14006 32628 15098
rect 32692 15026 32720 15506
rect 32680 15020 32732 15026
rect 32680 14962 32732 14968
rect 32692 14482 32720 14962
rect 32680 14476 32732 14482
rect 32680 14418 32732 14424
rect 32968 14006 32996 16594
rect 32588 14000 32640 14006
rect 32588 13942 32640 13948
rect 32956 14000 33008 14006
rect 32956 13942 33008 13948
rect 32404 13388 32456 13394
rect 32404 13330 32456 13336
rect 32416 12782 32444 13330
rect 32404 12776 32456 12782
rect 32404 12718 32456 12724
rect 32588 12300 32640 12306
rect 32588 12242 32640 12248
rect 32600 11694 32628 12242
rect 32680 12232 32732 12238
rect 32680 12174 32732 12180
rect 32772 12232 32824 12238
rect 32772 12174 32824 12180
rect 32692 11830 32720 12174
rect 32784 12102 32812 12174
rect 32772 12096 32824 12102
rect 32772 12038 32824 12044
rect 32680 11824 32732 11830
rect 32680 11766 32732 11772
rect 32784 11762 32812 12038
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32784 11354 32812 11698
rect 32772 11348 32824 11354
rect 32772 11290 32824 11296
rect 32220 11212 32272 11218
rect 32220 11154 32272 11160
rect 32232 10810 32260 11154
rect 32968 10810 32996 13942
rect 33060 13870 33088 18022
rect 33520 17678 33548 18838
rect 33690 18799 33746 18808
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33692 18760 33744 18766
rect 33692 18702 33744 18708
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 33612 18290 33640 18702
rect 33704 18630 33732 18702
rect 33692 18624 33744 18630
rect 33876 18624 33928 18630
rect 33692 18566 33744 18572
rect 33874 18592 33876 18601
rect 33928 18592 33930 18601
rect 33874 18527 33930 18536
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 33508 17672 33560 17678
rect 33508 17614 33560 17620
rect 33324 17536 33376 17542
rect 33324 17478 33376 17484
rect 33336 17338 33364 17478
rect 33324 17332 33376 17338
rect 33324 17274 33376 17280
rect 33232 17060 33284 17066
rect 33232 17002 33284 17008
rect 33244 15094 33272 17002
rect 33232 15088 33284 15094
rect 33232 15030 33284 15036
rect 33048 13864 33100 13870
rect 33048 13806 33100 13812
rect 33520 13326 33548 17614
rect 33600 17128 33652 17134
rect 33600 17070 33652 17076
rect 33612 16794 33640 17070
rect 33600 16788 33652 16794
rect 33600 16730 33652 16736
rect 33968 15972 34020 15978
rect 33968 15914 34020 15920
rect 33980 15706 34008 15914
rect 33968 15700 34020 15706
rect 33968 15642 34020 15648
rect 34060 14816 34112 14822
rect 34060 14758 34112 14764
rect 34072 14482 34100 14758
rect 34060 14476 34112 14482
rect 34060 14418 34112 14424
rect 34152 14408 34204 14414
rect 34152 14350 34204 14356
rect 34164 13870 34192 14350
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 34164 13462 34192 13806
rect 34152 13456 34204 13462
rect 34152 13398 34204 13404
rect 33968 13388 34020 13394
rect 33968 13330 34020 13336
rect 33232 13320 33284 13326
rect 33232 13262 33284 13268
rect 33508 13320 33560 13326
rect 33508 13262 33560 13268
rect 33244 11218 33272 13262
rect 33980 12850 34008 13330
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33416 12776 33468 12782
rect 33416 12718 33468 12724
rect 33324 12708 33376 12714
rect 33324 12650 33376 12656
rect 33336 11694 33364 12650
rect 33428 11898 33456 12718
rect 34348 12306 34376 18702
rect 34532 17649 34560 19314
rect 35622 18456 35678 18465
rect 34980 18420 35032 18426
rect 35622 18391 35678 18400
rect 34980 18362 35032 18368
rect 34992 18222 35020 18362
rect 35636 18222 35664 18391
rect 34980 18216 35032 18222
rect 34980 18158 35032 18164
rect 35164 18216 35216 18222
rect 35164 18158 35216 18164
rect 35624 18216 35676 18222
rect 35624 18158 35676 18164
rect 35716 18216 35768 18222
rect 35716 18158 35768 18164
rect 35176 18086 35204 18158
rect 35164 18080 35216 18086
rect 35164 18022 35216 18028
rect 35728 17746 35756 18158
rect 34612 17740 34664 17746
rect 34612 17682 34664 17688
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 34518 17640 34574 17649
rect 34518 17575 34574 17584
rect 34532 17202 34560 17575
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34428 15496 34480 15502
rect 34428 15438 34480 15444
rect 34440 15162 34468 15438
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34428 14340 34480 14346
rect 34428 14282 34480 14288
rect 34440 12986 34468 14282
rect 34520 13388 34572 13394
rect 34520 13330 34572 13336
rect 34428 12980 34480 12986
rect 34428 12922 34480 12928
rect 34336 12300 34388 12306
rect 34336 12242 34388 12248
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 33324 11688 33376 11694
rect 33324 11630 33376 11636
rect 33336 11354 33364 11630
rect 34348 11558 34376 12242
rect 34336 11552 34388 11558
rect 34336 11494 34388 11500
rect 34532 11354 34560 13330
rect 34624 12646 34652 17682
rect 35912 17610 35940 20198
rect 36188 20058 36216 20810
rect 36464 20806 36492 21082
rect 36452 20800 36504 20806
rect 36452 20742 36504 20748
rect 36817 20156 37113 20176
rect 36873 20154 36897 20156
rect 36953 20154 36977 20156
rect 37033 20154 37057 20156
rect 36895 20102 36897 20154
rect 36959 20102 36971 20154
rect 37033 20102 37035 20154
rect 36873 20100 36897 20102
rect 36953 20100 36977 20102
rect 37033 20100 37057 20102
rect 36817 20080 37113 20100
rect 36176 20052 36228 20058
rect 36176 19994 36228 20000
rect 36268 19304 36320 19310
rect 36820 19304 36872 19310
rect 36268 19246 36320 19252
rect 36648 19264 36820 19292
rect 36176 19236 36228 19242
rect 36176 19178 36228 19184
rect 36188 18970 36216 19178
rect 36280 18970 36308 19246
rect 36176 18964 36228 18970
rect 36176 18906 36228 18912
rect 36268 18964 36320 18970
rect 36268 18906 36320 18912
rect 36188 18834 36216 18906
rect 36176 18828 36228 18834
rect 36176 18770 36228 18776
rect 36452 18692 36504 18698
rect 36452 18634 36504 18640
rect 36464 18086 36492 18634
rect 36452 18080 36504 18086
rect 36452 18022 36504 18028
rect 36648 17814 36676 19264
rect 36820 19246 36872 19252
rect 36817 19068 37113 19088
rect 36873 19066 36897 19068
rect 36953 19066 36977 19068
rect 37033 19066 37057 19068
rect 36895 19014 36897 19066
rect 36959 19014 36971 19066
rect 37033 19014 37035 19066
rect 36873 19012 36897 19014
rect 36953 19012 36977 19014
rect 37033 19012 37057 19014
rect 36817 18992 37113 19012
rect 36726 18864 36782 18873
rect 36726 18799 36728 18808
rect 36780 18799 36782 18808
rect 36728 18770 36780 18776
rect 36817 17980 37113 18000
rect 36873 17978 36897 17980
rect 36953 17978 36977 17980
rect 37033 17978 37057 17980
rect 36895 17926 36897 17978
rect 36959 17926 36971 17978
rect 37033 17926 37035 17978
rect 36873 17924 36897 17926
rect 36953 17924 36977 17926
rect 37033 17924 37057 17926
rect 36817 17904 37113 17924
rect 37200 17814 37228 21354
rect 38120 20466 38148 23054
rect 38200 22976 38252 22982
rect 38200 22918 38252 22924
rect 38212 21894 38240 22918
rect 38200 21888 38252 21894
rect 38200 21830 38252 21836
rect 38212 21486 38240 21830
rect 38304 21554 38332 26400
rect 39040 24410 39068 26400
rect 39028 24404 39080 24410
rect 39028 24346 39080 24352
rect 38752 24200 38804 24206
rect 38752 24142 38804 24148
rect 38764 23866 38792 24142
rect 38752 23860 38804 23866
rect 38752 23802 38804 23808
rect 38844 23520 38896 23526
rect 38844 23462 38896 23468
rect 38752 23112 38804 23118
rect 38566 23080 38622 23089
rect 38622 23038 38700 23066
rect 38752 23054 38804 23060
rect 38566 23015 38622 23024
rect 38384 22772 38436 22778
rect 38384 22714 38436 22720
rect 38292 21548 38344 21554
rect 38292 21490 38344 21496
rect 38396 21486 38424 22714
rect 38672 22658 38700 23038
rect 38764 22778 38792 23054
rect 38752 22772 38804 22778
rect 38752 22714 38804 22720
rect 38672 22642 38792 22658
rect 38672 22636 38804 22642
rect 38672 22630 38752 22636
rect 38752 22578 38804 22584
rect 38856 22574 38884 23462
rect 39776 23186 39804 26400
rect 40512 24818 40540 26400
rect 41248 24834 41276 26400
rect 40500 24812 40552 24818
rect 41248 24806 41368 24834
rect 40500 24754 40552 24760
rect 40408 24744 40460 24750
rect 40408 24686 40460 24692
rect 41236 24744 41288 24750
rect 41236 24686 41288 24692
rect 39948 24608 40000 24614
rect 39948 24550 40000 24556
rect 39960 23730 39988 24550
rect 39948 23724 40000 23730
rect 39948 23666 40000 23672
rect 40040 23656 40092 23662
rect 40040 23598 40092 23604
rect 40132 23656 40184 23662
rect 40132 23598 40184 23604
rect 39764 23180 39816 23186
rect 39764 23122 39816 23128
rect 38844 22568 38896 22574
rect 38844 22510 38896 22516
rect 39488 22568 39540 22574
rect 39488 22510 39540 22516
rect 38200 21480 38252 21486
rect 38200 21422 38252 21428
rect 38384 21480 38436 21486
rect 38384 21422 38436 21428
rect 38752 21480 38804 21486
rect 38752 21422 38804 21428
rect 38292 20800 38344 20806
rect 38292 20742 38344 20748
rect 38108 20460 38160 20466
rect 38108 20402 38160 20408
rect 38304 20398 38332 20742
rect 38016 20392 38068 20398
rect 38016 20334 38068 20340
rect 38292 20392 38344 20398
rect 38292 20334 38344 20340
rect 37280 20324 37332 20330
rect 37280 20266 37332 20272
rect 37292 19310 37320 20266
rect 37372 19916 37424 19922
rect 37372 19858 37424 19864
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37280 19168 37332 19174
rect 37280 19110 37332 19116
rect 37292 18358 37320 19110
rect 37384 18630 37412 19858
rect 37648 19168 37700 19174
rect 37648 19110 37700 19116
rect 37660 18970 37688 19110
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 37372 18624 37424 18630
rect 37372 18566 37424 18572
rect 37280 18352 37332 18358
rect 37280 18294 37332 18300
rect 36636 17808 36688 17814
rect 36636 17750 36688 17756
rect 37188 17808 37240 17814
rect 37188 17750 37240 17756
rect 36360 17740 36412 17746
rect 36360 17682 36412 17688
rect 35900 17604 35952 17610
rect 35820 17564 35900 17592
rect 35624 17128 35676 17134
rect 35624 17070 35676 17076
rect 35636 16998 35664 17070
rect 35624 16992 35676 16998
rect 35624 16934 35676 16940
rect 35820 16658 35848 17564
rect 35900 17546 35952 17552
rect 36082 17368 36138 17377
rect 36082 17303 36138 17312
rect 36096 17270 36124 17303
rect 36084 17264 36136 17270
rect 36084 17206 36136 17212
rect 36084 17128 36136 17134
rect 36004 17076 36084 17082
rect 36004 17070 36136 17076
rect 35900 17060 35952 17066
rect 36004 17054 36124 17070
rect 36004 17048 36032 17054
rect 35952 17020 36032 17048
rect 35900 17002 35952 17008
rect 35808 16652 35860 16658
rect 35808 16594 35860 16600
rect 35820 16454 35848 16594
rect 35900 16584 35952 16590
rect 35900 16526 35952 16532
rect 35808 16448 35860 16454
rect 35808 16390 35860 16396
rect 35912 16250 35940 16526
rect 36372 16522 36400 17682
rect 36450 17368 36506 17377
rect 36450 17303 36506 17312
rect 36464 17134 36492 17303
rect 36452 17128 36504 17134
rect 36452 17070 36504 17076
rect 36360 16516 36412 16522
rect 36360 16458 36412 16464
rect 36452 16448 36504 16454
rect 36452 16390 36504 16396
rect 35900 16244 35952 16250
rect 35900 16186 35952 16192
rect 35532 16040 35584 16046
rect 35532 15982 35584 15988
rect 35808 16040 35860 16046
rect 35808 15982 35860 15988
rect 34980 15564 35032 15570
rect 34980 15506 35032 15512
rect 34992 14958 35020 15506
rect 34980 14952 35032 14958
rect 34980 14894 35032 14900
rect 35164 14476 35216 14482
rect 35440 14476 35492 14482
rect 35216 14436 35440 14464
rect 35164 14418 35216 14424
rect 35440 14418 35492 14424
rect 35348 14340 35400 14346
rect 35348 14282 35400 14288
rect 35360 14006 35388 14282
rect 35348 14000 35400 14006
rect 35348 13942 35400 13948
rect 35360 13462 35388 13942
rect 35452 13870 35480 14418
rect 35544 14346 35572 15982
rect 35624 15972 35676 15978
rect 35624 15914 35676 15920
rect 35636 15026 35664 15914
rect 35820 15570 35848 15982
rect 35808 15564 35860 15570
rect 35808 15506 35860 15512
rect 35624 15020 35676 15026
rect 35624 14962 35676 14968
rect 35716 14884 35768 14890
rect 35716 14826 35768 14832
rect 35728 14618 35756 14826
rect 35716 14612 35768 14618
rect 35716 14554 35768 14560
rect 35532 14340 35584 14346
rect 35532 14282 35584 14288
rect 35440 13864 35492 13870
rect 35440 13806 35492 13812
rect 35348 13456 35400 13462
rect 35348 13398 35400 13404
rect 34980 13320 35032 13326
rect 34980 13262 35032 13268
rect 34992 12850 35020 13262
rect 35544 13258 35572 14282
rect 35992 13864 36044 13870
rect 35992 13806 36044 13812
rect 36004 13394 36032 13806
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 34980 12844 35032 12850
rect 34980 12786 35032 12792
rect 36004 12782 36032 13330
rect 36464 12918 36492 16390
rect 36648 15570 36676 17750
rect 37200 17066 37228 17750
rect 37384 17746 37412 18566
rect 37924 17876 37976 17882
rect 37924 17818 37976 17824
rect 37372 17740 37424 17746
rect 37372 17682 37424 17688
rect 37936 17649 37964 17818
rect 37922 17640 37978 17649
rect 37922 17575 37978 17584
rect 38028 17202 38056 20334
rect 38476 20324 38528 20330
rect 38476 20266 38528 20272
rect 38488 20058 38516 20266
rect 38476 20052 38528 20058
rect 38476 19994 38528 20000
rect 38384 19984 38436 19990
rect 38384 19926 38436 19932
rect 38292 19848 38344 19854
rect 38292 19790 38344 19796
rect 38304 19310 38332 19790
rect 38396 19310 38424 19926
rect 38292 19304 38344 19310
rect 38292 19246 38344 19252
rect 38384 19304 38436 19310
rect 38384 19246 38436 19252
rect 38290 18728 38346 18737
rect 38290 18663 38292 18672
rect 38344 18663 38346 18672
rect 38292 18634 38344 18640
rect 38396 17762 38424 19246
rect 38764 19174 38792 21422
rect 38936 20936 38988 20942
rect 38936 20878 38988 20884
rect 38948 20534 38976 20878
rect 39120 20800 39172 20806
rect 39120 20742 39172 20748
rect 38936 20528 38988 20534
rect 38936 20470 38988 20476
rect 38752 19168 38804 19174
rect 38752 19110 38804 19116
rect 39026 19136 39082 19145
rect 38660 17808 38712 17814
rect 38396 17746 38608 17762
rect 38660 17750 38712 17756
rect 38108 17740 38160 17746
rect 38108 17682 38160 17688
rect 38384 17740 38620 17746
rect 38436 17734 38568 17740
rect 38384 17682 38436 17688
rect 38568 17682 38620 17688
rect 38016 17196 38068 17202
rect 38016 17138 38068 17144
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 37188 17060 37240 17066
rect 37188 17002 37240 17008
rect 36817 16892 37113 16912
rect 36873 16890 36897 16892
rect 36953 16890 36977 16892
rect 37033 16890 37057 16892
rect 36895 16838 36897 16890
rect 36959 16838 36971 16890
rect 37033 16838 37035 16890
rect 36873 16836 36897 16838
rect 36953 16836 36977 16838
rect 37033 16836 37057 16838
rect 36817 16816 37113 16836
rect 37188 16788 37240 16794
rect 37188 16730 37240 16736
rect 37200 16697 37228 16730
rect 37186 16688 37242 16697
rect 37186 16623 37242 16632
rect 36817 15804 37113 15824
rect 36873 15802 36897 15804
rect 36953 15802 36977 15804
rect 37033 15802 37057 15804
rect 36895 15750 36897 15802
rect 36959 15750 36971 15802
rect 37033 15750 37035 15802
rect 36873 15748 36897 15750
rect 36953 15748 36977 15750
rect 37033 15748 37057 15750
rect 36817 15728 37113 15748
rect 36636 15564 36688 15570
rect 36636 15506 36688 15512
rect 36648 15008 36676 15506
rect 36728 15020 36780 15026
rect 36648 14980 36728 15008
rect 36728 14962 36780 14968
rect 36817 14716 37113 14736
rect 36873 14714 36897 14716
rect 36953 14714 36977 14716
rect 37033 14714 37057 14716
rect 36895 14662 36897 14714
rect 36959 14662 36971 14714
rect 37033 14662 37035 14714
rect 36873 14660 36897 14662
rect 36953 14660 36977 14662
rect 37033 14660 37057 14662
rect 36817 14640 37113 14660
rect 37740 14544 37792 14550
rect 37740 14486 37792 14492
rect 37372 14340 37424 14346
rect 37372 14282 37424 14288
rect 37384 14006 37412 14282
rect 37556 14272 37608 14278
rect 37556 14214 37608 14220
rect 37372 14000 37424 14006
rect 37372 13942 37424 13948
rect 37568 13870 37596 14214
rect 37556 13864 37608 13870
rect 37556 13806 37608 13812
rect 37648 13864 37700 13870
rect 37648 13806 37700 13812
rect 36817 13628 37113 13648
rect 36873 13626 36897 13628
rect 36953 13626 36977 13628
rect 37033 13626 37057 13628
rect 36895 13574 36897 13626
rect 36959 13574 36971 13626
rect 37033 13574 37035 13626
rect 36873 13572 36897 13574
rect 36953 13572 36977 13574
rect 37033 13572 37057 13574
rect 36817 13552 37113 13572
rect 37660 13462 37688 13806
rect 37648 13456 37700 13462
rect 37648 13398 37700 13404
rect 37752 12918 37780 14486
rect 37844 14482 37872 17070
rect 38120 16998 38148 17682
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 38384 16584 38436 16590
rect 38672 16572 38700 17750
rect 38764 17066 38792 19110
rect 39026 19071 39082 19080
rect 38844 18828 38896 18834
rect 38844 18770 38896 18776
rect 38856 18630 38884 18770
rect 38934 18728 38990 18737
rect 38934 18663 38990 18672
rect 38844 18624 38896 18630
rect 38844 18566 38896 18572
rect 38948 18222 38976 18663
rect 39040 18290 39068 19071
rect 39132 18714 39160 20742
rect 39396 19372 39448 19378
rect 39396 19314 39448 19320
rect 39304 18828 39356 18834
rect 39304 18770 39356 18776
rect 39132 18686 39252 18714
rect 39120 18624 39172 18630
rect 39120 18566 39172 18572
rect 39132 18358 39160 18566
rect 39120 18352 39172 18358
rect 39120 18294 39172 18300
rect 39028 18284 39080 18290
rect 39028 18226 39080 18232
rect 38936 18216 38988 18222
rect 38936 18158 38988 18164
rect 38844 18148 38896 18154
rect 38844 18090 38896 18096
rect 38856 17882 38884 18090
rect 38844 17876 38896 17882
rect 38844 17818 38896 17824
rect 39028 17876 39080 17882
rect 39028 17818 39080 17824
rect 39040 17338 39068 17818
rect 39028 17332 39080 17338
rect 39028 17274 39080 17280
rect 39224 17270 39252 18686
rect 39316 18358 39344 18770
rect 39304 18352 39356 18358
rect 39304 18294 39356 18300
rect 39304 17536 39356 17542
rect 39304 17478 39356 17484
rect 39212 17264 39264 17270
rect 39212 17206 39264 17212
rect 39316 17202 39344 17478
rect 39304 17196 39356 17202
rect 39304 17138 39356 17144
rect 38752 17060 38804 17066
rect 38752 17002 38804 17008
rect 38752 16584 38804 16590
rect 38672 16544 38752 16572
rect 38384 16526 38436 16532
rect 38752 16526 38804 16532
rect 39120 16584 39172 16590
rect 39120 16526 39172 16532
rect 38396 15638 38424 16526
rect 39132 16046 39160 16526
rect 39408 16250 39436 19314
rect 39500 18834 39528 22510
rect 39856 22024 39908 22030
rect 39856 21966 39908 21972
rect 39868 21554 39896 21966
rect 39856 21548 39908 21554
rect 39856 21490 39908 21496
rect 40052 21078 40080 23598
rect 40144 22982 40172 23598
rect 40132 22976 40184 22982
rect 40132 22918 40184 22924
rect 40144 22098 40172 22918
rect 40420 22574 40448 24686
rect 41248 24274 41276 24686
rect 41236 24268 41288 24274
rect 41236 24210 41288 24216
rect 41052 23520 41104 23526
rect 41052 23462 41104 23468
rect 40592 23044 40644 23050
rect 40592 22986 40644 22992
rect 40604 22710 40632 22986
rect 40592 22704 40644 22710
rect 40592 22646 40644 22652
rect 40408 22568 40460 22574
rect 40408 22510 40460 22516
rect 40224 22500 40276 22506
rect 40224 22442 40276 22448
rect 40132 22092 40184 22098
rect 40132 22034 40184 22040
rect 40236 21146 40264 22442
rect 41064 21622 41092 23462
rect 41144 23180 41196 23186
rect 41144 23122 41196 23128
rect 41052 21616 41104 21622
rect 41052 21558 41104 21564
rect 41052 21480 41104 21486
rect 41052 21422 41104 21428
rect 40224 21140 40276 21146
rect 40224 21082 40276 21088
rect 40040 21072 40092 21078
rect 40040 21014 40092 21020
rect 40776 21072 40828 21078
rect 40776 21014 40828 21020
rect 40224 20936 40276 20942
rect 40224 20878 40276 20884
rect 40040 20392 40092 20398
rect 40040 20334 40092 20340
rect 39764 19916 39816 19922
rect 39764 19858 39816 19864
rect 39578 19816 39634 19825
rect 39776 19802 39804 19858
rect 39578 19751 39634 19760
rect 39684 19774 39804 19802
rect 39488 18828 39540 18834
rect 39488 18770 39540 18776
rect 39500 18068 39528 18770
rect 39592 18630 39620 19751
rect 39684 19378 39712 19774
rect 39672 19372 39724 19378
rect 39672 19314 39724 19320
rect 39764 19304 39816 19310
rect 39764 19246 39816 19252
rect 39776 19174 39804 19246
rect 39764 19168 39816 19174
rect 39764 19110 39816 19116
rect 40052 18902 40080 20334
rect 40132 19780 40184 19786
rect 40132 19722 40184 19728
rect 39856 18896 39908 18902
rect 39684 18844 39856 18850
rect 39684 18838 39908 18844
rect 40040 18896 40092 18902
rect 40040 18838 40092 18844
rect 39684 18822 39896 18838
rect 39580 18624 39632 18630
rect 39580 18566 39632 18572
rect 39592 18306 39620 18566
rect 39684 18426 39712 18822
rect 39946 18592 40002 18601
rect 39946 18527 40002 18536
rect 39960 18426 39988 18527
rect 39672 18420 39724 18426
rect 39672 18362 39724 18368
rect 39764 18420 39816 18426
rect 39764 18362 39816 18368
rect 39948 18420 40000 18426
rect 39948 18362 40000 18368
rect 39776 18306 39804 18362
rect 39592 18278 39804 18306
rect 40144 18290 40172 19722
rect 40236 18630 40264 20878
rect 40224 18624 40276 18630
rect 40224 18566 40276 18572
rect 40132 18284 40184 18290
rect 40132 18226 40184 18232
rect 40788 18222 40816 21014
rect 41064 19922 41092 21422
rect 41156 21350 41184 23122
rect 41236 22432 41288 22438
rect 41236 22374 41288 22380
rect 41248 21876 41276 22374
rect 41340 22166 41368 24806
rect 41788 23656 41840 23662
rect 41788 23598 41840 23604
rect 41604 23316 41656 23322
rect 41604 23258 41656 23264
rect 41616 22642 41644 23258
rect 41604 22636 41656 22642
rect 41604 22578 41656 22584
rect 41328 22160 41380 22166
rect 41328 22102 41380 22108
rect 41328 21888 41380 21894
rect 41248 21848 41328 21876
rect 41328 21830 41380 21836
rect 41144 21344 41196 21350
rect 41144 21286 41196 21292
rect 41052 19916 41104 19922
rect 41052 19858 41104 19864
rect 41064 19718 41092 19858
rect 41052 19712 41104 19718
rect 41052 19654 41104 19660
rect 41064 19514 41092 19654
rect 41052 19508 41104 19514
rect 41052 19450 41104 19456
rect 41340 19174 41368 21830
rect 41696 21140 41748 21146
rect 41696 21082 41748 21088
rect 41420 19712 41472 19718
rect 41420 19654 41472 19660
rect 41432 19310 41460 19654
rect 41420 19304 41472 19310
rect 41420 19246 41472 19252
rect 41602 19272 41658 19281
rect 41602 19207 41604 19216
rect 41656 19207 41658 19216
rect 41604 19178 41656 19184
rect 41328 19168 41380 19174
rect 41328 19110 41380 19116
rect 41340 18873 41368 19110
rect 41708 18970 41736 21082
rect 41800 20466 41828 23598
rect 41892 23322 41920 26400
rect 41972 24744 42024 24750
rect 41972 24686 42024 24692
rect 41984 23866 42012 24686
rect 41972 23860 42024 23866
rect 41972 23802 42024 23808
rect 41880 23316 41932 23322
rect 41880 23258 41932 23264
rect 41880 23180 41932 23186
rect 41880 23122 41932 23128
rect 42340 23180 42392 23186
rect 42340 23122 42392 23128
rect 41892 22778 41920 23122
rect 41880 22772 41932 22778
rect 41880 22714 41932 22720
rect 41892 22574 41920 22714
rect 42248 22636 42300 22642
rect 42248 22578 42300 22584
rect 41880 22568 41932 22574
rect 41880 22510 41932 22516
rect 41972 22500 42024 22506
rect 41972 22442 42024 22448
rect 41788 20460 41840 20466
rect 41788 20402 41840 20408
rect 41512 18964 41564 18970
rect 41512 18906 41564 18912
rect 41696 18964 41748 18970
rect 41696 18906 41748 18912
rect 41326 18864 41382 18873
rect 41326 18799 41382 18808
rect 41524 18630 41552 18906
rect 41708 18834 41736 18906
rect 41696 18828 41748 18834
rect 41696 18770 41748 18776
rect 41512 18624 41564 18630
rect 41512 18566 41564 18572
rect 41604 18420 41656 18426
rect 41604 18362 41656 18368
rect 41616 18329 41644 18362
rect 41602 18320 41658 18329
rect 41602 18255 41658 18264
rect 39948 18216 40000 18222
rect 39948 18158 40000 18164
rect 40776 18216 40828 18222
rect 40776 18158 40828 18164
rect 39960 18068 39988 18158
rect 39500 18040 39988 18068
rect 40040 18080 40092 18086
rect 40040 18022 40092 18028
rect 40052 17626 40080 18022
rect 40788 17746 40816 18158
rect 40880 17870 41368 17898
rect 40880 17746 40908 17870
rect 41050 17776 41106 17785
rect 40776 17740 40828 17746
rect 40776 17682 40828 17688
rect 40868 17740 40920 17746
rect 41340 17746 41368 17870
rect 41050 17711 41106 17720
rect 41328 17740 41380 17746
rect 40868 17682 40920 17688
rect 39960 17610 40080 17626
rect 39948 17604 40080 17610
rect 40000 17598 40080 17604
rect 40776 17604 40828 17610
rect 39948 17546 40000 17552
rect 40776 17546 40828 17552
rect 40038 17368 40094 17377
rect 40038 17303 40094 17312
rect 39948 17264 40000 17270
rect 39948 17206 40000 17212
rect 39488 17128 39540 17134
rect 39486 17096 39488 17105
rect 39540 17096 39542 17105
rect 39486 17031 39542 17040
rect 39672 17060 39724 17066
rect 39672 17002 39724 17008
rect 39684 16590 39712 17002
rect 39764 16992 39816 16998
rect 39764 16934 39816 16940
rect 39672 16584 39724 16590
rect 39672 16526 39724 16532
rect 39396 16244 39448 16250
rect 39396 16186 39448 16192
rect 39120 16040 39172 16046
rect 39120 15982 39172 15988
rect 38384 15632 38436 15638
rect 38384 15574 38436 15580
rect 39408 15570 39436 16186
rect 39028 15564 39080 15570
rect 39028 15506 39080 15512
rect 39396 15564 39448 15570
rect 39396 15506 39448 15512
rect 38752 15496 38804 15502
rect 38752 15438 38804 15444
rect 38764 15094 38792 15438
rect 38752 15088 38804 15094
rect 38752 15030 38804 15036
rect 39040 15026 39068 15506
rect 39408 15162 39436 15506
rect 39396 15156 39448 15162
rect 39396 15098 39448 15104
rect 39028 15020 39080 15026
rect 39028 14962 39080 14968
rect 39408 14958 39436 15098
rect 39396 14952 39448 14958
rect 39396 14894 39448 14900
rect 39396 14816 39448 14822
rect 39396 14758 39448 14764
rect 39672 14816 39724 14822
rect 39672 14758 39724 14764
rect 39408 14550 39436 14758
rect 39396 14544 39448 14550
rect 39396 14486 39448 14492
rect 37832 14476 37884 14482
rect 37832 14418 37884 14424
rect 38568 14476 38620 14482
rect 38568 14418 38620 14424
rect 38580 14278 38608 14418
rect 38568 14272 38620 14278
rect 38568 14214 38620 14220
rect 38580 13938 38608 14214
rect 38568 13932 38620 13938
rect 38568 13874 38620 13880
rect 38200 13796 38252 13802
rect 38200 13738 38252 13744
rect 38212 13394 38240 13738
rect 38200 13388 38252 13394
rect 38200 13330 38252 13336
rect 38580 13326 38608 13874
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 36452 12912 36504 12918
rect 36452 12854 36504 12860
rect 37740 12912 37792 12918
rect 37740 12854 37792 12860
rect 35992 12776 36044 12782
rect 35992 12718 36044 12724
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34612 11688 34664 11694
rect 34612 11630 34664 11636
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 34520 11348 34572 11354
rect 34520 11290 34572 11296
rect 34624 11218 34652 11630
rect 34716 11626 34744 12378
rect 35072 12300 35124 12306
rect 35072 12242 35124 12248
rect 35440 12300 35492 12306
rect 35440 12242 35492 12248
rect 34704 11620 34756 11626
rect 34704 11562 34756 11568
rect 34716 11218 34744 11562
rect 35084 11286 35112 12242
rect 35452 11830 35480 12242
rect 35624 12096 35676 12102
rect 35624 12038 35676 12044
rect 35440 11824 35492 11830
rect 35440 11766 35492 11772
rect 35636 11694 35664 12038
rect 36464 11898 36492 12854
rect 39684 12850 39712 14758
rect 39776 14414 39804 16934
rect 39960 16726 39988 17206
rect 39948 16720 40000 16726
rect 39948 16662 40000 16668
rect 39960 16454 39988 16662
rect 39948 16448 40000 16454
rect 39948 16390 40000 16396
rect 39764 14408 39816 14414
rect 39764 14350 39816 14356
rect 40052 12918 40080 17303
rect 40500 16720 40552 16726
rect 40500 16662 40552 16668
rect 40512 16590 40540 16662
rect 40788 16658 40816 17546
rect 40880 17377 40908 17682
rect 40866 17368 40922 17377
rect 40866 17303 40922 17312
rect 41064 16658 41092 17711
rect 41328 17682 41380 17688
rect 41708 17338 41736 18770
rect 41696 17332 41748 17338
rect 41696 17274 41748 17280
rect 41604 17196 41656 17202
rect 41800 17184 41828 20402
rect 41984 18086 42012 22442
rect 42154 22264 42210 22273
rect 42154 22199 42156 22208
rect 42208 22199 42210 22208
rect 42156 22170 42208 22176
rect 42260 22098 42288 22578
rect 42352 22234 42380 23122
rect 42628 22574 42656 26400
rect 43364 24818 43392 26400
rect 43352 24812 43404 24818
rect 43352 24754 43404 24760
rect 42892 24608 42944 24614
rect 42892 24550 42944 24556
rect 42984 24608 43036 24614
rect 42984 24550 43036 24556
rect 42904 24342 42932 24550
rect 42892 24336 42944 24342
rect 42892 24278 42944 24284
rect 42996 24274 43024 24550
rect 42984 24268 43036 24274
rect 42984 24210 43036 24216
rect 42800 22772 42852 22778
rect 42800 22714 42852 22720
rect 43076 22772 43128 22778
rect 43076 22714 43128 22720
rect 42616 22568 42668 22574
rect 42616 22510 42668 22516
rect 42340 22228 42392 22234
rect 42340 22170 42392 22176
rect 42812 22098 42840 22714
rect 43088 22574 43116 22714
rect 43076 22568 43128 22574
rect 43076 22510 43128 22516
rect 43536 22500 43588 22506
rect 43536 22442 43588 22448
rect 42248 22092 42300 22098
rect 42248 22034 42300 22040
rect 42616 22092 42668 22098
rect 42616 22034 42668 22040
rect 42800 22092 42852 22098
rect 42800 22034 42852 22040
rect 42628 21894 42656 22034
rect 42616 21888 42668 21894
rect 42616 21830 42668 21836
rect 42340 19304 42392 19310
rect 42340 19246 42392 19252
rect 42432 19304 42484 19310
rect 42432 19246 42484 19252
rect 42352 18986 42380 19246
rect 42444 19174 42472 19246
rect 42432 19168 42484 19174
rect 42432 19110 42484 19116
rect 42524 19168 42576 19174
rect 42524 19110 42576 19116
rect 42536 18986 42564 19110
rect 42352 18958 42564 18986
rect 41972 18080 42024 18086
rect 41972 18022 42024 18028
rect 42248 17332 42300 17338
rect 42248 17274 42300 17280
rect 41656 17156 41828 17184
rect 41604 17138 41656 17144
rect 41800 16658 41828 17156
rect 42260 17134 42288 17274
rect 42248 17128 42300 17134
rect 42248 17070 42300 17076
rect 42352 16794 42380 18958
rect 42628 18222 42656 21830
rect 42812 21146 42840 22034
rect 43548 21554 43576 22442
rect 43536 21548 43588 21554
rect 43536 21490 43588 21496
rect 42984 21344 43036 21350
rect 42984 21286 43036 21292
rect 43168 21344 43220 21350
rect 43168 21286 43220 21292
rect 42996 21146 43024 21286
rect 42800 21140 42852 21146
rect 42800 21082 42852 21088
rect 42984 21140 43036 21146
rect 42984 21082 43036 21088
rect 42892 20392 42944 20398
rect 42892 20334 42944 20340
rect 42904 19514 42932 20334
rect 42996 20262 43024 21082
rect 43180 21078 43208 21286
rect 43168 21072 43220 21078
rect 43168 21014 43220 21020
rect 42984 20256 43036 20262
rect 42984 20198 43036 20204
rect 42892 19508 42944 19514
rect 42892 19450 42944 19456
rect 44100 19242 44128 26400
rect 44272 24744 44324 24750
rect 44272 24686 44324 24692
rect 44284 23866 44312 24686
rect 44548 24608 44600 24614
rect 44548 24550 44600 24556
rect 44836 24562 44864 26400
rect 44560 24070 44588 24550
rect 44836 24534 45048 24562
rect 44548 24064 44600 24070
rect 44548 24006 44600 24012
rect 44272 23860 44324 23866
rect 44272 23802 44324 23808
rect 44180 23656 44232 23662
rect 44180 23598 44232 23604
rect 44192 19310 44220 23598
rect 44560 23254 44588 24006
rect 44548 23248 44600 23254
rect 44548 23190 44600 23196
rect 44560 23118 44588 23190
rect 44548 23112 44600 23118
rect 44548 23054 44600 23060
rect 44916 23112 44968 23118
rect 44916 23054 44968 23060
rect 44364 22976 44416 22982
rect 44364 22918 44416 22924
rect 44376 22642 44404 22918
rect 44364 22636 44416 22642
rect 44364 22578 44416 22584
rect 44824 22432 44876 22438
rect 44824 22374 44876 22380
rect 44836 22098 44864 22374
rect 44928 22166 44956 23054
rect 45020 22234 45048 24534
rect 45376 24064 45428 24070
rect 45376 24006 45428 24012
rect 45388 23798 45416 24006
rect 45376 23792 45428 23798
rect 45376 23734 45428 23740
rect 45008 22228 45060 22234
rect 45008 22170 45060 22176
rect 44916 22160 44968 22166
rect 44916 22102 44968 22108
rect 44272 22092 44324 22098
rect 44272 22034 44324 22040
rect 44824 22092 44876 22098
rect 44824 22034 44876 22040
rect 44284 20942 44312 22034
rect 45388 21894 45416 23734
rect 45480 23202 45508 26400
rect 45782 25052 46078 25072
rect 45838 25050 45862 25052
rect 45918 25050 45942 25052
rect 45998 25050 46022 25052
rect 45860 24998 45862 25050
rect 45924 24998 45936 25050
rect 45998 24998 46000 25050
rect 45838 24996 45862 24998
rect 45918 24996 45942 24998
rect 45998 24996 46022 24998
rect 45782 24976 46078 24996
rect 45560 24608 45612 24614
rect 45560 24550 45612 24556
rect 45572 23322 45600 24550
rect 45782 23964 46078 23984
rect 45838 23962 45862 23964
rect 45918 23962 45942 23964
rect 45998 23962 46022 23964
rect 45860 23910 45862 23962
rect 45924 23910 45936 23962
rect 45998 23910 46000 23962
rect 45838 23908 45862 23910
rect 45918 23908 45942 23910
rect 45998 23908 46022 23910
rect 45782 23888 46078 23908
rect 46216 23746 46244 26400
rect 46572 24200 46624 24206
rect 46572 24142 46624 24148
rect 46584 23866 46612 24142
rect 46664 24064 46716 24070
rect 46664 24006 46716 24012
rect 46572 23860 46624 23866
rect 46572 23802 46624 23808
rect 46124 23718 46244 23746
rect 46124 23322 46152 23718
rect 46204 23656 46256 23662
rect 46204 23598 46256 23604
rect 46388 23656 46440 23662
rect 46388 23598 46440 23604
rect 45560 23316 45612 23322
rect 45560 23258 45612 23264
rect 46112 23316 46164 23322
rect 46112 23258 46164 23264
rect 45480 23174 45600 23202
rect 45376 21888 45428 21894
rect 45376 21830 45428 21836
rect 45388 21146 45416 21830
rect 45376 21140 45428 21146
rect 45376 21082 45428 21088
rect 44456 21004 44508 21010
rect 44456 20946 44508 20952
rect 44272 20936 44324 20942
rect 44272 20878 44324 20884
rect 44468 20806 44496 20946
rect 44456 20800 44508 20806
rect 44456 20742 44508 20748
rect 44468 20602 44496 20742
rect 44456 20596 44508 20602
rect 44456 20538 44508 20544
rect 45572 20466 45600 23174
rect 46216 23118 46244 23598
rect 46400 23254 46428 23598
rect 46388 23248 46440 23254
rect 46388 23190 46440 23196
rect 46204 23112 46256 23118
rect 46204 23054 46256 23060
rect 45782 22876 46078 22896
rect 45838 22874 45862 22876
rect 45918 22874 45942 22876
rect 45998 22874 46022 22876
rect 45860 22822 45862 22874
rect 45924 22822 45936 22874
rect 45998 22822 46000 22874
rect 45838 22820 45862 22822
rect 45918 22820 45942 22822
rect 45998 22820 46022 22822
rect 45782 22800 46078 22820
rect 46400 22574 46428 23190
rect 46676 23186 46704 24006
rect 46664 23180 46716 23186
rect 46664 23122 46716 23128
rect 46388 22568 46440 22574
rect 46388 22510 46440 22516
rect 46296 22432 46348 22438
rect 46296 22374 46348 22380
rect 46308 22273 46336 22374
rect 46294 22264 46350 22273
rect 46294 22199 46350 22208
rect 46112 22092 46164 22098
rect 46112 22034 46164 22040
rect 46124 21894 46152 22034
rect 46296 22024 46348 22030
rect 46296 21966 46348 21972
rect 46112 21888 46164 21894
rect 46112 21830 46164 21836
rect 45782 21788 46078 21808
rect 45838 21786 45862 21788
rect 45918 21786 45942 21788
rect 45998 21786 46022 21788
rect 45860 21734 45862 21786
rect 45924 21734 45936 21786
rect 45998 21734 46000 21786
rect 45838 21732 45862 21734
rect 45918 21732 45942 21734
rect 45998 21732 46022 21734
rect 45782 21712 46078 21732
rect 46124 21690 46152 21830
rect 46308 21690 46336 21966
rect 46112 21684 46164 21690
rect 46112 21626 46164 21632
rect 46296 21684 46348 21690
rect 46296 21626 46348 21632
rect 46952 21146 46980 26400
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47400 23180 47452 23186
rect 47400 23122 47452 23128
rect 47412 22982 47440 23122
rect 47504 23050 47532 24754
rect 47492 23044 47544 23050
rect 47492 22986 47544 22992
rect 47400 22976 47452 22982
rect 47400 22918 47452 22924
rect 47688 22030 47716 26400
rect 47860 23180 47912 23186
rect 47860 23122 47912 23128
rect 47872 22982 47900 23122
rect 47860 22976 47912 22982
rect 47860 22918 47912 22924
rect 47676 22024 47728 22030
rect 47676 21966 47728 21972
rect 47032 21480 47084 21486
rect 47032 21422 47084 21428
rect 45652 21140 45704 21146
rect 45652 21082 45704 21088
rect 46940 21140 46992 21146
rect 46940 21082 46992 21088
rect 45560 20460 45612 20466
rect 45560 20402 45612 20408
rect 45664 20058 45692 21082
rect 47044 21078 47072 21422
rect 47872 21350 47900 22918
rect 47860 21344 47912 21350
rect 47860 21286 47912 21292
rect 47032 21072 47084 21078
rect 47032 21014 47084 21020
rect 45928 21004 45980 21010
rect 45928 20946 45980 20952
rect 46664 21004 46716 21010
rect 46664 20946 46716 20952
rect 45940 20890 45968 20946
rect 45940 20862 46152 20890
rect 45782 20700 46078 20720
rect 45838 20698 45862 20700
rect 45918 20698 45942 20700
rect 45998 20698 46022 20700
rect 45860 20646 45862 20698
rect 45924 20646 45936 20698
rect 45998 20646 46000 20698
rect 45838 20644 45862 20646
rect 45918 20644 45942 20646
rect 45998 20644 46022 20646
rect 45782 20624 46078 20644
rect 46124 20330 46152 20862
rect 46676 20806 46704 20946
rect 46664 20800 46716 20806
rect 46664 20742 46716 20748
rect 46112 20324 46164 20330
rect 46112 20266 46164 20272
rect 45560 20052 45612 20058
rect 45560 19994 45612 20000
rect 45652 20052 45704 20058
rect 45652 19994 45704 20000
rect 46020 20052 46072 20058
rect 46020 19994 46072 20000
rect 45572 19904 45600 19994
rect 45744 19916 45796 19922
rect 45572 19876 45744 19904
rect 45744 19858 45796 19864
rect 46032 19854 46060 19994
rect 46020 19848 46072 19854
rect 46020 19790 46072 19796
rect 45782 19612 46078 19632
rect 45838 19610 45862 19612
rect 45918 19610 45942 19612
rect 45998 19610 46022 19612
rect 45860 19558 45862 19610
rect 45924 19558 45936 19610
rect 45998 19558 46000 19610
rect 45838 19556 45862 19558
rect 45918 19556 45942 19558
rect 45998 19556 46022 19558
rect 45782 19536 46078 19556
rect 44824 19508 44876 19514
rect 44824 19450 44876 19456
rect 44836 19310 44864 19450
rect 46124 19394 46152 20266
rect 46296 20256 46348 20262
rect 46296 20198 46348 20204
rect 46308 19922 46336 20198
rect 46388 20052 46440 20058
rect 46388 19994 46440 20000
rect 46296 19916 46348 19922
rect 46296 19858 46348 19864
rect 46400 19825 46428 19994
rect 46386 19816 46442 19825
rect 46386 19751 46442 19760
rect 46032 19378 46152 19394
rect 46020 19372 46152 19378
rect 46072 19366 46152 19372
rect 46020 19314 46072 19320
rect 44180 19304 44232 19310
rect 44180 19246 44232 19252
rect 44824 19304 44876 19310
rect 46112 19304 46164 19310
rect 44824 19246 44876 19252
rect 46110 19272 46112 19281
rect 46164 19272 46166 19281
rect 44088 19236 44140 19242
rect 44088 19178 44140 19184
rect 44192 18766 44220 19246
rect 46110 19207 46166 19216
rect 46676 19174 46704 20742
rect 46756 20392 46808 20398
rect 46756 20334 46808 20340
rect 46768 19242 46796 20334
rect 46940 20324 46992 20330
rect 46940 20266 46992 20272
rect 46952 19718 46980 20266
rect 46940 19712 46992 19718
rect 46940 19654 46992 19660
rect 47400 19712 47452 19718
rect 47400 19654 47452 19660
rect 47412 19514 47440 19654
rect 47400 19508 47452 19514
rect 47400 19450 47452 19456
rect 47872 19310 47900 21286
rect 48424 21010 48452 26400
rect 48504 24812 48556 24818
rect 48504 24754 48556 24760
rect 48516 23254 48544 24754
rect 48596 24608 48648 24614
rect 48596 24550 48648 24556
rect 48608 23730 48636 24550
rect 49068 23866 49096 26400
rect 49056 23860 49108 23866
rect 49056 23802 49108 23808
rect 48596 23724 48648 23730
rect 48596 23666 48648 23672
rect 48504 23248 48556 23254
rect 48504 23190 48556 23196
rect 48608 22574 48636 23666
rect 48964 22636 49016 22642
rect 48964 22578 49016 22584
rect 48596 22568 48648 22574
rect 48596 22510 48648 22516
rect 48608 21690 48636 22510
rect 48976 22234 49004 22578
rect 48964 22228 49016 22234
rect 48964 22170 49016 22176
rect 49804 22098 49832 26400
rect 50540 24410 50568 26400
rect 50620 24744 50672 24750
rect 50620 24686 50672 24692
rect 50528 24404 50580 24410
rect 50528 24346 50580 24352
rect 50632 24342 50660 24686
rect 51080 24608 51132 24614
rect 51080 24550 51132 24556
rect 50620 24336 50672 24342
rect 50620 24278 50672 24284
rect 51092 23050 51120 24550
rect 52368 23656 52420 23662
rect 52368 23598 52420 23604
rect 51816 23520 51868 23526
rect 51816 23462 51868 23468
rect 51724 23180 51776 23186
rect 51724 23122 51776 23128
rect 51080 23044 51132 23050
rect 51080 22986 51132 22992
rect 51448 22976 51500 22982
rect 51448 22918 51500 22924
rect 51460 22778 51488 22918
rect 51448 22772 51500 22778
rect 51448 22714 51500 22720
rect 49976 22432 50028 22438
rect 49976 22374 50028 22380
rect 49792 22092 49844 22098
rect 49792 22034 49844 22040
rect 48596 21684 48648 21690
rect 48596 21626 48648 21632
rect 48412 21004 48464 21010
rect 48412 20946 48464 20952
rect 48412 20392 48464 20398
rect 48412 20334 48464 20340
rect 48424 19310 48452 20334
rect 48608 19922 48636 21626
rect 49240 20256 49292 20262
rect 49240 20198 49292 20204
rect 49252 19922 49280 20198
rect 48596 19916 48648 19922
rect 48596 19858 48648 19864
rect 49240 19916 49292 19922
rect 49240 19858 49292 19864
rect 48504 19848 48556 19854
rect 48504 19790 48556 19796
rect 48516 19378 48544 19790
rect 48504 19372 48556 19378
rect 48504 19314 48556 19320
rect 49240 19372 49292 19378
rect 49240 19314 49292 19320
rect 47860 19304 47912 19310
rect 47860 19246 47912 19252
rect 48412 19304 48464 19310
rect 48412 19246 48464 19252
rect 48596 19304 48648 19310
rect 48596 19246 48648 19252
rect 49056 19304 49108 19310
rect 49056 19246 49108 19252
rect 46756 19236 46808 19242
rect 46756 19178 46808 19184
rect 47124 19236 47176 19242
rect 47124 19178 47176 19184
rect 46112 19168 46164 19174
rect 46204 19168 46256 19174
rect 46112 19110 46164 19116
rect 46202 19136 46204 19145
rect 46664 19168 46716 19174
rect 46256 19136 46258 19145
rect 44730 18864 44786 18873
rect 44456 18828 44508 18834
rect 44640 18828 44692 18834
rect 44508 18788 44588 18816
rect 44456 18770 44508 18776
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 44456 18692 44508 18698
rect 44456 18634 44508 18640
rect 44362 18320 44418 18329
rect 44468 18290 44496 18634
rect 44362 18255 44418 18264
rect 44456 18284 44508 18290
rect 42524 18216 42576 18222
rect 42522 18184 42524 18193
rect 42616 18216 42668 18222
rect 42576 18184 42578 18193
rect 44272 18216 44324 18222
rect 42616 18158 42668 18164
rect 44192 18176 44272 18204
rect 42522 18119 42578 18128
rect 42984 18148 43036 18154
rect 42984 18090 43036 18096
rect 42708 17128 42760 17134
rect 42708 17070 42760 17076
rect 42340 16788 42392 16794
rect 42340 16730 42392 16736
rect 40776 16652 40828 16658
rect 40776 16594 40828 16600
rect 41052 16652 41104 16658
rect 41052 16594 41104 16600
rect 41788 16652 41840 16658
rect 41788 16594 41840 16600
rect 40500 16584 40552 16590
rect 40500 16526 40552 16532
rect 42064 16584 42116 16590
rect 42064 16526 42116 16532
rect 40316 16448 40368 16454
rect 40316 16390 40368 16396
rect 40328 15434 40356 16390
rect 41788 16108 41840 16114
rect 41788 16050 41840 16056
rect 41800 15638 41828 16050
rect 42076 16046 42104 16526
rect 42720 16454 42748 17070
rect 42996 17066 43024 18090
rect 44192 17882 44220 18176
rect 44272 18158 44324 18164
rect 44180 17876 44232 17882
rect 44180 17818 44232 17824
rect 44088 17672 44140 17678
rect 44088 17614 44140 17620
rect 43996 17536 44048 17542
rect 43996 17478 44048 17484
rect 44008 17270 44036 17478
rect 44100 17338 44128 17614
rect 44088 17332 44140 17338
rect 44088 17274 44140 17280
rect 43996 17264 44048 17270
rect 43996 17206 44048 17212
rect 42984 17060 43036 17066
rect 42984 17002 43036 17008
rect 42892 16516 42944 16522
rect 42892 16458 42944 16464
rect 42708 16448 42760 16454
rect 42708 16390 42760 16396
rect 42720 16114 42748 16390
rect 42708 16108 42760 16114
rect 42708 16050 42760 16056
rect 42064 16040 42116 16046
rect 42064 15982 42116 15988
rect 42800 16040 42852 16046
rect 42800 15982 42852 15988
rect 41880 15972 41932 15978
rect 41880 15914 41932 15920
rect 41788 15632 41840 15638
rect 41788 15574 41840 15580
rect 40408 15564 40460 15570
rect 40408 15506 40460 15512
rect 40420 15450 40448 15506
rect 40316 15428 40368 15434
rect 40420 15422 40540 15450
rect 40316 15370 40368 15376
rect 40512 14958 40540 15422
rect 41696 15360 41748 15366
rect 41696 15302 41748 15308
rect 41512 15020 41564 15026
rect 41512 14962 41564 14968
rect 40500 14952 40552 14958
rect 40500 14894 40552 14900
rect 40132 14884 40184 14890
rect 40132 14826 40184 14832
rect 40144 14482 40172 14826
rect 40512 14618 40540 14894
rect 40500 14612 40552 14618
rect 40500 14554 40552 14560
rect 40132 14476 40184 14482
rect 40132 14418 40184 14424
rect 40224 14272 40276 14278
rect 40224 14214 40276 14220
rect 40236 13938 40264 14214
rect 41236 14068 41288 14074
rect 41236 14010 41288 14016
rect 41248 13954 41276 14010
rect 40224 13932 40276 13938
rect 41248 13926 41460 13954
rect 40224 13874 40276 13880
rect 40868 13864 40920 13870
rect 40868 13806 40920 13812
rect 40880 13394 40908 13806
rect 41328 13728 41380 13734
rect 41328 13670 41380 13676
rect 41340 13462 41368 13670
rect 41328 13456 41380 13462
rect 41328 13398 41380 13404
rect 41432 13394 41460 13926
rect 41524 13734 41552 14962
rect 41708 14346 41736 15302
rect 41892 14958 41920 15914
rect 42156 15904 42208 15910
rect 42156 15846 42208 15852
rect 42168 15638 42196 15846
rect 42156 15632 42208 15638
rect 42156 15574 42208 15580
rect 42812 14958 42840 15982
rect 41880 14952 41932 14958
rect 41880 14894 41932 14900
rect 42524 14952 42576 14958
rect 42524 14894 42576 14900
rect 42800 14952 42852 14958
rect 42800 14894 42852 14900
rect 42536 14482 42564 14894
rect 42812 14550 42840 14894
rect 42800 14544 42852 14550
rect 42800 14486 42852 14492
rect 42904 14482 42932 16458
rect 43536 16040 43588 16046
rect 43536 15982 43588 15988
rect 43548 15026 43576 15982
rect 44008 15706 44036 17206
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 43996 15700 44048 15706
rect 43996 15642 44048 15648
rect 44008 15502 44036 15642
rect 43996 15496 44048 15502
rect 43996 15438 44048 15444
rect 43536 15020 43588 15026
rect 43536 14962 43588 14968
rect 43720 14952 43772 14958
rect 43720 14894 43772 14900
rect 42524 14476 42576 14482
rect 42524 14418 42576 14424
rect 42892 14476 42944 14482
rect 42892 14418 42944 14424
rect 41696 14340 41748 14346
rect 41696 14282 41748 14288
rect 42156 14340 42208 14346
rect 42156 14282 42208 14288
rect 41696 13796 41748 13802
rect 41696 13738 41748 13744
rect 41512 13728 41564 13734
rect 41512 13670 41564 13676
rect 40868 13388 40920 13394
rect 40868 13330 40920 13336
rect 41420 13388 41472 13394
rect 41420 13330 41472 13336
rect 40868 13184 40920 13190
rect 40868 13126 40920 13132
rect 41052 13184 41104 13190
rect 41052 13126 41104 13132
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 39672 12844 39724 12850
rect 39672 12786 39724 12792
rect 39120 12776 39172 12782
rect 39120 12718 39172 12724
rect 36817 12540 37113 12560
rect 36873 12538 36897 12540
rect 36953 12538 36977 12540
rect 37033 12538 37057 12540
rect 36895 12486 36897 12538
rect 36959 12486 36971 12538
rect 37033 12486 37035 12538
rect 36873 12484 36897 12486
rect 36953 12484 36977 12486
rect 37033 12484 37057 12486
rect 36817 12464 37113 12484
rect 39132 11898 39160 12718
rect 39684 12714 39712 12786
rect 39580 12708 39632 12714
rect 39580 12650 39632 12656
rect 39672 12708 39724 12714
rect 39672 12650 39724 12656
rect 39592 12238 39620 12650
rect 40052 12646 40080 12854
rect 40040 12640 40092 12646
rect 40040 12582 40092 12588
rect 40316 12640 40368 12646
rect 40316 12582 40368 12588
rect 40328 12442 40356 12582
rect 40880 12442 40908 13126
rect 41064 12782 41092 13126
rect 41708 12986 41736 13738
rect 42168 13530 42196 14282
rect 43732 14074 43760 14894
rect 43720 14068 43772 14074
rect 43720 14010 43772 14016
rect 42708 13932 42760 13938
rect 42708 13874 42760 13880
rect 42156 13524 42208 13530
rect 42156 13466 42208 13472
rect 42720 13394 42748 13874
rect 44008 13870 44036 15438
rect 44192 15094 44220 16934
rect 44180 15088 44232 15094
rect 44180 15030 44232 15036
rect 44192 14618 44220 15030
rect 44376 14958 44404 18255
rect 44456 18226 44508 18232
rect 44560 17882 44588 18788
rect 44730 18799 44786 18808
rect 44640 18770 44692 18776
rect 44548 17876 44600 17882
rect 44548 17818 44600 17824
rect 44560 17338 44588 17818
rect 44548 17332 44600 17338
rect 44548 17274 44600 17280
rect 44652 16658 44680 18770
rect 44744 18222 44772 18799
rect 45008 18692 45060 18698
rect 45008 18634 45060 18640
rect 45652 18692 45704 18698
rect 45652 18634 45704 18640
rect 45020 18426 45048 18634
rect 45008 18420 45060 18426
rect 45008 18362 45060 18368
rect 44732 18216 44784 18222
rect 44732 18158 44784 18164
rect 45664 18154 45692 18634
rect 45782 18524 46078 18544
rect 45838 18522 45862 18524
rect 45918 18522 45942 18524
rect 45998 18522 46022 18524
rect 45860 18470 45862 18522
rect 45924 18470 45936 18522
rect 45998 18470 46000 18522
rect 45838 18468 45862 18470
rect 45918 18468 45942 18470
rect 45998 18468 46022 18470
rect 45782 18448 46078 18468
rect 46124 18290 46152 19110
rect 46664 19110 46716 19116
rect 46202 19071 46258 19080
rect 46940 18760 46992 18766
rect 46940 18702 46992 18708
rect 46112 18284 46164 18290
rect 46112 18226 46164 18232
rect 46296 18216 46348 18222
rect 46952 18193 46980 18702
rect 46296 18158 46348 18164
rect 46938 18184 46994 18193
rect 45652 18148 45704 18154
rect 45652 18090 45704 18096
rect 46308 17814 46336 18158
rect 46938 18119 46994 18128
rect 45560 17808 45612 17814
rect 45560 17750 45612 17756
rect 46296 17808 46348 17814
rect 46296 17750 46348 17756
rect 45192 17536 45244 17542
rect 45192 17478 45244 17484
rect 45204 17338 45232 17478
rect 45192 17332 45244 17338
rect 45192 17274 45244 17280
rect 45572 17134 45600 17750
rect 45652 17740 45704 17746
rect 45652 17682 45704 17688
rect 45560 17128 45612 17134
rect 45560 17070 45612 17076
rect 44640 16652 44692 16658
rect 44640 16594 44692 16600
rect 45468 16652 45520 16658
rect 45468 16594 45520 16600
rect 45480 15706 45508 16594
rect 45468 15700 45520 15706
rect 45468 15642 45520 15648
rect 45664 15026 45692 17682
rect 46480 17536 46532 17542
rect 46480 17478 46532 17484
rect 45782 17436 46078 17456
rect 45838 17434 45862 17436
rect 45918 17434 45942 17436
rect 45998 17434 46022 17436
rect 45860 17382 45862 17434
rect 45924 17382 45936 17434
rect 45998 17382 46000 17434
rect 45838 17380 45862 17382
rect 45918 17380 45942 17382
rect 45998 17380 46022 17382
rect 45782 17360 46078 17380
rect 46492 17202 46520 17478
rect 46480 17196 46532 17202
rect 46480 17138 46532 17144
rect 45782 16348 46078 16368
rect 45838 16346 45862 16348
rect 45918 16346 45942 16348
rect 45998 16346 46022 16348
rect 45860 16294 45862 16346
rect 45924 16294 45936 16346
rect 45998 16294 46000 16346
rect 45838 16292 45862 16294
rect 45918 16292 45942 16294
rect 45998 16292 46022 16294
rect 45782 16272 46078 16292
rect 46952 15570 46980 18119
rect 47136 17678 47164 19178
rect 48608 18970 48636 19246
rect 48596 18964 48648 18970
rect 48596 18906 48648 18912
rect 49068 18834 49096 19246
rect 49252 19174 49280 19314
rect 49608 19236 49660 19242
rect 49608 19178 49660 19184
rect 49240 19168 49292 19174
rect 49240 19110 49292 19116
rect 49252 18834 49280 19110
rect 49620 18902 49648 19178
rect 49608 18896 49660 18902
rect 49608 18838 49660 18844
rect 49988 18834 50016 22374
rect 51460 22234 51488 22714
rect 51448 22228 51500 22234
rect 51448 22170 51500 22176
rect 51736 22166 51764 23122
rect 51828 22506 51856 23462
rect 52380 23254 52408 23598
rect 53472 23520 53524 23526
rect 53472 23462 53524 23468
rect 53484 23322 53512 23462
rect 53472 23316 53524 23322
rect 53472 23258 53524 23264
rect 52368 23248 52420 23254
rect 52368 23190 52420 23196
rect 52000 23180 52052 23186
rect 52000 23122 52052 23128
rect 51816 22500 51868 22506
rect 51816 22442 51868 22448
rect 51724 22160 51776 22166
rect 51724 22102 51776 22108
rect 50068 22092 50120 22098
rect 50068 22034 50120 22040
rect 50712 22092 50764 22098
rect 50712 22034 50764 22040
rect 50080 21078 50108 22034
rect 50068 21072 50120 21078
rect 50068 21014 50120 21020
rect 50160 21004 50212 21010
rect 50160 20946 50212 20952
rect 50172 20602 50200 20946
rect 50160 20596 50212 20602
rect 50160 20538 50212 20544
rect 50724 20534 50752 22034
rect 51724 21548 51776 21554
rect 51828 21536 51856 22442
rect 52012 21978 52040 23122
rect 52460 22568 52512 22574
rect 52460 22510 52512 22516
rect 52012 21950 52132 21978
rect 52000 21888 52052 21894
rect 52000 21830 52052 21836
rect 52012 21554 52040 21830
rect 52104 21554 52132 21950
rect 52276 21956 52328 21962
rect 52276 21898 52328 21904
rect 51776 21508 51856 21536
rect 52000 21548 52052 21554
rect 51724 21490 51776 21496
rect 52000 21490 52052 21496
rect 52092 21548 52144 21554
rect 52092 21490 52144 21496
rect 51736 21146 51764 21490
rect 52104 21434 52132 21490
rect 52012 21406 52132 21434
rect 51724 21140 51776 21146
rect 51724 21082 51776 21088
rect 50712 20528 50764 20534
rect 50710 20496 50712 20505
rect 50764 20496 50766 20505
rect 50710 20431 50766 20440
rect 50712 20392 50764 20398
rect 50712 20334 50764 20340
rect 50724 19990 50752 20334
rect 51356 20324 51408 20330
rect 51356 20266 51408 20272
rect 50712 19984 50764 19990
rect 50712 19926 50764 19932
rect 50724 19310 50752 19926
rect 50712 19304 50764 19310
rect 50712 19246 50764 19252
rect 51368 18834 51396 20266
rect 51736 19990 51764 21082
rect 52012 20330 52040 21406
rect 52288 20806 52316 21898
rect 52472 21894 52500 22510
rect 54128 22438 54156 26400
rect 54864 24274 54892 26400
rect 54852 24268 54904 24274
rect 54852 24210 54904 24216
rect 54116 22432 54168 22438
rect 54116 22374 54168 22380
rect 52460 21888 52512 21894
rect 52460 21830 52512 21836
rect 52276 20800 52328 20806
rect 52276 20742 52328 20748
rect 52090 20496 52146 20505
rect 52090 20431 52146 20440
rect 52104 20398 52132 20431
rect 52092 20392 52144 20398
rect 52092 20334 52144 20340
rect 52000 20324 52052 20330
rect 52000 20266 52052 20272
rect 52288 20262 52316 20742
rect 52366 20496 52422 20505
rect 52366 20431 52422 20440
rect 52276 20256 52328 20262
rect 52276 20198 52328 20204
rect 51724 19984 51776 19990
rect 51724 19926 51776 19932
rect 52380 19446 52408 20431
rect 53380 20392 53432 20398
rect 53380 20334 53432 20340
rect 52920 20256 52972 20262
rect 52920 20198 52972 20204
rect 52932 20058 52960 20198
rect 53392 20058 53420 20334
rect 52920 20052 52972 20058
rect 52920 19994 52972 20000
rect 53380 20052 53432 20058
rect 53380 19994 53432 20000
rect 52736 19848 52788 19854
rect 52736 19790 52788 19796
rect 52368 19440 52420 19446
rect 52368 19382 52420 19388
rect 52460 19372 52512 19378
rect 52460 19314 52512 19320
rect 52472 18834 52500 19314
rect 52644 19236 52696 19242
rect 52644 19178 52696 19184
rect 47860 18828 47912 18834
rect 47860 18770 47912 18776
rect 48872 18828 48924 18834
rect 48872 18770 48924 18776
rect 49056 18828 49108 18834
rect 49056 18770 49108 18776
rect 49240 18828 49292 18834
rect 49240 18770 49292 18776
rect 49976 18828 50028 18834
rect 49976 18770 50028 18776
rect 51356 18828 51408 18834
rect 51356 18770 51408 18776
rect 52460 18828 52512 18834
rect 52460 18770 52512 18776
rect 47872 18737 47900 18770
rect 47858 18728 47914 18737
rect 47858 18663 47914 18672
rect 47952 18624 48004 18630
rect 47952 18566 48004 18572
rect 47964 18426 47992 18566
rect 47952 18420 48004 18426
rect 47952 18362 48004 18368
rect 48320 18216 48372 18222
rect 48320 18158 48372 18164
rect 48596 18216 48648 18222
rect 48596 18158 48648 18164
rect 47308 18080 47360 18086
rect 47308 18022 47360 18028
rect 47124 17672 47176 17678
rect 47044 17632 47124 17660
rect 47044 16114 47072 17632
rect 47124 17614 47176 17620
rect 47320 16726 47348 18022
rect 48332 17746 48360 18158
rect 48608 17882 48636 18158
rect 48596 17876 48648 17882
rect 48596 17818 48648 17824
rect 48320 17740 48372 17746
rect 48320 17682 48372 17688
rect 47492 17128 47544 17134
rect 47492 17070 47544 17076
rect 47950 17096 48006 17105
rect 47504 16794 47532 17070
rect 47950 17031 47952 17040
rect 48004 17031 48006 17040
rect 47952 17002 48004 17008
rect 47492 16788 47544 16794
rect 47492 16730 47544 16736
rect 47308 16720 47360 16726
rect 47308 16662 47360 16668
rect 47400 16652 47452 16658
rect 47400 16594 47452 16600
rect 47412 16250 47440 16594
rect 47400 16244 47452 16250
rect 47400 16186 47452 16192
rect 47032 16108 47084 16114
rect 47032 16050 47084 16056
rect 48136 16108 48188 16114
rect 48136 16050 48188 16056
rect 46756 15564 46808 15570
rect 46756 15506 46808 15512
rect 46940 15564 46992 15570
rect 46940 15506 46992 15512
rect 45782 15260 46078 15280
rect 45838 15258 45862 15260
rect 45918 15258 45942 15260
rect 45998 15258 46022 15260
rect 45860 15206 45862 15258
rect 45924 15206 45936 15258
rect 45998 15206 46000 15258
rect 45838 15204 45862 15206
rect 45918 15204 45942 15206
rect 45998 15204 46022 15206
rect 45782 15184 46078 15204
rect 45284 15020 45336 15026
rect 45284 14962 45336 14968
rect 45652 15020 45704 15026
rect 45652 14962 45704 14968
rect 44364 14952 44416 14958
rect 44364 14894 44416 14900
rect 45192 14952 45244 14958
rect 45192 14894 45244 14900
rect 44180 14612 44232 14618
rect 44180 14554 44232 14560
rect 43076 13864 43128 13870
rect 43076 13806 43128 13812
rect 43996 13864 44048 13870
rect 43996 13806 44048 13812
rect 42708 13388 42760 13394
rect 42708 13330 42760 13336
rect 41696 12980 41748 12986
rect 41696 12922 41748 12928
rect 41052 12776 41104 12782
rect 41052 12718 41104 12724
rect 41972 12640 42024 12646
rect 41972 12582 42024 12588
rect 40316 12436 40368 12442
rect 40316 12378 40368 12384
rect 40868 12436 40920 12442
rect 40868 12378 40920 12384
rect 39580 12232 39632 12238
rect 39580 12174 39632 12180
rect 41984 12102 42012 12582
rect 43088 12442 43116 13806
rect 44192 13410 44220 14554
rect 44732 14476 44784 14482
rect 44732 14418 44784 14424
rect 44192 13382 44312 13410
rect 44284 13326 44312 13382
rect 44456 13388 44508 13394
rect 44456 13330 44508 13336
rect 43628 13320 43680 13326
rect 43628 13262 43680 13268
rect 44088 13320 44140 13326
rect 44088 13262 44140 13268
rect 44272 13320 44324 13326
rect 44272 13262 44324 13268
rect 43076 12436 43128 12442
rect 43076 12378 43128 12384
rect 43640 12306 43668 13262
rect 44100 12918 44128 13262
rect 44088 12912 44140 12918
rect 44088 12854 44140 12860
rect 44284 12782 44312 13262
rect 44468 12850 44496 13330
rect 44456 12844 44508 12850
rect 44456 12786 44508 12792
rect 44272 12776 44324 12782
rect 44272 12718 44324 12724
rect 44744 12442 44772 14418
rect 45204 14074 45232 14894
rect 44824 14068 44876 14074
rect 44824 14010 44876 14016
rect 45192 14068 45244 14074
rect 45192 14010 45244 14016
rect 44836 13870 44864 14010
rect 45296 14006 45324 14962
rect 45284 14000 45336 14006
rect 45284 13942 45336 13948
rect 44824 13864 44876 13870
rect 44824 13806 44876 13812
rect 44836 12986 44864 13806
rect 45664 13530 45692 14962
rect 45836 14884 45888 14890
rect 45836 14826 45888 14832
rect 45848 14482 45876 14826
rect 46204 14816 46256 14822
rect 46204 14758 46256 14764
rect 45836 14476 45888 14482
rect 45836 14418 45888 14424
rect 46216 14414 46244 14758
rect 46768 14482 46796 15506
rect 47044 15450 47072 16050
rect 47216 15564 47268 15570
rect 47216 15506 47268 15512
rect 46952 15422 47072 15450
rect 46952 15162 46980 15422
rect 47032 15360 47084 15366
rect 47032 15302 47084 15308
rect 47044 15162 47072 15302
rect 46940 15156 46992 15162
rect 46940 15098 46992 15104
rect 47032 15156 47084 15162
rect 47032 15098 47084 15104
rect 46940 14884 46992 14890
rect 46940 14826 46992 14832
rect 46952 14482 46980 14826
rect 47228 14482 47256 15506
rect 47584 14952 47636 14958
rect 47584 14894 47636 14900
rect 47596 14550 47624 14894
rect 48148 14618 48176 16050
rect 48332 15162 48360 17682
rect 48884 17270 48912 18770
rect 49068 18290 49096 18770
rect 49056 18284 49108 18290
rect 49056 18226 49108 18232
rect 49056 18148 49108 18154
rect 49056 18090 49108 18096
rect 49884 18148 49936 18154
rect 49884 18090 49936 18096
rect 48872 17264 48924 17270
rect 48872 17206 48924 17212
rect 48504 16992 48556 16998
rect 48504 16934 48556 16940
rect 48516 16658 48544 16934
rect 49068 16726 49096 18090
rect 49896 17814 49924 18090
rect 49988 18086 50016 18770
rect 51356 18216 51408 18222
rect 51356 18158 51408 18164
rect 49976 18080 50028 18086
rect 49976 18022 50028 18028
rect 49884 17808 49936 17814
rect 49884 17750 49936 17756
rect 50804 17740 50856 17746
rect 50804 17682 50856 17688
rect 50252 17604 50304 17610
rect 50252 17546 50304 17552
rect 50264 17134 50292 17546
rect 50436 17264 50488 17270
rect 50436 17206 50488 17212
rect 50448 17134 50476 17206
rect 50816 17202 50844 17682
rect 51368 17678 51396 18158
rect 51632 18148 51684 18154
rect 51632 18090 51684 18096
rect 51644 17746 51672 18090
rect 52472 17882 52500 18770
rect 52552 18624 52604 18630
rect 52552 18566 52604 18572
rect 52564 18154 52592 18566
rect 52656 18222 52684 19178
rect 52748 18426 52776 19790
rect 53392 19258 53420 19994
rect 53300 19230 53420 19258
rect 53300 18834 53328 19230
rect 53380 19168 53432 19174
rect 53380 19110 53432 19116
rect 53392 18970 53420 19110
rect 53380 18964 53432 18970
rect 53380 18906 53432 18912
rect 53288 18828 53340 18834
rect 53288 18770 53340 18776
rect 52736 18420 52788 18426
rect 52736 18362 52788 18368
rect 52644 18216 52696 18222
rect 52644 18158 52696 18164
rect 52552 18148 52604 18154
rect 52552 18090 52604 18096
rect 52460 17876 52512 17882
rect 52460 17818 52512 17824
rect 53300 17746 53328 18770
rect 51632 17740 51684 17746
rect 51632 17682 51684 17688
rect 53288 17740 53340 17746
rect 53288 17682 53340 17688
rect 51356 17672 51408 17678
rect 51356 17614 51408 17620
rect 52368 17672 52420 17678
rect 52368 17614 52420 17620
rect 50896 17332 50948 17338
rect 50896 17274 50948 17280
rect 50804 17196 50856 17202
rect 50804 17138 50856 17144
rect 50252 17128 50304 17134
rect 50252 17070 50304 17076
rect 50436 17128 50488 17134
rect 50436 17070 50488 17076
rect 49056 16720 49108 16726
rect 49056 16662 49108 16668
rect 48504 16652 48556 16658
rect 48504 16594 48556 16600
rect 48596 16448 48648 16454
rect 48596 16390 48648 16396
rect 48608 16046 48636 16390
rect 48596 16040 48648 16046
rect 48596 15982 48648 15988
rect 48608 15638 48636 15982
rect 48964 15972 49016 15978
rect 48964 15914 49016 15920
rect 48596 15632 48648 15638
rect 48596 15574 48648 15580
rect 48976 15570 49004 15914
rect 49068 15570 49096 16662
rect 50160 16652 50212 16658
rect 50160 16594 50212 16600
rect 50172 15978 50200 16594
rect 50908 16522 50936 17274
rect 50988 17196 51040 17202
rect 51080 17196 51132 17202
rect 51040 17156 51080 17184
rect 50988 17138 51040 17144
rect 51368 17184 51396 17614
rect 52380 17202 52408 17614
rect 52368 17196 52420 17202
rect 51368 17156 51488 17184
rect 51080 17138 51132 17144
rect 51356 17060 51408 17066
rect 51356 17002 51408 17008
rect 51264 16992 51316 16998
rect 51264 16934 51316 16940
rect 51276 16522 51304 16934
rect 51368 16522 51396 17002
rect 51460 16658 51488 17156
rect 52368 17138 52420 17144
rect 51448 16652 51500 16658
rect 51448 16594 51500 16600
rect 51724 16652 51776 16658
rect 51724 16594 51776 16600
rect 50896 16516 50948 16522
rect 50896 16458 50948 16464
rect 51264 16516 51316 16522
rect 51264 16458 51316 16464
rect 51356 16516 51408 16522
rect 51356 16458 51408 16464
rect 50620 16176 50672 16182
rect 50620 16118 50672 16124
rect 50160 15972 50212 15978
rect 50160 15914 50212 15920
rect 48964 15564 49016 15570
rect 48964 15506 49016 15512
rect 49056 15564 49108 15570
rect 49056 15506 49108 15512
rect 49608 15496 49660 15502
rect 49608 15438 49660 15444
rect 48320 15156 48372 15162
rect 48320 15098 48372 15104
rect 48136 14612 48188 14618
rect 48136 14554 48188 14560
rect 49620 14550 49648 15438
rect 50172 14958 50200 15914
rect 50632 15570 50660 16118
rect 51276 16046 51304 16458
rect 51264 16040 51316 16046
rect 51264 15982 51316 15988
rect 51368 15570 51396 16458
rect 50620 15564 50672 15570
rect 50620 15506 50672 15512
rect 51356 15564 51408 15570
rect 51356 15506 51408 15512
rect 50632 15162 50660 15506
rect 51460 15162 51488 16594
rect 51736 15638 51764 16594
rect 52368 16584 52420 16590
rect 52368 16526 52420 16532
rect 52380 16114 52408 16526
rect 53472 16516 53524 16522
rect 53472 16458 53524 16464
rect 53484 16250 53512 16458
rect 53472 16244 53524 16250
rect 53472 16186 53524 16192
rect 52368 16108 52420 16114
rect 52368 16050 52420 16056
rect 51816 15904 51868 15910
rect 51816 15846 51868 15852
rect 51724 15632 51776 15638
rect 51724 15574 51776 15580
rect 50620 15156 50672 15162
rect 50620 15098 50672 15104
rect 51448 15156 51500 15162
rect 51448 15098 51500 15104
rect 50160 14952 50212 14958
rect 50160 14894 50212 14900
rect 49700 14816 49752 14822
rect 49700 14758 49752 14764
rect 47584 14544 47636 14550
rect 47584 14486 47636 14492
rect 49608 14544 49660 14550
rect 49608 14486 49660 14492
rect 49712 14482 49740 14758
rect 46756 14476 46808 14482
rect 46756 14418 46808 14424
rect 46940 14476 46992 14482
rect 46940 14418 46992 14424
rect 47216 14476 47268 14482
rect 47216 14418 47268 14424
rect 49700 14476 49752 14482
rect 49700 14418 49752 14424
rect 46204 14408 46256 14414
rect 46204 14350 46256 14356
rect 45782 14172 46078 14192
rect 45838 14170 45862 14172
rect 45918 14170 45942 14172
rect 45998 14170 46022 14172
rect 45860 14118 45862 14170
rect 45924 14118 45936 14170
rect 45998 14118 46000 14170
rect 45838 14116 45862 14118
rect 45918 14116 45942 14118
rect 45998 14116 46022 14118
rect 45782 14096 46078 14116
rect 45652 13524 45704 13530
rect 45652 13466 45704 13472
rect 46216 13394 46244 14350
rect 47228 14346 47256 14418
rect 47216 14340 47268 14346
rect 47216 14282 47268 14288
rect 49608 14272 49660 14278
rect 49608 14214 49660 14220
rect 49620 13870 49648 14214
rect 49712 13938 49740 14418
rect 50712 14340 50764 14346
rect 50712 14282 50764 14288
rect 49792 14272 49844 14278
rect 49792 14214 49844 14220
rect 49804 14074 49832 14214
rect 50724 14074 50752 14282
rect 51460 14278 51488 15098
rect 51828 14278 51856 15846
rect 55600 15026 55628 26400
rect 55588 15020 55640 15026
rect 55588 14962 55640 14968
rect 52000 14952 52052 14958
rect 52000 14894 52052 14900
rect 51448 14272 51500 14278
rect 51448 14214 51500 14220
rect 51816 14272 51868 14278
rect 51816 14214 51868 14220
rect 49792 14068 49844 14074
rect 49792 14010 49844 14016
rect 50712 14068 50764 14074
rect 50712 14010 50764 14016
rect 49700 13932 49752 13938
rect 49700 13874 49752 13880
rect 47308 13864 47360 13870
rect 47308 13806 47360 13812
rect 49608 13864 49660 13870
rect 49608 13806 49660 13812
rect 51448 13864 51500 13870
rect 51448 13806 51500 13812
rect 47124 13796 47176 13802
rect 47124 13738 47176 13744
rect 46756 13456 46808 13462
rect 46756 13398 46808 13404
rect 46204 13388 46256 13394
rect 46204 13330 46256 13336
rect 46572 13388 46624 13394
rect 46572 13330 46624 13336
rect 45782 13084 46078 13104
rect 45838 13082 45862 13084
rect 45918 13082 45942 13084
rect 45998 13082 46022 13084
rect 45860 13030 45862 13082
rect 45924 13030 45936 13082
rect 45998 13030 46000 13082
rect 45838 13028 45862 13030
rect 45918 13028 45942 13030
rect 45998 13028 46022 13030
rect 45782 13008 46078 13028
rect 44824 12980 44876 12986
rect 44824 12922 44876 12928
rect 46584 12782 46612 13330
rect 46768 12782 46796 13398
rect 47136 12850 47164 13738
rect 47320 13394 47348 13806
rect 48228 13796 48280 13802
rect 48228 13738 48280 13744
rect 47308 13388 47360 13394
rect 47308 13330 47360 13336
rect 47860 13320 47912 13326
rect 47860 13262 47912 13268
rect 47872 12986 47900 13262
rect 47860 12980 47912 12986
rect 47860 12922 47912 12928
rect 48240 12850 48268 13738
rect 49700 13728 49752 13734
rect 49700 13670 49752 13676
rect 49712 13394 49740 13670
rect 51460 13530 51488 13806
rect 51448 13524 51500 13530
rect 51448 13466 51500 13472
rect 49700 13388 49752 13394
rect 49700 13330 49752 13336
rect 51828 13326 51856 14214
rect 52012 14074 52040 14894
rect 52276 14884 52328 14890
rect 52276 14826 52328 14832
rect 52288 14482 52316 14826
rect 52276 14476 52328 14482
rect 52276 14418 52328 14424
rect 52460 14272 52512 14278
rect 52460 14214 52512 14220
rect 52472 14074 52500 14214
rect 52000 14068 52052 14074
rect 52000 14010 52052 14016
rect 52460 14068 52512 14074
rect 52460 14010 52512 14016
rect 51816 13320 51868 13326
rect 51816 13262 51868 13268
rect 49332 13184 49384 13190
rect 49332 13126 49384 13132
rect 49344 12986 49372 13126
rect 49332 12980 49384 12986
rect 49332 12922 49384 12928
rect 47124 12844 47176 12850
rect 47124 12786 47176 12792
rect 48228 12844 48280 12850
rect 48228 12786 48280 12792
rect 46572 12776 46624 12782
rect 46572 12718 46624 12724
rect 46756 12776 46808 12782
rect 46756 12718 46808 12724
rect 44732 12436 44784 12442
rect 44732 12378 44784 12384
rect 43628 12300 43680 12306
rect 43628 12242 43680 12248
rect 41972 12096 42024 12102
rect 41972 12038 42024 12044
rect 45782 11996 46078 12016
rect 45838 11994 45862 11996
rect 45918 11994 45942 11996
rect 45998 11994 46022 11996
rect 45860 11942 45862 11994
rect 45924 11942 45936 11994
rect 45998 11942 46000 11994
rect 45838 11940 45862 11942
rect 45918 11940 45942 11942
rect 45998 11940 46022 11942
rect 45782 11920 46078 11940
rect 36452 11892 36504 11898
rect 36452 11834 36504 11840
rect 36820 11892 36872 11898
rect 36820 11834 36872 11840
rect 39120 11892 39172 11898
rect 39120 11834 39172 11840
rect 36832 11762 36860 11834
rect 36820 11756 36872 11762
rect 36820 11698 36872 11704
rect 35624 11688 35676 11694
rect 35624 11630 35676 11636
rect 36817 11452 37113 11472
rect 36873 11450 36897 11452
rect 36953 11450 36977 11452
rect 37033 11450 37057 11452
rect 36895 11398 36897 11450
rect 36959 11398 36971 11450
rect 37033 11398 37035 11450
rect 36873 11396 36897 11398
rect 36953 11396 36977 11398
rect 37033 11396 37057 11398
rect 36817 11376 37113 11396
rect 35072 11280 35124 11286
rect 35072 11222 35124 11228
rect 33232 11212 33284 11218
rect 33232 11154 33284 11160
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 34704 11212 34756 11218
rect 34704 11154 34756 11160
rect 45782 10908 46078 10928
rect 45838 10906 45862 10908
rect 45918 10906 45942 10908
rect 45998 10906 46022 10908
rect 45860 10854 45862 10906
rect 45924 10854 45936 10906
rect 45998 10854 46000 10906
rect 45838 10852 45862 10854
rect 45918 10852 45942 10854
rect 45998 10852 46022 10854
rect 45782 10832 46078 10852
rect 32220 10804 32272 10810
rect 32220 10746 32272 10752
rect 32956 10804 33008 10810
rect 32956 10746 33008 10752
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 31116 10600 31168 10606
rect 31116 10542 31168 10548
rect 34520 10600 34572 10606
rect 34520 10542 34572 10548
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 27436 10260 27488 10266
rect 27436 10202 27488 10208
rect 27436 10124 27488 10130
rect 27436 10066 27488 10072
rect 27528 10124 27580 10130
rect 27528 10066 27580 10072
rect 27448 9722 27476 10066
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27540 9178 27568 10066
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27632 9518 27660 9862
rect 27852 9820 28148 9840
rect 27908 9818 27932 9820
rect 27988 9818 28012 9820
rect 28068 9818 28092 9820
rect 27930 9766 27932 9818
rect 27994 9766 28006 9818
rect 28068 9766 28070 9818
rect 27908 9764 27932 9766
rect 27988 9764 28012 9766
rect 28068 9764 28092 9766
rect 27852 9744 28148 9764
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 28724 9512 28776 9518
rect 28724 9454 28776 9460
rect 28736 9178 28764 9454
rect 27528 9172 27580 9178
rect 27528 9114 27580 9120
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 27252 9104 27304 9110
rect 27252 9046 27304 9052
rect 27160 9036 27212 9042
rect 27160 8978 27212 8984
rect 27172 8634 27200 8978
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 27852 8732 28148 8752
rect 27908 8730 27932 8732
rect 27988 8730 28012 8732
rect 28068 8730 28092 8732
rect 27930 8678 27932 8730
rect 27994 8678 28006 8730
rect 28068 8678 28070 8730
rect 27908 8676 27932 8678
rect 27988 8676 28012 8678
rect 28068 8676 28092 8678
rect 27852 8656 28148 8676
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 27356 8090 27384 8366
rect 28368 8090 28396 8366
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28736 7954 28764 8774
rect 29012 8022 29040 10406
rect 29288 10266 29316 10542
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 29000 8016 29052 8022
rect 29000 7958 29052 7964
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 28724 7948 28776 7954
rect 28724 7890 28776 7896
rect 27356 7546 27384 7890
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27540 7342 27568 7686
rect 27852 7644 28148 7664
rect 27908 7642 27932 7644
rect 27988 7642 28012 7644
rect 28068 7642 28092 7644
rect 27930 7590 27932 7642
rect 27994 7590 28006 7642
rect 28068 7590 28070 7642
rect 27908 7588 27932 7590
rect 27988 7588 28012 7590
rect 28068 7588 28092 7590
rect 27852 7568 28148 7588
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 27632 6254 27660 6598
rect 27852 6556 28148 6576
rect 27908 6554 27932 6556
rect 27988 6554 28012 6556
rect 28068 6554 28092 6556
rect 27930 6502 27932 6554
rect 27994 6502 28006 6554
rect 28068 6502 28070 6554
rect 27908 6500 27932 6502
rect 27988 6500 28012 6502
rect 28068 6500 28092 6502
rect 27852 6480 28148 6500
rect 29380 6458 29408 10542
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 32864 10124 32916 10130
rect 32864 10066 32916 10072
rect 34244 10124 34296 10130
rect 34244 10066 34296 10072
rect 29472 9450 29500 10066
rect 29564 9654 29592 10066
rect 30748 9920 30800 9926
rect 30748 9862 30800 9868
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29460 9444 29512 9450
rect 29460 9386 29512 9392
rect 29748 9178 29776 9454
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 29552 9036 29604 9042
rect 29552 8978 29604 8984
rect 30564 9036 30616 9042
rect 30564 8978 30616 8984
rect 29564 8090 29592 8978
rect 30576 8634 30604 8978
rect 30564 8628 30616 8634
rect 30564 8570 30616 8576
rect 29736 8560 29788 8566
rect 29736 8502 29788 8508
rect 29552 8084 29604 8090
rect 29552 8026 29604 8032
rect 29748 6866 29776 8502
rect 30760 8430 30788 9862
rect 31760 9512 31812 9518
rect 31760 9454 31812 9460
rect 32128 9512 32180 9518
rect 32128 9454 32180 9460
rect 30932 9376 30984 9382
rect 30932 9318 30984 9324
rect 30944 9042 30972 9318
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 31208 8832 31260 8838
rect 31208 8774 31260 8780
rect 31220 8430 31248 8774
rect 31772 8634 31800 9454
rect 32140 9178 32168 9454
rect 32312 9376 32364 9382
rect 32312 9318 32364 9324
rect 32128 9172 32180 9178
rect 32128 9114 32180 9120
rect 31760 8628 31812 8634
rect 31760 8570 31812 8576
rect 30748 8424 30800 8430
rect 30748 8366 30800 8372
rect 31208 8424 31260 8430
rect 31208 8366 31260 8372
rect 30012 7948 30064 7954
rect 30012 7890 30064 7896
rect 30024 7546 30052 7890
rect 30012 7540 30064 7546
rect 30012 7482 30064 7488
rect 32324 7342 32352 9318
rect 32772 9036 32824 9042
rect 32772 8978 32824 8984
rect 32784 8634 32812 8978
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32876 7546 32904 10066
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 33324 9920 33376 9926
rect 33324 9862 33376 9868
rect 32968 8430 32996 9862
rect 33140 9512 33192 9518
rect 33140 9454 33192 9460
rect 33152 9178 33180 9454
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33336 9042 33364 9862
rect 34256 9654 34284 10066
rect 34244 9648 34296 9654
rect 34244 9590 34296 9596
rect 34532 9382 34560 10542
rect 37188 10464 37240 10470
rect 37188 10406 37240 10412
rect 36817 10364 37113 10384
rect 36873 10362 36897 10364
rect 36953 10362 36977 10364
rect 37033 10362 37057 10364
rect 36895 10310 36897 10362
rect 36959 10310 36971 10362
rect 37033 10310 37035 10362
rect 36873 10308 36897 10310
rect 36953 10308 36977 10310
rect 37033 10308 37057 10310
rect 36817 10288 37113 10308
rect 36176 10124 36228 10130
rect 36176 10066 36228 10072
rect 35992 9920 36044 9926
rect 35992 9862 36044 9868
rect 35808 9512 35860 9518
rect 35808 9454 35860 9460
rect 34520 9376 34572 9382
rect 34520 9318 34572 9324
rect 33324 9036 33376 9042
rect 33324 8978 33376 8984
rect 35348 9036 35400 9042
rect 35348 8978 35400 8984
rect 33968 8832 34020 8838
rect 33968 8774 34020 8780
rect 35164 8832 35216 8838
rect 35164 8774 35216 8780
rect 33980 8430 34008 8774
rect 34520 8560 34572 8566
rect 34520 8502 34572 8508
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 33968 8424 34020 8430
rect 33968 8366 34020 8372
rect 34532 7954 34560 8502
rect 34612 8424 34664 8430
rect 34612 8366 34664 8372
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 32864 7540 32916 7546
rect 32864 7482 32916 7488
rect 30196 7336 30248 7342
rect 30196 7278 30248 7284
rect 32312 7336 32364 7342
rect 32312 7278 32364 7284
rect 30208 7002 30236 7278
rect 30196 6996 30248 7002
rect 30196 6938 30248 6944
rect 34532 6934 34560 7686
rect 34624 7546 34652 8366
rect 34980 8288 35032 8294
rect 34980 8230 35032 8236
rect 34992 7954 35020 8230
rect 34980 7948 35032 7954
rect 34980 7890 35032 7896
rect 35072 7948 35124 7954
rect 35072 7890 35124 7896
rect 34612 7540 34664 7546
rect 34612 7482 34664 7488
rect 34520 6928 34572 6934
rect 34520 6870 34572 6876
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 34428 6792 34480 6798
rect 34612 6792 34664 6798
rect 34480 6740 34612 6746
rect 34428 6734 34664 6740
rect 34440 6718 34652 6734
rect 33968 6656 34020 6662
rect 33968 6598 34020 6604
rect 29368 6452 29420 6458
rect 29368 6394 29420 6400
rect 33980 6254 34008 6598
rect 35084 6458 35112 7890
rect 35176 7342 35204 8774
rect 35360 8090 35388 8978
rect 35820 8634 35848 9454
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 36004 8498 36032 9862
rect 36188 9654 36216 10066
rect 36820 9920 36872 9926
rect 36820 9862 36872 9868
rect 36176 9648 36228 9654
rect 36176 9590 36228 9596
rect 36832 9518 36860 9862
rect 36820 9512 36872 9518
rect 36820 9454 36872 9460
rect 36728 9376 36780 9382
rect 36728 9318 36780 9324
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 36740 8430 36768 9318
rect 36817 9276 37113 9296
rect 36873 9274 36897 9276
rect 36953 9274 36977 9276
rect 37033 9274 37057 9276
rect 36895 9222 36897 9274
rect 36959 9222 36971 9274
rect 37033 9222 37035 9274
rect 36873 9220 36897 9222
rect 36953 9220 36977 9222
rect 37033 9220 37057 9222
rect 36817 9200 37113 9220
rect 37200 9110 37228 10406
rect 37648 10124 37700 10130
rect 37648 10066 37700 10072
rect 37660 9654 37688 10066
rect 45782 9820 46078 9840
rect 45838 9818 45862 9820
rect 45918 9818 45942 9820
rect 45998 9818 46022 9820
rect 45860 9766 45862 9818
rect 45924 9766 45936 9818
rect 45998 9766 46000 9818
rect 45838 9764 45862 9766
rect 45918 9764 45942 9766
rect 45998 9764 46022 9766
rect 45782 9744 46078 9764
rect 37648 9648 37700 9654
rect 37648 9590 37700 9596
rect 38476 9512 38528 9518
rect 38476 9454 38528 9460
rect 38488 9178 38516 9454
rect 38476 9172 38528 9178
rect 38476 9114 38528 9120
rect 37188 9104 37240 9110
rect 37188 9046 37240 9052
rect 37648 9036 37700 9042
rect 37648 8978 37700 8984
rect 37660 8634 37688 8978
rect 45782 8732 46078 8752
rect 45838 8730 45862 8732
rect 45918 8730 45942 8732
rect 45998 8730 46022 8732
rect 45860 8678 45862 8730
rect 45924 8678 45936 8730
rect 45998 8678 46000 8730
rect 45838 8676 45862 8678
rect 45918 8676 45942 8678
rect 45998 8676 46022 8678
rect 45782 8656 46078 8676
rect 37648 8628 37700 8634
rect 37648 8570 37700 8576
rect 36728 8424 36780 8430
rect 36728 8366 36780 8372
rect 36817 8188 37113 8208
rect 36873 8186 36897 8188
rect 36953 8186 36977 8188
rect 37033 8186 37057 8188
rect 36895 8134 36897 8186
rect 36959 8134 36971 8186
rect 37033 8134 37035 8186
rect 36873 8132 36897 8134
rect 36953 8132 36977 8134
rect 37033 8132 37057 8134
rect 36817 8112 37113 8132
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 36084 7948 36136 7954
rect 36084 7890 36136 7896
rect 35808 7744 35860 7750
rect 35808 7686 35860 7692
rect 35900 7744 35952 7750
rect 35900 7686 35952 7692
rect 35820 7342 35848 7686
rect 35164 7336 35216 7342
rect 35164 7278 35216 7284
rect 35808 7336 35860 7342
rect 35808 7278 35860 7284
rect 35808 7200 35860 7206
rect 35808 7142 35860 7148
rect 35820 6866 35848 7142
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35072 6452 35124 6458
rect 35072 6394 35124 6400
rect 35912 6254 35940 7686
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 30196 6248 30248 6254
rect 30196 6190 30248 6196
rect 33968 6248 34020 6254
rect 33968 6190 34020 6196
rect 35900 6248 35952 6254
rect 35900 6190 35952 6196
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 26528 4758 26556 6054
rect 29092 5772 29144 5778
rect 29092 5714 29144 5720
rect 26608 5568 26660 5574
rect 26608 5510 26660 5516
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 26620 5166 26648 5510
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26516 4752 26568 4758
rect 26516 4694 26568 4700
rect 26620 4078 26648 4966
rect 27356 4690 27384 5510
rect 27852 5468 28148 5488
rect 27908 5466 27932 5468
rect 27988 5466 28012 5468
rect 28068 5466 28092 5468
rect 27930 5414 27932 5466
rect 27994 5414 28006 5466
rect 28068 5414 28070 5466
rect 27908 5412 27932 5414
rect 27988 5412 28012 5414
rect 28068 5412 28092 5414
rect 27852 5392 28148 5412
rect 27712 5160 27764 5166
rect 27712 5102 27764 5108
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27540 4690 27568 4966
rect 27344 4684 27396 4690
rect 27344 4626 27396 4632
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27632 4078 27660 4422
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27724 3942 27752 5102
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 27852 4380 28148 4400
rect 27908 4378 27932 4380
rect 27988 4378 28012 4380
rect 28068 4378 28092 4380
rect 27930 4326 27932 4378
rect 27994 4326 28006 4378
rect 28068 4326 28070 4378
rect 27908 4324 27932 4326
rect 27988 4324 28012 4326
rect 28068 4324 28092 4326
rect 27852 4304 28148 4324
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 28276 3738 28304 4014
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26804 3194 26832 3538
rect 27852 3292 28148 3312
rect 27908 3290 27932 3292
rect 27988 3290 28012 3292
rect 28068 3290 28092 3292
rect 27930 3238 27932 3290
rect 27994 3238 28006 3290
rect 28068 3238 28070 3290
rect 27908 3236 27932 3238
rect 27988 3236 28012 3238
rect 28068 3236 28092 3238
rect 27852 3216 28148 3236
rect 26792 3188 26844 3194
rect 26792 3130 26844 3136
rect 28368 3058 28396 4422
rect 29012 3942 29040 4626
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 28448 3596 28500 3602
rect 28448 3538 28500 3544
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 24952 2984 25004 2990
rect 24952 2926 25004 2932
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 22940 2650 22968 2926
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 23492 2310 23520 2518
rect 23860 2514 23888 2790
rect 27816 2514 27844 2790
rect 28460 2650 28488 3538
rect 29104 3126 29132 5714
rect 29276 5568 29328 5574
rect 29276 5510 29328 5516
rect 29288 5234 29316 5510
rect 29840 5234 29868 6054
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 29092 3120 29144 3126
rect 29092 3062 29144 3068
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 27804 2508 27856 2514
rect 27804 2450 27856 2456
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 9921 2204 10217 2224
rect 9977 2202 10001 2204
rect 10057 2202 10081 2204
rect 10137 2202 10161 2204
rect 9999 2150 10001 2202
rect 10063 2150 10075 2202
rect 10137 2150 10139 2202
rect 9977 2148 10001 2150
rect 10057 2148 10081 2150
rect 10137 2148 10161 2150
rect 9921 2128 10217 2148
rect 19812 2106 19840 2246
rect 27852 2204 28148 2224
rect 27908 2202 27932 2204
rect 27988 2202 28012 2204
rect 28068 2202 28092 2204
rect 27930 2150 27932 2202
rect 27994 2150 28006 2202
rect 28068 2150 28070 2202
rect 27908 2148 27932 2150
rect 27988 2148 28012 2150
rect 28068 2148 28092 2150
rect 27852 2128 28148 2148
rect 29196 2106 29224 5102
rect 29460 4480 29512 4486
rect 29460 4422 29512 4428
rect 29472 3602 29500 4422
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 29288 2990 29316 3334
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 30208 2650 30236 6190
rect 34336 6180 34388 6186
rect 34336 6122 34388 6128
rect 31484 6112 31536 6118
rect 31484 6054 31536 6060
rect 30472 5772 30524 5778
rect 30472 5714 30524 5720
rect 30380 5024 30432 5030
rect 30380 4966 30432 4972
rect 30196 2644 30248 2650
rect 30196 2586 30248 2592
rect 30392 2582 30420 4966
rect 30484 4826 30512 5714
rect 30472 4820 30524 4826
rect 30472 4762 30524 4768
rect 31496 4690 31524 6054
rect 33508 5296 33560 5302
rect 33508 5238 33560 5244
rect 30472 4684 30524 4690
rect 30472 4626 30524 4632
rect 31484 4684 31536 4690
rect 31484 4626 31536 4632
rect 33048 4684 33100 4690
rect 33048 4626 33100 4632
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 30484 2378 30512 4626
rect 33060 4282 33088 4626
rect 33048 4276 33100 4282
rect 33048 4218 33100 4224
rect 31852 4072 31904 4078
rect 31852 4014 31904 4020
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 30564 3596 30616 3602
rect 30564 3538 30616 3544
rect 30576 3194 30604 3538
rect 31208 3392 31260 3398
rect 31208 3334 31260 3340
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 31220 2990 31248 3334
rect 31312 2990 31340 3878
rect 31680 3602 31708 3878
rect 31668 3596 31720 3602
rect 31668 3538 31720 3544
rect 31864 3466 31892 4014
rect 33048 4004 33100 4010
rect 33048 3946 33100 3952
rect 31852 3460 31904 3466
rect 31852 3402 31904 3408
rect 33060 3194 33088 3946
rect 33232 3392 33284 3398
rect 33232 3334 33284 3340
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 33244 2990 33272 3334
rect 31024 2984 31076 2990
rect 31024 2926 31076 2932
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 30656 2848 30708 2854
rect 30656 2790 30708 2796
rect 30668 2514 30696 2790
rect 31036 2650 31064 2926
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 31680 2514 31708 2790
rect 33520 2514 33548 5238
rect 34060 4480 34112 4486
rect 34060 4422 34112 4428
rect 33692 4072 33744 4078
rect 33692 4014 33744 4020
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33704 3466 33732 4014
rect 33888 3738 33916 4014
rect 33876 3732 33928 3738
rect 33876 3674 33928 3680
rect 34072 3602 34100 4422
rect 34244 3936 34296 3942
rect 34244 3878 34296 3884
rect 34060 3596 34112 3602
rect 34060 3538 34112 3544
rect 33692 3460 33744 3466
rect 33692 3402 33744 3408
rect 34256 2990 34284 3878
rect 34244 2984 34296 2990
rect 34244 2926 34296 2932
rect 34348 2650 34376 6122
rect 36004 5778 36032 7142
rect 36096 6730 36124 7890
rect 45782 7644 46078 7664
rect 45838 7642 45862 7644
rect 45918 7642 45942 7644
rect 45998 7642 46022 7644
rect 45860 7590 45862 7642
rect 45924 7590 45936 7642
rect 45998 7590 46000 7642
rect 45838 7588 45862 7590
rect 45918 7588 45942 7590
rect 45998 7588 46022 7590
rect 45782 7568 46078 7588
rect 36176 7336 36228 7342
rect 36176 7278 36228 7284
rect 38016 7336 38068 7342
rect 38016 7278 38068 7284
rect 36084 6724 36136 6730
rect 36084 6666 36136 6672
rect 36188 6458 36216 7278
rect 36817 7100 37113 7120
rect 36873 7098 36897 7100
rect 36953 7098 36977 7100
rect 37033 7098 37057 7100
rect 36895 7046 36897 7098
rect 36959 7046 36971 7098
rect 37033 7046 37035 7098
rect 36873 7044 36897 7046
rect 36953 7044 36977 7046
rect 37033 7044 37057 7046
rect 36817 7024 37113 7044
rect 36268 6860 36320 6866
rect 36268 6802 36320 6808
rect 36176 6452 36228 6458
rect 36176 6394 36228 6400
rect 36280 5914 36308 6802
rect 38028 6730 38056 7278
rect 39856 7200 39908 7206
rect 39856 7142 39908 7148
rect 38660 6860 38712 6866
rect 38660 6802 38712 6808
rect 38016 6724 38068 6730
rect 38016 6666 38068 6672
rect 38672 6458 38700 6802
rect 38844 6656 38896 6662
rect 38844 6598 38896 6604
rect 38936 6656 38988 6662
rect 38936 6598 38988 6604
rect 38660 6452 38712 6458
rect 38660 6394 38712 6400
rect 37188 6248 37240 6254
rect 37188 6190 37240 6196
rect 36817 6012 37113 6032
rect 36873 6010 36897 6012
rect 36953 6010 36977 6012
rect 37033 6010 37057 6012
rect 36895 5958 36897 6010
rect 36959 5958 36971 6010
rect 37033 5958 37035 6010
rect 36873 5956 36897 5958
rect 36953 5956 36977 5958
rect 37033 5956 37057 5958
rect 36817 5936 37113 5956
rect 37200 5914 37228 6190
rect 38568 6180 38620 6186
rect 38568 6122 38620 6128
rect 37280 6112 37332 6118
rect 37280 6054 37332 6060
rect 36268 5908 36320 5914
rect 36268 5850 36320 5856
rect 37188 5908 37240 5914
rect 37188 5850 37240 5856
rect 35992 5772 36044 5778
rect 35992 5714 36044 5720
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34336 2644 34388 2650
rect 34336 2586 34388 2592
rect 34532 2514 34560 5510
rect 37292 5166 37320 6054
rect 37372 5772 37424 5778
rect 37372 5714 37424 5720
rect 37384 5370 37412 5714
rect 37556 5568 37608 5574
rect 37556 5510 37608 5516
rect 37372 5364 37424 5370
rect 37372 5306 37424 5312
rect 37568 5166 37596 5510
rect 38580 5370 38608 6122
rect 38568 5364 38620 5370
rect 38568 5306 38620 5312
rect 37280 5160 37332 5166
rect 37280 5102 37332 5108
rect 37556 5160 37608 5166
rect 37556 5102 37608 5108
rect 38752 5160 38804 5166
rect 38752 5102 38804 5108
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 36817 4924 37113 4944
rect 36873 4922 36897 4924
rect 36953 4922 36977 4924
rect 37033 4922 37057 4924
rect 36895 4870 36897 4922
rect 36959 4870 36971 4922
rect 37033 4870 37035 4922
rect 36873 4868 36897 4870
rect 36953 4868 36977 4870
rect 37033 4868 37057 4870
rect 36817 4848 37113 4868
rect 37568 4690 37596 4966
rect 38764 4826 38792 5102
rect 38752 4820 38804 4826
rect 38752 4762 38804 4768
rect 38856 4758 38884 6598
rect 38948 6254 38976 6598
rect 38936 6248 38988 6254
rect 38936 6190 38988 6196
rect 39868 5846 39896 7142
rect 51078 6896 51134 6905
rect 40500 6860 40552 6866
rect 51078 6831 51134 6840
rect 40500 6802 40552 6808
rect 40040 6112 40092 6118
rect 40040 6054 40092 6060
rect 39856 5840 39908 5846
rect 39856 5782 39908 5788
rect 40052 5166 40080 6054
rect 40512 5914 40540 6802
rect 51092 6798 51120 6831
rect 51080 6792 51132 6798
rect 51080 6734 51132 6740
rect 45782 6556 46078 6576
rect 45838 6554 45862 6556
rect 45918 6554 45942 6556
rect 45998 6554 46022 6556
rect 45860 6502 45862 6554
rect 45924 6502 45936 6554
rect 45998 6502 46000 6554
rect 45838 6500 45862 6502
rect 45918 6500 45942 6502
rect 45998 6500 46022 6502
rect 45782 6480 46078 6500
rect 40500 5908 40552 5914
rect 40500 5850 40552 5856
rect 40592 5772 40644 5778
rect 40592 5714 40644 5720
rect 40040 5160 40092 5166
rect 40040 5102 40092 5108
rect 39396 5024 39448 5030
rect 39396 4966 39448 4972
rect 38844 4752 38896 4758
rect 38844 4694 38896 4700
rect 36176 4684 36228 4690
rect 36176 4626 36228 4632
rect 37556 4684 37608 4690
rect 37556 4626 37608 4632
rect 35624 4072 35676 4078
rect 35624 4014 35676 4020
rect 35072 3596 35124 3602
rect 35072 3538 35124 3544
rect 35084 3194 35112 3538
rect 35636 3194 35664 4014
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 36096 3602 36124 3878
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 35072 3188 35124 3194
rect 35072 3130 35124 3136
rect 35624 3188 35676 3194
rect 35624 3130 35676 3136
rect 36004 2990 36032 3334
rect 35992 2984 36044 2990
rect 35992 2926 36044 2932
rect 36188 2650 36216 4626
rect 36544 4480 36596 4486
rect 36544 4422 36596 4428
rect 36556 2990 36584 4422
rect 39408 4078 39436 4966
rect 40604 4826 40632 5714
rect 45782 5468 46078 5488
rect 45838 5466 45862 5468
rect 45918 5466 45942 5468
rect 45998 5466 46022 5468
rect 45860 5414 45862 5466
rect 45924 5414 45936 5466
rect 45998 5414 46000 5466
rect 45838 5412 45862 5414
rect 45918 5412 45942 5414
rect 45998 5412 46022 5414
rect 45782 5392 46078 5412
rect 40592 4820 40644 4826
rect 40592 4762 40644 4768
rect 40684 4684 40736 4690
rect 40684 4626 40736 4632
rect 40592 4480 40644 4486
rect 40592 4422 40644 4428
rect 40604 4078 40632 4422
rect 36728 4072 36780 4078
rect 36728 4014 36780 4020
rect 39396 4072 39448 4078
rect 39396 4014 39448 4020
rect 40408 4072 40460 4078
rect 40408 4014 40460 4020
rect 40592 4072 40644 4078
rect 40592 4014 40644 4020
rect 36636 3936 36688 3942
rect 36636 3878 36688 3884
rect 36648 3602 36676 3878
rect 36636 3596 36688 3602
rect 36636 3538 36688 3544
rect 36740 3194 36768 4014
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 40316 3936 40368 3942
rect 40316 3878 40368 3884
rect 36817 3836 37113 3856
rect 36873 3834 36897 3836
rect 36953 3834 36977 3836
rect 37033 3834 37057 3836
rect 36895 3782 36897 3834
rect 36959 3782 36971 3834
rect 37033 3782 37035 3834
rect 36873 3780 36897 3782
rect 36953 3780 36977 3782
rect 37033 3780 37057 3782
rect 36817 3760 37113 3780
rect 38396 3670 38424 3878
rect 38384 3664 38436 3670
rect 38384 3606 38436 3612
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 38672 3194 38700 3538
rect 39212 3392 39264 3398
rect 39212 3334 39264 3340
rect 40224 3392 40276 3398
rect 40224 3334 40276 3340
rect 36728 3188 36780 3194
rect 36728 3130 36780 3136
rect 38660 3188 38712 3194
rect 38660 3130 38712 3136
rect 36544 2984 36596 2990
rect 36544 2926 36596 2932
rect 37832 2984 37884 2990
rect 37832 2926 37884 2932
rect 38844 2984 38896 2990
rect 38844 2926 38896 2932
rect 37280 2848 37332 2854
rect 37280 2790 37332 2796
rect 36817 2748 37113 2768
rect 36873 2746 36897 2748
rect 36953 2746 36977 2748
rect 37033 2746 37057 2748
rect 36895 2694 36897 2746
rect 36959 2694 36971 2746
rect 37033 2694 37035 2746
rect 36873 2692 36897 2694
rect 36953 2692 36977 2694
rect 37033 2692 37057 2694
rect 36817 2672 37113 2692
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 37292 2514 37320 2790
rect 37844 2650 37872 2926
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 38672 2514 38700 2790
rect 38856 2650 38884 2926
rect 38844 2644 38896 2650
rect 38844 2586 38896 2592
rect 39224 2514 39252 3334
rect 40040 2984 40092 2990
rect 40040 2926 40092 2932
rect 40052 2650 40080 2926
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40236 2514 40264 3334
rect 40328 2990 40356 3878
rect 40316 2984 40368 2990
rect 40316 2926 40368 2932
rect 30656 2508 30708 2514
rect 30656 2450 30708 2456
rect 31668 2508 31720 2514
rect 31668 2450 31720 2456
rect 33508 2508 33560 2514
rect 33508 2450 33560 2456
rect 34520 2508 34572 2514
rect 34520 2450 34572 2456
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 38660 2508 38712 2514
rect 38660 2450 38712 2456
rect 39212 2508 39264 2514
rect 39212 2450 39264 2456
rect 40224 2508 40276 2514
rect 40224 2450 40276 2456
rect 40420 2378 40448 4014
rect 40696 3738 40724 4626
rect 45782 4380 46078 4400
rect 45838 4378 45862 4380
rect 45918 4378 45942 4380
rect 45998 4378 46022 4380
rect 45860 4326 45862 4378
rect 45924 4326 45936 4378
rect 45998 4326 46000 4378
rect 45838 4324 45862 4326
rect 45918 4324 45942 4326
rect 45998 4324 46022 4326
rect 45782 4304 46078 4324
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 40684 3732 40736 3738
rect 40684 3674 40736 3680
rect 40592 3596 40644 3602
rect 40592 3538 40644 3544
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 42248 3596 42300 3602
rect 42248 3538 42300 3544
rect 40604 2650 40632 3538
rect 41248 3194 41276 3538
rect 41420 3392 41472 3398
rect 41420 3334 41472 3340
rect 41236 3188 41288 3194
rect 41236 3130 41288 3136
rect 40592 2644 40644 2650
rect 40592 2586 40644 2592
rect 41432 2514 41460 3334
rect 42260 3194 42288 3538
rect 42248 3188 42300 3194
rect 42248 3130 42300 3136
rect 42444 2990 42472 3878
rect 43076 3460 43128 3466
rect 43076 3402 43128 3408
rect 42432 2984 42484 2990
rect 42432 2926 42484 2932
rect 43088 2514 43116 3402
rect 45782 3292 46078 3312
rect 45838 3290 45862 3292
rect 45918 3290 45942 3292
rect 45998 3290 46022 3292
rect 45860 3238 45862 3290
rect 45924 3238 45936 3290
rect 45998 3238 46000 3290
rect 45838 3236 45862 3238
rect 45918 3236 45942 3238
rect 45998 3236 46022 3238
rect 45782 3216 46078 3236
rect 41420 2508 41472 2514
rect 41420 2450 41472 2456
rect 43076 2508 43128 2514
rect 43076 2450 43128 2456
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 40408 2372 40460 2378
rect 40408 2314 40460 2320
rect 45782 2204 46078 2224
rect 45838 2202 45862 2204
rect 45918 2202 45942 2204
rect 45998 2202 46022 2204
rect 45860 2150 45862 2202
rect 45924 2150 45936 2202
rect 45998 2150 46000 2202
rect 45838 2148 45862 2150
rect 45918 2148 45942 2150
rect 45998 2148 46022 2150
rect 45782 2128 46078 2148
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 29184 2100 29236 2106
rect 29184 2042 29236 2048
<< via2 >>
rect 2502 21936 2558 21992
rect 7286 21956 7342 21992
rect 7286 21936 7288 21956
rect 7288 21936 7340 21956
rect 7340 21936 7342 21956
rect 9921 25050 9977 25052
rect 10001 25050 10057 25052
rect 10081 25050 10137 25052
rect 10161 25050 10217 25052
rect 9921 24998 9947 25050
rect 9947 24998 9977 25050
rect 10001 24998 10011 25050
rect 10011 24998 10057 25050
rect 10081 24998 10127 25050
rect 10127 24998 10137 25050
rect 10161 24998 10191 25050
rect 10191 24998 10217 25050
rect 9921 24996 9977 24998
rect 10001 24996 10057 24998
rect 10081 24996 10137 24998
rect 10161 24996 10217 24998
rect 8298 19252 8300 19272
rect 8300 19252 8352 19272
rect 8352 19252 8354 19272
rect 8298 19216 8354 19252
rect 9921 23962 9977 23964
rect 10001 23962 10057 23964
rect 10081 23962 10137 23964
rect 10161 23962 10217 23964
rect 9921 23910 9947 23962
rect 9947 23910 9977 23962
rect 10001 23910 10011 23962
rect 10011 23910 10057 23962
rect 10081 23910 10127 23962
rect 10127 23910 10137 23962
rect 10161 23910 10191 23962
rect 10191 23910 10217 23962
rect 9921 23908 9977 23910
rect 10001 23908 10057 23910
rect 10081 23908 10137 23910
rect 10161 23908 10217 23910
rect 9921 22874 9977 22876
rect 10001 22874 10057 22876
rect 10081 22874 10137 22876
rect 10161 22874 10217 22876
rect 9921 22822 9947 22874
rect 9947 22822 9977 22874
rect 10001 22822 10011 22874
rect 10011 22822 10057 22874
rect 10081 22822 10127 22874
rect 10127 22822 10137 22874
rect 10161 22822 10191 22874
rect 10191 22822 10217 22874
rect 9921 22820 9977 22822
rect 10001 22820 10057 22822
rect 10081 22820 10137 22822
rect 10161 22820 10217 22822
rect 9494 19216 9550 19272
rect 9921 21786 9977 21788
rect 10001 21786 10057 21788
rect 10081 21786 10137 21788
rect 10161 21786 10217 21788
rect 9921 21734 9947 21786
rect 9947 21734 9977 21786
rect 10001 21734 10011 21786
rect 10011 21734 10057 21786
rect 10081 21734 10127 21786
rect 10127 21734 10137 21786
rect 10161 21734 10191 21786
rect 10191 21734 10217 21786
rect 9921 21732 9977 21734
rect 10001 21732 10057 21734
rect 10081 21732 10137 21734
rect 10161 21732 10217 21734
rect 9921 20698 9977 20700
rect 10001 20698 10057 20700
rect 10081 20698 10137 20700
rect 10161 20698 10217 20700
rect 9921 20646 9947 20698
rect 9947 20646 9977 20698
rect 10001 20646 10011 20698
rect 10011 20646 10057 20698
rect 10081 20646 10127 20698
rect 10127 20646 10137 20698
rect 10161 20646 10191 20698
rect 10191 20646 10217 20698
rect 9921 20644 9977 20646
rect 10001 20644 10057 20646
rect 10081 20644 10137 20646
rect 10161 20644 10217 20646
rect 9921 19610 9977 19612
rect 10001 19610 10057 19612
rect 10081 19610 10137 19612
rect 10161 19610 10217 19612
rect 9921 19558 9947 19610
rect 9947 19558 9977 19610
rect 10001 19558 10011 19610
rect 10011 19558 10057 19610
rect 10081 19558 10127 19610
rect 10127 19558 10137 19610
rect 10161 19558 10191 19610
rect 10191 19558 10217 19610
rect 9921 19556 9977 19558
rect 10001 19556 10057 19558
rect 10081 19556 10137 19558
rect 10161 19556 10217 19558
rect 9921 18522 9977 18524
rect 10001 18522 10057 18524
rect 10081 18522 10137 18524
rect 10161 18522 10217 18524
rect 9921 18470 9947 18522
rect 9947 18470 9977 18522
rect 10001 18470 10011 18522
rect 10011 18470 10057 18522
rect 10081 18470 10127 18522
rect 10127 18470 10137 18522
rect 10161 18470 10191 18522
rect 10191 18470 10217 18522
rect 9921 18468 9977 18470
rect 10001 18468 10057 18470
rect 10081 18468 10137 18470
rect 10161 18468 10217 18470
rect 9921 17434 9977 17436
rect 10001 17434 10057 17436
rect 10081 17434 10137 17436
rect 10161 17434 10217 17436
rect 9921 17382 9947 17434
rect 9947 17382 9977 17434
rect 10001 17382 10011 17434
rect 10011 17382 10057 17434
rect 10081 17382 10127 17434
rect 10127 17382 10137 17434
rect 10161 17382 10191 17434
rect 10191 17382 10217 17434
rect 9921 17380 9977 17382
rect 10001 17380 10057 17382
rect 10081 17380 10137 17382
rect 10161 17380 10217 17382
rect 12254 21548 12310 21584
rect 12254 21528 12256 21548
rect 12256 21528 12308 21548
rect 12308 21528 12310 21548
rect 9921 16346 9977 16348
rect 10001 16346 10057 16348
rect 10081 16346 10137 16348
rect 10161 16346 10217 16348
rect 9921 16294 9947 16346
rect 9947 16294 9977 16346
rect 10001 16294 10011 16346
rect 10011 16294 10057 16346
rect 10081 16294 10127 16346
rect 10127 16294 10137 16346
rect 10161 16294 10191 16346
rect 10191 16294 10217 16346
rect 9921 16292 9977 16294
rect 10001 16292 10057 16294
rect 10081 16292 10137 16294
rect 10161 16292 10217 16294
rect 9770 15408 9826 15464
rect 9921 15258 9977 15260
rect 10001 15258 10057 15260
rect 10081 15258 10137 15260
rect 10161 15258 10217 15260
rect 9921 15206 9947 15258
rect 9947 15206 9977 15258
rect 10001 15206 10011 15258
rect 10011 15206 10057 15258
rect 10081 15206 10127 15258
rect 10127 15206 10137 15258
rect 10161 15206 10191 15258
rect 10191 15206 10217 15258
rect 9921 15204 9977 15206
rect 10001 15204 10057 15206
rect 10081 15204 10137 15206
rect 10161 15204 10217 15206
rect 10322 15000 10378 15056
rect 9921 14170 9977 14172
rect 10001 14170 10057 14172
rect 10081 14170 10137 14172
rect 10161 14170 10217 14172
rect 9921 14118 9947 14170
rect 9947 14118 9977 14170
rect 10001 14118 10011 14170
rect 10011 14118 10057 14170
rect 10081 14118 10127 14170
rect 10127 14118 10137 14170
rect 10161 14118 10191 14170
rect 10191 14118 10217 14170
rect 9921 14116 9977 14118
rect 10001 14116 10057 14118
rect 10081 14116 10137 14118
rect 10161 14116 10217 14118
rect 9921 13082 9977 13084
rect 10001 13082 10057 13084
rect 10081 13082 10137 13084
rect 10161 13082 10217 13084
rect 9921 13030 9947 13082
rect 9947 13030 9977 13082
rect 10001 13030 10011 13082
rect 10011 13030 10057 13082
rect 10081 13030 10127 13082
rect 10127 13030 10137 13082
rect 10161 13030 10191 13082
rect 10191 13030 10217 13082
rect 9921 13028 9977 13030
rect 10001 13028 10057 13030
rect 10081 13028 10137 13030
rect 10161 13028 10217 13030
rect 9921 11994 9977 11996
rect 10001 11994 10057 11996
rect 10081 11994 10137 11996
rect 10161 11994 10217 11996
rect 9921 11942 9947 11994
rect 9947 11942 9977 11994
rect 10001 11942 10011 11994
rect 10011 11942 10057 11994
rect 10081 11942 10127 11994
rect 10127 11942 10137 11994
rect 10161 11942 10191 11994
rect 10191 11942 10217 11994
rect 9921 11940 9977 11942
rect 10001 11940 10057 11942
rect 10081 11940 10137 11942
rect 10161 11940 10217 11942
rect 9921 10906 9977 10908
rect 10001 10906 10057 10908
rect 10081 10906 10137 10908
rect 10161 10906 10217 10908
rect 9921 10854 9947 10906
rect 9947 10854 9977 10906
rect 10001 10854 10011 10906
rect 10011 10854 10057 10906
rect 10081 10854 10127 10906
rect 10127 10854 10137 10906
rect 10161 10854 10191 10906
rect 10191 10854 10217 10906
rect 9921 10852 9977 10854
rect 10001 10852 10057 10854
rect 10081 10852 10137 10854
rect 10161 10852 10217 10854
rect 9921 9818 9977 9820
rect 10001 9818 10057 9820
rect 10081 9818 10137 9820
rect 10161 9818 10217 9820
rect 9921 9766 9947 9818
rect 9947 9766 9977 9818
rect 10001 9766 10011 9818
rect 10011 9766 10057 9818
rect 10081 9766 10127 9818
rect 10127 9766 10137 9818
rect 10161 9766 10191 9818
rect 10191 9766 10217 9818
rect 9921 9764 9977 9766
rect 10001 9764 10057 9766
rect 10081 9764 10137 9766
rect 10161 9764 10217 9766
rect 12714 21548 12770 21584
rect 12714 21528 12716 21548
rect 12716 21528 12768 21548
rect 12768 21528 12770 21548
rect 12530 15408 12586 15464
rect 13082 15000 13138 15056
rect 9921 8730 9977 8732
rect 10001 8730 10057 8732
rect 10081 8730 10137 8732
rect 10161 8730 10217 8732
rect 9921 8678 9947 8730
rect 9947 8678 9977 8730
rect 10001 8678 10011 8730
rect 10011 8678 10057 8730
rect 10081 8678 10127 8730
rect 10127 8678 10137 8730
rect 10161 8678 10191 8730
rect 10191 8678 10217 8730
rect 9921 8676 9977 8678
rect 10001 8676 10057 8678
rect 10081 8676 10137 8678
rect 10161 8676 10217 8678
rect 9921 7642 9977 7644
rect 10001 7642 10057 7644
rect 10081 7642 10137 7644
rect 10161 7642 10217 7644
rect 9921 7590 9947 7642
rect 9947 7590 9977 7642
rect 10001 7590 10011 7642
rect 10011 7590 10057 7642
rect 10081 7590 10127 7642
rect 10127 7590 10137 7642
rect 10161 7590 10191 7642
rect 10191 7590 10217 7642
rect 9921 7588 9977 7590
rect 10001 7588 10057 7590
rect 10081 7588 10137 7590
rect 10161 7588 10217 7590
rect 9921 6554 9977 6556
rect 10001 6554 10057 6556
rect 10081 6554 10137 6556
rect 10161 6554 10217 6556
rect 9921 6502 9947 6554
rect 9947 6502 9977 6554
rect 10001 6502 10011 6554
rect 10011 6502 10057 6554
rect 10081 6502 10127 6554
rect 10127 6502 10137 6554
rect 10161 6502 10191 6554
rect 10191 6502 10217 6554
rect 9921 6500 9977 6502
rect 10001 6500 10057 6502
rect 10081 6500 10137 6502
rect 10161 6500 10217 6502
rect 11242 8900 11298 8936
rect 11242 8880 11244 8900
rect 11244 8880 11296 8900
rect 11296 8880 11298 8900
rect 9921 5466 9977 5468
rect 10001 5466 10057 5468
rect 10081 5466 10137 5468
rect 10161 5466 10217 5468
rect 9921 5414 9947 5466
rect 9947 5414 9977 5466
rect 10001 5414 10011 5466
rect 10011 5414 10057 5466
rect 10081 5414 10127 5466
rect 10127 5414 10137 5466
rect 10161 5414 10191 5466
rect 10191 5414 10217 5466
rect 9921 5412 9977 5414
rect 10001 5412 10057 5414
rect 10081 5412 10137 5414
rect 10161 5412 10217 5414
rect 9921 4378 9977 4380
rect 10001 4378 10057 4380
rect 10081 4378 10137 4380
rect 10161 4378 10217 4380
rect 9921 4326 9947 4378
rect 9947 4326 9977 4378
rect 10001 4326 10011 4378
rect 10011 4326 10057 4378
rect 10081 4326 10127 4378
rect 10127 4326 10137 4378
rect 10161 4326 10191 4378
rect 10191 4326 10217 4378
rect 9921 4324 9977 4326
rect 10001 4324 10057 4326
rect 10081 4324 10137 4326
rect 10161 4324 10217 4326
rect 15382 15000 15438 15056
rect 18886 24506 18942 24508
rect 18966 24506 19022 24508
rect 19046 24506 19102 24508
rect 19126 24506 19182 24508
rect 18886 24454 18912 24506
rect 18912 24454 18942 24506
rect 18966 24454 18976 24506
rect 18976 24454 19022 24506
rect 19046 24454 19092 24506
rect 19092 24454 19102 24506
rect 19126 24454 19156 24506
rect 19156 24454 19182 24506
rect 18886 24452 18942 24454
rect 18966 24452 19022 24454
rect 19046 24452 19102 24454
rect 19126 24452 19182 24454
rect 18886 23418 18942 23420
rect 18966 23418 19022 23420
rect 19046 23418 19102 23420
rect 19126 23418 19182 23420
rect 18886 23366 18912 23418
rect 18912 23366 18942 23418
rect 18966 23366 18976 23418
rect 18976 23366 19022 23418
rect 19046 23366 19092 23418
rect 19092 23366 19102 23418
rect 19126 23366 19156 23418
rect 19156 23366 19182 23418
rect 18886 23364 18942 23366
rect 18966 23364 19022 23366
rect 19046 23364 19102 23366
rect 19126 23364 19182 23366
rect 18886 22330 18942 22332
rect 18966 22330 19022 22332
rect 19046 22330 19102 22332
rect 19126 22330 19182 22332
rect 18886 22278 18912 22330
rect 18912 22278 18942 22330
rect 18966 22278 18976 22330
rect 18976 22278 19022 22330
rect 19046 22278 19092 22330
rect 19092 22278 19102 22330
rect 19126 22278 19156 22330
rect 19156 22278 19182 22330
rect 18886 22276 18942 22278
rect 18966 22276 19022 22278
rect 19046 22276 19102 22278
rect 19126 22276 19182 22278
rect 18886 21242 18942 21244
rect 18966 21242 19022 21244
rect 19046 21242 19102 21244
rect 19126 21242 19182 21244
rect 18886 21190 18912 21242
rect 18912 21190 18942 21242
rect 18966 21190 18976 21242
rect 18976 21190 19022 21242
rect 19046 21190 19092 21242
rect 19092 21190 19102 21242
rect 19126 21190 19156 21242
rect 19156 21190 19182 21242
rect 18886 21188 18942 21190
rect 18966 21188 19022 21190
rect 19046 21188 19102 21190
rect 19126 21188 19182 21190
rect 18886 20154 18942 20156
rect 18966 20154 19022 20156
rect 19046 20154 19102 20156
rect 19126 20154 19182 20156
rect 18886 20102 18912 20154
rect 18912 20102 18942 20154
rect 18966 20102 18976 20154
rect 18976 20102 19022 20154
rect 19046 20102 19092 20154
rect 19092 20102 19102 20154
rect 19126 20102 19156 20154
rect 19156 20102 19182 20154
rect 18886 20100 18942 20102
rect 18966 20100 19022 20102
rect 19046 20100 19102 20102
rect 19126 20100 19182 20102
rect 18886 19066 18942 19068
rect 18966 19066 19022 19068
rect 19046 19066 19102 19068
rect 19126 19066 19182 19068
rect 18886 19014 18912 19066
rect 18912 19014 18942 19066
rect 18966 19014 18976 19066
rect 18976 19014 19022 19066
rect 19046 19014 19092 19066
rect 19092 19014 19102 19066
rect 19126 19014 19156 19066
rect 19156 19014 19182 19066
rect 18886 19012 18942 19014
rect 18966 19012 19022 19014
rect 19046 19012 19102 19014
rect 19126 19012 19182 19014
rect 18886 17978 18942 17980
rect 18966 17978 19022 17980
rect 19046 17978 19102 17980
rect 19126 17978 19182 17980
rect 18886 17926 18912 17978
rect 18912 17926 18942 17978
rect 18966 17926 18976 17978
rect 18976 17926 19022 17978
rect 19046 17926 19092 17978
rect 19092 17926 19102 17978
rect 19126 17926 19156 17978
rect 19156 17926 19182 17978
rect 18886 17924 18942 17926
rect 18966 17924 19022 17926
rect 19046 17924 19102 17926
rect 19126 17924 19182 17926
rect 22006 19372 22062 19408
rect 22006 19352 22008 19372
rect 22008 19352 22060 19372
rect 22060 19352 22062 19372
rect 24030 22516 24032 22536
rect 24032 22516 24084 22536
rect 24084 22516 24086 22536
rect 24030 22480 24086 22516
rect 24306 22516 24308 22536
rect 24308 22516 24360 22536
rect 24360 22516 24362 22536
rect 24306 22480 24362 22516
rect 24030 20476 24032 20496
rect 24032 20476 24084 20496
rect 24084 20476 24086 20496
rect 24030 20440 24086 20476
rect 18886 16890 18942 16892
rect 18966 16890 19022 16892
rect 19046 16890 19102 16892
rect 19126 16890 19182 16892
rect 18886 16838 18912 16890
rect 18912 16838 18942 16890
rect 18966 16838 18976 16890
rect 18976 16838 19022 16890
rect 19046 16838 19092 16890
rect 19092 16838 19102 16890
rect 19126 16838 19156 16890
rect 19156 16838 19182 16890
rect 18886 16836 18942 16838
rect 18966 16836 19022 16838
rect 19046 16836 19102 16838
rect 19126 16836 19182 16838
rect 17038 8900 17094 8936
rect 17038 8880 17040 8900
rect 17040 8880 17092 8900
rect 17092 8880 17094 8900
rect 18886 15802 18942 15804
rect 18966 15802 19022 15804
rect 19046 15802 19102 15804
rect 19126 15802 19182 15804
rect 18886 15750 18912 15802
rect 18912 15750 18942 15802
rect 18966 15750 18976 15802
rect 18976 15750 19022 15802
rect 19046 15750 19092 15802
rect 19092 15750 19102 15802
rect 19126 15750 19156 15802
rect 19156 15750 19182 15802
rect 18886 15748 18942 15750
rect 18966 15748 19022 15750
rect 19046 15748 19102 15750
rect 19126 15748 19182 15750
rect 19522 15952 19578 16008
rect 18886 14714 18942 14716
rect 18966 14714 19022 14716
rect 19046 14714 19102 14716
rect 19126 14714 19182 14716
rect 18886 14662 18912 14714
rect 18912 14662 18942 14714
rect 18966 14662 18976 14714
rect 18976 14662 19022 14714
rect 19046 14662 19092 14714
rect 19092 14662 19102 14714
rect 19126 14662 19156 14714
rect 19156 14662 19182 14714
rect 18886 14660 18942 14662
rect 18966 14660 19022 14662
rect 19046 14660 19102 14662
rect 19126 14660 19182 14662
rect 18886 13626 18942 13628
rect 18966 13626 19022 13628
rect 19046 13626 19102 13628
rect 19126 13626 19182 13628
rect 18886 13574 18912 13626
rect 18912 13574 18942 13626
rect 18966 13574 18976 13626
rect 18976 13574 19022 13626
rect 19046 13574 19092 13626
rect 19092 13574 19102 13626
rect 19126 13574 19156 13626
rect 19156 13574 19182 13626
rect 18886 13572 18942 13574
rect 18966 13572 19022 13574
rect 19046 13572 19102 13574
rect 19126 13572 19182 13574
rect 18886 12538 18942 12540
rect 18966 12538 19022 12540
rect 19046 12538 19102 12540
rect 19126 12538 19182 12540
rect 18886 12486 18912 12538
rect 18912 12486 18942 12538
rect 18966 12486 18976 12538
rect 18976 12486 19022 12538
rect 19046 12486 19092 12538
rect 19092 12486 19102 12538
rect 19126 12486 19156 12538
rect 19156 12486 19182 12538
rect 18886 12484 18942 12486
rect 18966 12484 19022 12486
rect 19046 12484 19102 12486
rect 19126 12484 19182 12486
rect 22098 15988 22100 16008
rect 22100 15988 22152 16008
rect 22152 15988 22154 16008
rect 22098 15952 22154 15988
rect 27852 25050 27908 25052
rect 27932 25050 27988 25052
rect 28012 25050 28068 25052
rect 28092 25050 28148 25052
rect 27852 24998 27878 25050
rect 27878 24998 27908 25050
rect 27932 24998 27942 25050
rect 27942 24998 27988 25050
rect 28012 24998 28058 25050
rect 28058 24998 28068 25050
rect 28092 24998 28122 25050
rect 28122 24998 28148 25050
rect 27852 24996 27908 24998
rect 27932 24996 27988 24998
rect 28012 24996 28068 24998
rect 28092 24996 28148 24998
rect 27852 23962 27908 23964
rect 27932 23962 27988 23964
rect 28012 23962 28068 23964
rect 28092 23962 28148 23964
rect 27852 23910 27878 23962
rect 27878 23910 27908 23962
rect 27932 23910 27942 23962
rect 27942 23910 27988 23962
rect 28012 23910 28058 23962
rect 28058 23910 28068 23962
rect 28092 23910 28122 23962
rect 28122 23910 28148 23962
rect 27852 23908 27908 23910
rect 27932 23908 27988 23910
rect 28012 23908 28068 23910
rect 28092 23908 28148 23910
rect 27852 22874 27908 22876
rect 27932 22874 27988 22876
rect 28012 22874 28068 22876
rect 28092 22874 28148 22876
rect 27852 22822 27878 22874
rect 27878 22822 27908 22874
rect 27932 22822 27942 22874
rect 27942 22822 27988 22874
rect 28012 22822 28058 22874
rect 28058 22822 28068 22874
rect 28092 22822 28122 22874
rect 28122 22822 28148 22874
rect 27852 22820 27908 22822
rect 27932 22820 27988 22822
rect 28012 22820 28068 22822
rect 28092 22820 28148 22822
rect 28262 22500 28318 22536
rect 28262 22480 28264 22500
rect 28264 22480 28316 22500
rect 28316 22480 28318 22500
rect 27852 21786 27908 21788
rect 27932 21786 27988 21788
rect 28012 21786 28068 21788
rect 28092 21786 28148 21788
rect 27852 21734 27878 21786
rect 27878 21734 27908 21786
rect 27932 21734 27942 21786
rect 27942 21734 27988 21786
rect 28012 21734 28058 21786
rect 28058 21734 28068 21786
rect 28092 21734 28122 21786
rect 28122 21734 28148 21786
rect 27852 21732 27908 21734
rect 27932 21732 27988 21734
rect 28012 21732 28068 21734
rect 28092 21732 28148 21734
rect 28354 21392 28410 21448
rect 25778 17756 25780 17776
rect 25780 17756 25832 17776
rect 25832 17756 25834 17776
rect 25778 17720 25834 17756
rect 24398 16496 24454 16552
rect 25962 16496 26018 16552
rect 26882 21004 26938 21040
rect 26882 20984 26884 21004
rect 26884 20984 26936 21004
rect 26936 20984 26938 21004
rect 28722 21020 28724 21040
rect 28724 21020 28776 21040
rect 28776 21020 28778 21040
rect 28722 20984 28778 21020
rect 27852 20698 27908 20700
rect 27932 20698 27988 20700
rect 28012 20698 28068 20700
rect 28092 20698 28148 20700
rect 27852 20646 27878 20698
rect 27878 20646 27908 20698
rect 27932 20646 27942 20698
rect 27942 20646 27988 20698
rect 28012 20646 28058 20698
rect 28058 20646 28068 20698
rect 28092 20646 28122 20698
rect 28122 20646 28148 20698
rect 27852 20644 27908 20646
rect 27932 20644 27988 20646
rect 28012 20644 28068 20646
rect 28092 20644 28148 20646
rect 26974 20440 27030 20496
rect 27852 19610 27908 19612
rect 27932 19610 27988 19612
rect 28012 19610 28068 19612
rect 28092 19610 28148 19612
rect 27852 19558 27878 19610
rect 27878 19558 27908 19610
rect 27932 19558 27942 19610
rect 27942 19558 27988 19610
rect 28012 19558 28058 19610
rect 28058 19558 28068 19610
rect 28092 19558 28122 19610
rect 28122 19558 28148 19610
rect 27852 19556 27908 19558
rect 27932 19556 27988 19558
rect 28012 19556 28068 19558
rect 28092 19556 28148 19558
rect 27802 19388 27804 19408
rect 27804 19388 27856 19408
rect 27856 19388 27858 19408
rect 27802 19352 27858 19388
rect 18886 11450 18942 11452
rect 18966 11450 19022 11452
rect 19046 11450 19102 11452
rect 19126 11450 19182 11452
rect 18886 11398 18912 11450
rect 18912 11398 18942 11450
rect 18966 11398 18976 11450
rect 18976 11398 19022 11450
rect 19046 11398 19092 11450
rect 19092 11398 19102 11450
rect 19126 11398 19156 11450
rect 19156 11398 19182 11450
rect 18886 11396 18942 11398
rect 18966 11396 19022 11398
rect 19046 11396 19102 11398
rect 19126 11396 19182 11398
rect 18886 10362 18942 10364
rect 18966 10362 19022 10364
rect 19046 10362 19102 10364
rect 19126 10362 19182 10364
rect 18886 10310 18912 10362
rect 18912 10310 18942 10362
rect 18966 10310 18976 10362
rect 18976 10310 19022 10362
rect 19046 10310 19092 10362
rect 19092 10310 19102 10362
rect 19126 10310 19156 10362
rect 19156 10310 19182 10362
rect 18886 10308 18942 10310
rect 18966 10308 19022 10310
rect 19046 10308 19102 10310
rect 19126 10308 19182 10310
rect 18886 9274 18942 9276
rect 18966 9274 19022 9276
rect 19046 9274 19102 9276
rect 19126 9274 19182 9276
rect 18886 9222 18912 9274
rect 18912 9222 18942 9274
rect 18966 9222 18976 9274
rect 18976 9222 19022 9274
rect 19046 9222 19092 9274
rect 19092 9222 19102 9274
rect 19126 9222 19156 9274
rect 19156 9222 19182 9274
rect 18886 9220 18942 9222
rect 18966 9220 19022 9222
rect 19046 9220 19102 9222
rect 19126 9220 19182 9222
rect 18886 8186 18942 8188
rect 18966 8186 19022 8188
rect 19046 8186 19102 8188
rect 19126 8186 19182 8188
rect 18886 8134 18912 8186
rect 18912 8134 18942 8186
rect 18966 8134 18976 8186
rect 18976 8134 19022 8186
rect 19046 8134 19092 8186
rect 19092 8134 19102 8186
rect 19126 8134 19156 8186
rect 19156 8134 19182 8186
rect 18886 8132 18942 8134
rect 18966 8132 19022 8134
rect 19046 8132 19102 8134
rect 19126 8132 19182 8134
rect 18886 7098 18942 7100
rect 18966 7098 19022 7100
rect 19046 7098 19102 7100
rect 19126 7098 19182 7100
rect 18886 7046 18912 7098
rect 18912 7046 18942 7098
rect 18966 7046 18976 7098
rect 18976 7046 19022 7098
rect 19046 7046 19092 7098
rect 19092 7046 19102 7098
rect 19126 7046 19156 7098
rect 19156 7046 19182 7098
rect 18886 7044 18942 7046
rect 18966 7044 19022 7046
rect 19046 7044 19102 7046
rect 19126 7044 19182 7046
rect 18886 6010 18942 6012
rect 18966 6010 19022 6012
rect 19046 6010 19102 6012
rect 19126 6010 19182 6012
rect 18886 5958 18912 6010
rect 18912 5958 18942 6010
rect 18966 5958 18976 6010
rect 18976 5958 19022 6010
rect 19046 5958 19092 6010
rect 19092 5958 19102 6010
rect 19126 5958 19156 6010
rect 19156 5958 19182 6010
rect 18886 5956 18942 5958
rect 18966 5956 19022 5958
rect 19046 5956 19102 5958
rect 19126 5956 19182 5958
rect 18886 4922 18942 4924
rect 18966 4922 19022 4924
rect 19046 4922 19102 4924
rect 19126 4922 19182 4924
rect 18886 4870 18912 4922
rect 18912 4870 18942 4922
rect 18966 4870 18976 4922
rect 18976 4870 19022 4922
rect 19046 4870 19092 4922
rect 19092 4870 19102 4922
rect 19126 4870 19156 4922
rect 19156 4870 19182 4922
rect 18886 4868 18942 4870
rect 18966 4868 19022 4870
rect 19046 4868 19102 4870
rect 19126 4868 19182 4870
rect 18886 3834 18942 3836
rect 18966 3834 19022 3836
rect 19046 3834 19102 3836
rect 19126 3834 19182 3836
rect 18886 3782 18912 3834
rect 18912 3782 18942 3834
rect 18966 3782 18976 3834
rect 18976 3782 19022 3834
rect 19046 3782 19092 3834
rect 19092 3782 19102 3834
rect 19126 3782 19156 3834
rect 19156 3782 19182 3834
rect 18886 3780 18942 3782
rect 18966 3780 19022 3782
rect 19046 3780 19102 3782
rect 19126 3780 19182 3782
rect 9921 3290 9977 3292
rect 10001 3290 10057 3292
rect 10081 3290 10137 3292
rect 10161 3290 10217 3292
rect 9921 3238 9947 3290
rect 9947 3238 9977 3290
rect 10001 3238 10011 3290
rect 10011 3238 10057 3290
rect 10081 3238 10127 3290
rect 10127 3238 10137 3290
rect 10161 3238 10191 3290
rect 10191 3238 10217 3290
rect 9921 3236 9977 3238
rect 10001 3236 10057 3238
rect 10081 3236 10137 3238
rect 10161 3236 10217 3238
rect 18886 2746 18942 2748
rect 18966 2746 19022 2748
rect 19046 2746 19102 2748
rect 19126 2746 19182 2748
rect 18886 2694 18912 2746
rect 18912 2694 18942 2746
rect 18966 2694 18976 2746
rect 18976 2694 19022 2746
rect 19046 2694 19092 2746
rect 19092 2694 19102 2746
rect 19126 2694 19156 2746
rect 19156 2694 19182 2746
rect 18886 2692 18942 2694
rect 18966 2692 19022 2694
rect 19046 2692 19102 2694
rect 19126 2692 19182 2694
rect 27852 18522 27908 18524
rect 27932 18522 27988 18524
rect 28012 18522 28068 18524
rect 28092 18522 28148 18524
rect 27852 18470 27878 18522
rect 27878 18470 27908 18522
rect 27932 18470 27942 18522
rect 27942 18470 27988 18522
rect 28012 18470 28058 18522
rect 28058 18470 28068 18522
rect 28092 18470 28122 18522
rect 28122 18470 28148 18522
rect 27852 18468 27908 18470
rect 27932 18468 27988 18470
rect 28012 18468 28068 18470
rect 28092 18468 28148 18470
rect 27852 17434 27908 17436
rect 27932 17434 27988 17436
rect 28012 17434 28068 17436
rect 28092 17434 28148 17436
rect 27852 17382 27878 17434
rect 27878 17382 27908 17434
rect 27932 17382 27942 17434
rect 27942 17382 27988 17434
rect 28012 17382 28058 17434
rect 28058 17382 28068 17434
rect 28092 17382 28122 17434
rect 28122 17382 28148 17434
rect 27852 17380 27908 17382
rect 27932 17380 27988 17382
rect 28012 17380 28068 17382
rect 28092 17380 28148 17382
rect 28906 21412 28962 21448
rect 28906 21392 28908 21412
rect 28908 21392 28960 21412
rect 28960 21392 28962 21412
rect 32494 23024 32550 23080
rect 29366 18672 29422 18728
rect 30010 18400 30066 18456
rect 28630 17484 28632 17504
rect 28632 17484 28684 17504
rect 28684 17484 28686 17504
rect 28630 17448 28686 17484
rect 28906 17484 28908 17504
rect 28908 17484 28960 17504
rect 28960 17484 28962 17504
rect 28906 17448 28962 17484
rect 27852 16346 27908 16348
rect 27932 16346 27988 16348
rect 28012 16346 28068 16348
rect 28092 16346 28148 16348
rect 27852 16294 27878 16346
rect 27878 16294 27908 16346
rect 27932 16294 27942 16346
rect 27942 16294 27988 16346
rect 28012 16294 28058 16346
rect 28058 16294 28068 16346
rect 28092 16294 28122 16346
rect 28122 16294 28148 16346
rect 27852 16292 27908 16294
rect 27932 16292 27988 16294
rect 28012 16292 28068 16294
rect 28092 16292 28148 16294
rect 29826 17332 29882 17368
rect 29826 17312 29828 17332
rect 29828 17312 29880 17332
rect 29880 17312 29882 17332
rect 31758 18536 31814 18592
rect 36817 24506 36873 24508
rect 36897 24506 36953 24508
rect 36977 24506 37033 24508
rect 37057 24506 37113 24508
rect 36817 24454 36843 24506
rect 36843 24454 36873 24506
rect 36897 24454 36907 24506
rect 36907 24454 36953 24506
rect 36977 24454 37023 24506
rect 37023 24454 37033 24506
rect 37057 24454 37087 24506
rect 37087 24454 37113 24506
rect 36817 24452 36873 24454
rect 36897 24452 36953 24454
rect 36977 24452 37033 24454
rect 37057 24452 37113 24454
rect 36817 23418 36873 23420
rect 36897 23418 36953 23420
rect 36977 23418 37033 23420
rect 37057 23418 37113 23420
rect 36817 23366 36843 23418
rect 36843 23366 36873 23418
rect 36897 23366 36907 23418
rect 36907 23366 36953 23418
rect 36977 23366 37023 23418
rect 37023 23366 37033 23418
rect 37057 23366 37087 23418
rect 37087 23366 37113 23418
rect 36817 23364 36873 23366
rect 36897 23364 36953 23366
rect 36977 23364 37033 23366
rect 37057 23364 37113 23366
rect 36817 22330 36873 22332
rect 36897 22330 36953 22332
rect 36977 22330 37033 22332
rect 37057 22330 37113 22332
rect 36817 22278 36843 22330
rect 36843 22278 36873 22330
rect 36897 22278 36907 22330
rect 36907 22278 36953 22330
rect 36977 22278 37023 22330
rect 37023 22278 37033 22330
rect 37057 22278 37087 22330
rect 37087 22278 37113 22330
rect 36817 22276 36873 22278
rect 36897 22276 36953 22278
rect 36977 22276 37033 22278
rect 37057 22276 37113 22278
rect 36817 21242 36873 21244
rect 36897 21242 36953 21244
rect 36977 21242 37033 21244
rect 37057 21242 37113 21244
rect 36817 21190 36843 21242
rect 36843 21190 36873 21242
rect 36897 21190 36907 21242
rect 36907 21190 36953 21242
rect 36977 21190 37023 21242
rect 37023 21190 37033 21242
rect 37057 21190 37087 21242
rect 37087 21190 37113 21242
rect 36817 21188 36873 21190
rect 36897 21188 36953 21190
rect 36977 21188 37033 21190
rect 37057 21188 37113 21190
rect 32402 18828 32458 18864
rect 32402 18808 32404 18828
rect 32404 18808 32456 18828
rect 32456 18808 32458 18828
rect 32310 18536 32366 18592
rect 30470 16652 30526 16688
rect 30470 16632 30472 16652
rect 30472 16632 30524 16652
rect 30524 16632 30526 16652
rect 27852 15258 27908 15260
rect 27932 15258 27988 15260
rect 28012 15258 28068 15260
rect 28092 15258 28148 15260
rect 27852 15206 27878 15258
rect 27878 15206 27908 15258
rect 27932 15206 27942 15258
rect 27942 15206 27988 15258
rect 28012 15206 28058 15258
rect 28058 15206 28068 15258
rect 28092 15206 28122 15258
rect 28122 15206 28148 15258
rect 27852 15204 27908 15206
rect 27932 15204 27988 15206
rect 28012 15204 28068 15206
rect 28092 15204 28148 15206
rect 27852 14170 27908 14172
rect 27932 14170 27988 14172
rect 28012 14170 28068 14172
rect 28092 14170 28148 14172
rect 27852 14118 27878 14170
rect 27878 14118 27908 14170
rect 27932 14118 27942 14170
rect 27942 14118 27988 14170
rect 28012 14118 28058 14170
rect 28058 14118 28068 14170
rect 28092 14118 28122 14170
rect 28122 14118 28148 14170
rect 27852 14116 27908 14118
rect 27932 14116 27988 14118
rect 28012 14116 28068 14118
rect 28092 14116 28148 14118
rect 27852 13082 27908 13084
rect 27932 13082 27988 13084
rect 28012 13082 28068 13084
rect 28092 13082 28148 13084
rect 27852 13030 27878 13082
rect 27878 13030 27908 13082
rect 27932 13030 27942 13082
rect 27942 13030 27988 13082
rect 28012 13030 28058 13082
rect 28058 13030 28068 13082
rect 28092 13030 28122 13082
rect 28122 13030 28148 13082
rect 27852 13028 27908 13030
rect 27932 13028 27988 13030
rect 28012 13028 28068 13030
rect 28092 13028 28148 13030
rect 27852 11994 27908 11996
rect 27932 11994 27988 11996
rect 28012 11994 28068 11996
rect 28092 11994 28148 11996
rect 27852 11942 27878 11994
rect 27878 11942 27908 11994
rect 27932 11942 27942 11994
rect 27942 11942 27988 11994
rect 28012 11942 28058 11994
rect 28058 11942 28068 11994
rect 28092 11942 28122 11994
rect 28122 11942 28148 11994
rect 27852 11940 27908 11942
rect 27932 11940 27988 11942
rect 28012 11940 28068 11942
rect 28092 11940 28148 11942
rect 27852 10906 27908 10908
rect 27932 10906 27988 10908
rect 28012 10906 28068 10908
rect 28092 10906 28148 10908
rect 27852 10854 27878 10906
rect 27878 10854 27908 10906
rect 27932 10854 27942 10906
rect 27942 10854 27988 10906
rect 28012 10854 28058 10906
rect 28058 10854 28068 10906
rect 28092 10854 28122 10906
rect 28122 10854 28148 10906
rect 27852 10852 27908 10854
rect 27932 10852 27988 10854
rect 28012 10852 28068 10854
rect 28092 10852 28148 10854
rect 32954 18536 33010 18592
rect 33690 18808 33746 18864
rect 33874 18572 33876 18592
rect 33876 18572 33928 18592
rect 33928 18572 33930 18592
rect 33874 18536 33930 18572
rect 35622 18400 35678 18456
rect 34518 17584 34574 17640
rect 36817 20154 36873 20156
rect 36897 20154 36953 20156
rect 36977 20154 37033 20156
rect 37057 20154 37113 20156
rect 36817 20102 36843 20154
rect 36843 20102 36873 20154
rect 36897 20102 36907 20154
rect 36907 20102 36953 20154
rect 36977 20102 37023 20154
rect 37023 20102 37033 20154
rect 37057 20102 37087 20154
rect 37087 20102 37113 20154
rect 36817 20100 36873 20102
rect 36897 20100 36953 20102
rect 36977 20100 37033 20102
rect 37057 20100 37113 20102
rect 36817 19066 36873 19068
rect 36897 19066 36953 19068
rect 36977 19066 37033 19068
rect 37057 19066 37113 19068
rect 36817 19014 36843 19066
rect 36843 19014 36873 19066
rect 36897 19014 36907 19066
rect 36907 19014 36953 19066
rect 36977 19014 37023 19066
rect 37023 19014 37033 19066
rect 37057 19014 37087 19066
rect 37087 19014 37113 19066
rect 36817 19012 36873 19014
rect 36897 19012 36953 19014
rect 36977 19012 37033 19014
rect 37057 19012 37113 19014
rect 36726 18828 36782 18864
rect 36726 18808 36728 18828
rect 36728 18808 36780 18828
rect 36780 18808 36782 18828
rect 36817 17978 36873 17980
rect 36897 17978 36953 17980
rect 36977 17978 37033 17980
rect 37057 17978 37113 17980
rect 36817 17926 36843 17978
rect 36843 17926 36873 17978
rect 36897 17926 36907 17978
rect 36907 17926 36953 17978
rect 36977 17926 37023 17978
rect 37023 17926 37033 17978
rect 37057 17926 37087 17978
rect 37087 17926 37113 17978
rect 36817 17924 36873 17926
rect 36897 17924 36953 17926
rect 36977 17924 37033 17926
rect 37057 17924 37113 17926
rect 38566 23024 38622 23080
rect 36082 17312 36138 17368
rect 36450 17312 36506 17368
rect 37922 17584 37978 17640
rect 38290 18692 38346 18728
rect 38290 18672 38292 18692
rect 38292 18672 38344 18692
rect 38344 18672 38346 18692
rect 36817 16890 36873 16892
rect 36897 16890 36953 16892
rect 36977 16890 37033 16892
rect 37057 16890 37113 16892
rect 36817 16838 36843 16890
rect 36843 16838 36873 16890
rect 36897 16838 36907 16890
rect 36907 16838 36953 16890
rect 36977 16838 37023 16890
rect 37023 16838 37033 16890
rect 37057 16838 37087 16890
rect 37087 16838 37113 16890
rect 36817 16836 36873 16838
rect 36897 16836 36953 16838
rect 36977 16836 37033 16838
rect 37057 16836 37113 16838
rect 37186 16632 37242 16688
rect 36817 15802 36873 15804
rect 36897 15802 36953 15804
rect 36977 15802 37033 15804
rect 37057 15802 37113 15804
rect 36817 15750 36843 15802
rect 36843 15750 36873 15802
rect 36897 15750 36907 15802
rect 36907 15750 36953 15802
rect 36977 15750 37023 15802
rect 37023 15750 37033 15802
rect 37057 15750 37087 15802
rect 37087 15750 37113 15802
rect 36817 15748 36873 15750
rect 36897 15748 36953 15750
rect 36977 15748 37033 15750
rect 37057 15748 37113 15750
rect 36817 14714 36873 14716
rect 36897 14714 36953 14716
rect 36977 14714 37033 14716
rect 37057 14714 37113 14716
rect 36817 14662 36843 14714
rect 36843 14662 36873 14714
rect 36897 14662 36907 14714
rect 36907 14662 36953 14714
rect 36977 14662 37023 14714
rect 37023 14662 37033 14714
rect 37057 14662 37087 14714
rect 37087 14662 37113 14714
rect 36817 14660 36873 14662
rect 36897 14660 36953 14662
rect 36977 14660 37033 14662
rect 37057 14660 37113 14662
rect 36817 13626 36873 13628
rect 36897 13626 36953 13628
rect 36977 13626 37033 13628
rect 37057 13626 37113 13628
rect 36817 13574 36843 13626
rect 36843 13574 36873 13626
rect 36897 13574 36907 13626
rect 36907 13574 36953 13626
rect 36977 13574 37023 13626
rect 37023 13574 37033 13626
rect 37057 13574 37087 13626
rect 37087 13574 37113 13626
rect 36817 13572 36873 13574
rect 36897 13572 36953 13574
rect 36977 13572 37033 13574
rect 37057 13572 37113 13574
rect 39026 19080 39082 19136
rect 38934 18672 38990 18728
rect 39578 19760 39634 19816
rect 39946 18536 40002 18592
rect 41602 19236 41658 19272
rect 41602 19216 41604 19236
rect 41604 19216 41656 19236
rect 41656 19216 41658 19236
rect 41326 18808 41382 18864
rect 41602 18264 41658 18320
rect 41050 17720 41106 17776
rect 40038 17312 40094 17368
rect 39486 17076 39488 17096
rect 39488 17076 39540 17096
rect 39540 17076 39542 17096
rect 39486 17040 39542 17076
rect 40866 17312 40922 17368
rect 42154 22228 42210 22264
rect 42154 22208 42156 22228
rect 42156 22208 42208 22228
rect 42208 22208 42210 22228
rect 45782 25050 45838 25052
rect 45862 25050 45918 25052
rect 45942 25050 45998 25052
rect 46022 25050 46078 25052
rect 45782 24998 45808 25050
rect 45808 24998 45838 25050
rect 45862 24998 45872 25050
rect 45872 24998 45918 25050
rect 45942 24998 45988 25050
rect 45988 24998 45998 25050
rect 46022 24998 46052 25050
rect 46052 24998 46078 25050
rect 45782 24996 45838 24998
rect 45862 24996 45918 24998
rect 45942 24996 45998 24998
rect 46022 24996 46078 24998
rect 45782 23962 45838 23964
rect 45862 23962 45918 23964
rect 45942 23962 45998 23964
rect 46022 23962 46078 23964
rect 45782 23910 45808 23962
rect 45808 23910 45838 23962
rect 45862 23910 45872 23962
rect 45872 23910 45918 23962
rect 45942 23910 45988 23962
rect 45988 23910 45998 23962
rect 46022 23910 46052 23962
rect 46052 23910 46078 23962
rect 45782 23908 45838 23910
rect 45862 23908 45918 23910
rect 45942 23908 45998 23910
rect 46022 23908 46078 23910
rect 45782 22874 45838 22876
rect 45862 22874 45918 22876
rect 45942 22874 45998 22876
rect 46022 22874 46078 22876
rect 45782 22822 45808 22874
rect 45808 22822 45838 22874
rect 45862 22822 45872 22874
rect 45872 22822 45918 22874
rect 45942 22822 45988 22874
rect 45988 22822 45998 22874
rect 46022 22822 46052 22874
rect 46052 22822 46078 22874
rect 45782 22820 45838 22822
rect 45862 22820 45918 22822
rect 45942 22820 45998 22822
rect 46022 22820 46078 22822
rect 46294 22208 46350 22264
rect 45782 21786 45838 21788
rect 45862 21786 45918 21788
rect 45942 21786 45998 21788
rect 46022 21786 46078 21788
rect 45782 21734 45808 21786
rect 45808 21734 45838 21786
rect 45862 21734 45872 21786
rect 45872 21734 45918 21786
rect 45942 21734 45988 21786
rect 45988 21734 45998 21786
rect 46022 21734 46052 21786
rect 46052 21734 46078 21786
rect 45782 21732 45838 21734
rect 45862 21732 45918 21734
rect 45942 21732 45998 21734
rect 46022 21732 46078 21734
rect 45782 20698 45838 20700
rect 45862 20698 45918 20700
rect 45942 20698 45998 20700
rect 46022 20698 46078 20700
rect 45782 20646 45808 20698
rect 45808 20646 45838 20698
rect 45862 20646 45872 20698
rect 45872 20646 45918 20698
rect 45942 20646 45988 20698
rect 45988 20646 45998 20698
rect 46022 20646 46052 20698
rect 46052 20646 46078 20698
rect 45782 20644 45838 20646
rect 45862 20644 45918 20646
rect 45942 20644 45998 20646
rect 46022 20644 46078 20646
rect 45782 19610 45838 19612
rect 45862 19610 45918 19612
rect 45942 19610 45998 19612
rect 46022 19610 46078 19612
rect 45782 19558 45808 19610
rect 45808 19558 45838 19610
rect 45862 19558 45872 19610
rect 45872 19558 45918 19610
rect 45942 19558 45988 19610
rect 45988 19558 45998 19610
rect 46022 19558 46052 19610
rect 46052 19558 46078 19610
rect 45782 19556 45838 19558
rect 45862 19556 45918 19558
rect 45942 19556 45998 19558
rect 46022 19556 46078 19558
rect 46386 19760 46442 19816
rect 46110 19252 46112 19272
rect 46112 19252 46164 19272
rect 46164 19252 46166 19272
rect 46110 19216 46166 19252
rect 46202 19116 46204 19136
rect 46204 19116 46256 19136
rect 46256 19116 46258 19136
rect 44362 18264 44418 18320
rect 42522 18164 42524 18184
rect 42524 18164 42576 18184
rect 42576 18164 42578 18184
rect 42522 18128 42578 18164
rect 36817 12538 36873 12540
rect 36897 12538 36953 12540
rect 36977 12538 37033 12540
rect 37057 12538 37113 12540
rect 36817 12486 36843 12538
rect 36843 12486 36873 12538
rect 36897 12486 36907 12538
rect 36907 12486 36953 12538
rect 36977 12486 37023 12538
rect 37023 12486 37033 12538
rect 37057 12486 37087 12538
rect 37087 12486 37113 12538
rect 36817 12484 36873 12486
rect 36897 12484 36953 12486
rect 36977 12484 37033 12486
rect 37057 12484 37113 12486
rect 44730 18808 44786 18864
rect 45782 18522 45838 18524
rect 45862 18522 45918 18524
rect 45942 18522 45998 18524
rect 46022 18522 46078 18524
rect 45782 18470 45808 18522
rect 45808 18470 45838 18522
rect 45862 18470 45872 18522
rect 45872 18470 45918 18522
rect 45942 18470 45988 18522
rect 45988 18470 45998 18522
rect 46022 18470 46052 18522
rect 46052 18470 46078 18522
rect 45782 18468 45838 18470
rect 45862 18468 45918 18470
rect 45942 18468 45998 18470
rect 46022 18468 46078 18470
rect 46202 19080 46258 19116
rect 46938 18128 46994 18184
rect 45782 17434 45838 17436
rect 45862 17434 45918 17436
rect 45942 17434 45998 17436
rect 46022 17434 46078 17436
rect 45782 17382 45808 17434
rect 45808 17382 45838 17434
rect 45862 17382 45872 17434
rect 45872 17382 45918 17434
rect 45942 17382 45988 17434
rect 45988 17382 45998 17434
rect 46022 17382 46052 17434
rect 46052 17382 46078 17434
rect 45782 17380 45838 17382
rect 45862 17380 45918 17382
rect 45942 17380 45998 17382
rect 46022 17380 46078 17382
rect 45782 16346 45838 16348
rect 45862 16346 45918 16348
rect 45942 16346 45998 16348
rect 46022 16346 46078 16348
rect 45782 16294 45808 16346
rect 45808 16294 45838 16346
rect 45862 16294 45872 16346
rect 45872 16294 45918 16346
rect 45942 16294 45988 16346
rect 45988 16294 45998 16346
rect 46022 16294 46052 16346
rect 46052 16294 46078 16346
rect 45782 16292 45838 16294
rect 45862 16292 45918 16294
rect 45942 16292 45998 16294
rect 46022 16292 46078 16294
rect 50710 20476 50712 20496
rect 50712 20476 50764 20496
rect 50764 20476 50766 20496
rect 50710 20440 50766 20476
rect 52090 20440 52146 20496
rect 52366 20440 52422 20496
rect 47858 18672 47914 18728
rect 47950 17060 48006 17096
rect 47950 17040 47952 17060
rect 47952 17040 48004 17060
rect 48004 17040 48006 17060
rect 45782 15258 45838 15260
rect 45862 15258 45918 15260
rect 45942 15258 45998 15260
rect 46022 15258 46078 15260
rect 45782 15206 45808 15258
rect 45808 15206 45838 15258
rect 45862 15206 45872 15258
rect 45872 15206 45918 15258
rect 45942 15206 45988 15258
rect 45988 15206 45998 15258
rect 46022 15206 46052 15258
rect 46052 15206 46078 15258
rect 45782 15204 45838 15206
rect 45862 15204 45918 15206
rect 45942 15204 45998 15206
rect 46022 15204 46078 15206
rect 45782 14170 45838 14172
rect 45862 14170 45918 14172
rect 45942 14170 45998 14172
rect 46022 14170 46078 14172
rect 45782 14118 45808 14170
rect 45808 14118 45838 14170
rect 45862 14118 45872 14170
rect 45872 14118 45918 14170
rect 45942 14118 45988 14170
rect 45988 14118 45998 14170
rect 46022 14118 46052 14170
rect 46052 14118 46078 14170
rect 45782 14116 45838 14118
rect 45862 14116 45918 14118
rect 45942 14116 45998 14118
rect 46022 14116 46078 14118
rect 45782 13082 45838 13084
rect 45862 13082 45918 13084
rect 45942 13082 45998 13084
rect 46022 13082 46078 13084
rect 45782 13030 45808 13082
rect 45808 13030 45838 13082
rect 45862 13030 45872 13082
rect 45872 13030 45918 13082
rect 45942 13030 45988 13082
rect 45988 13030 45998 13082
rect 46022 13030 46052 13082
rect 46052 13030 46078 13082
rect 45782 13028 45838 13030
rect 45862 13028 45918 13030
rect 45942 13028 45998 13030
rect 46022 13028 46078 13030
rect 45782 11994 45838 11996
rect 45862 11994 45918 11996
rect 45942 11994 45998 11996
rect 46022 11994 46078 11996
rect 45782 11942 45808 11994
rect 45808 11942 45838 11994
rect 45862 11942 45872 11994
rect 45872 11942 45918 11994
rect 45942 11942 45988 11994
rect 45988 11942 45998 11994
rect 46022 11942 46052 11994
rect 46052 11942 46078 11994
rect 45782 11940 45838 11942
rect 45862 11940 45918 11942
rect 45942 11940 45998 11942
rect 46022 11940 46078 11942
rect 36817 11450 36873 11452
rect 36897 11450 36953 11452
rect 36977 11450 37033 11452
rect 37057 11450 37113 11452
rect 36817 11398 36843 11450
rect 36843 11398 36873 11450
rect 36897 11398 36907 11450
rect 36907 11398 36953 11450
rect 36977 11398 37023 11450
rect 37023 11398 37033 11450
rect 37057 11398 37087 11450
rect 37087 11398 37113 11450
rect 36817 11396 36873 11398
rect 36897 11396 36953 11398
rect 36977 11396 37033 11398
rect 37057 11396 37113 11398
rect 45782 10906 45838 10908
rect 45862 10906 45918 10908
rect 45942 10906 45998 10908
rect 46022 10906 46078 10908
rect 45782 10854 45808 10906
rect 45808 10854 45838 10906
rect 45862 10854 45872 10906
rect 45872 10854 45918 10906
rect 45942 10854 45988 10906
rect 45988 10854 45998 10906
rect 46022 10854 46052 10906
rect 46052 10854 46078 10906
rect 45782 10852 45838 10854
rect 45862 10852 45918 10854
rect 45942 10852 45998 10854
rect 46022 10852 46078 10854
rect 27852 9818 27908 9820
rect 27932 9818 27988 9820
rect 28012 9818 28068 9820
rect 28092 9818 28148 9820
rect 27852 9766 27878 9818
rect 27878 9766 27908 9818
rect 27932 9766 27942 9818
rect 27942 9766 27988 9818
rect 28012 9766 28058 9818
rect 28058 9766 28068 9818
rect 28092 9766 28122 9818
rect 28122 9766 28148 9818
rect 27852 9764 27908 9766
rect 27932 9764 27988 9766
rect 28012 9764 28068 9766
rect 28092 9764 28148 9766
rect 27852 8730 27908 8732
rect 27932 8730 27988 8732
rect 28012 8730 28068 8732
rect 28092 8730 28148 8732
rect 27852 8678 27878 8730
rect 27878 8678 27908 8730
rect 27932 8678 27942 8730
rect 27942 8678 27988 8730
rect 28012 8678 28058 8730
rect 28058 8678 28068 8730
rect 28092 8678 28122 8730
rect 28122 8678 28148 8730
rect 27852 8676 27908 8678
rect 27932 8676 27988 8678
rect 28012 8676 28068 8678
rect 28092 8676 28148 8678
rect 27852 7642 27908 7644
rect 27932 7642 27988 7644
rect 28012 7642 28068 7644
rect 28092 7642 28148 7644
rect 27852 7590 27878 7642
rect 27878 7590 27908 7642
rect 27932 7590 27942 7642
rect 27942 7590 27988 7642
rect 28012 7590 28058 7642
rect 28058 7590 28068 7642
rect 28092 7590 28122 7642
rect 28122 7590 28148 7642
rect 27852 7588 27908 7590
rect 27932 7588 27988 7590
rect 28012 7588 28068 7590
rect 28092 7588 28148 7590
rect 27852 6554 27908 6556
rect 27932 6554 27988 6556
rect 28012 6554 28068 6556
rect 28092 6554 28148 6556
rect 27852 6502 27878 6554
rect 27878 6502 27908 6554
rect 27932 6502 27942 6554
rect 27942 6502 27988 6554
rect 28012 6502 28058 6554
rect 28058 6502 28068 6554
rect 28092 6502 28122 6554
rect 28122 6502 28148 6554
rect 27852 6500 27908 6502
rect 27932 6500 27988 6502
rect 28012 6500 28068 6502
rect 28092 6500 28148 6502
rect 36817 10362 36873 10364
rect 36897 10362 36953 10364
rect 36977 10362 37033 10364
rect 37057 10362 37113 10364
rect 36817 10310 36843 10362
rect 36843 10310 36873 10362
rect 36897 10310 36907 10362
rect 36907 10310 36953 10362
rect 36977 10310 37023 10362
rect 37023 10310 37033 10362
rect 37057 10310 37087 10362
rect 37087 10310 37113 10362
rect 36817 10308 36873 10310
rect 36897 10308 36953 10310
rect 36977 10308 37033 10310
rect 37057 10308 37113 10310
rect 36817 9274 36873 9276
rect 36897 9274 36953 9276
rect 36977 9274 37033 9276
rect 37057 9274 37113 9276
rect 36817 9222 36843 9274
rect 36843 9222 36873 9274
rect 36897 9222 36907 9274
rect 36907 9222 36953 9274
rect 36977 9222 37023 9274
rect 37023 9222 37033 9274
rect 37057 9222 37087 9274
rect 37087 9222 37113 9274
rect 36817 9220 36873 9222
rect 36897 9220 36953 9222
rect 36977 9220 37033 9222
rect 37057 9220 37113 9222
rect 45782 9818 45838 9820
rect 45862 9818 45918 9820
rect 45942 9818 45998 9820
rect 46022 9818 46078 9820
rect 45782 9766 45808 9818
rect 45808 9766 45838 9818
rect 45862 9766 45872 9818
rect 45872 9766 45918 9818
rect 45942 9766 45988 9818
rect 45988 9766 45998 9818
rect 46022 9766 46052 9818
rect 46052 9766 46078 9818
rect 45782 9764 45838 9766
rect 45862 9764 45918 9766
rect 45942 9764 45998 9766
rect 46022 9764 46078 9766
rect 45782 8730 45838 8732
rect 45862 8730 45918 8732
rect 45942 8730 45998 8732
rect 46022 8730 46078 8732
rect 45782 8678 45808 8730
rect 45808 8678 45838 8730
rect 45862 8678 45872 8730
rect 45872 8678 45918 8730
rect 45942 8678 45988 8730
rect 45988 8678 45998 8730
rect 46022 8678 46052 8730
rect 46052 8678 46078 8730
rect 45782 8676 45838 8678
rect 45862 8676 45918 8678
rect 45942 8676 45998 8678
rect 46022 8676 46078 8678
rect 36817 8186 36873 8188
rect 36897 8186 36953 8188
rect 36977 8186 37033 8188
rect 37057 8186 37113 8188
rect 36817 8134 36843 8186
rect 36843 8134 36873 8186
rect 36897 8134 36907 8186
rect 36907 8134 36953 8186
rect 36977 8134 37023 8186
rect 37023 8134 37033 8186
rect 37057 8134 37087 8186
rect 37087 8134 37113 8186
rect 36817 8132 36873 8134
rect 36897 8132 36953 8134
rect 36977 8132 37033 8134
rect 37057 8132 37113 8134
rect 27852 5466 27908 5468
rect 27932 5466 27988 5468
rect 28012 5466 28068 5468
rect 28092 5466 28148 5468
rect 27852 5414 27878 5466
rect 27878 5414 27908 5466
rect 27932 5414 27942 5466
rect 27942 5414 27988 5466
rect 28012 5414 28058 5466
rect 28058 5414 28068 5466
rect 28092 5414 28122 5466
rect 28122 5414 28148 5466
rect 27852 5412 27908 5414
rect 27932 5412 27988 5414
rect 28012 5412 28068 5414
rect 28092 5412 28148 5414
rect 27852 4378 27908 4380
rect 27932 4378 27988 4380
rect 28012 4378 28068 4380
rect 28092 4378 28148 4380
rect 27852 4326 27878 4378
rect 27878 4326 27908 4378
rect 27932 4326 27942 4378
rect 27942 4326 27988 4378
rect 28012 4326 28058 4378
rect 28058 4326 28068 4378
rect 28092 4326 28122 4378
rect 28122 4326 28148 4378
rect 27852 4324 27908 4326
rect 27932 4324 27988 4326
rect 28012 4324 28068 4326
rect 28092 4324 28148 4326
rect 27852 3290 27908 3292
rect 27932 3290 27988 3292
rect 28012 3290 28068 3292
rect 28092 3290 28148 3292
rect 27852 3238 27878 3290
rect 27878 3238 27908 3290
rect 27932 3238 27942 3290
rect 27942 3238 27988 3290
rect 28012 3238 28058 3290
rect 28058 3238 28068 3290
rect 28092 3238 28122 3290
rect 28122 3238 28148 3290
rect 27852 3236 27908 3238
rect 27932 3236 27988 3238
rect 28012 3236 28068 3238
rect 28092 3236 28148 3238
rect 9921 2202 9977 2204
rect 10001 2202 10057 2204
rect 10081 2202 10137 2204
rect 10161 2202 10217 2204
rect 9921 2150 9947 2202
rect 9947 2150 9977 2202
rect 10001 2150 10011 2202
rect 10011 2150 10057 2202
rect 10081 2150 10127 2202
rect 10127 2150 10137 2202
rect 10161 2150 10191 2202
rect 10191 2150 10217 2202
rect 9921 2148 9977 2150
rect 10001 2148 10057 2150
rect 10081 2148 10137 2150
rect 10161 2148 10217 2150
rect 27852 2202 27908 2204
rect 27932 2202 27988 2204
rect 28012 2202 28068 2204
rect 28092 2202 28148 2204
rect 27852 2150 27878 2202
rect 27878 2150 27908 2202
rect 27932 2150 27942 2202
rect 27942 2150 27988 2202
rect 28012 2150 28058 2202
rect 28058 2150 28068 2202
rect 28092 2150 28122 2202
rect 28122 2150 28148 2202
rect 27852 2148 27908 2150
rect 27932 2148 27988 2150
rect 28012 2148 28068 2150
rect 28092 2148 28148 2150
rect 45782 7642 45838 7644
rect 45862 7642 45918 7644
rect 45942 7642 45998 7644
rect 46022 7642 46078 7644
rect 45782 7590 45808 7642
rect 45808 7590 45838 7642
rect 45862 7590 45872 7642
rect 45872 7590 45918 7642
rect 45942 7590 45988 7642
rect 45988 7590 45998 7642
rect 46022 7590 46052 7642
rect 46052 7590 46078 7642
rect 45782 7588 45838 7590
rect 45862 7588 45918 7590
rect 45942 7588 45998 7590
rect 46022 7588 46078 7590
rect 36817 7098 36873 7100
rect 36897 7098 36953 7100
rect 36977 7098 37033 7100
rect 37057 7098 37113 7100
rect 36817 7046 36843 7098
rect 36843 7046 36873 7098
rect 36897 7046 36907 7098
rect 36907 7046 36953 7098
rect 36977 7046 37023 7098
rect 37023 7046 37033 7098
rect 37057 7046 37087 7098
rect 37087 7046 37113 7098
rect 36817 7044 36873 7046
rect 36897 7044 36953 7046
rect 36977 7044 37033 7046
rect 37057 7044 37113 7046
rect 36817 6010 36873 6012
rect 36897 6010 36953 6012
rect 36977 6010 37033 6012
rect 37057 6010 37113 6012
rect 36817 5958 36843 6010
rect 36843 5958 36873 6010
rect 36897 5958 36907 6010
rect 36907 5958 36953 6010
rect 36977 5958 37023 6010
rect 37023 5958 37033 6010
rect 37057 5958 37087 6010
rect 37087 5958 37113 6010
rect 36817 5956 36873 5958
rect 36897 5956 36953 5958
rect 36977 5956 37033 5958
rect 37057 5956 37113 5958
rect 36817 4922 36873 4924
rect 36897 4922 36953 4924
rect 36977 4922 37033 4924
rect 37057 4922 37113 4924
rect 36817 4870 36843 4922
rect 36843 4870 36873 4922
rect 36897 4870 36907 4922
rect 36907 4870 36953 4922
rect 36977 4870 37023 4922
rect 37023 4870 37033 4922
rect 37057 4870 37087 4922
rect 37087 4870 37113 4922
rect 36817 4868 36873 4870
rect 36897 4868 36953 4870
rect 36977 4868 37033 4870
rect 37057 4868 37113 4870
rect 51078 6840 51134 6896
rect 45782 6554 45838 6556
rect 45862 6554 45918 6556
rect 45942 6554 45998 6556
rect 46022 6554 46078 6556
rect 45782 6502 45808 6554
rect 45808 6502 45838 6554
rect 45862 6502 45872 6554
rect 45872 6502 45918 6554
rect 45942 6502 45988 6554
rect 45988 6502 45998 6554
rect 46022 6502 46052 6554
rect 46052 6502 46078 6554
rect 45782 6500 45838 6502
rect 45862 6500 45918 6502
rect 45942 6500 45998 6502
rect 46022 6500 46078 6502
rect 45782 5466 45838 5468
rect 45862 5466 45918 5468
rect 45942 5466 45998 5468
rect 46022 5466 46078 5468
rect 45782 5414 45808 5466
rect 45808 5414 45838 5466
rect 45862 5414 45872 5466
rect 45872 5414 45918 5466
rect 45942 5414 45988 5466
rect 45988 5414 45998 5466
rect 46022 5414 46052 5466
rect 46052 5414 46078 5466
rect 45782 5412 45838 5414
rect 45862 5412 45918 5414
rect 45942 5412 45998 5414
rect 46022 5412 46078 5414
rect 36817 3834 36873 3836
rect 36897 3834 36953 3836
rect 36977 3834 37033 3836
rect 37057 3834 37113 3836
rect 36817 3782 36843 3834
rect 36843 3782 36873 3834
rect 36897 3782 36907 3834
rect 36907 3782 36953 3834
rect 36977 3782 37023 3834
rect 37023 3782 37033 3834
rect 37057 3782 37087 3834
rect 37087 3782 37113 3834
rect 36817 3780 36873 3782
rect 36897 3780 36953 3782
rect 36977 3780 37033 3782
rect 37057 3780 37113 3782
rect 36817 2746 36873 2748
rect 36897 2746 36953 2748
rect 36977 2746 37033 2748
rect 37057 2746 37113 2748
rect 36817 2694 36843 2746
rect 36843 2694 36873 2746
rect 36897 2694 36907 2746
rect 36907 2694 36953 2746
rect 36977 2694 37023 2746
rect 37023 2694 37033 2746
rect 37057 2694 37087 2746
rect 37087 2694 37113 2746
rect 36817 2692 36873 2694
rect 36897 2692 36953 2694
rect 36977 2692 37033 2694
rect 37057 2692 37113 2694
rect 45782 4378 45838 4380
rect 45862 4378 45918 4380
rect 45942 4378 45998 4380
rect 46022 4378 46078 4380
rect 45782 4326 45808 4378
rect 45808 4326 45838 4378
rect 45862 4326 45872 4378
rect 45872 4326 45918 4378
rect 45942 4326 45988 4378
rect 45988 4326 45998 4378
rect 46022 4326 46052 4378
rect 46052 4326 46078 4378
rect 45782 4324 45838 4326
rect 45862 4324 45918 4326
rect 45942 4324 45998 4326
rect 46022 4324 46078 4326
rect 45782 3290 45838 3292
rect 45862 3290 45918 3292
rect 45942 3290 45998 3292
rect 46022 3290 46078 3292
rect 45782 3238 45808 3290
rect 45808 3238 45838 3290
rect 45862 3238 45872 3290
rect 45872 3238 45918 3290
rect 45942 3238 45988 3290
rect 45988 3238 45998 3290
rect 46022 3238 46052 3290
rect 46052 3238 46078 3290
rect 45782 3236 45838 3238
rect 45862 3236 45918 3238
rect 45942 3236 45998 3238
rect 46022 3236 46078 3238
rect 45782 2202 45838 2204
rect 45862 2202 45918 2204
rect 45942 2202 45998 2204
rect 46022 2202 46078 2204
rect 45782 2150 45808 2202
rect 45808 2150 45838 2202
rect 45862 2150 45872 2202
rect 45872 2150 45918 2202
rect 45942 2150 45988 2202
rect 45988 2150 45998 2202
rect 46022 2150 46052 2202
rect 46052 2150 46078 2202
rect 45782 2148 45838 2150
rect 45862 2148 45918 2150
rect 45942 2148 45998 2150
rect 46022 2148 46078 2150
<< metal3 >>
rect 9909 25056 10229 25057
rect 9909 24992 9917 25056
rect 9981 24992 9997 25056
rect 10061 24992 10077 25056
rect 10141 24992 10157 25056
rect 10221 24992 10229 25056
rect 9909 24991 10229 24992
rect 27840 25056 28160 25057
rect 27840 24992 27848 25056
rect 27912 24992 27928 25056
rect 27992 24992 28008 25056
rect 28072 24992 28088 25056
rect 28152 24992 28160 25056
rect 27840 24991 28160 24992
rect 45770 25056 46090 25057
rect 45770 24992 45778 25056
rect 45842 24992 45858 25056
rect 45922 24992 45938 25056
rect 46002 24992 46018 25056
rect 46082 24992 46090 25056
rect 45770 24991 46090 24992
rect 18874 24512 19194 24513
rect 18874 24448 18882 24512
rect 18946 24448 18962 24512
rect 19026 24448 19042 24512
rect 19106 24448 19122 24512
rect 19186 24448 19194 24512
rect 18874 24447 19194 24448
rect 36805 24512 37125 24513
rect 36805 24448 36813 24512
rect 36877 24448 36893 24512
rect 36957 24448 36973 24512
rect 37037 24448 37053 24512
rect 37117 24448 37125 24512
rect 36805 24447 37125 24448
rect 9909 23968 10229 23969
rect 9909 23904 9917 23968
rect 9981 23904 9997 23968
rect 10061 23904 10077 23968
rect 10141 23904 10157 23968
rect 10221 23904 10229 23968
rect 9909 23903 10229 23904
rect 27840 23968 28160 23969
rect 27840 23904 27848 23968
rect 27912 23904 27928 23968
rect 27992 23904 28008 23968
rect 28072 23904 28088 23968
rect 28152 23904 28160 23968
rect 27840 23903 28160 23904
rect 45770 23968 46090 23969
rect 45770 23904 45778 23968
rect 45842 23904 45858 23968
rect 45922 23904 45938 23968
rect 46002 23904 46018 23968
rect 46082 23904 46090 23968
rect 45770 23903 46090 23904
rect 18874 23424 19194 23425
rect 18874 23360 18882 23424
rect 18946 23360 18962 23424
rect 19026 23360 19042 23424
rect 19106 23360 19122 23424
rect 19186 23360 19194 23424
rect 18874 23359 19194 23360
rect 36805 23424 37125 23425
rect 36805 23360 36813 23424
rect 36877 23360 36893 23424
rect 36957 23360 36973 23424
rect 37037 23360 37053 23424
rect 37117 23360 37125 23424
rect 36805 23359 37125 23360
rect 32489 23082 32555 23085
rect 38561 23082 38627 23085
rect 32489 23080 38627 23082
rect 32489 23024 32494 23080
rect 32550 23024 38566 23080
rect 38622 23024 38627 23080
rect 32489 23022 38627 23024
rect 32489 23019 32555 23022
rect 38561 23019 38627 23022
rect 9909 22880 10229 22881
rect 9909 22816 9917 22880
rect 9981 22816 9997 22880
rect 10061 22816 10077 22880
rect 10141 22816 10157 22880
rect 10221 22816 10229 22880
rect 9909 22815 10229 22816
rect 27840 22880 28160 22881
rect 27840 22816 27848 22880
rect 27912 22816 27928 22880
rect 27992 22816 28008 22880
rect 28072 22816 28088 22880
rect 28152 22816 28160 22880
rect 27840 22815 28160 22816
rect 45770 22880 46090 22881
rect 45770 22816 45778 22880
rect 45842 22816 45858 22880
rect 45922 22816 45938 22880
rect 46002 22816 46018 22880
rect 46082 22816 46090 22880
rect 45770 22815 46090 22816
rect 24025 22538 24091 22541
rect 24301 22538 24367 22541
rect 28257 22538 28323 22541
rect 24025 22536 28323 22538
rect 24025 22480 24030 22536
rect 24086 22480 24306 22536
rect 24362 22480 28262 22536
rect 28318 22480 28323 22536
rect 24025 22478 28323 22480
rect 24025 22475 24091 22478
rect 24301 22475 24367 22478
rect 28257 22475 28323 22478
rect 18874 22336 19194 22337
rect 18874 22272 18882 22336
rect 18946 22272 18962 22336
rect 19026 22272 19042 22336
rect 19106 22272 19122 22336
rect 19186 22272 19194 22336
rect 18874 22271 19194 22272
rect 36805 22336 37125 22337
rect 36805 22272 36813 22336
rect 36877 22272 36893 22336
rect 36957 22272 36973 22336
rect 37037 22272 37053 22336
rect 37117 22272 37125 22336
rect 36805 22271 37125 22272
rect 42149 22266 42215 22269
rect 46289 22266 46355 22269
rect 42149 22264 46355 22266
rect 42149 22208 42154 22264
rect 42210 22208 46294 22264
rect 46350 22208 46355 22264
rect 42149 22206 46355 22208
rect 42149 22203 42215 22206
rect 46289 22203 46355 22206
rect 2497 21994 2563 21997
rect 7281 21994 7347 21997
rect 2497 21992 7347 21994
rect 2497 21936 2502 21992
rect 2558 21936 7286 21992
rect 7342 21936 7347 21992
rect 2497 21934 7347 21936
rect 2497 21931 2563 21934
rect 7281 21931 7347 21934
rect 9909 21792 10229 21793
rect 9909 21728 9917 21792
rect 9981 21728 9997 21792
rect 10061 21728 10077 21792
rect 10141 21728 10157 21792
rect 10221 21728 10229 21792
rect 9909 21727 10229 21728
rect 27840 21792 28160 21793
rect 27840 21728 27848 21792
rect 27912 21728 27928 21792
rect 27992 21728 28008 21792
rect 28072 21728 28088 21792
rect 28152 21728 28160 21792
rect 27840 21727 28160 21728
rect 45770 21792 46090 21793
rect 45770 21728 45778 21792
rect 45842 21728 45858 21792
rect 45922 21728 45938 21792
rect 46002 21728 46018 21792
rect 46082 21728 46090 21792
rect 45770 21727 46090 21728
rect 12249 21586 12315 21589
rect 12709 21586 12775 21589
rect 12249 21584 12775 21586
rect 12249 21528 12254 21584
rect 12310 21528 12714 21584
rect 12770 21528 12775 21584
rect 12249 21526 12775 21528
rect 12249 21523 12315 21526
rect 12709 21523 12775 21526
rect 28349 21450 28415 21453
rect 28901 21450 28967 21453
rect 28349 21448 28967 21450
rect 28349 21392 28354 21448
rect 28410 21392 28906 21448
rect 28962 21392 28967 21448
rect 28349 21390 28967 21392
rect 28349 21387 28415 21390
rect 28901 21387 28967 21390
rect 18874 21248 19194 21249
rect 18874 21184 18882 21248
rect 18946 21184 18962 21248
rect 19026 21184 19042 21248
rect 19106 21184 19122 21248
rect 19186 21184 19194 21248
rect 18874 21183 19194 21184
rect 36805 21248 37125 21249
rect 36805 21184 36813 21248
rect 36877 21184 36893 21248
rect 36957 21184 36973 21248
rect 37037 21184 37053 21248
rect 37117 21184 37125 21248
rect 36805 21183 37125 21184
rect 26877 21042 26943 21045
rect 28717 21042 28783 21045
rect 26877 21040 28783 21042
rect 26877 20984 26882 21040
rect 26938 20984 28722 21040
rect 28778 20984 28783 21040
rect 26877 20982 28783 20984
rect 26877 20979 26943 20982
rect 28717 20979 28783 20982
rect 9909 20704 10229 20705
rect 9909 20640 9917 20704
rect 9981 20640 9997 20704
rect 10061 20640 10077 20704
rect 10141 20640 10157 20704
rect 10221 20640 10229 20704
rect 9909 20639 10229 20640
rect 27840 20704 28160 20705
rect 27840 20640 27848 20704
rect 27912 20640 27928 20704
rect 27992 20640 28008 20704
rect 28072 20640 28088 20704
rect 28152 20640 28160 20704
rect 27840 20639 28160 20640
rect 45770 20704 46090 20705
rect 45770 20640 45778 20704
rect 45842 20640 45858 20704
rect 45922 20640 45938 20704
rect 46002 20640 46018 20704
rect 46082 20640 46090 20704
rect 45770 20639 46090 20640
rect 24025 20498 24091 20501
rect 26969 20498 27035 20501
rect 24025 20496 27035 20498
rect 24025 20440 24030 20496
rect 24086 20440 26974 20496
rect 27030 20440 27035 20496
rect 24025 20438 27035 20440
rect 24025 20435 24091 20438
rect 26969 20435 27035 20438
rect 50705 20498 50771 20501
rect 52085 20498 52151 20501
rect 50705 20496 52151 20498
rect 50705 20440 50710 20496
rect 50766 20440 52090 20496
rect 52146 20440 52151 20496
rect 50705 20438 52151 20440
rect 50705 20435 50771 20438
rect 52085 20435 52151 20438
rect 52361 20498 52427 20501
rect 55200 20498 56000 20528
rect 52361 20496 56000 20498
rect 52361 20440 52366 20496
rect 52422 20440 56000 20496
rect 52361 20438 56000 20440
rect 52361 20435 52427 20438
rect 55200 20408 56000 20438
rect 18874 20160 19194 20161
rect 18874 20096 18882 20160
rect 18946 20096 18962 20160
rect 19026 20096 19042 20160
rect 19106 20096 19122 20160
rect 19186 20096 19194 20160
rect 18874 20095 19194 20096
rect 36805 20160 37125 20161
rect 36805 20096 36813 20160
rect 36877 20096 36893 20160
rect 36957 20096 36973 20160
rect 37037 20096 37053 20160
rect 37117 20096 37125 20160
rect 36805 20095 37125 20096
rect 39573 19818 39639 19821
rect 46381 19818 46447 19821
rect 39573 19816 46447 19818
rect 39573 19760 39578 19816
rect 39634 19760 46386 19816
rect 46442 19760 46447 19816
rect 39573 19758 46447 19760
rect 39573 19755 39639 19758
rect 46381 19755 46447 19758
rect 9909 19616 10229 19617
rect 9909 19552 9917 19616
rect 9981 19552 9997 19616
rect 10061 19552 10077 19616
rect 10141 19552 10157 19616
rect 10221 19552 10229 19616
rect 9909 19551 10229 19552
rect 27840 19616 28160 19617
rect 27840 19552 27848 19616
rect 27912 19552 27928 19616
rect 27992 19552 28008 19616
rect 28072 19552 28088 19616
rect 28152 19552 28160 19616
rect 27840 19551 28160 19552
rect 45770 19616 46090 19617
rect 45770 19552 45778 19616
rect 45842 19552 45858 19616
rect 45922 19552 45938 19616
rect 46002 19552 46018 19616
rect 46082 19552 46090 19616
rect 45770 19551 46090 19552
rect 22001 19410 22067 19413
rect 27797 19410 27863 19413
rect 22001 19408 27863 19410
rect 22001 19352 22006 19408
rect 22062 19352 27802 19408
rect 27858 19352 27863 19408
rect 22001 19350 27863 19352
rect 22001 19347 22067 19350
rect 27797 19347 27863 19350
rect 8293 19274 8359 19277
rect 9489 19274 9555 19277
rect 8293 19272 9555 19274
rect 8293 19216 8298 19272
rect 8354 19216 9494 19272
rect 9550 19216 9555 19272
rect 8293 19214 9555 19216
rect 8293 19211 8359 19214
rect 9489 19211 9555 19214
rect 41597 19274 41663 19277
rect 46105 19274 46171 19277
rect 41597 19272 46171 19274
rect 41597 19216 41602 19272
rect 41658 19216 46110 19272
rect 46166 19216 46171 19272
rect 41597 19214 46171 19216
rect 41597 19211 41663 19214
rect 46105 19211 46171 19214
rect 39021 19138 39087 19141
rect 46197 19138 46263 19141
rect 39021 19136 46263 19138
rect 39021 19080 39026 19136
rect 39082 19080 46202 19136
rect 46258 19080 46263 19136
rect 39021 19078 46263 19080
rect 39021 19075 39087 19078
rect 46197 19075 46263 19078
rect 18874 19072 19194 19073
rect 18874 19008 18882 19072
rect 18946 19008 18962 19072
rect 19026 19008 19042 19072
rect 19106 19008 19122 19072
rect 19186 19008 19194 19072
rect 18874 19007 19194 19008
rect 36805 19072 37125 19073
rect 36805 19008 36813 19072
rect 36877 19008 36893 19072
rect 36957 19008 36973 19072
rect 37037 19008 37053 19072
rect 37117 19008 37125 19072
rect 36805 19007 37125 19008
rect 32397 18866 32463 18869
rect 33685 18866 33751 18869
rect 36721 18866 36787 18869
rect 32397 18864 36787 18866
rect 32397 18808 32402 18864
rect 32458 18808 33690 18864
rect 33746 18808 36726 18864
rect 36782 18808 36787 18864
rect 32397 18806 36787 18808
rect 32397 18803 32463 18806
rect 33685 18803 33751 18806
rect 36721 18803 36787 18806
rect 41321 18866 41387 18869
rect 44725 18866 44791 18869
rect 41321 18864 44791 18866
rect 41321 18808 41326 18864
rect 41382 18808 44730 18864
rect 44786 18808 44791 18864
rect 41321 18806 44791 18808
rect 41321 18803 41387 18806
rect 44725 18803 44791 18806
rect 29361 18730 29427 18733
rect 38285 18730 38351 18733
rect 29361 18728 38351 18730
rect 29361 18672 29366 18728
rect 29422 18672 38290 18728
rect 38346 18672 38351 18728
rect 29361 18670 38351 18672
rect 29361 18667 29427 18670
rect 38285 18667 38351 18670
rect 38929 18730 38995 18733
rect 47853 18730 47919 18733
rect 38929 18728 47919 18730
rect 38929 18672 38934 18728
rect 38990 18672 47858 18728
rect 47914 18672 47919 18728
rect 38929 18670 47919 18672
rect 38929 18667 38995 18670
rect 47853 18667 47919 18670
rect 31753 18594 31819 18597
rect 32305 18594 32371 18597
rect 32949 18594 33015 18597
rect 33869 18594 33935 18597
rect 39941 18594 40007 18597
rect 31753 18592 40007 18594
rect 31753 18536 31758 18592
rect 31814 18536 32310 18592
rect 32366 18536 32954 18592
rect 33010 18536 33874 18592
rect 33930 18536 39946 18592
rect 40002 18536 40007 18592
rect 31753 18534 40007 18536
rect 31753 18531 31819 18534
rect 32305 18531 32371 18534
rect 32949 18531 33015 18534
rect 33869 18531 33935 18534
rect 39941 18531 40007 18534
rect 9909 18528 10229 18529
rect 9909 18464 9917 18528
rect 9981 18464 9997 18528
rect 10061 18464 10077 18528
rect 10141 18464 10157 18528
rect 10221 18464 10229 18528
rect 9909 18463 10229 18464
rect 27840 18528 28160 18529
rect 27840 18464 27848 18528
rect 27912 18464 27928 18528
rect 27992 18464 28008 18528
rect 28072 18464 28088 18528
rect 28152 18464 28160 18528
rect 27840 18463 28160 18464
rect 45770 18528 46090 18529
rect 45770 18464 45778 18528
rect 45842 18464 45858 18528
rect 45922 18464 45938 18528
rect 46002 18464 46018 18528
rect 46082 18464 46090 18528
rect 45770 18463 46090 18464
rect 30005 18458 30071 18461
rect 35617 18458 35683 18461
rect 30005 18456 35683 18458
rect 30005 18400 30010 18456
rect 30066 18400 35622 18456
rect 35678 18400 35683 18456
rect 30005 18398 35683 18400
rect 30005 18395 30071 18398
rect 35617 18395 35683 18398
rect 41597 18322 41663 18325
rect 44357 18322 44423 18325
rect 41597 18320 44423 18322
rect 41597 18264 41602 18320
rect 41658 18264 44362 18320
rect 44418 18264 44423 18320
rect 41597 18262 44423 18264
rect 41597 18259 41663 18262
rect 44357 18259 44423 18262
rect 42517 18186 42583 18189
rect 46933 18186 46999 18189
rect 42517 18184 46999 18186
rect 42517 18128 42522 18184
rect 42578 18128 46938 18184
rect 46994 18128 46999 18184
rect 42517 18126 46999 18128
rect 42517 18123 42583 18126
rect 46933 18123 46999 18126
rect 18874 17984 19194 17985
rect 18874 17920 18882 17984
rect 18946 17920 18962 17984
rect 19026 17920 19042 17984
rect 19106 17920 19122 17984
rect 19186 17920 19194 17984
rect 18874 17919 19194 17920
rect 36805 17984 37125 17985
rect 36805 17920 36813 17984
rect 36877 17920 36893 17984
rect 36957 17920 36973 17984
rect 37037 17920 37053 17984
rect 37117 17920 37125 17984
rect 36805 17919 37125 17920
rect 25773 17778 25839 17781
rect 41045 17778 41111 17781
rect 25773 17776 41111 17778
rect 25773 17720 25778 17776
rect 25834 17720 41050 17776
rect 41106 17720 41111 17776
rect 25773 17718 41111 17720
rect 25773 17715 25839 17718
rect 41045 17715 41111 17718
rect 34513 17642 34579 17645
rect 37917 17642 37983 17645
rect 34513 17640 37983 17642
rect 34513 17584 34518 17640
rect 34574 17584 37922 17640
rect 37978 17584 37983 17640
rect 34513 17582 37983 17584
rect 34513 17579 34579 17582
rect 37917 17579 37983 17582
rect 28625 17506 28691 17509
rect 28901 17506 28967 17509
rect 28625 17504 28967 17506
rect 28625 17448 28630 17504
rect 28686 17448 28906 17504
rect 28962 17448 28967 17504
rect 28625 17446 28967 17448
rect 28625 17443 28691 17446
rect 28901 17443 28967 17446
rect 9909 17440 10229 17441
rect 9909 17376 9917 17440
rect 9981 17376 9997 17440
rect 10061 17376 10077 17440
rect 10141 17376 10157 17440
rect 10221 17376 10229 17440
rect 9909 17375 10229 17376
rect 27840 17440 28160 17441
rect 27840 17376 27848 17440
rect 27912 17376 27928 17440
rect 27992 17376 28008 17440
rect 28072 17376 28088 17440
rect 28152 17376 28160 17440
rect 27840 17375 28160 17376
rect 45770 17440 46090 17441
rect 45770 17376 45778 17440
rect 45842 17376 45858 17440
rect 45922 17376 45938 17440
rect 46002 17376 46018 17440
rect 46082 17376 46090 17440
rect 45770 17375 46090 17376
rect 29821 17370 29887 17373
rect 36077 17370 36143 17373
rect 29821 17368 36143 17370
rect 29821 17312 29826 17368
rect 29882 17312 36082 17368
rect 36138 17312 36143 17368
rect 29821 17310 36143 17312
rect 29821 17307 29887 17310
rect 36077 17307 36143 17310
rect 36445 17370 36511 17373
rect 40033 17370 40099 17373
rect 40861 17370 40927 17373
rect 36445 17368 40927 17370
rect 36445 17312 36450 17368
rect 36506 17312 40038 17368
rect 40094 17312 40866 17368
rect 40922 17312 40927 17368
rect 36445 17310 40927 17312
rect 36445 17307 36511 17310
rect 40033 17307 40099 17310
rect 40861 17307 40927 17310
rect 39481 17098 39547 17101
rect 47945 17098 48011 17101
rect 39481 17096 48011 17098
rect 39481 17040 39486 17096
rect 39542 17040 47950 17096
rect 48006 17040 48011 17096
rect 39481 17038 48011 17040
rect 39481 17035 39547 17038
rect 47945 17035 48011 17038
rect 18874 16896 19194 16897
rect 18874 16832 18882 16896
rect 18946 16832 18962 16896
rect 19026 16832 19042 16896
rect 19106 16832 19122 16896
rect 19186 16832 19194 16896
rect 18874 16831 19194 16832
rect 36805 16896 37125 16897
rect 36805 16832 36813 16896
rect 36877 16832 36893 16896
rect 36957 16832 36973 16896
rect 37037 16832 37053 16896
rect 37117 16832 37125 16896
rect 36805 16831 37125 16832
rect 30465 16690 30531 16693
rect 37181 16690 37247 16693
rect 30465 16688 37247 16690
rect 30465 16632 30470 16688
rect 30526 16632 37186 16688
rect 37242 16632 37247 16688
rect 30465 16630 37247 16632
rect 30465 16627 30531 16630
rect 37181 16627 37247 16630
rect 24393 16554 24459 16557
rect 25957 16554 26023 16557
rect 24393 16552 26023 16554
rect 24393 16496 24398 16552
rect 24454 16496 25962 16552
rect 26018 16496 26023 16552
rect 24393 16494 26023 16496
rect 24393 16491 24459 16494
rect 25957 16491 26023 16494
rect 9909 16352 10229 16353
rect 9909 16288 9917 16352
rect 9981 16288 9997 16352
rect 10061 16288 10077 16352
rect 10141 16288 10157 16352
rect 10221 16288 10229 16352
rect 9909 16287 10229 16288
rect 27840 16352 28160 16353
rect 27840 16288 27848 16352
rect 27912 16288 27928 16352
rect 27992 16288 28008 16352
rect 28072 16288 28088 16352
rect 28152 16288 28160 16352
rect 27840 16287 28160 16288
rect 45770 16352 46090 16353
rect 45770 16288 45778 16352
rect 45842 16288 45858 16352
rect 45922 16288 45938 16352
rect 46002 16288 46018 16352
rect 46082 16288 46090 16352
rect 45770 16287 46090 16288
rect 19517 16010 19583 16013
rect 22093 16010 22159 16013
rect 19517 16008 22159 16010
rect 19517 15952 19522 16008
rect 19578 15952 22098 16008
rect 22154 15952 22159 16008
rect 19517 15950 22159 15952
rect 19517 15947 19583 15950
rect 22093 15947 22159 15950
rect 18874 15808 19194 15809
rect 18874 15744 18882 15808
rect 18946 15744 18962 15808
rect 19026 15744 19042 15808
rect 19106 15744 19122 15808
rect 19186 15744 19194 15808
rect 18874 15743 19194 15744
rect 36805 15808 37125 15809
rect 36805 15744 36813 15808
rect 36877 15744 36893 15808
rect 36957 15744 36973 15808
rect 37037 15744 37053 15808
rect 37117 15744 37125 15808
rect 36805 15743 37125 15744
rect 9765 15466 9831 15469
rect 12525 15466 12591 15469
rect 9765 15464 12591 15466
rect 9765 15408 9770 15464
rect 9826 15408 12530 15464
rect 12586 15408 12591 15464
rect 9765 15406 12591 15408
rect 9765 15403 9831 15406
rect 12525 15403 12591 15406
rect 9909 15264 10229 15265
rect 9909 15200 9917 15264
rect 9981 15200 9997 15264
rect 10061 15200 10077 15264
rect 10141 15200 10157 15264
rect 10221 15200 10229 15264
rect 9909 15199 10229 15200
rect 27840 15264 28160 15265
rect 27840 15200 27848 15264
rect 27912 15200 27928 15264
rect 27992 15200 28008 15264
rect 28072 15200 28088 15264
rect 28152 15200 28160 15264
rect 27840 15199 28160 15200
rect 45770 15264 46090 15265
rect 45770 15200 45778 15264
rect 45842 15200 45858 15264
rect 45922 15200 45938 15264
rect 46002 15200 46018 15264
rect 46082 15200 46090 15264
rect 45770 15199 46090 15200
rect 10317 15058 10383 15061
rect 13077 15058 13143 15061
rect 15377 15058 15443 15061
rect 10317 15056 15443 15058
rect 10317 15000 10322 15056
rect 10378 15000 13082 15056
rect 13138 15000 15382 15056
rect 15438 15000 15443 15056
rect 10317 14998 15443 15000
rect 10317 14995 10383 14998
rect 13077 14995 13143 14998
rect 15377 14995 15443 14998
rect 18874 14720 19194 14721
rect 18874 14656 18882 14720
rect 18946 14656 18962 14720
rect 19026 14656 19042 14720
rect 19106 14656 19122 14720
rect 19186 14656 19194 14720
rect 18874 14655 19194 14656
rect 36805 14720 37125 14721
rect 36805 14656 36813 14720
rect 36877 14656 36893 14720
rect 36957 14656 36973 14720
rect 37037 14656 37053 14720
rect 37117 14656 37125 14720
rect 36805 14655 37125 14656
rect 9909 14176 10229 14177
rect 9909 14112 9917 14176
rect 9981 14112 9997 14176
rect 10061 14112 10077 14176
rect 10141 14112 10157 14176
rect 10221 14112 10229 14176
rect 9909 14111 10229 14112
rect 27840 14176 28160 14177
rect 27840 14112 27848 14176
rect 27912 14112 27928 14176
rect 27992 14112 28008 14176
rect 28072 14112 28088 14176
rect 28152 14112 28160 14176
rect 27840 14111 28160 14112
rect 45770 14176 46090 14177
rect 45770 14112 45778 14176
rect 45842 14112 45858 14176
rect 45922 14112 45938 14176
rect 46002 14112 46018 14176
rect 46082 14112 46090 14176
rect 45770 14111 46090 14112
rect 18874 13632 19194 13633
rect 18874 13568 18882 13632
rect 18946 13568 18962 13632
rect 19026 13568 19042 13632
rect 19106 13568 19122 13632
rect 19186 13568 19194 13632
rect 18874 13567 19194 13568
rect 36805 13632 37125 13633
rect 36805 13568 36813 13632
rect 36877 13568 36893 13632
rect 36957 13568 36973 13632
rect 37037 13568 37053 13632
rect 37117 13568 37125 13632
rect 36805 13567 37125 13568
rect 9909 13088 10229 13089
rect 9909 13024 9917 13088
rect 9981 13024 9997 13088
rect 10061 13024 10077 13088
rect 10141 13024 10157 13088
rect 10221 13024 10229 13088
rect 9909 13023 10229 13024
rect 27840 13088 28160 13089
rect 27840 13024 27848 13088
rect 27912 13024 27928 13088
rect 27992 13024 28008 13088
rect 28072 13024 28088 13088
rect 28152 13024 28160 13088
rect 27840 13023 28160 13024
rect 45770 13088 46090 13089
rect 45770 13024 45778 13088
rect 45842 13024 45858 13088
rect 45922 13024 45938 13088
rect 46002 13024 46018 13088
rect 46082 13024 46090 13088
rect 45770 13023 46090 13024
rect 18874 12544 19194 12545
rect 18874 12480 18882 12544
rect 18946 12480 18962 12544
rect 19026 12480 19042 12544
rect 19106 12480 19122 12544
rect 19186 12480 19194 12544
rect 18874 12479 19194 12480
rect 36805 12544 37125 12545
rect 36805 12480 36813 12544
rect 36877 12480 36893 12544
rect 36957 12480 36973 12544
rect 37037 12480 37053 12544
rect 37117 12480 37125 12544
rect 36805 12479 37125 12480
rect 9909 12000 10229 12001
rect 9909 11936 9917 12000
rect 9981 11936 9997 12000
rect 10061 11936 10077 12000
rect 10141 11936 10157 12000
rect 10221 11936 10229 12000
rect 9909 11935 10229 11936
rect 27840 12000 28160 12001
rect 27840 11936 27848 12000
rect 27912 11936 27928 12000
rect 27992 11936 28008 12000
rect 28072 11936 28088 12000
rect 28152 11936 28160 12000
rect 27840 11935 28160 11936
rect 45770 12000 46090 12001
rect 45770 11936 45778 12000
rect 45842 11936 45858 12000
rect 45922 11936 45938 12000
rect 46002 11936 46018 12000
rect 46082 11936 46090 12000
rect 45770 11935 46090 11936
rect 18874 11456 19194 11457
rect 18874 11392 18882 11456
rect 18946 11392 18962 11456
rect 19026 11392 19042 11456
rect 19106 11392 19122 11456
rect 19186 11392 19194 11456
rect 18874 11391 19194 11392
rect 36805 11456 37125 11457
rect 36805 11392 36813 11456
rect 36877 11392 36893 11456
rect 36957 11392 36973 11456
rect 37037 11392 37053 11456
rect 37117 11392 37125 11456
rect 36805 11391 37125 11392
rect 9909 10912 10229 10913
rect 9909 10848 9917 10912
rect 9981 10848 9997 10912
rect 10061 10848 10077 10912
rect 10141 10848 10157 10912
rect 10221 10848 10229 10912
rect 9909 10847 10229 10848
rect 27840 10912 28160 10913
rect 27840 10848 27848 10912
rect 27912 10848 27928 10912
rect 27992 10848 28008 10912
rect 28072 10848 28088 10912
rect 28152 10848 28160 10912
rect 27840 10847 28160 10848
rect 45770 10912 46090 10913
rect 45770 10848 45778 10912
rect 45842 10848 45858 10912
rect 45922 10848 45938 10912
rect 46002 10848 46018 10912
rect 46082 10848 46090 10912
rect 45770 10847 46090 10848
rect 18874 10368 19194 10369
rect 18874 10304 18882 10368
rect 18946 10304 18962 10368
rect 19026 10304 19042 10368
rect 19106 10304 19122 10368
rect 19186 10304 19194 10368
rect 18874 10303 19194 10304
rect 36805 10368 37125 10369
rect 36805 10304 36813 10368
rect 36877 10304 36893 10368
rect 36957 10304 36973 10368
rect 37037 10304 37053 10368
rect 37117 10304 37125 10368
rect 36805 10303 37125 10304
rect 9909 9824 10229 9825
rect 9909 9760 9917 9824
rect 9981 9760 9997 9824
rect 10061 9760 10077 9824
rect 10141 9760 10157 9824
rect 10221 9760 10229 9824
rect 9909 9759 10229 9760
rect 27840 9824 28160 9825
rect 27840 9760 27848 9824
rect 27912 9760 27928 9824
rect 27992 9760 28008 9824
rect 28072 9760 28088 9824
rect 28152 9760 28160 9824
rect 27840 9759 28160 9760
rect 45770 9824 46090 9825
rect 45770 9760 45778 9824
rect 45842 9760 45858 9824
rect 45922 9760 45938 9824
rect 46002 9760 46018 9824
rect 46082 9760 46090 9824
rect 45770 9759 46090 9760
rect 18874 9280 19194 9281
rect 18874 9216 18882 9280
rect 18946 9216 18962 9280
rect 19026 9216 19042 9280
rect 19106 9216 19122 9280
rect 19186 9216 19194 9280
rect 18874 9215 19194 9216
rect 36805 9280 37125 9281
rect 36805 9216 36813 9280
rect 36877 9216 36893 9280
rect 36957 9216 36973 9280
rect 37037 9216 37053 9280
rect 37117 9216 37125 9280
rect 36805 9215 37125 9216
rect 11237 8938 11303 8941
rect 17033 8938 17099 8941
rect 11237 8936 17099 8938
rect 11237 8880 11242 8936
rect 11298 8880 17038 8936
rect 17094 8880 17099 8936
rect 11237 8878 17099 8880
rect 11237 8875 11303 8878
rect 17033 8875 17099 8878
rect 9909 8736 10229 8737
rect 9909 8672 9917 8736
rect 9981 8672 9997 8736
rect 10061 8672 10077 8736
rect 10141 8672 10157 8736
rect 10221 8672 10229 8736
rect 9909 8671 10229 8672
rect 27840 8736 28160 8737
rect 27840 8672 27848 8736
rect 27912 8672 27928 8736
rect 27992 8672 28008 8736
rect 28072 8672 28088 8736
rect 28152 8672 28160 8736
rect 27840 8671 28160 8672
rect 45770 8736 46090 8737
rect 45770 8672 45778 8736
rect 45842 8672 45858 8736
rect 45922 8672 45938 8736
rect 46002 8672 46018 8736
rect 46082 8672 46090 8736
rect 45770 8671 46090 8672
rect 18874 8192 19194 8193
rect 18874 8128 18882 8192
rect 18946 8128 18962 8192
rect 19026 8128 19042 8192
rect 19106 8128 19122 8192
rect 19186 8128 19194 8192
rect 18874 8127 19194 8128
rect 36805 8192 37125 8193
rect 36805 8128 36813 8192
rect 36877 8128 36893 8192
rect 36957 8128 36973 8192
rect 37037 8128 37053 8192
rect 37117 8128 37125 8192
rect 36805 8127 37125 8128
rect 9909 7648 10229 7649
rect 9909 7584 9917 7648
rect 9981 7584 9997 7648
rect 10061 7584 10077 7648
rect 10141 7584 10157 7648
rect 10221 7584 10229 7648
rect 9909 7583 10229 7584
rect 27840 7648 28160 7649
rect 27840 7584 27848 7648
rect 27912 7584 27928 7648
rect 27992 7584 28008 7648
rect 28072 7584 28088 7648
rect 28152 7584 28160 7648
rect 27840 7583 28160 7584
rect 45770 7648 46090 7649
rect 45770 7584 45778 7648
rect 45842 7584 45858 7648
rect 45922 7584 45938 7648
rect 46002 7584 46018 7648
rect 46082 7584 46090 7648
rect 45770 7583 46090 7584
rect 18874 7104 19194 7105
rect 18874 7040 18882 7104
rect 18946 7040 18962 7104
rect 19026 7040 19042 7104
rect 19106 7040 19122 7104
rect 19186 7040 19194 7104
rect 18874 7039 19194 7040
rect 36805 7104 37125 7105
rect 36805 7040 36813 7104
rect 36877 7040 36893 7104
rect 36957 7040 36973 7104
rect 37037 7040 37053 7104
rect 37117 7040 37125 7104
rect 36805 7039 37125 7040
rect 51073 6898 51139 6901
rect 55200 6898 56000 6928
rect 51073 6896 56000 6898
rect 51073 6840 51078 6896
rect 51134 6840 56000 6896
rect 51073 6838 56000 6840
rect 51073 6835 51139 6838
rect 55200 6808 56000 6838
rect 9909 6560 10229 6561
rect 9909 6496 9917 6560
rect 9981 6496 9997 6560
rect 10061 6496 10077 6560
rect 10141 6496 10157 6560
rect 10221 6496 10229 6560
rect 9909 6495 10229 6496
rect 27840 6560 28160 6561
rect 27840 6496 27848 6560
rect 27912 6496 27928 6560
rect 27992 6496 28008 6560
rect 28072 6496 28088 6560
rect 28152 6496 28160 6560
rect 27840 6495 28160 6496
rect 45770 6560 46090 6561
rect 45770 6496 45778 6560
rect 45842 6496 45858 6560
rect 45922 6496 45938 6560
rect 46002 6496 46018 6560
rect 46082 6496 46090 6560
rect 45770 6495 46090 6496
rect 18874 6016 19194 6017
rect 18874 5952 18882 6016
rect 18946 5952 18962 6016
rect 19026 5952 19042 6016
rect 19106 5952 19122 6016
rect 19186 5952 19194 6016
rect 18874 5951 19194 5952
rect 36805 6016 37125 6017
rect 36805 5952 36813 6016
rect 36877 5952 36893 6016
rect 36957 5952 36973 6016
rect 37037 5952 37053 6016
rect 37117 5952 37125 6016
rect 36805 5951 37125 5952
rect 9909 5472 10229 5473
rect 9909 5408 9917 5472
rect 9981 5408 9997 5472
rect 10061 5408 10077 5472
rect 10141 5408 10157 5472
rect 10221 5408 10229 5472
rect 9909 5407 10229 5408
rect 27840 5472 28160 5473
rect 27840 5408 27848 5472
rect 27912 5408 27928 5472
rect 27992 5408 28008 5472
rect 28072 5408 28088 5472
rect 28152 5408 28160 5472
rect 27840 5407 28160 5408
rect 45770 5472 46090 5473
rect 45770 5408 45778 5472
rect 45842 5408 45858 5472
rect 45922 5408 45938 5472
rect 46002 5408 46018 5472
rect 46082 5408 46090 5472
rect 45770 5407 46090 5408
rect 18874 4928 19194 4929
rect 18874 4864 18882 4928
rect 18946 4864 18962 4928
rect 19026 4864 19042 4928
rect 19106 4864 19122 4928
rect 19186 4864 19194 4928
rect 18874 4863 19194 4864
rect 36805 4928 37125 4929
rect 36805 4864 36813 4928
rect 36877 4864 36893 4928
rect 36957 4864 36973 4928
rect 37037 4864 37053 4928
rect 37117 4864 37125 4928
rect 36805 4863 37125 4864
rect 9909 4384 10229 4385
rect 9909 4320 9917 4384
rect 9981 4320 9997 4384
rect 10061 4320 10077 4384
rect 10141 4320 10157 4384
rect 10221 4320 10229 4384
rect 9909 4319 10229 4320
rect 27840 4384 28160 4385
rect 27840 4320 27848 4384
rect 27912 4320 27928 4384
rect 27992 4320 28008 4384
rect 28072 4320 28088 4384
rect 28152 4320 28160 4384
rect 27840 4319 28160 4320
rect 45770 4384 46090 4385
rect 45770 4320 45778 4384
rect 45842 4320 45858 4384
rect 45922 4320 45938 4384
rect 46002 4320 46018 4384
rect 46082 4320 46090 4384
rect 45770 4319 46090 4320
rect 18874 3840 19194 3841
rect 18874 3776 18882 3840
rect 18946 3776 18962 3840
rect 19026 3776 19042 3840
rect 19106 3776 19122 3840
rect 19186 3776 19194 3840
rect 18874 3775 19194 3776
rect 36805 3840 37125 3841
rect 36805 3776 36813 3840
rect 36877 3776 36893 3840
rect 36957 3776 36973 3840
rect 37037 3776 37053 3840
rect 37117 3776 37125 3840
rect 36805 3775 37125 3776
rect 9909 3296 10229 3297
rect 9909 3232 9917 3296
rect 9981 3232 9997 3296
rect 10061 3232 10077 3296
rect 10141 3232 10157 3296
rect 10221 3232 10229 3296
rect 9909 3231 10229 3232
rect 27840 3296 28160 3297
rect 27840 3232 27848 3296
rect 27912 3232 27928 3296
rect 27992 3232 28008 3296
rect 28072 3232 28088 3296
rect 28152 3232 28160 3296
rect 27840 3231 28160 3232
rect 45770 3296 46090 3297
rect 45770 3232 45778 3296
rect 45842 3232 45858 3296
rect 45922 3232 45938 3296
rect 46002 3232 46018 3296
rect 46082 3232 46090 3296
rect 45770 3231 46090 3232
rect 18874 2752 19194 2753
rect 18874 2688 18882 2752
rect 18946 2688 18962 2752
rect 19026 2688 19042 2752
rect 19106 2688 19122 2752
rect 19186 2688 19194 2752
rect 18874 2687 19194 2688
rect 36805 2752 37125 2753
rect 36805 2688 36813 2752
rect 36877 2688 36893 2752
rect 36957 2688 36973 2752
rect 37037 2688 37053 2752
rect 37117 2688 37125 2752
rect 36805 2687 37125 2688
rect 9909 2208 10229 2209
rect 9909 2144 9917 2208
rect 9981 2144 9997 2208
rect 10061 2144 10077 2208
rect 10141 2144 10157 2208
rect 10221 2144 10229 2208
rect 9909 2143 10229 2144
rect 27840 2208 28160 2209
rect 27840 2144 27848 2208
rect 27912 2144 27928 2208
rect 27992 2144 28008 2208
rect 28072 2144 28088 2208
rect 28152 2144 28160 2208
rect 27840 2143 28160 2144
rect 45770 2208 46090 2209
rect 45770 2144 45778 2208
rect 45842 2144 45858 2208
rect 45922 2144 45938 2208
rect 46002 2144 46018 2208
rect 46082 2144 46090 2208
rect 45770 2143 46090 2144
<< via3 >>
rect 9917 25052 9981 25056
rect 9917 24996 9921 25052
rect 9921 24996 9977 25052
rect 9977 24996 9981 25052
rect 9917 24992 9981 24996
rect 9997 25052 10061 25056
rect 9997 24996 10001 25052
rect 10001 24996 10057 25052
rect 10057 24996 10061 25052
rect 9997 24992 10061 24996
rect 10077 25052 10141 25056
rect 10077 24996 10081 25052
rect 10081 24996 10137 25052
rect 10137 24996 10141 25052
rect 10077 24992 10141 24996
rect 10157 25052 10221 25056
rect 10157 24996 10161 25052
rect 10161 24996 10217 25052
rect 10217 24996 10221 25052
rect 10157 24992 10221 24996
rect 27848 25052 27912 25056
rect 27848 24996 27852 25052
rect 27852 24996 27908 25052
rect 27908 24996 27912 25052
rect 27848 24992 27912 24996
rect 27928 25052 27992 25056
rect 27928 24996 27932 25052
rect 27932 24996 27988 25052
rect 27988 24996 27992 25052
rect 27928 24992 27992 24996
rect 28008 25052 28072 25056
rect 28008 24996 28012 25052
rect 28012 24996 28068 25052
rect 28068 24996 28072 25052
rect 28008 24992 28072 24996
rect 28088 25052 28152 25056
rect 28088 24996 28092 25052
rect 28092 24996 28148 25052
rect 28148 24996 28152 25052
rect 28088 24992 28152 24996
rect 45778 25052 45842 25056
rect 45778 24996 45782 25052
rect 45782 24996 45838 25052
rect 45838 24996 45842 25052
rect 45778 24992 45842 24996
rect 45858 25052 45922 25056
rect 45858 24996 45862 25052
rect 45862 24996 45918 25052
rect 45918 24996 45922 25052
rect 45858 24992 45922 24996
rect 45938 25052 46002 25056
rect 45938 24996 45942 25052
rect 45942 24996 45998 25052
rect 45998 24996 46002 25052
rect 45938 24992 46002 24996
rect 46018 25052 46082 25056
rect 46018 24996 46022 25052
rect 46022 24996 46078 25052
rect 46078 24996 46082 25052
rect 46018 24992 46082 24996
rect 18882 24508 18946 24512
rect 18882 24452 18886 24508
rect 18886 24452 18942 24508
rect 18942 24452 18946 24508
rect 18882 24448 18946 24452
rect 18962 24508 19026 24512
rect 18962 24452 18966 24508
rect 18966 24452 19022 24508
rect 19022 24452 19026 24508
rect 18962 24448 19026 24452
rect 19042 24508 19106 24512
rect 19042 24452 19046 24508
rect 19046 24452 19102 24508
rect 19102 24452 19106 24508
rect 19042 24448 19106 24452
rect 19122 24508 19186 24512
rect 19122 24452 19126 24508
rect 19126 24452 19182 24508
rect 19182 24452 19186 24508
rect 19122 24448 19186 24452
rect 36813 24508 36877 24512
rect 36813 24452 36817 24508
rect 36817 24452 36873 24508
rect 36873 24452 36877 24508
rect 36813 24448 36877 24452
rect 36893 24508 36957 24512
rect 36893 24452 36897 24508
rect 36897 24452 36953 24508
rect 36953 24452 36957 24508
rect 36893 24448 36957 24452
rect 36973 24508 37037 24512
rect 36973 24452 36977 24508
rect 36977 24452 37033 24508
rect 37033 24452 37037 24508
rect 36973 24448 37037 24452
rect 37053 24508 37117 24512
rect 37053 24452 37057 24508
rect 37057 24452 37113 24508
rect 37113 24452 37117 24508
rect 37053 24448 37117 24452
rect 9917 23964 9981 23968
rect 9917 23908 9921 23964
rect 9921 23908 9977 23964
rect 9977 23908 9981 23964
rect 9917 23904 9981 23908
rect 9997 23964 10061 23968
rect 9997 23908 10001 23964
rect 10001 23908 10057 23964
rect 10057 23908 10061 23964
rect 9997 23904 10061 23908
rect 10077 23964 10141 23968
rect 10077 23908 10081 23964
rect 10081 23908 10137 23964
rect 10137 23908 10141 23964
rect 10077 23904 10141 23908
rect 10157 23964 10221 23968
rect 10157 23908 10161 23964
rect 10161 23908 10217 23964
rect 10217 23908 10221 23964
rect 10157 23904 10221 23908
rect 27848 23964 27912 23968
rect 27848 23908 27852 23964
rect 27852 23908 27908 23964
rect 27908 23908 27912 23964
rect 27848 23904 27912 23908
rect 27928 23964 27992 23968
rect 27928 23908 27932 23964
rect 27932 23908 27988 23964
rect 27988 23908 27992 23964
rect 27928 23904 27992 23908
rect 28008 23964 28072 23968
rect 28008 23908 28012 23964
rect 28012 23908 28068 23964
rect 28068 23908 28072 23964
rect 28008 23904 28072 23908
rect 28088 23964 28152 23968
rect 28088 23908 28092 23964
rect 28092 23908 28148 23964
rect 28148 23908 28152 23964
rect 28088 23904 28152 23908
rect 45778 23964 45842 23968
rect 45778 23908 45782 23964
rect 45782 23908 45838 23964
rect 45838 23908 45842 23964
rect 45778 23904 45842 23908
rect 45858 23964 45922 23968
rect 45858 23908 45862 23964
rect 45862 23908 45918 23964
rect 45918 23908 45922 23964
rect 45858 23904 45922 23908
rect 45938 23964 46002 23968
rect 45938 23908 45942 23964
rect 45942 23908 45998 23964
rect 45998 23908 46002 23964
rect 45938 23904 46002 23908
rect 46018 23964 46082 23968
rect 46018 23908 46022 23964
rect 46022 23908 46078 23964
rect 46078 23908 46082 23964
rect 46018 23904 46082 23908
rect 18882 23420 18946 23424
rect 18882 23364 18886 23420
rect 18886 23364 18942 23420
rect 18942 23364 18946 23420
rect 18882 23360 18946 23364
rect 18962 23420 19026 23424
rect 18962 23364 18966 23420
rect 18966 23364 19022 23420
rect 19022 23364 19026 23420
rect 18962 23360 19026 23364
rect 19042 23420 19106 23424
rect 19042 23364 19046 23420
rect 19046 23364 19102 23420
rect 19102 23364 19106 23420
rect 19042 23360 19106 23364
rect 19122 23420 19186 23424
rect 19122 23364 19126 23420
rect 19126 23364 19182 23420
rect 19182 23364 19186 23420
rect 19122 23360 19186 23364
rect 36813 23420 36877 23424
rect 36813 23364 36817 23420
rect 36817 23364 36873 23420
rect 36873 23364 36877 23420
rect 36813 23360 36877 23364
rect 36893 23420 36957 23424
rect 36893 23364 36897 23420
rect 36897 23364 36953 23420
rect 36953 23364 36957 23420
rect 36893 23360 36957 23364
rect 36973 23420 37037 23424
rect 36973 23364 36977 23420
rect 36977 23364 37033 23420
rect 37033 23364 37037 23420
rect 36973 23360 37037 23364
rect 37053 23420 37117 23424
rect 37053 23364 37057 23420
rect 37057 23364 37113 23420
rect 37113 23364 37117 23420
rect 37053 23360 37117 23364
rect 9917 22876 9981 22880
rect 9917 22820 9921 22876
rect 9921 22820 9977 22876
rect 9977 22820 9981 22876
rect 9917 22816 9981 22820
rect 9997 22876 10061 22880
rect 9997 22820 10001 22876
rect 10001 22820 10057 22876
rect 10057 22820 10061 22876
rect 9997 22816 10061 22820
rect 10077 22876 10141 22880
rect 10077 22820 10081 22876
rect 10081 22820 10137 22876
rect 10137 22820 10141 22876
rect 10077 22816 10141 22820
rect 10157 22876 10221 22880
rect 10157 22820 10161 22876
rect 10161 22820 10217 22876
rect 10217 22820 10221 22876
rect 10157 22816 10221 22820
rect 27848 22876 27912 22880
rect 27848 22820 27852 22876
rect 27852 22820 27908 22876
rect 27908 22820 27912 22876
rect 27848 22816 27912 22820
rect 27928 22876 27992 22880
rect 27928 22820 27932 22876
rect 27932 22820 27988 22876
rect 27988 22820 27992 22876
rect 27928 22816 27992 22820
rect 28008 22876 28072 22880
rect 28008 22820 28012 22876
rect 28012 22820 28068 22876
rect 28068 22820 28072 22876
rect 28008 22816 28072 22820
rect 28088 22876 28152 22880
rect 28088 22820 28092 22876
rect 28092 22820 28148 22876
rect 28148 22820 28152 22876
rect 28088 22816 28152 22820
rect 45778 22876 45842 22880
rect 45778 22820 45782 22876
rect 45782 22820 45838 22876
rect 45838 22820 45842 22876
rect 45778 22816 45842 22820
rect 45858 22876 45922 22880
rect 45858 22820 45862 22876
rect 45862 22820 45918 22876
rect 45918 22820 45922 22876
rect 45858 22816 45922 22820
rect 45938 22876 46002 22880
rect 45938 22820 45942 22876
rect 45942 22820 45998 22876
rect 45998 22820 46002 22876
rect 45938 22816 46002 22820
rect 46018 22876 46082 22880
rect 46018 22820 46022 22876
rect 46022 22820 46078 22876
rect 46078 22820 46082 22876
rect 46018 22816 46082 22820
rect 18882 22332 18946 22336
rect 18882 22276 18886 22332
rect 18886 22276 18942 22332
rect 18942 22276 18946 22332
rect 18882 22272 18946 22276
rect 18962 22332 19026 22336
rect 18962 22276 18966 22332
rect 18966 22276 19022 22332
rect 19022 22276 19026 22332
rect 18962 22272 19026 22276
rect 19042 22332 19106 22336
rect 19042 22276 19046 22332
rect 19046 22276 19102 22332
rect 19102 22276 19106 22332
rect 19042 22272 19106 22276
rect 19122 22332 19186 22336
rect 19122 22276 19126 22332
rect 19126 22276 19182 22332
rect 19182 22276 19186 22332
rect 19122 22272 19186 22276
rect 36813 22332 36877 22336
rect 36813 22276 36817 22332
rect 36817 22276 36873 22332
rect 36873 22276 36877 22332
rect 36813 22272 36877 22276
rect 36893 22332 36957 22336
rect 36893 22276 36897 22332
rect 36897 22276 36953 22332
rect 36953 22276 36957 22332
rect 36893 22272 36957 22276
rect 36973 22332 37037 22336
rect 36973 22276 36977 22332
rect 36977 22276 37033 22332
rect 37033 22276 37037 22332
rect 36973 22272 37037 22276
rect 37053 22332 37117 22336
rect 37053 22276 37057 22332
rect 37057 22276 37113 22332
rect 37113 22276 37117 22332
rect 37053 22272 37117 22276
rect 9917 21788 9981 21792
rect 9917 21732 9921 21788
rect 9921 21732 9977 21788
rect 9977 21732 9981 21788
rect 9917 21728 9981 21732
rect 9997 21788 10061 21792
rect 9997 21732 10001 21788
rect 10001 21732 10057 21788
rect 10057 21732 10061 21788
rect 9997 21728 10061 21732
rect 10077 21788 10141 21792
rect 10077 21732 10081 21788
rect 10081 21732 10137 21788
rect 10137 21732 10141 21788
rect 10077 21728 10141 21732
rect 10157 21788 10221 21792
rect 10157 21732 10161 21788
rect 10161 21732 10217 21788
rect 10217 21732 10221 21788
rect 10157 21728 10221 21732
rect 27848 21788 27912 21792
rect 27848 21732 27852 21788
rect 27852 21732 27908 21788
rect 27908 21732 27912 21788
rect 27848 21728 27912 21732
rect 27928 21788 27992 21792
rect 27928 21732 27932 21788
rect 27932 21732 27988 21788
rect 27988 21732 27992 21788
rect 27928 21728 27992 21732
rect 28008 21788 28072 21792
rect 28008 21732 28012 21788
rect 28012 21732 28068 21788
rect 28068 21732 28072 21788
rect 28008 21728 28072 21732
rect 28088 21788 28152 21792
rect 28088 21732 28092 21788
rect 28092 21732 28148 21788
rect 28148 21732 28152 21788
rect 28088 21728 28152 21732
rect 45778 21788 45842 21792
rect 45778 21732 45782 21788
rect 45782 21732 45838 21788
rect 45838 21732 45842 21788
rect 45778 21728 45842 21732
rect 45858 21788 45922 21792
rect 45858 21732 45862 21788
rect 45862 21732 45918 21788
rect 45918 21732 45922 21788
rect 45858 21728 45922 21732
rect 45938 21788 46002 21792
rect 45938 21732 45942 21788
rect 45942 21732 45998 21788
rect 45998 21732 46002 21788
rect 45938 21728 46002 21732
rect 46018 21788 46082 21792
rect 46018 21732 46022 21788
rect 46022 21732 46078 21788
rect 46078 21732 46082 21788
rect 46018 21728 46082 21732
rect 18882 21244 18946 21248
rect 18882 21188 18886 21244
rect 18886 21188 18942 21244
rect 18942 21188 18946 21244
rect 18882 21184 18946 21188
rect 18962 21244 19026 21248
rect 18962 21188 18966 21244
rect 18966 21188 19022 21244
rect 19022 21188 19026 21244
rect 18962 21184 19026 21188
rect 19042 21244 19106 21248
rect 19042 21188 19046 21244
rect 19046 21188 19102 21244
rect 19102 21188 19106 21244
rect 19042 21184 19106 21188
rect 19122 21244 19186 21248
rect 19122 21188 19126 21244
rect 19126 21188 19182 21244
rect 19182 21188 19186 21244
rect 19122 21184 19186 21188
rect 36813 21244 36877 21248
rect 36813 21188 36817 21244
rect 36817 21188 36873 21244
rect 36873 21188 36877 21244
rect 36813 21184 36877 21188
rect 36893 21244 36957 21248
rect 36893 21188 36897 21244
rect 36897 21188 36953 21244
rect 36953 21188 36957 21244
rect 36893 21184 36957 21188
rect 36973 21244 37037 21248
rect 36973 21188 36977 21244
rect 36977 21188 37033 21244
rect 37033 21188 37037 21244
rect 36973 21184 37037 21188
rect 37053 21244 37117 21248
rect 37053 21188 37057 21244
rect 37057 21188 37113 21244
rect 37113 21188 37117 21244
rect 37053 21184 37117 21188
rect 9917 20700 9981 20704
rect 9917 20644 9921 20700
rect 9921 20644 9977 20700
rect 9977 20644 9981 20700
rect 9917 20640 9981 20644
rect 9997 20700 10061 20704
rect 9997 20644 10001 20700
rect 10001 20644 10057 20700
rect 10057 20644 10061 20700
rect 9997 20640 10061 20644
rect 10077 20700 10141 20704
rect 10077 20644 10081 20700
rect 10081 20644 10137 20700
rect 10137 20644 10141 20700
rect 10077 20640 10141 20644
rect 10157 20700 10221 20704
rect 10157 20644 10161 20700
rect 10161 20644 10217 20700
rect 10217 20644 10221 20700
rect 10157 20640 10221 20644
rect 27848 20700 27912 20704
rect 27848 20644 27852 20700
rect 27852 20644 27908 20700
rect 27908 20644 27912 20700
rect 27848 20640 27912 20644
rect 27928 20700 27992 20704
rect 27928 20644 27932 20700
rect 27932 20644 27988 20700
rect 27988 20644 27992 20700
rect 27928 20640 27992 20644
rect 28008 20700 28072 20704
rect 28008 20644 28012 20700
rect 28012 20644 28068 20700
rect 28068 20644 28072 20700
rect 28008 20640 28072 20644
rect 28088 20700 28152 20704
rect 28088 20644 28092 20700
rect 28092 20644 28148 20700
rect 28148 20644 28152 20700
rect 28088 20640 28152 20644
rect 45778 20700 45842 20704
rect 45778 20644 45782 20700
rect 45782 20644 45838 20700
rect 45838 20644 45842 20700
rect 45778 20640 45842 20644
rect 45858 20700 45922 20704
rect 45858 20644 45862 20700
rect 45862 20644 45918 20700
rect 45918 20644 45922 20700
rect 45858 20640 45922 20644
rect 45938 20700 46002 20704
rect 45938 20644 45942 20700
rect 45942 20644 45998 20700
rect 45998 20644 46002 20700
rect 45938 20640 46002 20644
rect 46018 20700 46082 20704
rect 46018 20644 46022 20700
rect 46022 20644 46078 20700
rect 46078 20644 46082 20700
rect 46018 20640 46082 20644
rect 18882 20156 18946 20160
rect 18882 20100 18886 20156
rect 18886 20100 18942 20156
rect 18942 20100 18946 20156
rect 18882 20096 18946 20100
rect 18962 20156 19026 20160
rect 18962 20100 18966 20156
rect 18966 20100 19022 20156
rect 19022 20100 19026 20156
rect 18962 20096 19026 20100
rect 19042 20156 19106 20160
rect 19042 20100 19046 20156
rect 19046 20100 19102 20156
rect 19102 20100 19106 20156
rect 19042 20096 19106 20100
rect 19122 20156 19186 20160
rect 19122 20100 19126 20156
rect 19126 20100 19182 20156
rect 19182 20100 19186 20156
rect 19122 20096 19186 20100
rect 36813 20156 36877 20160
rect 36813 20100 36817 20156
rect 36817 20100 36873 20156
rect 36873 20100 36877 20156
rect 36813 20096 36877 20100
rect 36893 20156 36957 20160
rect 36893 20100 36897 20156
rect 36897 20100 36953 20156
rect 36953 20100 36957 20156
rect 36893 20096 36957 20100
rect 36973 20156 37037 20160
rect 36973 20100 36977 20156
rect 36977 20100 37033 20156
rect 37033 20100 37037 20156
rect 36973 20096 37037 20100
rect 37053 20156 37117 20160
rect 37053 20100 37057 20156
rect 37057 20100 37113 20156
rect 37113 20100 37117 20156
rect 37053 20096 37117 20100
rect 9917 19612 9981 19616
rect 9917 19556 9921 19612
rect 9921 19556 9977 19612
rect 9977 19556 9981 19612
rect 9917 19552 9981 19556
rect 9997 19612 10061 19616
rect 9997 19556 10001 19612
rect 10001 19556 10057 19612
rect 10057 19556 10061 19612
rect 9997 19552 10061 19556
rect 10077 19612 10141 19616
rect 10077 19556 10081 19612
rect 10081 19556 10137 19612
rect 10137 19556 10141 19612
rect 10077 19552 10141 19556
rect 10157 19612 10221 19616
rect 10157 19556 10161 19612
rect 10161 19556 10217 19612
rect 10217 19556 10221 19612
rect 10157 19552 10221 19556
rect 27848 19612 27912 19616
rect 27848 19556 27852 19612
rect 27852 19556 27908 19612
rect 27908 19556 27912 19612
rect 27848 19552 27912 19556
rect 27928 19612 27992 19616
rect 27928 19556 27932 19612
rect 27932 19556 27988 19612
rect 27988 19556 27992 19612
rect 27928 19552 27992 19556
rect 28008 19612 28072 19616
rect 28008 19556 28012 19612
rect 28012 19556 28068 19612
rect 28068 19556 28072 19612
rect 28008 19552 28072 19556
rect 28088 19612 28152 19616
rect 28088 19556 28092 19612
rect 28092 19556 28148 19612
rect 28148 19556 28152 19612
rect 28088 19552 28152 19556
rect 45778 19612 45842 19616
rect 45778 19556 45782 19612
rect 45782 19556 45838 19612
rect 45838 19556 45842 19612
rect 45778 19552 45842 19556
rect 45858 19612 45922 19616
rect 45858 19556 45862 19612
rect 45862 19556 45918 19612
rect 45918 19556 45922 19612
rect 45858 19552 45922 19556
rect 45938 19612 46002 19616
rect 45938 19556 45942 19612
rect 45942 19556 45998 19612
rect 45998 19556 46002 19612
rect 45938 19552 46002 19556
rect 46018 19612 46082 19616
rect 46018 19556 46022 19612
rect 46022 19556 46078 19612
rect 46078 19556 46082 19612
rect 46018 19552 46082 19556
rect 18882 19068 18946 19072
rect 18882 19012 18886 19068
rect 18886 19012 18942 19068
rect 18942 19012 18946 19068
rect 18882 19008 18946 19012
rect 18962 19068 19026 19072
rect 18962 19012 18966 19068
rect 18966 19012 19022 19068
rect 19022 19012 19026 19068
rect 18962 19008 19026 19012
rect 19042 19068 19106 19072
rect 19042 19012 19046 19068
rect 19046 19012 19102 19068
rect 19102 19012 19106 19068
rect 19042 19008 19106 19012
rect 19122 19068 19186 19072
rect 19122 19012 19126 19068
rect 19126 19012 19182 19068
rect 19182 19012 19186 19068
rect 19122 19008 19186 19012
rect 36813 19068 36877 19072
rect 36813 19012 36817 19068
rect 36817 19012 36873 19068
rect 36873 19012 36877 19068
rect 36813 19008 36877 19012
rect 36893 19068 36957 19072
rect 36893 19012 36897 19068
rect 36897 19012 36953 19068
rect 36953 19012 36957 19068
rect 36893 19008 36957 19012
rect 36973 19068 37037 19072
rect 36973 19012 36977 19068
rect 36977 19012 37033 19068
rect 37033 19012 37037 19068
rect 36973 19008 37037 19012
rect 37053 19068 37117 19072
rect 37053 19012 37057 19068
rect 37057 19012 37113 19068
rect 37113 19012 37117 19068
rect 37053 19008 37117 19012
rect 9917 18524 9981 18528
rect 9917 18468 9921 18524
rect 9921 18468 9977 18524
rect 9977 18468 9981 18524
rect 9917 18464 9981 18468
rect 9997 18524 10061 18528
rect 9997 18468 10001 18524
rect 10001 18468 10057 18524
rect 10057 18468 10061 18524
rect 9997 18464 10061 18468
rect 10077 18524 10141 18528
rect 10077 18468 10081 18524
rect 10081 18468 10137 18524
rect 10137 18468 10141 18524
rect 10077 18464 10141 18468
rect 10157 18524 10221 18528
rect 10157 18468 10161 18524
rect 10161 18468 10217 18524
rect 10217 18468 10221 18524
rect 10157 18464 10221 18468
rect 27848 18524 27912 18528
rect 27848 18468 27852 18524
rect 27852 18468 27908 18524
rect 27908 18468 27912 18524
rect 27848 18464 27912 18468
rect 27928 18524 27992 18528
rect 27928 18468 27932 18524
rect 27932 18468 27988 18524
rect 27988 18468 27992 18524
rect 27928 18464 27992 18468
rect 28008 18524 28072 18528
rect 28008 18468 28012 18524
rect 28012 18468 28068 18524
rect 28068 18468 28072 18524
rect 28008 18464 28072 18468
rect 28088 18524 28152 18528
rect 28088 18468 28092 18524
rect 28092 18468 28148 18524
rect 28148 18468 28152 18524
rect 28088 18464 28152 18468
rect 45778 18524 45842 18528
rect 45778 18468 45782 18524
rect 45782 18468 45838 18524
rect 45838 18468 45842 18524
rect 45778 18464 45842 18468
rect 45858 18524 45922 18528
rect 45858 18468 45862 18524
rect 45862 18468 45918 18524
rect 45918 18468 45922 18524
rect 45858 18464 45922 18468
rect 45938 18524 46002 18528
rect 45938 18468 45942 18524
rect 45942 18468 45998 18524
rect 45998 18468 46002 18524
rect 45938 18464 46002 18468
rect 46018 18524 46082 18528
rect 46018 18468 46022 18524
rect 46022 18468 46078 18524
rect 46078 18468 46082 18524
rect 46018 18464 46082 18468
rect 18882 17980 18946 17984
rect 18882 17924 18886 17980
rect 18886 17924 18942 17980
rect 18942 17924 18946 17980
rect 18882 17920 18946 17924
rect 18962 17980 19026 17984
rect 18962 17924 18966 17980
rect 18966 17924 19022 17980
rect 19022 17924 19026 17980
rect 18962 17920 19026 17924
rect 19042 17980 19106 17984
rect 19042 17924 19046 17980
rect 19046 17924 19102 17980
rect 19102 17924 19106 17980
rect 19042 17920 19106 17924
rect 19122 17980 19186 17984
rect 19122 17924 19126 17980
rect 19126 17924 19182 17980
rect 19182 17924 19186 17980
rect 19122 17920 19186 17924
rect 36813 17980 36877 17984
rect 36813 17924 36817 17980
rect 36817 17924 36873 17980
rect 36873 17924 36877 17980
rect 36813 17920 36877 17924
rect 36893 17980 36957 17984
rect 36893 17924 36897 17980
rect 36897 17924 36953 17980
rect 36953 17924 36957 17980
rect 36893 17920 36957 17924
rect 36973 17980 37037 17984
rect 36973 17924 36977 17980
rect 36977 17924 37033 17980
rect 37033 17924 37037 17980
rect 36973 17920 37037 17924
rect 37053 17980 37117 17984
rect 37053 17924 37057 17980
rect 37057 17924 37113 17980
rect 37113 17924 37117 17980
rect 37053 17920 37117 17924
rect 9917 17436 9981 17440
rect 9917 17380 9921 17436
rect 9921 17380 9977 17436
rect 9977 17380 9981 17436
rect 9917 17376 9981 17380
rect 9997 17436 10061 17440
rect 9997 17380 10001 17436
rect 10001 17380 10057 17436
rect 10057 17380 10061 17436
rect 9997 17376 10061 17380
rect 10077 17436 10141 17440
rect 10077 17380 10081 17436
rect 10081 17380 10137 17436
rect 10137 17380 10141 17436
rect 10077 17376 10141 17380
rect 10157 17436 10221 17440
rect 10157 17380 10161 17436
rect 10161 17380 10217 17436
rect 10217 17380 10221 17436
rect 10157 17376 10221 17380
rect 27848 17436 27912 17440
rect 27848 17380 27852 17436
rect 27852 17380 27908 17436
rect 27908 17380 27912 17436
rect 27848 17376 27912 17380
rect 27928 17436 27992 17440
rect 27928 17380 27932 17436
rect 27932 17380 27988 17436
rect 27988 17380 27992 17436
rect 27928 17376 27992 17380
rect 28008 17436 28072 17440
rect 28008 17380 28012 17436
rect 28012 17380 28068 17436
rect 28068 17380 28072 17436
rect 28008 17376 28072 17380
rect 28088 17436 28152 17440
rect 28088 17380 28092 17436
rect 28092 17380 28148 17436
rect 28148 17380 28152 17436
rect 28088 17376 28152 17380
rect 45778 17436 45842 17440
rect 45778 17380 45782 17436
rect 45782 17380 45838 17436
rect 45838 17380 45842 17436
rect 45778 17376 45842 17380
rect 45858 17436 45922 17440
rect 45858 17380 45862 17436
rect 45862 17380 45918 17436
rect 45918 17380 45922 17436
rect 45858 17376 45922 17380
rect 45938 17436 46002 17440
rect 45938 17380 45942 17436
rect 45942 17380 45998 17436
rect 45998 17380 46002 17436
rect 45938 17376 46002 17380
rect 46018 17436 46082 17440
rect 46018 17380 46022 17436
rect 46022 17380 46078 17436
rect 46078 17380 46082 17436
rect 46018 17376 46082 17380
rect 18882 16892 18946 16896
rect 18882 16836 18886 16892
rect 18886 16836 18942 16892
rect 18942 16836 18946 16892
rect 18882 16832 18946 16836
rect 18962 16892 19026 16896
rect 18962 16836 18966 16892
rect 18966 16836 19022 16892
rect 19022 16836 19026 16892
rect 18962 16832 19026 16836
rect 19042 16892 19106 16896
rect 19042 16836 19046 16892
rect 19046 16836 19102 16892
rect 19102 16836 19106 16892
rect 19042 16832 19106 16836
rect 19122 16892 19186 16896
rect 19122 16836 19126 16892
rect 19126 16836 19182 16892
rect 19182 16836 19186 16892
rect 19122 16832 19186 16836
rect 36813 16892 36877 16896
rect 36813 16836 36817 16892
rect 36817 16836 36873 16892
rect 36873 16836 36877 16892
rect 36813 16832 36877 16836
rect 36893 16892 36957 16896
rect 36893 16836 36897 16892
rect 36897 16836 36953 16892
rect 36953 16836 36957 16892
rect 36893 16832 36957 16836
rect 36973 16892 37037 16896
rect 36973 16836 36977 16892
rect 36977 16836 37033 16892
rect 37033 16836 37037 16892
rect 36973 16832 37037 16836
rect 37053 16892 37117 16896
rect 37053 16836 37057 16892
rect 37057 16836 37113 16892
rect 37113 16836 37117 16892
rect 37053 16832 37117 16836
rect 9917 16348 9981 16352
rect 9917 16292 9921 16348
rect 9921 16292 9977 16348
rect 9977 16292 9981 16348
rect 9917 16288 9981 16292
rect 9997 16348 10061 16352
rect 9997 16292 10001 16348
rect 10001 16292 10057 16348
rect 10057 16292 10061 16348
rect 9997 16288 10061 16292
rect 10077 16348 10141 16352
rect 10077 16292 10081 16348
rect 10081 16292 10137 16348
rect 10137 16292 10141 16348
rect 10077 16288 10141 16292
rect 10157 16348 10221 16352
rect 10157 16292 10161 16348
rect 10161 16292 10217 16348
rect 10217 16292 10221 16348
rect 10157 16288 10221 16292
rect 27848 16348 27912 16352
rect 27848 16292 27852 16348
rect 27852 16292 27908 16348
rect 27908 16292 27912 16348
rect 27848 16288 27912 16292
rect 27928 16348 27992 16352
rect 27928 16292 27932 16348
rect 27932 16292 27988 16348
rect 27988 16292 27992 16348
rect 27928 16288 27992 16292
rect 28008 16348 28072 16352
rect 28008 16292 28012 16348
rect 28012 16292 28068 16348
rect 28068 16292 28072 16348
rect 28008 16288 28072 16292
rect 28088 16348 28152 16352
rect 28088 16292 28092 16348
rect 28092 16292 28148 16348
rect 28148 16292 28152 16348
rect 28088 16288 28152 16292
rect 45778 16348 45842 16352
rect 45778 16292 45782 16348
rect 45782 16292 45838 16348
rect 45838 16292 45842 16348
rect 45778 16288 45842 16292
rect 45858 16348 45922 16352
rect 45858 16292 45862 16348
rect 45862 16292 45918 16348
rect 45918 16292 45922 16348
rect 45858 16288 45922 16292
rect 45938 16348 46002 16352
rect 45938 16292 45942 16348
rect 45942 16292 45998 16348
rect 45998 16292 46002 16348
rect 45938 16288 46002 16292
rect 46018 16348 46082 16352
rect 46018 16292 46022 16348
rect 46022 16292 46078 16348
rect 46078 16292 46082 16348
rect 46018 16288 46082 16292
rect 18882 15804 18946 15808
rect 18882 15748 18886 15804
rect 18886 15748 18942 15804
rect 18942 15748 18946 15804
rect 18882 15744 18946 15748
rect 18962 15804 19026 15808
rect 18962 15748 18966 15804
rect 18966 15748 19022 15804
rect 19022 15748 19026 15804
rect 18962 15744 19026 15748
rect 19042 15804 19106 15808
rect 19042 15748 19046 15804
rect 19046 15748 19102 15804
rect 19102 15748 19106 15804
rect 19042 15744 19106 15748
rect 19122 15804 19186 15808
rect 19122 15748 19126 15804
rect 19126 15748 19182 15804
rect 19182 15748 19186 15804
rect 19122 15744 19186 15748
rect 36813 15804 36877 15808
rect 36813 15748 36817 15804
rect 36817 15748 36873 15804
rect 36873 15748 36877 15804
rect 36813 15744 36877 15748
rect 36893 15804 36957 15808
rect 36893 15748 36897 15804
rect 36897 15748 36953 15804
rect 36953 15748 36957 15804
rect 36893 15744 36957 15748
rect 36973 15804 37037 15808
rect 36973 15748 36977 15804
rect 36977 15748 37033 15804
rect 37033 15748 37037 15804
rect 36973 15744 37037 15748
rect 37053 15804 37117 15808
rect 37053 15748 37057 15804
rect 37057 15748 37113 15804
rect 37113 15748 37117 15804
rect 37053 15744 37117 15748
rect 9917 15260 9981 15264
rect 9917 15204 9921 15260
rect 9921 15204 9977 15260
rect 9977 15204 9981 15260
rect 9917 15200 9981 15204
rect 9997 15260 10061 15264
rect 9997 15204 10001 15260
rect 10001 15204 10057 15260
rect 10057 15204 10061 15260
rect 9997 15200 10061 15204
rect 10077 15260 10141 15264
rect 10077 15204 10081 15260
rect 10081 15204 10137 15260
rect 10137 15204 10141 15260
rect 10077 15200 10141 15204
rect 10157 15260 10221 15264
rect 10157 15204 10161 15260
rect 10161 15204 10217 15260
rect 10217 15204 10221 15260
rect 10157 15200 10221 15204
rect 27848 15260 27912 15264
rect 27848 15204 27852 15260
rect 27852 15204 27908 15260
rect 27908 15204 27912 15260
rect 27848 15200 27912 15204
rect 27928 15260 27992 15264
rect 27928 15204 27932 15260
rect 27932 15204 27988 15260
rect 27988 15204 27992 15260
rect 27928 15200 27992 15204
rect 28008 15260 28072 15264
rect 28008 15204 28012 15260
rect 28012 15204 28068 15260
rect 28068 15204 28072 15260
rect 28008 15200 28072 15204
rect 28088 15260 28152 15264
rect 28088 15204 28092 15260
rect 28092 15204 28148 15260
rect 28148 15204 28152 15260
rect 28088 15200 28152 15204
rect 45778 15260 45842 15264
rect 45778 15204 45782 15260
rect 45782 15204 45838 15260
rect 45838 15204 45842 15260
rect 45778 15200 45842 15204
rect 45858 15260 45922 15264
rect 45858 15204 45862 15260
rect 45862 15204 45918 15260
rect 45918 15204 45922 15260
rect 45858 15200 45922 15204
rect 45938 15260 46002 15264
rect 45938 15204 45942 15260
rect 45942 15204 45998 15260
rect 45998 15204 46002 15260
rect 45938 15200 46002 15204
rect 46018 15260 46082 15264
rect 46018 15204 46022 15260
rect 46022 15204 46078 15260
rect 46078 15204 46082 15260
rect 46018 15200 46082 15204
rect 18882 14716 18946 14720
rect 18882 14660 18886 14716
rect 18886 14660 18942 14716
rect 18942 14660 18946 14716
rect 18882 14656 18946 14660
rect 18962 14716 19026 14720
rect 18962 14660 18966 14716
rect 18966 14660 19022 14716
rect 19022 14660 19026 14716
rect 18962 14656 19026 14660
rect 19042 14716 19106 14720
rect 19042 14660 19046 14716
rect 19046 14660 19102 14716
rect 19102 14660 19106 14716
rect 19042 14656 19106 14660
rect 19122 14716 19186 14720
rect 19122 14660 19126 14716
rect 19126 14660 19182 14716
rect 19182 14660 19186 14716
rect 19122 14656 19186 14660
rect 36813 14716 36877 14720
rect 36813 14660 36817 14716
rect 36817 14660 36873 14716
rect 36873 14660 36877 14716
rect 36813 14656 36877 14660
rect 36893 14716 36957 14720
rect 36893 14660 36897 14716
rect 36897 14660 36953 14716
rect 36953 14660 36957 14716
rect 36893 14656 36957 14660
rect 36973 14716 37037 14720
rect 36973 14660 36977 14716
rect 36977 14660 37033 14716
rect 37033 14660 37037 14716
rect 36973 14656 37037 14660
rect 37053 14716 37117 14720
rect 37053 14660 37057 14716
rect 37057 14660 37113 14716
rect 37113 14660 37117 14716
rect 37053 14656 37117 14660
rect 9917 14172 9981 14176
rect 9917 14116 9921 14172
rect 9921 14116 9977 14172
rect 9977 14116 9981 14172
rect 9917 14112 9981 14116
rect 9997 14172 10061 14176
rect 9997 14116 10001 14172
rect 10001 14116 10057 14172
rect 10057 14116 10061 14172
rect 9997 14112 10061 14116
rect 10077 14172 10141 14176
rect 10077 14116 10081 14172
rect 10081 14116 10137 14172
rect 10137 14116 10141 14172
rect 10077 14112 10141 14116
rect 10157 14172 10221 14176
rect 10157 14116 10161 14172
rect 10161 14116 10217 14172
rect 10217 14116 10221 14172
rect 10157 14112 10221 14116
rect 27848 14172 27912 14176
rect 27848 14116 27852 14172
rect 27852 14116 27908 14172
rect 27908 14116 27912 14172
rect 27848 14112 27912 14116
rect 27928 14172 27992 14176
rect 27928 14116 27932 14172
rect 27932 14116 27988 14172
rect 27988 14116 27992 14172
rect 27928 14112 27992 14116
rect 28008 14172 28072 14176
rect 28008 14116 28012 14172
rect 28012 14116 28068 14172
rect 28068 14116 28072 14172
rect 28008 14112 28072 14116
rect 28088 14172 28152 14176
rect 28088 14116 28092 14172
rect 28092 14116 28148 14172
rect 28148 14116 28152 14172
rect 28088 14112 28152 14116
rect 45778 14172 45842 14176
rect 45778 14116 45782 14172
rect 45782 14116 45838 14172
rect 45838 14116 45842 14172
rect 45778 14112 45842 14116
rect 45858 14172 45922 14176
rect 45858 14116 45862 14172
rect 45862 14116 45918 14172
rect 45918 14116 45922 14172
rect 45858 14112 45922 14116
rect 45938 14172 46002 14176
rect 45938 14116 45942 14172
rect 45942 14116 45998 14172
rect 45998 14116 46002 14172
rect 45938 14112 46002 14116
rect 46018 14172 46082 14176
rect 46018 14116 46022 14172
rect 46022 14116 46078 14172
rect 46078 14116 46082 14172
rect 46018 14112 46082 14116
rect 18882 13628 18946 13632
rect 18882 13572 18886 13628
rect 18886 13572 18942 13628
rect 18942 13572 18946 13628
rect 18882 13568 18946 13572
rect 18962 13628 19026 13632
rect 18962 13572 18966 13628
rect 18966 13572 19022 13628
rect 19022 13572 19026 13628
rect 18962 13568 19026 13572
rect 19042 13628 19106 13632
rect 19042 13572 19046 13628
rect 19046 13572 19102 13628
rect 19102 13572 19106 13628
rect 19042 13568 19106 13572
rect 19122 13628 19186 13632
rect 19122 13572 19126 13628
rect 19126 13572 19182 13628
rect 19182 13572 19186 13628
rect 19122 13568 19186 13572
rect 36813 13628 36877 13632
rect 36813 13572 36817 13628
rect 36817 13572 36873 13628
rect 36873 13572 36877 13628
rect 36813 13568 36877 13572
rect 36893 13628 36957 13632
rect 36893 13572 36897 13628
rect 36897 13572 36953 13628
rect 36953 13572 36957 13628
rect 36893 13568 36957 13572
rect 36973 13628 37037 13632
rect 36973 13572 36977 13628
rect 36977 13572 37033 13628
rect 37033 13572 37037 13628
rect 36973 13568 37037 13572
rect 37053 13628 37117 13632
rect 37053 13572 37057 13628
rect 37057 13572 37113 13628
rect 37113 13572 37117 13628
rect 37053 13568 37117 13572
rect 9917 13084 9981 13088
rect 9917 13028 9921 13084
rect 9921 13028 9977 13084
rect 9977 13028 9981 13084
rect 9917 13024 9981 13028
rect 9997 13084 10061 13088
rect 9997 13028 10001 13084
rect 10001 13028 10057 13084
rect 10057 13028 10061 13084
rect 9997 13024 10061 13028
rect 10077 13084 10141 13088
rect 10077 13028 10081 13084
rect 10081 13028 10137 13084
rect 10137 13028 10141 13084
rect 10077 13024 10141 13028
rect 10157 13084 10221 13088
rect 10157 13028 10161 13084
rect 10161 13028 10217 13084
rect 10217 13028 10221 13084
rect 10157 13024 10221 13028
rect 27848 13084 27912 13088
rect 27848 13028 27852 13084
rect 27852 13028 27908 13084
rect 27908 13028 27912 13084
rect 27848 13024 27912 13028
rect 27928 13084 27992 13088
rect 27928 13028 27932 13084
rect 27932 13028 27988 13084
rect 27988 13028 27992 13084
rect 27928 13024 27992 13028
rect 28008 13084 28072 13088
rect 28008 13028 28012 13084
rect 28012 13028 28068 13084
rect 28068 13028 28072 13084
rect 28008 13024 28072 13028
rect 28088 13084 28152 13088
rect 28088 13028 28092 13084
rect 28092 13028 28148 13084
rect 28148 13028 28152 13084
rect 28088 13024 28152 13028
rect 45778 13084 45842 13088
rect 45778 13028 45782 13084
rect 45782 13028 45838 13084
rect 45838 13028 45842 13084
rect 45778 13024 45842 13028
rect 45858 13084 45922 13088
rect 45858 13028 45862 13084
rect 45862 13028 45918 13084
rect 45918 13028 45922 13084
rect 45858 13024 45922 13028
rect 45938 13084 46002 13088
rect 45938 13028 45942 13084
rect 45942 13028 45998 13084
rect 45998 13028 46002 13084
rect 45938 13024 46002 13028
rect 46018 13084 46082 13088
rect 46018 13028 46022 13084
rect 46022 13028 46078 13084
rect 46078 13028 46082 13084
rect 46018 13024 46082 13028
rect 18882 12540 18946 12544
rect 18882 12484 18886 12540
rect 18886 12484 18942 12540
rect 18942 12484 18946 12540
rect 18882 12480 18946 12484
rect 18962 12540 19026 12544
rect 18962 12484 18966 12540
rect 18966 12484 19022 12540
rect 19022 12484 19026 12540
rect 18962 12480 19026 12484
rect 19042 12540 19106 12544
rect 19042 12484 19046 12540
rect 19046 12484 19102 12540
rect 19102 12484 19106 12540
rect 19042 12480 19106 12484
rect 19122 12540 19186 12544
rect 19122 12484 19126 12540
rect 19126 12484 19182 12540
rect 19182 12484 19186 12540
rect 19122 12480 19186 12484
rect 36813 12540 36877 12544
rect 36813 12484 36817 12540
rect 36817 12484 36873 12540
rect 36873 12484 36877 12540
rect 36813 12480 36877 12484
rect 36893 12540 36957 12544
rect 36893 12484 36897 12540
rect 36897 12484 36953 12540
rect 36953 12484 36957 12540
rect 36893 12480 36957 12484
rect 36973 12540 37037 12544
rect 36973 12484 36977 12540
rect 36977 12484 37033 12540
rect 37033 12484 37037 12540
rect 36973 12480 37037 12484
rect 37053 12540 37117 12544
rect 37053 12484 37057 12540
rect 37057 12484 37113 12540
rect 37113 12484 37117 12540
rect 37053 12480 37117 12484
rect 9917 11996 9981 12000
rect 9917 11940 9921 11996
rect 9921 11940 9977 11996
rect 9977 11940 9981 11996
rect 9917 11936 9981 11940
rect 9997 11996 10061 12000
rect 9997 11940 10001 11996
rect 10001 11940 10057 11996
rect 10057 11940 10061 11996
rect 9997 11936 10061 11940
rect 10077 11996 10141 12000
rect 10077 11940 10081 11996
rect 10081 11940 10137 11996
rect 10137 11940 10141 11996
rect 10077 11936 10141 11940
rect 10157 11996 10221 12000
rect 10157 11940 10161 11996
rect 10161 11940 10217 11996
rect 10217 11940 10221 11996
rect 10157 11936 10221 11940
rect 27848 11996 27912 12000
rect 27848 11940 27852 11996
rect 27852 11940 27908 11996
rect 27908 11940 27912 11996
rect 27848 11936 27912 11940
rect 27928 11996 27992 12000
rect 27928 11940 27932 11996
rect 27932 11940 27988 11996
rect 27988 11940 27992 11996
rect 27928 11936 27992 11940
rect 28008 11996 28072 12000
rect 28008 11940 28012 11996
rect 28012 11940 28068 11996
rect 28068 11940 28072 11996
rect 28008 11936 28072 11940
rect 28088 11996 28152 12000
rect 28088 11940 28092 11996
rect 28092 11940 28148 11996
rect 28148 11940 28152 11996
rect 28088 11936 28152 11940
rect 45778 11996 45842 12000
rect 45778 11940 45782 11996
rect 45782 11940 45838 11996
rect 45838 11940 45842 11996
rect 45778 11936 45842 11940
rect 45858 11996 45922 12000
rect 45858 11940 45862 11996
rect 45862 11940 45918 11996
rect 45918 11940 45922 11996
rect 45858 11936 45922 11940
rect 45938 11996 46002 12000
rect 45938 11940 45942 11996
rect 45942 11940 45998 11996
rect 45998 11940 46002 11996
rect 45938 11936 46002 11940
rect 46018 11996 46082 12000
rect 46018 11940 46022 11996
rect 46022 11940 46078 11996
rect 46078 11940 46082 11996
rect 46018 11936 46082 11940
rect 18882 11452 18946 11456
rect 18882 11396 18886 11452
rect 18886 11396 18942 11452
rect 18942 11396 18946 11452
rect 18882 11392 18946 11396
rect 18962 11452 19026 11456
rect 18962 11396 18966 11452
rect 18966 11396 19022 11452
rect 19022 11396 19026 11452
rect 18962 11392 19026 11396
rect 19042 11452 19106 11456
rect 19042 11396 19046 11452
rect 19046 11396 19102 11452
rect 19102 11396 19106 11452
rect 19042 11392 19106 11396
rect 19122 11452 19186 11456
rect 19122 11396 19126 11452
rect 19126 11396 19182 11452
rect 19182 11396 19186 11452
rect 19122 11392 19186 11396
rect 36813 11452 36877 11456
rect 36813 11396 36817 11452
rect 36817 11396 36873 11452
rect 36873 11396 36877 11452
rect 36813 11392 36877 11396
rect 36893 11452 36957 11456
rect 36893 11396 36897 11452
rect 36897 11396 36953 11452
rect 36953 11396 36957 11452
rect 36893 11392 36957 11396
rect 36973 11452 37037 11456
rect 36973 11396 36977 11452
rect 36977 11396 37033 11452
rect 37033 11396 37037 11452
rect 36973 11392 37037 11396
rect 37053 11452 37117 11456
rect 37053 11396 37057 11452
rect 37057 11396 37113 11452
rect 37113 11396 37117 11452
rect 37053 11392 37117 11396
rect 9917 10908 9981 10912
rect 9917 10852 9921 10908
rect 9921 10852 9977 10908
rect 9977 10852 9981 10908
rect 9917 10848 9981 10852
rect 9997 10908 10061 10912
rect 9997 10852 10001 10908
rect 10001 10852 10057 10908
rect 10057 10852 10061 10908
rect 9997 10848 10061 10852
rect 10077 10908 10141 10912
rect 10077 10852 10081 10908
rect 10081 10852 10137 10908
rect 10137 10852 10141 10908
rect 10077 10848 10141 10852
rect 10157 10908 10221 10912
rect 10157 10852 10161 10908
rect 10161 10852 10217 10908
rect 10217 10852 10221 10908
rect 10157 10848 10221 10852
rect 27848 10908 27912 10912
rect 27848 10852 27852 10908
rect 27852 10852 27908 10908
rect 27908 10852 27912 10908
rect 27848 10848 27912 10852
rect 27928 10908 27992 10912
rect 27928 10852 27932 10908
rect 27932 10852 27988 10908
rect 27988 10852 27992 10908
rect 27928 10848 27992 10852
rect 28008 10908 28072 10912
rect 28008 10852 28012 10908
rect 28012 10852 28068 10908
rect 28068 10852 28072 10908
rect 28008 10848 28072 10852
rect 28088 10908 28152 10912
rect 28088 10852 28092 10908
rect 28092 10852 28148 10908
rect 28148 10852 28152 10908
rect 28088 10848 28152 10852
rect 45778 10908 45842 10912
rect 45778 10852 45782 10908
rect 45782 10852 45838 10908
rect 45838 10852 45842 10908
rect 45778 10848 45842 10852
rect 45858 10908 45922 10912
rect 45858 10852 45862 10908
rect 45862 10852 45918 10908
rect 45918 10852 45922 10908
rect 45858 10848 45922 10852
rect 45938 10908 46002 10912
rect 45938 10852 45942 10908
rect 45942 10852 45998 10908
rect 45998 10852 46002 10908
rect 45938 10848 46002 10852
rect 46018 10908 46082 10912
rect 46018 10852 46022 10908
rect 46022 10852 46078 10908
rect 46078 10852 46082 10908
rect 46018 10848 46082 10852
rect 18882 10364 18946 10368
rect 18882 10308 18886 10364
rect 18886 10308 18942 10364
rect 18942 10308 18946 10364
rect 18882 10304 18946 10308
rect 18962 10364 19026 10368
rect 18962 10308 18966 10364
rect 18966 10308 19022 10364
rect 19022 10308 19026 10364
rect 18962 10304 19026 10308
rect 19042 10364 19106 10368
rect 19042 10308 19046 10364
rect 19046 10308 19102 10364
rect 19102 10308 19106 10364
rect 19042 10304 19106 10308
rect 19122 10364 19186 10368
rect 19122 10308 19126 10364
rect 19126 10308 19182 10364
rect 19182 10308 19186 10364
rect 19122 10304 19186 10308
rect 36813 10364 36877 10368
rect 36813 10308 36817 10364
rect 36817 10308 36873 10364
rect 36873 10308 36877 10364
rect 36813 10304 36877 10308
rect 36893 10364 36957 10368
rect 36893 10308 36897 10364
rect 36897 10308 36953 10364
rect 36953 10308 36957 10364
rect 36893 10304 36957 10308
rect 36973 10364 37037 10368
rect 36973 10308 36977 10364
rect 36977 10308 37033 10364
rect 37033 10308 37037 10364
rect 36973 10304 37037 10308
rect 37053 10364 37117 10368
rect 37053 10308 37057 10364
rect 37057 10308 37113 10364
rect 37113 10308 37117 10364
rect 37053 10304 37117 10308
rect 9917 9820 9981 9824
rect 9917 9764 9921 9820
rect 9921 9764 9977 9820
rect 9977 9764 9981 9820
rect 9917 9760 9981 9764
rect 9997 9820 10061 9824
rect 9997 9764 10001 9820
rect 10001 9764 10057 9820
rect 10057 9764 10061 9820
rect 9997 9760 10061 9764
rect 10077 9820 10141 9824
rect 10077 9764 10081 9820
rect 10081 9764 10137 9820
rect 10137 9764 10141 9820
rect 10077 9760 10141 9764
rect 10157 9820 10221 9824
rect 10157 9764 10161 9820
rect 10161 9764 10217 9820
rect 10217 9764 10221 9820
rect 10157 9760 10221 9764
rect 27848 9820 27912 9824
rect 27848 9764 27852 9820
rect 27852 9764 27908 9820
rect 27908 9764 27912 9820
rect 27848 9760 27912 9764
rect 27928 9820 27992 9824
rect 27928 9764 27932 9820
rect 27932 9764 27988 9820
rect 27988 9764 27992 9820
rect 27928 9760 27992 9764
rect 28008 9820 28072 9824
rect 28008 9764 28012 9820
rect 28012 9764 28068 9820
rect 28068 9764 28072 9820
rect 28008 9760 28072 9764
rect 28088 9820 28152 9824
rect 28088 9764 28092 9820
rect 28092 9764 28148 9820
rect 28148 9764 28152 9820
rect 28088 9760 28152 9764
rect 45778 9820 45842 9824
rect 45778 9764 45782 9820
rect 45782 9764 45838 9820
rect 45838 9764 45842 9820
rect 45778 9760 45842 9764
rect 45858 9820 45922 9824
rect 45858 9764 45862 9820
rect 45862 9764 45918 9820
rect 45918 9764 45922 9820
rect 45858 9760 45922 9764
rect 45938 9820 46002 9824
rect 45938 9764 45942 9820
rect 45942 9764 45998 9820
rect 45998 9764 46002 9820
rect 45938 9760 46002 9764
rect 46018 9820 46082 9824
rect 46018 9764 46022 9820
rect 46022 9764 46078 9820
rect 46078 9764 46082 9820
rect 46018 9760 46082 9764
rect 18882 9276 18946 9280
rect 18882 9220 18886 9276
rect 18886 9220 18942 9276
rect 18942 9220 18946 9276
rect 18882 9216 18946 9220
rect 18962 9276 19026 9280
rect 18962 9220 18966 9276
rect 18966 9220 19022 9276
rect 19022 9220 19026 9276
rect 18962 9216 19026 9220
rect 19042 9276 19106 9280
rect 19042 9220 19046 9276
rect 19046 9220 19102 9276
rect 19102 9220 19106 9276
rect 19042 9216 19106 9220
rect 19122 9276 19186 9280
rect 19122 9220 19126 9276
rect 19126 9220 19182 9276
rect 19182 9220 19186 9276
rect 19122 9216 19186 9220
rect 36813 9276 36877 9280
rect 36813 9220 36817 9276
rect 36817 9220 36873 9276
rect 36873 9220 36877 9276
rect 36813 9216 36877 9220
rect 36893 9276 36957 9280
rect 36893 9220 36897 9276
rect 36897 9220 36953 9276
rect 36953 9220 36957 9276
rect 36893 9216 36957 9220
rect 36973 9276 37037 9280
rect 36973 9220 36977 9276
rect 36977 9220 37033 9276
rect 37033 9220 37037 9276
rect 36973 9216 37037 9220
rect 37053 9276 37117 9280
rect 37053 9220 37057 9276
rect 37057 9220 37113 9276
rect 37113 9220 37117 9276
rect 37053 9216 37117 9220
rect 9917 8732 9981 8736
rect 9917 8676 9921 8732
rect 9921 8676 9977 8732
rect 9977 8676 9981 8732
rect 9917 8672 9981 8676
rect 9997 8732 10061 8736
rect 9997 8676 10001 8732
rect 10001 8676 10057 8732
rect 10057 8676 10061 8732
rect 9997 8672 10061 8676
rect 10077 8732 10141 8736
rect 10077 8676 10081 8732
rect 10081 8676 10137 8732
rect 10137 8676 10141 8732
rect 10077 8672 10141 8676
rect 10157 8732 10221 8736
rect 10157 8676 10161 8732
rect 10161 8676 10217 8732
rect 10217 8676 10221 8732
rect 10157 8672 10221 8676
rect 27848 8732 27912 8736
rect 27848 8676 27852 8732
rect 27852 8676 27908 8732
rect 27908 8676 27912 8732
rect 27848 8672 27912 8676
rect 27928 8732 27992 8736
rect 27928 8676 27932 8732
rect 27932 8676 27988 8732
rect 27988 8676 27992 8732
rect 27928 8672 27992 8676
rect 28008 8732 28072 8736
rect 28008 8676 28012 8732
rect 28012 8676 28068 8732
rect 28068 8676 28072 8732
rect 28008 8672 28072 8676
rect 28088 8732 28152 8736
rect 28088 8676 28092 8732
rect 28092 8676 28148 8732
rect 28148 8676 28152 8732
rect 28088 8672 28152 8676
rect 45778 8732 45842 8736
rect 45778 8676 45782 8732
rect 45782 8676 45838 8732
rect 45838 8676 45842 8732
rect 45778 8672 45842 8676
rect 45858 8732 45922 8736
rect 45858 8676 45862 8732
rect 45862 8676 45918 8732
rect 45918 8676 45922 8732
rect 45858 8672 45922 8676
rect 45938 8732 46002 8736
rect 45938 8676 45942 8732
rect 45942 8676 45998 8732
rect 45998 8676 46002 8732
rect 45938 8672 46002 8676
rect 46018 8732 46082 8736
rect 46018 8676 46022 8732
rect 46022 8676 46078 8732
rect 46078 8676 46082 8732
rect 46018 8672 46082 8676
rect 18882 8188 18946 8192
rect 18882 8132 18886 8188
rect 18886 8132 18942 8188
rect 18942 8132 18946 8188
rect 18882 8128 18946 8132
rect 18962 8188 19026 8192
rect 18962 8132 18966 8188
rect 18966 8132 19022 8188
rect 19022 8132 19026 8188
rect 18962 8128 19026 8132
rect 19042 8188 19106 8192
rect 19042 8132 19046 8188
rect 19046 8132 19102 8188
rect 19102 8132 19106 8188
rect 19042 8128 19106 8132
rect 19122 8188 19186 8192
rect 19122 8132 19126 8188
rect 19126 8132 19182 8188
rect 19182 8132 19186 8188
rect 19122 8128 19186 8132
rect 36813 8188 36877 8192
rect 36813 8132 36817 8188
rect 36817 8132 36873 8188
rect 36873 8132 36877 8188
rect 36813 8128 36877 8132
rect 36893 8188 36957 8192
rect 36893 8132 36897 8188
rect 36897 8132 36953 8188
rect 36953 8132 36957 8188
rect 36893 8128 36957 8132
rect 36973 8188 37037 8192
rect 36973 8132 36977 8188
rect 36977 8132 37033 8188
rect 37033 8132 37037 8188
rect 36973 8128 37037 8132
rect 37053 8188 37117 8192
rect 37053 8132 37057 8188
rect 37057 8132 37113 8188
rect 37113 8132 37117 8188
rect 37053 8128 37117 8132
rect 9917 7644 9981 7648
rect 9917 7588 9921 7644
rect 9921 7588 9977 7644
rect 9977 7588 9981 7644
rect 9917 7584 9981 7588
rect 9997 7644 10061 7648
rect 9997 7588 10001 7644
rect 10001 7588 10057 7644
rect 10057 7588 10061 7644
rect 9997 7584 10061 7588
rect 10077 7644 10141 7648
rect 10077 7588 10081 7644
rect 10081 7588 10137 7644
rect 10137 7588 10141 7644
rect 10077 7584 10141 7588
rect 10157 7644 10221 7648
rect 10157 7588 10161 7644
rect 10161 7588 10217 7644
rect 10217 7588 10221 7644
rect 10157 7584 10221 7588
rect 27848 7644 27912 7648
rect 27848 7588 27852 7644
rect 27852 7588 27908 7644
rect 27908 7588 27912 7644
rect 27848 7584 27912 7588
rect 27928 7644 27992 7648
rect 27928 7588 27932 7644
rect 27932 7588 27988 7644
rect 27988 7588 27992 7644
rect 27928 7584 27992 7588
rect 28008 7644 28072 7648
rect 28008 7588 28012 7644
rect 28012 7588 28068 7644
rect 28068 7588 28072 7644
rect 28008 7584 28072 7588
rect 28088 7644 28152 7648
rect 28088 7588 28092 7644
rect 28092 7588 28148 7644
rect 28148 7588 28152 7644
rect 28088 7584 28152 7588
rect 45778 7644 45842 7648
rect 45778 7588 45782 7644
rect 45782 7588 45838 7644
rect 45838 7588 45842 7644
rect 45778 7584 45842 7588
rect 45858 7644 45922 7648
rect 45858 7588 45862 7644
rect 45862 7588 45918 7644
rect 45918 7588 45922 7644
rect 45858 7584 45922 7588
rect 45938 7644 46002 7648
rect 45938 7588 45942 7644
rect 45942 7588 45998 7644
rect 45998 7588 46002 7644
rect 45938 7584 46002 7588
rect 46018 7644 46082 7648
rect 46018 7588 46022 7644
rect 46022 7588 46078 7644
rect 46078 7588 46082 7644
rect 46018 7584 46082 7588
rect 18882 7100 18946 7104
rect 18882 7044 18886 7100
rect 18886 7044 18942 7100
rect 18942 7044 18946 7100
rect 18882 7040 18946 7044
rect 18962 7100 19026 7104
rect 18962 7044 18966 7100
rect 18966 7044 19022 7100
rect 19022 7044 19026 7100
rect 18962 7040 19026 7044
rect 19042 7100 19106 7104
rect 19042 7044 19046 7100
rect 19046 7044 19102 7100
rect 19102 7044 19106 7100
rect 19042 7040 19106 7044
rect 19122 7100 19186 7104
rect 19122 7044 19126 7100
rect 19126 7044 19182 7100
rect 19182 7044 19186 7100
rect 19122 7040 19186 7044
rect 36813 7100 36877 7104
rect 36813 7044 36817 7100
rect 36817 7044 36873 7100
rect 36873 7044 36877 7100
rect 36813 7040 36877 7044
rect 36893 7100 36957 7104
rect 36893 7044 36897 7100
rect 36897 7044 36953 7100
rect 36953 7044 36957 7100
rect 36893 7040 36957 7044
rect 36973 7100 37037 7104
rect 36973 7044 36977 7100
rect 36977 7044 37033 7100
rect 37033 7044 37037 7100
rect 36973 7040 37037 7044
rect 37053 7100 37117 7104
rect 37053 7044 37057 7100
rect 37057 7044 37113 7100
rect 37113 7044 37117 7100
rect 37053 7040 37117 7044
rect 9917 6556 9981 6560
rect 9917 6500 9921 6556
rect 9921 6500 9977 6556
rect 9977 6500 9981 6556
rect 9917 6496 9981 6500
rect 9997 6556 10061 6560
rect 9997 6500 10001 6556
rect 10001 6500 10057 6556
rect 10057 6500 10061 6556
rect 9997 6496 10061 6500
rect 10077 6556 10141 6560
rect 10077 6500 10081 6556
rect 10081 6500 10137 6556
rect 10137 6500 10141 6556
rect 10077 6496 10141 6500
rect 10157 6556 10221 6560
rect 10157 6500 10161 6556
rect 10161 6500 10217 6556
rect 10217 6500 10221 6556
rect 10157 6496 10221 6500
rect 27848 6556 27912 6560
rect 27848 6500 27852 6556
rect 27852 6500 27908 6556
rect 27908 6500 27912 6556
rect 27848 6496 27912 6500
rect 27928 6556 27992 6560
rect 27928 6500 27932 6556
rect 27932 6500 27988 6556
rect 27988 6500 27992 6556
rect 27928 6496 27992 6500
rect 28008 6556 28072 6560
rect 28008 6500 28012 6556
rect 28012 6500 28068 6556
rect 28068 6500 28072 6556
rect 28008 6496 28072 6500
rect 28088 6556 28152 6560
rect 28088 6500 28092 6556
rect 28092 6500 28148 6556
rect 28148 6500 28152 6556
rect 28088 6496 28152 6500
rect 45778 6556 45842 6560
rect 45778 6500 45782 6556
rect 45782 6500 45838 6556
rect 45838 6500 45842 6556
rect 45778 6496 45842 6500
rect 45858 6556 45922 6560
rect 45858 6500 45862 6556
rect 45862 6500 45918 6556
rect 45918 6500 45922 6556
rect 45858 6496 45922 6500
rect 45938 6556 46002 6560
rect 45938 6500 45942 6556
rect 45942 6500 45998 6556
rect 45998 6500 46002 6556
rect 45938 6496 46002 6500
rect 46018 6556 46082 6560
rect 46018 6500 46022 6556
rect 46022 6500 46078 6556
rect 46078 6500 46082 6556
rect 46018 6496 46082 6500
rect 18882 6012 18946 6016
rect 18882 5956 18886 6012
rect 18886 5956 18942 6012
rect 18942 5956 18946 6012
rect 18882 5952 18946 5956
rect 18962 6012 19026 6016
rect 18962 5956 18966 6012
rect 18966 5956 19022 6012
rect 19022 5956 19026 6012
rect 18962 5952 19026 5956
rect 19042 6012 19106 6016
rect 19042 5956 19046 6012
rect 19046 5956 19102 6012
rect 19102 5956 19106 6012
rect 19042 5952 19106 5956
rect 19122 6012 19186 6016
rect 19122 5956 19126 6012
rect 19126 5956 19182 6012
rect 19182 5956 19186 6012
rect 19122 5952 19186 5956
rect 36813 6012 36877 6016
rect 36813 5956 36817 6012
rect 36817 5956 36873 6012
rect 36873 5956 36877 6012
rect 36813 5952 36877 5956
rect 36893 6012 36957 6016
rect 36893 5956 36897 6012
rect 36897 5956 36953 6012
rect 36953 5956 36957 6012
rect 36893 5952 36957 5956
rect 36973 6012 37037 6016
rect 36973 5956 36977 6012
rect 36977 5956 37033 6012
rect 37033 5956 37037 6012
rect 36973 5952 37037 5956
rect 37053 6012 37117 6016
rect 37053 5956 37057 6012
rect 37057 5956 37113 6012
rect 37113 5956 37117 6012
rect 37053 5952 37117 5956
rect 9917 5468 9981 5472
rect 9917 5412 9921 5468
rect 9921 5412 9977 5468
rect 9977 5412 9981 5468
rect 9917 5408 9981 5412
rect 9997 5468 10061 5472
rect 9997 5412 10001 5468
rect 10001 5412 10057 5468
rect 10057 5412 10061 5468
rect 9997 5408 10061 5412
rect 10077 5468 10141 5472
rect 10077 5412 10081 5468
rect 10081 5412 10137 5468
rect 10137 5412 10141 5468
rect 10077 5408 10141 5412
rect 10157 5468 10221 5472
rect 10157 5412 10161 5468
rect 10161 5412 10217 5468
rect 10217 5412 10221 5468
rect 10157 5408 10221 5412
rect 27848 5468 27912 5472
rect 27848 5412 27852 5468
rect 27852 5412 27908 5468
rect 27908 5412 27912 5468
rect 27848 5408 27912 5412
rect 27928 5468 27992 5472
rect 27928 5412 27932 5468
rect 27932 5412 27988 5468
rect 27988 5412 27992 5468
rect 27928 5408 27992 5412
rect 28008 5468 28072 5472
rect 28008 5412 28012 5468
rect 28012 5412 28068 5468
rect 28068 5412 28072 5468
rect 28008 5408 28072 5412
rect 28088 5468 28152 5472
rect 28088 5412 28092 5468
rect 28092 5412 28148 5468
rect 28148 5412 28152 5468
rect 28088 5408 28152 5412
rect 45778 5468 45842 5472
rect 45778 5412 45782 5468
rect 45782 5412 45838 5468
rect 45838 5412 45842 5468
rect 45778 5408 45842 5412
rect 45858 5468 45922 5472
rect 45858 5412 45862 5468
rect 45862 5412 45918 5468
rect 45918 5412 45922 5468
rect 45858 5408 45922 5412
rect 45938 5468 46002 5472
rect 45938 5412 45942 5468
rect 45942 5412 45998 5468
rect 45998 5412 46002 5468
rect 45938 5408 46002 5412
rect 46018 5468 46082 5472
rect 46018 5412 46022 5468
rect 46022 5412 46078 5468
rect 46078 5412 46082 5468
rect 46018 5408 46082 5412
rect 18882 4924 18946 4928
rect 18882 4868 18886 4924
rect 18886 4868 18942 4924
rect 18942 4868 18946 4924
rect 18882 4864 18946 4868
rect 18962 4924 19026 4928
rect 18962 4868 18966 4924
rect 18966 4868 19022 4924
rect 19022 4868 19026 4924
rect 18962 4864 19026 4868
rect 19042 4924 19106 4928
rect 19042 4868 19046 4924
rect 19046 4868 19102 4924
rect 19102 4868 19106 4924
rect 19042 4864 19106 4868
rect 19122 4924 19186 4928
rect 19122 4868 19126 4924
rect 19126 4868 19182 4924
rect 19182 4868 19186 4924
rect 19122 4864 19186 4868
rect 36813 4924 36877 4928
rect 36813 4868 36817 4924
rect 36817 4868 36873 4924
rect 36873 4868 36877 4924
rect 36813 4864 36877 4868
rect 36893 4924 36957 4928
rect 36893 4868 36897 4924
rect 36897 4868 36953 4924
rect 36953 4868 36957 4924
rect 36893 4864 36957 4868
rect 36973 4924 37037 4928
rect 36973 4868 36977 4924
rect 36977 4868 37033 4924
rect 37033 4868 37037 4924
rect 36973 4864 37037 4868
rect 37053 4924 37117 4928
rect 37053 4868 37057 4924
rect 37057 4868 37113 4924
rect 37113 4868 37117 4924
rect 37053 4864 37117 4868
rect 9917 4380 9981 4384
rect 9917 4324 9921 4380
rect 9921 4324 9977 4380
rect 9977 4324 9981 4380
rect 9917 4320 9981 4324
rect 9997 4380 10061 4384
rect 9997 4324 10001 4380
rect 10001 4324 10057 4380
rect 10057 4324 10061 4380
rect 9997 4320 10061 4324
rect 10077 4380 10141 4384
rect 10077 4324 10081 4380
rect 10081 4324 10137 4380
rect 10137 4324 10141 4380
rect 10077 4320 10141 4324
rect 10157 4380 10221 4384
rect 10157 4324 10161 4380
rect 10161 4324 10217 4380
rect 10217 4324 10221 4380
rect 10157 4320 10221 4324
rect 27848 4380 27912 4384
rect 27848 4324 27852 4380
rect 27852 4324 27908 4380
rect 27908 4324 27912 4380
rect 27848 4320 27912 4324
rect 27928 4380 27992 4384
rect 27928 4324 27932 4380
rect 27932 4324 27988 4380
rect 27988 4324 27992 4380
rect 27928 4320 27992 4324
rect 28008 4380 28072 4384
rect 28008 4324 28012 4380
rect 28012 4324 28068 4380
rect 28068 4324 28072 4380
rect 28008 4320 28072 4324
rect 28088 4380 28152 4384
rect 28088 4324 28092 4380
rect 28092 4324 28148 4380
rect 28148 4324 28152 4380
rect 28088 4320 28152 4324
rect 45778 4380 45842 4384
rect 45778 4324 45782 4380
rect 45782 4324 45838 4380
rect 45838 4324 45842 4380
rect 45778 4320 45842 4324
rect 45858 4380 45922 4384
rect 45858 4324 45862 4380
rect 45862 4324 45918 4380
rect 45918 4324 45922 4380
rect 45858 4320 45922 4324
rect 45938 4380 46002 4384
rect 45938 4324 45942 4380
rect 45942 4324 45998 4380
rect 45998 4324 46002 4380
rect 45938 4320 46002 4324
rect 46018 4380 46082 4384
rect 46018 4324 46022 4380
rect 46022 4324 46078 4380
rect 46078 4324 46082 4380
rect 46018 4320 46082 4324
rect 18882 3836 18946 3840
rect 18882 3780 18886 3836
rect 18886 3780 18942 3836
rect 18942 3780 18946 3836
rect 18882 3776 18946 3780
rect 18962 3836 19026 3840
rect 18962 3780 18966 3836
rect 18966 3780 19022 3836
rect 19022 3780 19026 3836
rect 18962 3776 19026 3780
rect 19042 3836 19106 3840
rect 19042 3780 19046 3836
rect 19046 3780 19102 3836
rect 19102 3780 19106 3836
rect 19042 3776 19106 3780
rect 19122 3836 19186 3840
rect 19122 3780 19126 3836
rect 19126 3780 19182 3836
rect 19182 3780 19186 3836
rect 19122 3776 19186 3780
rect 36813 3836 36877 3840
rect 36813 3780 36817 3836
rect 36817 3780 36873 3836
rect 36873 3780 36877 3836
rect 36813 3776 36877 3780
rect 36893 3836 36957 3840
rect 36893 3780 36897 3836
rect 36897 3780 36953 3836
rect 36953 3780 36957 3836
rect 36893 3776 36957 3780
rect 36973 3836 37037 3840
rect 36973 3780 36977 3836
rect 36977 3780 37033 3836
rect 37033 3780 37037 3836
rect 36973 3776 37037 3780
rect 37053 3836 37117 3840
rect 37053 3780 37057 3836
rect 37057 3780 37113 3836
rect 37113 3780 37117 3836
rect 37053 3776 37117 3780
rect 9917 3292 9981 3296
rect 9917 3236 9921 3292
rect 9921 3236 9977 3292
rect 9977 3236 9981 3292
rect 9917 3232 9981 3236
rect 9997 3292 10061 3296
rect 9997 3236 10001 3292
rect 10001 3236 10057 3292
rect 10057 3236 10061 3292
rect 9997 3232 10061 3236
rect 10077 3292 10141 3296
rect 10077 3236 10081 3292
rect 10081 3236 10137 3292
rect 10137 3236 10141 3292
rect 10077 3232 10141 3236
rect 10157 3292 10221 3296
rect 10157 3236 10161 3292
rect 10161 3236 10217 3292
rect 10217 3236 10221 3292
rect 10157 3232 10221 3236
rect 27848 3292 27912 3296
rect 27848 3236 27852 3292
rect 27852 3236 27908 3292
rect 27908 3236 27912 3292
rect 27848 3232 27912 3236
rect 27928 3292 27992 3296
rect 27928 3236 27932 3292
rect 27932 3236 27988 3292
rect 27988 3236 27992 3292
rect 27928 3232 27992 3236
rect 28008 3292 28072 3296
rect 28008 3236 28012 3292
rect 28012 3236 28068 3292
rect 28068 3236 28072 3292
rect 28008 3232 28072 3236
rect 28088 3292 28152 3296
rect 28088 3236 28092 3292
rect 28092 3236 28148 3292
rect 28148 3236 28152 3292
rect 28088 3232 28152 3236
rect 45778 3292 45842 3296
rect 45778 3236 45782 3292
rect 45782 3236 45838 3292
rect 45838 3236 45842 3292
rect 45778 3232 45842 3236
rect 45858 3292 45922 3296
rect 45858 3236 45862 3292
rect 45862 3236 45918 3292
rect 45918 3236 45922 3292
rect 45858 3232 45922 3236
rect 45938 3292 46002 3296
rect 45938 3236 45942 3292
rect 45942 3236 45998 3292
rect 45998 3236 46002 3292
rect 45938 3232 46002 3236
rect 46018 3292 46082 3296
rect 46018 3236 46022 3292
rect 46022 3236 46078 3292
rect 46078 3236 46082 3292
rect 46018 3232 46082 3236
rect 18882 2748 18946 2752
rect 18882 2692 18886 2748
rect 18886 2692 18942 2748
rect 18942 2692 18946 2748
rect 18882 2688 18946 2692
rect 18962 2748 19026 2752
rect 18962 2692 18966 2748
rect 18966 2692 19022 2748
rect 19022 2692 19026 2748
rect 18962 2688 19026 2692
rect 19042 2748 19106 2752
rect 19042 2692 19046 2748
rect 19046 2692 19102 2748
rect 19102 2692 19106 2748
rect 19042 2688 19106 2692
rect 19122 2748 19186 2752
rect 19122 2692 19126 2748
rect 19126 2692 19182 2748
rect 19182 2692 19186 2748
rect 19122 2688 19186 2692
rect 36813 2748 36877 2752
rect 36813 2692 36817 2748
rect 36817 2692 36873 2748
rect 36873 2692 36877 2748
rect 36813 2688 36877 2692
rect 36893 2748 36957 2752
rect 36893 2692 36897 2748
rect 36897 2692 36953 2748
rect 36953 2692 36957 2748
rect 36893 2688 36957 2692
rect 36973 2748 37037 2752
rect 36973 2692 36977 2748
rect 36977 2692 37033 2748
rect 37033 2692 37037 2748
rect 36973 2688 37037 2692
rect 37053 2748 37117 2752
rect 37053 2692 37057 2748
rect 37057 2692 37113 2748
rect 37113 2692 37117 2748
rect 37053 2688 37117 2692
rect 9917 2204 9981 2208
rect 9917 2148 9921 2204
rect 9921 2148 9977 2204
rect 9977 2148 9981 2204
rect 9917 2144 9981 2148
rect 9997 2204 10061 2208
rect 9997 2148 10001 2204
rect 10001 2148 10057 2204
rect 10057 2148 10061 2204
rect 9997 2144 10061 2148
rect 10077 2204 10141 2208
rect 10077 2148 10081 2204
rect 10081 2148 10137 2204
rect 10137 2148 10141 2204
rect 10077 2144 10141 2148
rect 10157 2204 10221 2208
rect 10157 2148 10161 2204
rect 10161 2148 10217 2204
rect 10217 2148 10221 2204
rect 10157 2144 10221 2148
rect 27848 2204 27912 2208
rect 27848 2148 27852 2204
rect 27852 2148 27908 2204
rect 27908 2148 27912 2204
rect 27848 2144 27912 2148
rect 27928 2204 27992 2208
rect 27928 2148 27932 2204
rect 27932 2148 27988 2204
rect 27988 2148 27992 2204
rect 27928 2144 27992 2148
rect 28008 2204 28072 2208
rect 28008 2148 28012 2204
rect 28012 2148 28068 2204
rect 28068 2148 28072 2204
rect 28008 2144 28072 2148
rect 28088 2204 28152 2208
rect 28088 2148 28092 2204
rect 28092 2148 28148 2204
rect 28148 2148 28152 2204
rect 28088 2144 28152 2148
rect 45778 2204 45842 2208
rect 45778 2148 45782 2204
rect 45782 2148 45838 2204
rect 45838 2148 45842 2204
rect 45778 2144 45842 2148
rect 45858 2204 45922 2208
rect 45858 2148 45862 2204
rect 45862 2148 45918 2204
rect 45918 2148 45922 2204
rect 45858 2144 45922 2148
rect 45938 2204 46002 2208
rect 45938 2148 45942 2204
rect 45942 2148 45998 2204
rect 45998 2148 46002 2204
rect 45938 2144 46002 2148
rect 46018 2204 46082 2208
rect 46018 2148 46022 2204
rect 46022 2148 46078 2204
rect 46078 2148 46082 2204
rect 46018 2144 46082 2148
<< metal4 >>
rect 9909 25056 10229 25072
rect 9909 24992 9917 25056
rect 9981 24992 9997 25056
rect 10061 24992 10077 25056
rect 10141 24992 10157 25056
rect 10221 24992 10229 25056
rect 9909 23968 10229 24992
rect 9909 23904 9917 23968
rect 9981 23904 9997 23968
rect 10061 23904 10077 23968
rect 10141 23904 10157 23968
rect 10221 23904 10229 23968
rect 9909 22880 10229 23904
rect 9909 22816 9917 22880
rect 9981 22816 9997 22880
rect 10061 22816 10077 22880
rect 10141 22816 10157 22880
rect 10221 22816 10229 22880
rect 9909 21792 10229 22816
rect 9909 21728 9917 21792
rect 9981 21728 9997 21792
rect 10061 21728 10077 21792
rect 10141 21728 10157 21792
rect 10221 21728 10229 21792
rect 9909 20704 10229 21728
rect 9909 20640 9917 20704
rect 9981 20640 9997 20704
rect 10061 20640 10077 20704
rect 10141 20640 10157 20704
rect 10221 20640 10229 20704
rect 9909 19616 10229 20640
rect 9909 19552 9917 19616
rect 9981 19552 9997 19616
rect 10061 19552 10077 19616
rect 10141 19552 10157 19616
rect 10221 19552 10229 19616
rect 9909 18528 10229 19552
rect 9909 18464 9917 18528
rect 9981 18464 9997 18528
rect 10061 18464 10077 18528
rect 10141 18464 10157 18528
rect 10221 18464 10229 18528
rect 9909 17440 10229 18464
rect 9909 17376 9917 17440
rect 9981 17376 9997 17440
rect 10061 17376 10077 17440
rect 10141 17376 10157 17440
rect 10221 17376 10229 17440
rect 9909 16352 10229 17376
rect 9909 16288 9917 16352
rect 9981 16288 9997 16352
rect 10061 16288 10077 16352
rect 10141 16288 10157 16352
rect 10221 16288 10229 16352
rect 9909 15264 10229 16288
rect 9909 15200 9917 15264
rect 9981 15200 9997 15264
rect 10061 15200 10077 15264
rect 10141 15200 10157 15264
rect 10221 15200 10229 15264
rect 9909 14176 10229 15200
rect 9909 14112 9917 14176
rect 9981 14112 9997 14176
rect 10061 14112 10077 14176
rect 10141 14112 10157 14176
rect 10221 14112 10229 14176
rect 9909 13088 10229 14112
rect 9909 13024 9917 13088
rect 9981 13024 9997 13088
rect 10061 13024 10077 13088
rect 10141 13024 10157 13088
rect 10221 13024 10229 13088
rect 9909 12000 10229 13024
rect 9909 11936 9917 12000
rect 9981 11936 9997 12000
rect 10061 11936 10077 12000
rect 10141 11936 10157 12000
rect 10221 11936 10229 12000
rect 9909 10912 10229 11936
rect 9909 10848 9917 10912
rect 9981 10848 9997 10912
rect 10061 10848 10077 10912
rect 10141 10848 10157 10912
rect 10221 10848 10229 10912
rect 9909 9824 10229 10848
rect 9909 9760 9917 9824
rect 9981 9760 9997 9824
rect 10061 9760 10077 9824
rect 10141 9760 10157 9824
rect 10221 9760 10229 9824
rect 9909 8736 10229 9760
rect 9909 8672 9917 8736
rect 9981 8672 9997 8736
rect 10061 8672 10077 8736
rect 10141 8672 10157 8736
rect 10221 8672 10229 8736
rect 9909 7648 10229 8672
rect 9909 7584 9917 7648
rect 9981 7584 9997 7648
rect 10061 7584 10077 7648
rect 10141 7584 10157 7648
rect 10221 7584 10229 7648
rect 9909 6560 10229 7584
rect 9909 6496 9917 6560
rect 9981 6496 9997 6560
rect 10061 6496 10077 6560
rect 10141 6496 10157 6560
rect 10221 6496 10229 6560
rect 9909 5472 10229 6496
rect 9909 5408 9917 5472
rect 9981 5408 9997 5472
rect 10061 5408 10077 5472
rect 10141 5408 10157 5472
rect 10221 5408 10229 5472
rect 9909 4384 10229 5408
rect 9909 4320 9917 4384
rect 9981 4320 9997 4384
rect 10061 4320 10077 4384
rect 10141 4320 10157 4384
rect 10221 4320 10229 4384
rect 9909 3296 10229 4320
rect 9909 3232 9917 3296
rect 9981 3232 9997 3296
rect 10061 3232 10077 3296
rect 10141 3232 10157 3296
rect 10221 3232 10229 3296
rect 9909 2208 10229 3232
rect 9909 2144 9917 2208
rect 9981 2144 9997 2208
rect 10061 2144 10077 2208
rect 10141 2144 10157 2208
rect 10221 2144 10229 2208
rect 9909 2128 10229 2144
rect 18874 24512 19195 25072
rect 18874 24448 18882 24512
rect 18946 24448 18962 24512
rect 19026 24448 19042 24512
rect 19106 24448 19122 24512
rect 19186 24448 19195 24512
rect 18874 23424 19195 24448
rect 18874 23360 18882 23424
rect 18946 23360 18962 23424
rect 19026 23360 19042 23424
rect 19106 23360 19122 23424
rect 19186 23360 19195 23424
rect 18874 22336 19195 23360
rect 18874 22272 18882 22336
rect 18946 22272 18962 22336
rect 19026 22272 19042 22336
rect 19106 22272 19122 22336
rect 19186 22272 19195 22336
rect 18874 21248 19195 22272
rect 18874 21184 18882 21248
rect 18946 21184 18962 21248
rect 19026 21184 19042 21248
rect 19106 21184 19122 21248
rect 19186 21184 19195 21248
rect 18874 20160 19195 21184
rect 18874 20096 18882 20160
rect 18946 20096 18962 20160
rect 19026 20096 19042 20160
rect 19106 20096 19122 20160
rect 19186 20096 19195 20160
rect 18874 19072 19195 20096
rect 18874 19008 18882 19072
rect 18946 19008 18962 19072
rect 19026 19008 19042 19072
rect 19106 19008 19122 19072
rect 19186 19008 19195 19072
rect 18874 17984 19195 19008
rect 18874 17920 18882 17984
rect 18946 17920 18962 17984
rect 19026 17920 19042 17984
rect 19106 17920 19122 17984
rect 19186 17920 19195 17984
rect 18874 16896 19195 17920
rect 18874 16832 18882 16896
rect 18946 16832 18962 16896
rect 19026 16832 19042 16896
rect 19106 16832 19122 16896
rect 19186 16832 19195 16896
rect 18874 15808 19195 16832
rect 18874 15744 18882 15808
rect 18946 15744 18962 15808
rect 19026 15744 19042 15808
rect 19106 15744 19122 15808
rect 19186 15744 19195 15808
rect 18874 14720 19195 15744
rect 18874 14656 18882 14720
rect 18946 14656 18962 14720
rect 19026 14656 19042 14720
rect 19106 14656 19122 14720
rect 19186 14656 19195 14720
rect 18874 13632 19195 14656
rect 18874 13568 18882 13632
rect 18946 13568 18962 13632
rect 19026 13568 19042 13632
rect 19106 13568 19122 13632
rect 19186 13568 19195 13632
rect 18874 12544 19195 13568
rect 18874 12480 18882 12544
rect 18946 12480 18962 12544
rect 19026 12480 19042 12544
rect 19106 12480 19122 12544
rect 19186 12480 19195 12544
rect 18874 11456 19195 12480
rect 18874 11392 18882 11456
rect 18946 11392 18962 11456
rect 19026 11392 19042 11456
rect 19106 11392 19122 11456
rect 19186 11392 19195 11456
rect 18874 10368 19195 11392
rect 18874 10304 18882 10368
rect 18946 10304 18962 10368
rect 19026 10304 19042 10368
rect 19106 10304 19122 10368
rect 19186 10304 19195 10368
rect 18874 9280 19195 10304
rect 18874 9216 18882 9280
rect 18946 9216 18962 9280
rect 19026 9216 19042 9280
rect 19106 9216 19122 9280
rect 19186 9216 19195 9280
rect 18874 8192 19195 9216
rect 18874 8128 18882 8192
rect 18946 8128 18962 8192
rect 19026 8128 19042 8192
rect 19106 8128 19122 8192
rect 19186 8128 19195 8192
rect 18874 7104 19195 8128
rect 18874 7040 18882 7104
rect 18946 7040 18962 7104
rect 19026 7040 19042 7104
rect 19106 7040 19122 7104
rect 19186 7040 19195 7104
rect 18874 6016 19195 7040
rect 18874 5952 18882 6016
rect 18946 5952 18962 6016
rect 19026 5952 19042 6016
rect 19106 5952 19122 6016
rect 19186 5952 19195 6016
rect 18874 4928 19195 5952
rect 18874 4864 18882 4928
rect 18946 4864 18962 4928
rect 19026 4864 19042 4928
rect 19106 4864 19122 4928
rect 19186 4864 19195 4928
rect 18874 3840 19195 4864
rect 18874 3776 18882 3840
rect 18946 3776 18962 3840
rect 19026 3776 19042 3840
rect 19106 3776 19122 3840
rect 19186 3776 19195 3840
rect 18874 2752 19195 3776
rect 18874 2688 18882 2752
rect 18946 2688 18962 2752
rect 19026 2688 19042 2752
rect 19106 2688 19122 2752
rect 19186 2688 19195 2752
rect 18874 2128 19195 2688
rect 27840 25056 28160 25072
rect 27840 24992 27848 25056
rect 27912 24992 27928 25056
rect 27992 24992 28008 25056
rect 28072 24992 28088 25056
rect 28152 24992 28160 25056
rect 27840 23968 28160 24992
rect 27840 23904 27848 23968
rect 27912 23904 27928 23968
rect 27992 23904 28008 23968
rect 28072 23904 28088 23968
rect 28152 23904 28160 23968
rect 27840 22880 28160 23904
rect 27840 22816 27848 22880
rect 27912 22816 27928 22880
rect 27992 22816 28008 22880
rect 28072 22816 28088 22880
rect 28152 22816 28160 22880
rect 27840 21792 28160 22816
rect 27840 21728 27848 21792
rect 27912 21728 27928 21792
rect 27992 21728 28008 21792
rect 28072 21728 28088 21792
rect 28152 21728 28160 21792
rect 27840 20704 28160 21728
rect 27840 20640 27848 20704
rect 27912 20640 27928 20704
rect 27992 20640 28008 20704
rect 28072 20640 28088 20704
rect 28152 20640 28160 20704
rect 27840 19616 28160 20640
rect 27840 19552 27848 19616
rect 27912 19552 27928 19616
rect 27992 19552 28008 19616
rect 28072 19552 28088 19616
rect 28152 19552 28160 19616
rect 27840 18528 28160 19552
rect 27840 18464 27848 18528
rect 27912 18464 27928 18528
rect 27992 18464 28008 18528
rect 28072 18464 28088 18528
rect 28152 18464 28160 18528
rect 27840 17440 28160 18464
rect 27840 17376 27848 17440
rect 27912 17376 27928 17440
rect 27992 17376 28008 17440
rect 28072 17376 28088 17440
rect 28152 17376 28160 17440
rect 27840 16352 28160 17376
rect 27840 16288 27848 16352
rect 27912 16288 27928 16352
rect 27992 16288 28008 16352
rect 28072 16288 28088 16352
rect 28152 16288 28160 16352
rect 27840 15264 28160 16288
rect 27840 15200 27848 15264
rect 27912 15200 27928 15264
rect 27992 15200 28008 15264
rect 28072 15200 28088 15264
rect 28152 15200 28160 15264
rect 27840 14176 28160 15200
rect 27840 14112 27848 14176
rect 27912 14112 27928 14176
rect 27992 14112 28008 14176
rect 28072 14112 28088 14176
rect 28152 14112 28160 14176
rect 27840 13088 28160 14112
rect 27840 13024 27848 13088
rect 27912 13024 27928 13088
rect 27992 13024 28008 13088
rect 28072 13024 28088 13088
rect 28152 13024 28160 13088
rect 27840 12000 28160 13024
rect 27840 11936 27848 12000
rect 27912 11936 27928 12000
rect 27992 11936 28008 12000
rect 28072 11936 28088 12000
rect 28152 11936 28160 12000
rect 27840 10912 28160 11936
rect 27840 10848 27848 10912
rect 27912 10848 27928 10912
rect 27992 10848 28008 10912
rect 28072 10848 28088 10912
rect 28152 10848 28160 10912
rect 27840 9824 28160 10848
rect 27840 9760 27848 9824
rect 27912 9760 27928 9824
rect 27992 9760 28008 9824
rect 28072 9760 28088 9824
rect 28152 9760 28160 9824
rect 27840 8736 28160 9760
rect 27840 8672 27848 8736
rect 27912 8672 27928 8736
rect 27992 8672 28008 8736
rect 28072 8672 28088 8736
rect 28152 8672 28160 8736
rect 27840 7648 28160 8672
rect 27840 7584 27848 7648
rect 27912 7584 27928 7648
rect 27992 7584 28008 7648
rect 28072 7584 28088 7648
rect 28152 7584 28160 7648
rect 27840 6560 28160 7584
rect 27840 6496 27848 6560
rect 27912 6496 27928 6560
rect 27992 6496 28008 6560
rect 28072 6496 28088 6560
rect 28152 6496 28160 6560
rect 27840 5472 28160 6496
rect 27840 5408 27848 5472
rect 27912 5408 27928 5472
rect 27992 5408 28008 5472
rect 28072 5408 28088 5472
rect 28152 5408 28160 5472
rect 27840 4384 28160 5408
rect 27840 4320 27848 4384
rect 27912 4320 27928 4384
rect 27992 4320 28008 4384
rect 28072 4320 28088 4384
rect 28152 4320 28160 4384
rect 27840 3296 28160 4320
rect 27840 3232 27848 3296
rect 27912 3232 27928 3296
rect 27992 3232 28008 3296
rect 28072 3232 28088 3296
rect 28152 3232 28160 3296
rect 27840 2208 28160 3232
rect 27840 2144 27848 2208
rect 27912 2144 27928 2208
rect 27992 2144 28008 2208
rect 28072 2144 28088 2208
rect 28152 2144 28160 2208
rect 27840 2128 28160 2144
rect 36805 24512 37125 25072
rect 36805 24448 36813 24512
rect 36877 24448 36893 24512
rect 36957 24448 36973 24512
rect 37037 24448 37053 24512
rect 37117 24448 37125 24512
rect 36805 23424 37125 24448
rect 36805 23360 36813 23424
rect 36877 23360 36893 23424
rect 36957 23360 36973 23424
rect 37037 23360 37053 23424
rect 37117 23360 37125 23424
rect 36805 22336 37125 23360
rect 36805 22272 36813 22336
rect 36877 22272 36893 22336
rect 36957 22272 36973 22336
rect 37037 22272 37053 22336
rect 37117 22272 37125 22336
rect 36805 21248 37125 22272
rect 36805 21184 36813 21248
rect 36877 21184 36893 21248
rect 36957 21184 36973 21248
rect 37037 21184 37053 21248
rect 37117 21184 37125 21248
rect 36805 20160 37125 21184
rect 36805 20096 36813 20160
rect 36877 20096 36893 20160
rect 36957 20096 36973 20160
rect 37037 20096 37053 20160
rect 37117 20096 37125 20160
rect 36805 19072 37125 20096
rect 36805 19008 36813 19072
rect 36877 19008 36893 19072
rect 36957 19008 36973 19072
rect 37037 19008 37053 19072
rect 37117 19008 37125 19072
rect 36805 17984 37125 19008
rect 36805 17920 36813 17984
rect 36877 17920 36893 17984
rect 36957 17920 36973 17984
rect 37037 17920 37053 17984
rect 37117 17920 37125 17984
rect 36805 16896 37125 17920
rect 36805 16832 36813 16896
rect 36877 16832 36893 16896
rect 36957 16832 36973 16896
rect 37037 16832 37053 16896
rect 37117 16832 37125 16896
rect 36805 15808 37125 16832
rect 36805 15744 36813 15808
rect 36877 15744 36893 15808
rect 36957 15744 36973 15808
rect 37037 15744 37053 15808
rect 37117 15744 37125 15808
rect 36805 14720 37125 15744
rect 36805 14656 36813 14720
rect 36877 14656 36893 14720
rect 36957 14656 36973 14720
rect 37037 14656 37053 14720
rect 37117 14656 37125 14720
rect 36805 13632 37125 14656
rect 36805 13568 36813 13632
rect 36877 13568 36893 13632
rect 36957 13568 36973 13632
rect 37037 13568 37053 13632
rect 37117 13568 37125 13632
rect 36805 12544 37125 13568
rect 36805 12480 36813 12544
rect 36877 12480 36893 12544
rect 36957 12480 36973 12544
rect 37037 12480 37053 12544
rect 37117 12480 37125 12544
rect 36805 11456 37125 12480
rect 36805 11392 36813 11456
rect 36877 11392 36893 11456
rect 36957 11392 36973 11456
rect 37037 11392 37053 11456
rect 37117 11392 37125 11456
rect 36805 10368 37125 11392
rect 36805 10304 36813 10368
rect 36877 10304 36893 10368
rect 36957 10304 36973 10368
rect 37037 10304 37053 10368
rect 37117 10304 37125 10368
rect 36805 9280 37125 10304
rect 36805 9216 36813 9280
rect 36877 9216 36893 9280
rect 36957 9216 36973 9280
rect 37037 9216 37053 9280
rect 37117 9216 37125 9280
rect 36805 8192 37125 9216
rect 36805 8128 36813 8192
rect 36877 8128 36893 8192
rect 36957 8128 36973 8192
rect 37037 8128 37053 8192
rect 37117 8128 37125 8192
rect 36805 7104 37125 8128
rect 36805 7040 36813 7104
rect 36877 7040 36893 7104
rect 36957 7040 36973 7104
rect 37037 7040 37053 7104
rect 37117 7040 37125 7104
rect 36805 6016 37125 7040
rect 36805 5952 36813 6016
rect 36877 5952 36893 6016
rect 36957 5952 36973 6016
rect 37037 5952 37053 6016
rect 37117 5952 37125 6016
rect 36805 4928 37125 5952
rect 36805 4864 36813 4928
rect 36877 4864 36893 4928
rect 36957 4864 36973 4928
rect 37037 4864 37053 4928
rect 37117 4864 37125 4928
rect 36805 3840 37125 4864
rect 36805 3776 36813 3840
rect 36877 3776 36893 3840
rect 36957 3776 36973 3840
rect 37037 3776 37053 3840
rect 37117 3776 37125 3840
rect 36805 2752 37125 3776
rect 36805 2688 36813 2752
rect 36877 2688 36893 2752
rect 36957 2688 36973 2752
rect 37037 2688 37053 2752
rect 37117 2688 37125 2752
rect 36805 2128 37125 2688
rect 45770 25056 46090 25072
rect 45770 24992 45778 25056
rect 45842 24992 45858 25056
rect 45922 24992 45938 25056
rect 46002 24992 46018 25056
rect 46082 24992 46090 25056
rect 45770 23968 46090 24992
rect 45770 23904 45778 23968
rect 45842 23904 45858 23968
rect 45922 23904 45938 23968
rect 46002 23904 46018 23968
rect 46082 23904 46090 23968
rect 45770 22880 46090 23904
rect 45770 22816 45778 22880
rect 45842 22816 45858 22880
rect 45922 22816 45938 22880
rect 46002 22816 46018 22880
rect 46082 22816 46090 22880
rect 45770 21792 46090 22816
rect 45770 21728 45778 21792
rect 45842 21728 45858 21792
rect 45922 21728 45938 21792
rect 46002 21728 46018 21792
rect 46082 21728 46090 21792
rect 45770 20704 46090 21728
rect 45770 20640 45778 20704
rect 45842 20640 45858 20704
rect 45922 20640 45938 20704
rect 46002 20640 46018 20704
rect 46082 20640 46090 20704
rect 45770 19616 46090 20640
rect 45770 19552 45778 19616
rect 45842 19552 45858 19616
rect 45922 19552 45938 19616
rect 46002 19552 46018 19616
rect 46082 19552 46090 19616
rect 45770 18528 46090 19552
rect 45770 18464 45778 18528
rect 45842 18464 45858 18528
rect 45922 18464 45938 18528
rect 46002 18464 46018 18528
rect 46082 18464 46090 18528
rect 45770 17440 46090 18464
rect 45770 17376 45778 17440
rect 45842 17376 45858 17440
rect 45922 17376 45938 17440
rect 46002 17376 46018 17440
rect 46082 17376 46090 17440
rect 45770 16352 46090 17376
rect 45770 16288 45778 16352
rect 45842 16288 45858 16352
rect 45922 16288 45938 16352
rect 46002 16288 46018 16352
rect 46082 16288 46090 16352
rect 45770 15264 46090 16288
rect 45770 15200 45778 15264
rect 45842 15200 45858 15264
rect 45922 15200 45938 15264
rect 46002 15200 46018 15264
rect 46082 15200 46090 15264
rect 45770 14176 46090 15200
rect 45770 14112 45778 14176
rect 45842 14112 45858 14176
rect 45922 14112 45938 14176
rect 46002 14112 46018 14176
rect 46082 14112 46090 14176
rect 45770 13088 46090 14112
rect 45770 13024 45778 13088
rect 45842 13024 45858 13088
rect 45922 13024 45938 13088
rect 46002 13024 46018 13088
rect 46082 13024 46090 13088
rect 45770 12000 46090 13024
rect 45770 11936 45778 12000
rect 45842 11936 45858 12000
rect 45922 11936 45938 12000
rect 46002 11936 46018 12000
rect 46082 11936 46090 12000
rect 45770 10912 46090 11936
rect 45770 10848 45778 10912
rect 45842 10848 45858 10912
rect 45922 10848 45938 10912
rect 46002 10848 46018 10912
rect 46082 10848 46090 10912
rect 45770 9824 46090 10848
rect 45770 9760 45778 9824
rect 45842 9760 45858 9824
rect 45922 9760 45938 9824
rect 46002 9760 46018 9824
rect 46082 9760 46090 9824
rect 45770 8736 46090 9760
rect 45770 8672 45778 8736
rect 45842 8672 45858 8736
rect 45922 8672 45938 8736
rect 46002 8672 46018 8736
rect 46082 8672 46090 8736
rect 45770 7648 46090 8672
rect 45770 7584 45778 7648
rect 45842 7584 45858 7648
rect 45922 7584 45938 7648
rect 46002 7584 46018 7648
rect 46082 7584 46090 7648
rect 45770 6560 46090 7584
rect 45770 6496 45778 6560
rect 45842 6496 45858 6560
rect 45922 6496 45938 6560
rect 46002 6496 46018 6560
rect 46082 6496 46090 6560
rect 45770 5472 46090 6496
rect 45770 5408 45778 5472
rect 45842 5408 45858 5472
rect 45922 5408 45938 5472
rect 46002 5408 46018 5472
rect 46082 5408 46090 5472
rect 45770 4384 46090 5408
rect 45770 4320 45778 4384
rect 45842 4320 45858 4384
rect 45922 4320 45938 4384
rect 46002 4320 46018 4384
rect 46082 4320 46090 4384
rect 45770 3296 46090 4320
rect 45770 3232 45778 3296
rect 45842 3232 45858 3296
rect 45922 3232 45938 3296
rect 46002 3232 46018 3296
rect 46082 3232 46090 3296
rect 45770 2208 46090 3232
rect 45770 2144 45778 2208
rect 45842 2144 45858 2208
rect 45922 2144 45938 2208
rect 46002 2144 46018 2208
rect 46082 2144 46090 2208
rect 45770 2128 46090 2144
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607194113
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607194113
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1607194113
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1607194113
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607194113
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1607194113
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1607194113
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1607194113
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1607194113
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607194113
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607194113
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1607194113
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1607194113
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1607194113
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1607194113
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1607194113
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607194113
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1607194113
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1607194113
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1607194113
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1607194113
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607194113
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1607194113
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1607194113
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1607194113
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1607194113
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1607194113
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1607194113
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1607194113
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1607194113
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1607194113
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1607194113
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1607194113
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1607194113
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1607194113
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1607194113
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1607194113
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1607194113
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1607194113
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1607194113
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:93.inst_tap.g_clkbuf_1.dly $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 19780 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1607194113
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_206
timestamp 1607194113
transform 1 0 20056 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1607194113
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1607194113
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:55.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21712 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:89.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20700 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:90.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1607194113
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1607194113
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_212 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 20608 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1607194113
transform 1 0 20976 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_227
timestamp 1607194113
transform 1 0 21988 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_238
timestamp 1607194113
transform 1 0 23000 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_237
timestamp 1607194113
transform 1 0 22908 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1607194113
transform 1 0 22264 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:88.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22632 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:87.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_249
timestamp 1607194113
transform 1 0 24012 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1607194113
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1607194113
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:86.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23644 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1607194113
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:68.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24748 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:74.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:84.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25760 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:85.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24748 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_260
timestamp 1607194113
transform 1 0 25024 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_260
timestamp 1607194113
transform 1 0 25024 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:76.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26772 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:80.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27600 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:81.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27784 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1607194113
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 1607194113
transform 1 0 26036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_280
timestamp 1607194113
transform 1 0 26864 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_291
timestamp 1607194113
transform 1 0 27876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1607194113
transform 1 0 26036 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_282
timestamp 1607194113
transform 1 0 27048 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:100.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1607194113
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1607194113
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_302
timestamp 1607194113
transform 1 0 28888 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_311
timestamp 1607194113
transform 1 0 29716 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1607194113
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_306
timestamp 1607194113
transform 1 0 29256 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:101.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:102.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29992 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:103.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31464 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:104.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_322
timestamp 1607194113
transform 1 0 30728 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_333
timestamp 1607194113
transform 1 0 31740 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_317
timestamp 1607194113
transform 1 0 30268 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_328
timestamp 1607194113
transform 1 0 31280 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:106.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 32016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:108.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:91.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1607194113
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_342
timestamp 1607194113
transform 1 0 32568 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1607194113
transform 1 0 33580 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_339
timestamp 1607194113
transform 1 0 32292 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_350
timestamp 1607194113
transform 1 0 33304 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1607194113
transform 1 0 34316 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:96.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 34316 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:115.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 34040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_367
timestamp 1607194113
transform 1 0 34868 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_365
timestamp 1607194113
transform 1 0 34684 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_364
timestamp 1607194113
transform 1 0 34592 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1607194113
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_373
timestamp 1607194113
transform 1 0 35420 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1607194113
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:119.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:122.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36616 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:124.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36156 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:126.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37168 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1607194113
transform 1 0 36432 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_395
timestamp 1607194113
transform 1 0 37444 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_378
timestamp 1607194113
transform 1 0 35880 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_389
timestamp 1607194113
transform 1 0 36892 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:125.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:127.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38640 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:128.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1607194113
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_404
timestamp 1607194113
transform 1 0 38272 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_415
timestamp 1607194113
transform 1 0 39284 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_400
timestamp 1607194113
transform 1 0 37904 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_411
timestamp 1607194113
transform 1 0 38916 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_422
timestamp 1607194113
transform 1 0 39928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:131.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 40020 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:130.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39652 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_428
timestamp 1607194113
transform 1 0 40480 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_426
timestamp 1607194113
transform 1 0 40296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_426
timestamp 1607194113
transform 1 0 40296 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1607194113
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1607194113
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_435
timestamp 1607194113
transform 1 0 41124 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:135.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 41216 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:133.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 41860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:137.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 42872 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:139.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 42228 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_446
timestamp 1607194113
transform 1 0 42136 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_457
timestamp 1607194113
transform 1 0 43148 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_439
timestamp 1607194113
transform 1 0 41492 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_450
timestamp 1607194113
transform 1 0 42504 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1607194113
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_466
timestamp 1607194113
transform 1 0 43976 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_478
timestamp 1607194113
transform 1 0 45080 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_462
timestamp 1607194113
transform 1 0 43608 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_474
timestamp 1607194113
transform 1 0 44712 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1607194113
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1607194113
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_490
timestamp 1607194113
transform 1 0 46184 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_497
timestamp 1607194113
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_486
timestamp 1607194113
transform 1 0 45816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_489
timestamp 1607194113
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_509
timestamp 1607194113
transform 1 0 47932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_501
timestamp 1607194113
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_513
timestamp 1607194113
transform 1 0 48300 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1607194113
transform 1 0 49588 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_521
timestamp 1607194113
transform 1 0 49036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_528
timestamp 1607194113
transform 1 0 49680 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_540
timestamp 1607194113
transform 1 0 50784 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_525
timestamp 1607194113
transform 1 0 49404 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_537
timestamp 1607194113
transform 1 0 50508 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1607194113
transform 1 0 52440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1607194113
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_552
timestamp 1607194113
transform 1 0 51888 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_559
timestamp 1607194113
transform 1 0 52532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_550
timestamp 1607194113
transform 1 0 51704 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_562
timestamp 1607194113
transform 1 0 52808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607194113
transform -1 0 54832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607194113
transform -1 0 54832 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_571
timestamp 1607194113
transform 1 0 53636 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_579
timestamp 1607194113
transform 1 0 54372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_574
timestamp 1607194113
transform 1 0 53912 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_580
timestamp 1607194113
transform 1 0 54464 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607194113
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607194113
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607194113
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1607194113
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607194113
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607194113
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607194113
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607194113
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607194113
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1607194113
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1607194113
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607194113
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1607194113
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1607194113
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:97.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13984 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1607194113
transform 1 0 12972 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1607194113
transform 1 0 13708 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_143
timestamp 1607194113
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:9.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1607194113
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1607194113
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1607194113
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_169
timestamp 1607194113
transform 1 0 16652 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_181
timestamp 1607194113
transform 1 0 17756 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:35.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18676 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_189
timestamp 1607194113
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_194
timestamp 1607194113
transform 1 0 18952 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1607194113
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:49.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1607194113
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1607194113
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_226
timestamp 1607194113
transform 1 0 21896 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:59.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22724 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:60.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23736 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_234
timestamp 1607194113
transform 1 0 22632 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_238
timestamp 1607194113
transform 1 0 23000 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_249
timestamp 1607194113
transform 1 0 24012 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:64.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24748 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:69.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_260
timestamp 1607194113
transform 1 0 25024 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:75.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27232 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1607194113
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1607194113
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_276
timestamp 1607194113
transform 1 0 26496 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_287
timestamp 1607194113
transform 1 0 27508 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:79.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28244 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:82.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1607194113
transform 1 0 28520 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1607194113
transform 1 0 29532 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:105.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_317
timestamp 1607194113
transform 1 0 30268 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1607194113
transform 1 0 30636 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_333
timestamp 1607194113
transform 1 0 31740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:109.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 32844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1607194113
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_337
timestamp 1607194113
transform 1 0 32108 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_348
timestamp 1607194113
transform 1 0 33120 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:111.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:114.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 34868 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_359
timestamp 1607194113
transform 1 0 34132 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_370
timestamp 1607194113
transform 1 0 35144 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:117.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35880 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:120.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_381
timestamp 1607194113
transform 1 0 36156 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_392
timestamp 1607194113
transform 1 0 37168 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:129.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38456 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1607194113
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_396
timestamp 1607194113
transform 1 0 37536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1607194113
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_409
timestamp 1607194113
transform 1 0 38732 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:132.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39468 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:134.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 40480 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_420
timestamp 1607194113
transform 1 0 39744 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_431
timestamp 1607194113
transform 1 0 40756 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:138.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 41492 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:142.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 42504 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1607194113
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_442
timestamp 1607194113
transform 1 0 41768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1607194113
transform 1 0 42780 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_457
timestamp 1607194113
transform 1 0 43148 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_459
timestamp 1607194113
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_471
timestamp 1607194113
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_483
timestamp 1607194113
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_495
timestamp 1607194113
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1607194113
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_507
timestamp 1607194113
transform 1 0 47748 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_520
timestamp 1607194113
transform 1 0 48944 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_532
timestamp 1607194113
transform 1 0 50048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_544
timestamp 1607194113
transform 1 0 51152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_556
timestamp 1607194113
transform 1 0 52256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607194113
transform -1 0 54832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1607194113
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_568
timestamp 1607194113
transform 1 0 53360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607194113
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607194113
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1607194113
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1607194113
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1607194113
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:9.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1607194113
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1607194113
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1607194113
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1607194113
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:6.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7820 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_70
timestamp 1607194113
transform 1 0 7544 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_76
timestamp 1607194113
transform 1 0 8096 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_88
timestamp 1607194113
transform 1 0 9200 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_100
timestamp 1607194113
transform 1 0 10304 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1607194113
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_112
timestamp 1607194113
transform 1 0 11408 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1607194113
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_123
timestamp 1607194113
transform 1 0 12420 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:96.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:99.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_134
timestamp 1607194113
transform 1 0 13432 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_145
timestamp 1607194113
transform 1 0 14444 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:7.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:8.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16376 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_153
timestamp 1607194113
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_158
timestamp 1607194113
transform 1 0 15640 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1607194113
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1607194113
transform 1 0 16652 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1607194113
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1607194113
transform 1 0 18032 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:29.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:36.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19780 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_195
timestamp 1607194113
transform 1 0 19044 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_206
timestamp 1607194113
transform 1 0 20056 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:39.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20792 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_217
timestamp 1607194113
transform 1 0 21068 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_229
timestamp 1607194113
transform 1 0 22172 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:45.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22448 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1607194113
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_235
timestamp 1607194113
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1607194113
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1607194113
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:56.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:61.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25392 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_256
timestamp 1607194113
transform 1 0 24656 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_267
timestamp 1607194113
transform 1 0 25668 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:65.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26404 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:72.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_278
timestamp 1607194113
transform 1 0 26680 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_289
timestamp 1607194113
transform 1 0 27692 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:78.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1607194113
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1607194113
transform 1 0 28704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_304
timestamp 1607194113
transform 1 0 29072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1607194113
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:107.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30636 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:110.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_318
timestamp 1607194113
transform 1 0 30360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_324
timestamp 1607194113
transform 1 0 30912 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:113.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 32660 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:116.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_335
timestamp 1607194113
transform 1 0 31924 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_346
timestamp 1607194113
transform 1 0 32936 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:118.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1607194113
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_357
timestamp 1607194113
transform 1 0 33948 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_365
timestamp 1607194113
transform 1 0 34684 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_367
timestamp 1607194113
transform 1 0 34868 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:121.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36616 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_378
timestamp 1607194113
transform 1 0 35880 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_389
timestamp 1607194113
transform 1 0 36892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:136.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39376 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:143.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_401
timestamp 1607194113
transform 1 0 37996 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_408
timestamp 1607194113
transform 1 0 38640 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:140.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 41216 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1607194113
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_419
timestamp 1607194113
transform 1 0 39652 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_428
timestamp 1607194113
transform 1 0 40480 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_439
timestamp 1607194113
transform 1 0 41492 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_451
timestamp 1607194113
transform 1 0 42596 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_463
timestamp 1607194113
transform 1 0 43700 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_475
timestamp 1607194113
transform 1 0 44804 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1607194113
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_487
timestamp 1607194113
transform 1 0 45908 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_489
timestamp 1607194113
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_501
timestamp 1607194113
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_513
timestamp 1607194113
transform 1 0 48300 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_525
timestamp 1607194113
transform 1 0 49404 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_537
timestamp 1607194113
transform 1 0 50508 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1607194113
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_550
timestamp 1607194113
transform 1 0 51704 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_562
timestamp 1607194113
transform 1 0 52808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607194113
transform -1 0 54832 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_574
timestamp 1607194113
transform 1 0 53912 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_580
timestamp 1607194113
transform 1 0 54464 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607194113
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607194113
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607194113
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1607194113
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607194113
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607194113
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:29.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:31.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_44
timestamp 1607194113
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_49
timestamp 1607194113
transform 1 0 5612 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_60
timestamp 1607194113
transform 1 0 6624 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:35.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:39.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_71
timestamp 1607194113
transform 1 0 7636 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_82
timestamp 1607194113
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1607194113
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1607194113
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1607194113
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1607194113
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1607194113
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:95.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14076 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:98.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_129
timestamp 1607194113
transform 1 0 12972 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_133
timestamp 1607194113
transform 1 0 13340 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_144
timestamp 1607194113
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:5.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1607194113
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_delay_line.g_taps:8.g_subtaps:5.inst_tap.g_clkbuf_1.dly_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1607194113
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_154
timestamp 1607194113
transform 1 0 15272 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1607194113
transform 1 0 16284 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:31.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17848 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_177
timestamp 1607194113
transform 1 0 17388 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1607194113
transform 1 0 17756 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_185
timestamp 1607194113
transform 1 0 18124 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:28.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1607194113
transform 1 0 19136 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_208
timestamp 1607194113
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:32.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20424 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:37.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1607194113
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1607194113
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1607194113
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_226
timestamp 1607194113
transform 1 0 21896 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:44.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22632 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:50.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23644 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_237
timestamp 1607194113
transform 1 0 22908 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_248
timestamp 1607194113
transform 1 0 23920 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:52.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24932 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:62.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25944 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_256
timestamp 1607194113
transform 1 0 24656 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_262
timestamp 1607194113
transform 1 0 25208 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:70.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27232 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1607194113
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_273
timestamp 1607194113
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_276
timestamp 1607194113
transform 1 0 26496 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_287
timestamp 1607194113
transform 1 0 27508 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:73.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28244 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:77.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29256 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_298
timestamp 1607194113
transform 1 0 28520 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_309
timestamp 1607194113
transform 1 0 29532 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:83.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30268 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:98.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31280 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_320
timestamp 1607194113
transform 1 0 30544 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1607194113
transform 1 0 31556 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:112.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 32844 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1607194113
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1607194113
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_337
timestamp 1607194113
transform 1 0 32108 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_348
timestamp 1607194113
transform 1 0 33120 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:123.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_360
timestamp 1607194113
transform 1 0 34224 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_372
timestamp 1607194113
transform 1 0 35328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:146.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37352 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_378
timestamp 1607194113
transform 1 0 35880 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_390
timestamp 1607194113
transform 1 0 36984 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:145.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38732 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1607194113
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_398
timestamp 1607194113
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_406
timestamp 1607194113
transform 1 0 38456 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_412
timestamp 1607194113
transform 1 0 39008 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:141.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39744 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:155.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 40756 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_423
timestamp 1607194113
transform 1 0 40020 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_434
timestamp 1607194113
transform 1 0 41032 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1607194113
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_446
timestamp 1607194113
transform 1 0 42136 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_459
timestamp 1607194113
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_471
timestamp 1607194113
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_483
timestamp 1607194113
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_495
timestamp 1607194113
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1607194113
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_507
timestamp 1607194113
transform 1 0 47748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_520
timestamp 1607194113
transform 1 0 48944 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_532
timestamp 1607194113
transform 1 0 50048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_544
timestamp 1607194113
transform 1 0 51152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_556
timestamp 1607194113
transform 1 0 52256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607194113
transform -1 0 54832 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1607194113
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_568
timestamp 1607194113
transform 1 0 53360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:8.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607194113
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1607194113
transform 1 0 1380 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_14
timestamp 1607194113
transform 1 0 2392 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_26
timestamp 1607194113
transform 1 0 3496 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_38
timestamp 1607194113
transform 1 0 4600 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:26.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5152 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1607194113
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_47
timestamp 1607194113
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1607194113
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1607194113
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:30.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:33.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_73
timestamp 1607194113
transform 1 0 7820 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:36.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 9568 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:41.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10580 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1607194113
transform 1 0 8832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_95
timestamp 1607194113
transform 1 0 9844 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:44.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11592 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1607194113
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1607194113
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1607194113
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1607194113
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_123
timestamp 1607194113
transform 1 0 12420 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:50.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_134
timestamp 1607194113
transform 1 0 13432 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:65.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:94.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15088 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_146
timestamp 1607194113
transform 1 0 14536 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_155
timestamp 1607194113
transform 1 0 15364 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1607194113
transform 1 0 16376 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1607194113
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1607194113
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1607194113
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 1607194113
transform 1 0 18032 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:71.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:26.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19780 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_195
timestamp 1607194113
transform 1 0 19044 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_206
timestamp 1607194113
transform 1 0 20056 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:25.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:27.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22080 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_214
timestamp 1607194113
transform 1 0 20792 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_220
timestamp 1607194113
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:38.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1607194113
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_231
timestamp 1607194113
transform 1 0 22356 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_242
timestamp 1607194113
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_245
timestamp 1607194113
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:48.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:51.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25392 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_256
timestamp 1607194113
transform 1 0 24656 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_267
timestamp 1607194113
transform 1 0 25668 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:57.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26404 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:66.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_278
timestamp 1607194113
transform 1 0 26680 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_289
timestamp 1607194113
transform 1 0 27692 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:71.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1607194113
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_300
timestamp 1607194113
transform 1 0 28704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_304
timestamp 1607194113
transform 1 0 29072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_306
timestamp 1607194113
transform 1 0 29256 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:92.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:94.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31004 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_317
timestamp 1607194113
transform 1 0 30268 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_328
timestamp 1607194113
transform 1 0 31280 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_340
timestamp 1607194113
transform 1 0 32384 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_352
timestamp 1607194113
transform 1 0 33488 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1607194113
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_364
timestamp 1607194113
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1607194113
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:148.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37352 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:151.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36340 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_379
timestamp 1607194113
transform 1 0 35972 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_386
timestamp 1607194113
transform 1 0 36616 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:144.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39376 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:147.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_397
timestamp 1607194113
transform 1 0 37628 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_408
timestamp 1607194113
transform 1 0 38640 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:158.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 41216 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1607194113
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_419
timestamp 1607194113
transform 1 0 39652 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_428
timestamp 1607194113
transform 1 0 40480 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_439
timestamp 1607194113
transform 1 0 41492 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_451
timestamp 1607194113
transform 1 0 42596 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_463
timestamp 1607194113
transform 1 0 43700 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_475
timestamp 1607194113
transform 1 0 44804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1607194113
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_487
timestamp 1607194113
transform 1 0 45908 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_489
timestamp 1607194113
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_501
timestamp 1607194113
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_513
timestamp 1607194113
transform 1 0 48300 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_525
timestamp 1607194113
transform 1 0 49404 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_537
timestamp 1607194113
transform 1 0 50508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1607194113
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_550
timestamp 1607194113
transform 1 0 51704 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_562
timestamp 1607194113
transform 1 0 52808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607194113
transform -1 0 54832 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_574
timestamp 1607194113
transform 1 0 53912 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_580
timestamp 1607194113
transform 1 0 54464 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:27.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:5.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607194113
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607194113
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1607194113
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_14
timestamp 1607194113
transform 1 0 2392 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607194113
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1607194113
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_20
timestamp 1607194113
transform 1 0 2944 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:15.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:21.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4784 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:22.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3680 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1607194113
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_26
timestamp 1607194113
transform 1 0 3496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1607194113
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1607194113
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_31
timestamp 1607194113
transform 1 0 3956 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:17.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:24.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:25.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1607194113
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_43
timestamp 1607194113
transform 1 0 5060 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_54
timestamp 1607194113
transform 1 0 6072 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_42
timestamp 1607194113
transform 1 0 4968 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1607194113
transform 1 0 5980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1607194113
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:28.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8188 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:28.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7820 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1607194113
transform 1 0 7084 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1607194113
transform 1 0 8096 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_74
timestamp 1607194113
transform 1 0 7912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_80
timestamp 1607194113
transform 1 0 8464 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_91
timestamp 1607194113
transform 1 0 9476 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1607194113
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1607194113
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1607194113
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:32.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8832 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:3.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 9200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_93
timestamp 1607194113
transform 1 0 9660 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:38.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:37.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10212 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1607194113
transform 1 0 10488 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_104
timestamp 1607194113
transform 1 0 10672 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:40.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:42.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:45.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 12420 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1607194113
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_115
timestamp 1607194113
transform 1 0 11684 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1607194113
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1607194113
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_123
timestamp 1607194113
transform 1 0 12420 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:43.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:47.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13432 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:48.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:53.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_126
timestamp 1607194113
transform 1 0 12696 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_137
timestamp 1607194113
transform 1 0 13708 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_134
timestamp 1607194113
transform 1 0 13432 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_145
timestamp 1607194113
transform 1 0 14444 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:52.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15180 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:57.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16192 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:59.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1607194113
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1607194113
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1607194113
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_154
timestamp 1607194113
transform 1 0 15272 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1607194113
transform 1 0 16284 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_156
timestamp 1607194113
transform 1 0 15456 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_167
timestamp 1607194113
transform 1 0 16468 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:63.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17020 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:60.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17204 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_184
timestamp 1607194113
transform 1 0 18032 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1607194113
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1607194113
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_176
timestamp 1607194113
transform 1 0 17296 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1607194113
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:67.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18032 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_187
timestamp 1607194113
transform 1 0 18308 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:66.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:68.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:69.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19780 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:74.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20056 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_198
timestamp 1607194113
transform 1 0 19320 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_195
timestamp 1607194113
transform 1 0 19044 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_206
timestamp 1607194113
transform 1 0 20056 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:72.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20792 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:245.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1607194113
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1607194113
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1607194113
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1607194113
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_226
timestamp 1607194113
transform 1 0 21896 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_217
timestamp 1607194113
transform 1 0 21068 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_229
timestamp 1607194113
transform 1 0 22172 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:242.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:252.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22632 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:33.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23644 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1607194113
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_237
timestamp 1607194113
transform 1 0 22908 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_248
timestamp 1607194113
transform 1 0 23920 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_236
timestamp 1607194113
transform 1 0 22816 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_245
timestamp 1607194113
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:40.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:41.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25392 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:42.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24656 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:46.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25668 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_259
timestamp 1607194113
transform 1 0 24932 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1607194113
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_256
timestamp 1607194113
transform 1 0 24656 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_267
timestamp 1607194113
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:47.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:53.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:58.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1607194113
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1607194113
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_276
timestamp 1607194113
transform 1 0 26496 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_287
timestamp 1607194113
transform 1 0 27508 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_278
timestamp 1607194113
transform 1 0 26680 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_289
timestamp 1607194113
transform 1 0 27692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:63.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28244 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:67.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:95.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1607194113
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_298
timestamp 1607194113
transform 1 0 28520 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1607194113
transform 1 0 29532 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_300
timestamp 1607194113
transform 1 0 28704 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_304
timestamp 1607194113
transform 1 0 29072 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_306
timestamp 1607194113
transform 1 0 29256 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:97.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30268 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:99.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29992 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_320
timestamp 1607194113
transform 1 0 30544 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_332
timestamp 1607194113
transform 1 0 31648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1607194113
transform 1 0 30268 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_329
timestamp 1607194113
transform 1 0 31372 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1607194113
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_337
timestamp 1607194113
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_349
timestamp 1607194113
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_341
timestamp 1607194113
transform 1 0 32476 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_353
timestamp 1607194113
transform 1 0 33580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:164.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:166.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:171.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33764 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1607194113
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_361
timestamp 1607194113
transform 1 0 34316 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_369
timestamp 1607194113
transform 1 0 35052 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_375
timestamp 1607194113
transform 1 0 35604 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_358
timestamp 1607194113
transform 1 0 34040 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_367
timestamp 1607194113
transform 1 0 34868 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:150.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37352 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:153.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36340 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:157.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36616 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_386
timestamp 1607194113
transform 1 0 36616 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_378
timestamp 1607194113
transform 1 0 35880 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_389
timestamp 1607194113
transform 1 0 36892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:149.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:152.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37720 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:159.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38732 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1607194113
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_398
timestamp 1607194113
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_409
timestamp 1607194113
transform 1 0 38732 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_397
timestamp 1607194113
transform 1 0 37628 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_401
timestamp 1607194113
transform 1 0 37996 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_412
timestamp 1607194113
transform 1 0 39008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:154.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39468 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:161.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 40480 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1607194113
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_420
timestamp 1607194113
transform 1 0 39744 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_431
timestamp 1607194113
transform 1 0 40756 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_424
timestamp 1607194113
transform 1 0 40112 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_428
timestamp 1607194113
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1607194113
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_443
timestamp 1607194113
transform 1 0 41860 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_455
timestamp 1607194113
transform 1 0 42964 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_440
timestamp 1607194113
transform 1 0 41584 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_452
timestamp 1607194113
transform 1 0 42688 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_459
timestamp 1607194113
transform 1 0 43332 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_471
timestamp 1607194113
transform 1 0 44436 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_464
timestamp 1607194113
transform 1 0 43792 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_476
timestamp 1607194113
transform 1 0 44896 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1607194113
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_483
timestamp 1607194113
transform 1 0 45540 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_495
timestamp 1607194113
transform 1 0 46644 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_489
timestamp 1607194113
transform 1 0 46092 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1607194113
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_507
timestamp 1607194113
transform 1 0 47748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_520
timestamp 1607194113
transform 1 0 48944 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_501
timestamp 1607194113
transform 1 0 47196 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_513
timestamp 1607194113
transform 1 0 48300 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_532
timestamp 1607194113
transform 1 0 50048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_525
timestamp 1607194113
transform 1 0 49404 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_537
timestamp 1607194113
transform 1 0 50508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1607194113
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_544
timestamp 1607194113
transform 1 0 51152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_556
timestamp 1607194113
transform 1 0 52256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_550
timestamp 1607194113
transform 1 0 51704 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_562
timestamp 1607194113
transform 1 0 52808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607194113
transform -1 0 54832 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607194113
transform -1 0 54832 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1607194113
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_568
timestamp 1607194113
transform 1 0 53360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_574
timestamp 1607194113
transform 1 0 53912 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_580
timestamp 1607194113
transform 1 0 54464 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:23.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2668 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607194113
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607194113
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_15
timestamp 1607194113
transform 1 0 2484 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1607194113
transform 1 0 2944 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:16.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607194113
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1607194113
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:13.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5612 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1607194113
transform 1 0 5152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_48
timestamp 1607194113
transform 1 0 5520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_52
timestamp 1607194113
transform 1 0 5888 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:23.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7452 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:26.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_64
timestamp 1607194113
transform 1 0 6992 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_68
timestamp 1607194113
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_72
timestamp 1607194113
transform 1 0 7728 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_83
timestamp 1607194113
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:29.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607194113
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1607194113
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1607194113
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_104
timestamp 1607194113
transform 1 0 10672 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:120.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 12512 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:34.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11408 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_115
timestamp 1607194113
transform 1 0 11684 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_123
timestamp 1607194113
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:46.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13524 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_127
timestamp 1607194113
transform 1 0 12788 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_138
timestamp 1607194113
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:56.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607194113
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1607194113
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1607194113
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_165
timestamp 1607194113
transform 1 0 16284 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:58.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:61.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18032 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_176
timestamp 1607194113
transform 1 0 17296 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_187
timestamp 1607194113
transform 1 0 18308 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:64.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19044 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:73.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20056 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_198
timestamp 1607194113
transform 1 0 19320 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:78.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607194113
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1607194113
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1607194113
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1607194113
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_226
timestamp 1607194113
transform 1 0 21896 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:241.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22724 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:243.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23736 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_234
timestamp 1607194113
transform 1 0 22632 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_238
timestamp 1607194113
transform 1 0 23000 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_249
timestamp 1607194113
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:247.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:43.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_260
timestamp 1607194113
transform 1 0 25024 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:54.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27232 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607194113
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_271
timestamp 1607194113
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_276
timestamp 1607194113
transform 1 0 26496 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_287
timestamp 1607194113
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:210.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_299
timestamp 1607194113
transform 1 0 28612 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_307
timestamp 1607194113
transform 1 0 29348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_312
timestamp 1607194113
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_324
timestamp 1607194113
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:173.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607194113
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_337
timestamp 1607194113
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_349
timestamp 1607194113
transform 1 0 33212 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:168.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:172.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 34592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_356
timestamp 1607194113
transform 1 0 33856 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_367
timestamp 1607194113
transform 1 0 34868 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:163.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36708 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_378
timestamp 1607194113
transform 1 0 35880 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_386
timestamp 1607194113
transform 1 0 36616 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_390
timestamp 1607194113
transform 1 0 36984 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:156.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607194113
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_396
timestamp 1607194113
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1607194113
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_409
timestamp 1607194113
transform 1 0 38732 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:160.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 39468 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_420
timestamp 1607194113
transform 1 0 39744 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_432
timestamp 1607194113
transform 1 0 40848 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607194113
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_444
timestamp 1607194113
transform 1 0 41952 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_456
timestamp 1607194113
transform 1 0 43056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_459
timestamp 1607194113
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_471
timestamp 1607194113
transform 1 0 44436 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_483
timestamp 1607194113
transform 1 0 45540 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_495
timestamp 1607194113
transform 1 0 46644 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607194113
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_507
timestamp 1607194113
transform 1 0 47748 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_520
timestamp 1607194113
transform 1 0 48944 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_532
timestamp 1607194113
transform 1 0 50048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_544
timestamp 1607194113
transform 1 0 51152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_556
timestamp 1607194113
transform 1 0 52256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607194113
transform -1 0 54832 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607194113
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_568
timestamp 1607194113
transform 1 0 53360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:20.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607194113
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1607194113
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_14
timestamp 1607194113
transform 1 0 2392 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:14.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:19.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3496 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_29
timestamp 1607194113
transform 1 0 3772 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_40
timestamp 1607194113
transform 1 0 4784 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:12.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607194113
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1607194113
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1607194113
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1607194113
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:20.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:24.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_73
timestamp 1607194113
transform 1 0 7820 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:27.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 9568 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:30.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_84
timestamp 1607194113
transform 1 0 8832 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_95
timestamp 1607194113
transform 1 0 9844 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607194113
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_106
timestamp 1607194113
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1607194113
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_123
timestamp 1607194113
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:115.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:49.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_134
timestamp 1607194113
transform 1 0 13432 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_145
timestamp 1607194113
transform 1 0 14444 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:51.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:54.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16192 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_156
timestamp 1607194113
transform 1 0 15456 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:79.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17572 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607194113
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_167
timestamp 1607194113
transform 1 0 16468 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1607194113
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1607194113
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:70.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:75.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19780 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_195
timestamp 1607194113
transform 1 0 19044 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_206
timestamp 1607194113
transform 1 0 20056 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:77.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20792 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_217
timestamp 1607194113
transform 1 0 21068 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_229
timestamp 1607194113
transform 1 0 22172 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:240.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22540 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607194113
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_236
timestamp 1607194113
transform 1 0 22816 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_245
timestamp 1607194113
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:246.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:34.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25392 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_256
timestamp 1607194113
transform 1 0 24656 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_267
timestamp 1607194113
transform 1 0 25668 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:216.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_279
timestamp 1607194113
transform 1 0 26772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_288
timestamp 1607194113
transform 1 0 27600 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607194113
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_300
timestamp 1607194113
transform 1 0 28704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_304
timestamp 1607194113
transform 1 0 29072 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_306
timestamp 1607194113
transform 1 0 29256 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:209.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29992 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1607194113
transform 1 0 30268 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_329
timestamp 1607194113
transform 1 0 31372 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:198.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 32752 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_341
timestamp 1607194113
transform 1 0 32476 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_347
timestamp 1607194113
transform 1 0 33028 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:169.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:176.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607194113
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_358
timestamp 1607194113
transform 1 0 34040 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_367
timestamp 1607194113
transform 1 0 34868 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:165.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36616 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_378
timestamp 1607194113
transform 1 0 35880 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_389
timestamp 1607194113
transform 1 0 36892 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:162.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_397
timestamp 1607194113
transform 1 0 37628 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_402
timestamp 1607194113
transform 1 0 38088 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_414
timestamp 1607194113
transform 1 0 39192 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607194113
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_426
timestamp 1607194113
transform 1 0 40296 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_428
timestamp 1607194113
transform 1 0 40480 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_440
timestamp 1607194113
transform 1 0 41584 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_452
timestamp 1607194113
transform 1 0 42688 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_464
timestamp 1607194113
transform 1 0 43792 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_476
timestamp 1607194113
transform 1 0 44896 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607194113
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_489
timestamp 1607194113
transform 1 0 46092 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_501
timestamp 1607194113
transform 1 0 47196 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_513
timestamp 1607194113
transform 1 0 48300 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_525
timestamp 1607194113
transform 1 0 49404 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_537
timestamp 1607194113
transform 1 0 50508 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607194113
transform 1 0 51612 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_550
timestamp 1607194113
transform 1 0 51704 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_562
timestamp 1607194113
transform 1 0 52808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607194113
transform -1 0 54832 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_574
timestamp 1607194113
transform 1 0 53912 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_580
timestamp 1607194113
transform 1 0 54464 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:6.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607194113
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1607194113
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_14
timestamp 1607194113
transform 1 0 2392 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:18.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607194113
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1607194113
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1607194113
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:21.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:11.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5520 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_44
timestamp 1607194113
transform 1 0 5152 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1607194113
transform 1 0 5796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_62
timestamp 1607194113
transform 1 0 6808 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:17.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:22.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_73
timestamp 1607194113
transform 1 0 7820 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:25.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607194113
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1607194113
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1607194113
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_104
timestamp 1607194113
transform 1 0 10672 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:32.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11408 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:34.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 12420 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_115
timestamp 1607194113
transform 1 0 11684 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:101.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13432 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_126
timestamp 1607194113
transform 1 0 12696 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_137
timestamp 1607194113
transform 1 0 13708 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:55.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:85.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607194113
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_149
timestamp 1607194113
transform 1 0 14812 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_154
timestamp 1607194113
transform 1 0 15272 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_165
timestamp 1607194113
transform 1 0 16284 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:62.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17020 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_176
timestamp 1607194113
transform 1 0 17296 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:76.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18584 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:84.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19596 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1607194113
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_193
timestamp 1607194113
transform 1 0 18860 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1607194113
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:24.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607194113
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1607194113
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1607194113
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_226
timestamp 1607194113
transform 1 0 21896 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:236.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:238.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23092 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_238
timestamp 1607194113
transform 1 0 23000 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_242
timestamp 1607194113
transform 1 0 23368 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:250.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25116 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1607194113
transform 1 0 24380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_264
timestamp 1607194113
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:215.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27508 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:217.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607194113
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_276
timestamp 1607194113
transform 1 0 26496 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_284
timestamp 1607194113
transform 1 0 27232 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_290
timestamp 1607194113
transform 1 0 27784 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:208.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29532 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:212.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28520 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_301
timestamp 1607194113
transform 1 0 28796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_312
timestamp 1607194113
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_324
timestamp 1607194113
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607194113
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_337
timestamp 1607194113
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_349
timestamp 1607194113
transform 1 0 33212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:174.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 34776 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:178.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33764 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_358
timestamp 1607194113
transform 1 0 34040 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_369
timestamp 1607194113
transform 1 0 35052 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:167.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36800 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:170.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35788 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_380
timestamp 1607194113
transform 1 0 36064 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_391
timestamp 1607194113
transform 1 0 37076 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607194113
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_398
timestamp 1607194113
transform 1 0 37720 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_410
timestamp 1607194113
transform 1 0 38824 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_422
timestamp 1607194113
transform 1 0 39928 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_434
timestamp 1607194113
transform 1 0 41032 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607194113
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_446
timestamp 1607194113
transform 1 0 42136 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_459
timestamp 1607194113
transform 1 0 43332 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_471
timestamp 1607194113
transform 1 0 44436 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_483
timestamp 1607194113
transform 1 0 45540 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_495
timestamp 1607194113
transform 1 0 46644 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607194113
transform 1 0 48852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_507
timestamp 1607194113
transform 1 0 47748 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_520
timestamp 1607194113
transform 1 0 48944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_532
timestamp 1607194113
transform 1 0 50048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_544
timestamp 1607194113
transform 1 0 51152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_556
timestamp 1607194113
transform 1 0 52256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607194113
transform -1 0 54832 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607194113
transform 1 0 54464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_568
timestamp 1607194113
transform 1 0 53360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:5.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607194113
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607194113
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1607194113
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:10.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_22
timestamp 1607194113
transform 1 0 3128 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1607194113
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 1607194113
transform 1 0 4692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:7.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:8.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607194113
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_50
timestamp 1607194113
transform 1 0 5704 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1607194113
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:15.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:19.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_73
timestamp 1607194113
transform 1 0 7820 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:31.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:33.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10580 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_84
timestamp 1607194113
transform 1 0 8832 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_95
timestamp 1607194113
transform 1 0 9844 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607194113
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_106
timestamp 1607194113
transform 1 0 10856 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1607194113
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_123
timestamp 1607194113
transform 1 0 12420 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:39.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:100.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_134
timestamp 1607194113
transform 1 0 13432 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_145
timestamp 1607194113
transform 1 0 14444 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:110.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_156
timestamp 1607194113
transform 1 0 15456 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:82.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16928 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607194113
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_168
timestamp 1607194113
transform 1 0 16560 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1607194113
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_184
timestamp 1607194113
transform 1 0 18032 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:80.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:83.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19780 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_195
timestamp 1607194113
transform 1 0 19044 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_206
timestamp 1607194113
transform 1 0 20056 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:88.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20792 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:92.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21804 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_217
timestamp 1607194113
transform 1 0 21068 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_228
timestamp 1607194113
transform 1 0 22080 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:239.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22816 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607194113
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1607194113
transform 1 0 23092 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1607194113
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1607194113
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:221.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25116 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1607194113
transform 1 0 24748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_264
timestamp 1607194113
transform 1 0 25392 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:214.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27140 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:218.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26128 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_275
timestamp 1607194113
transform 1 0 26404 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_286
timestamp 1607194113
transform 1 0 27416 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:211.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607194113
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_297
timestamp 1607194113
transform 1 0 28428 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_306
timestamp 1607194113
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:200.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31740 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:204.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_318
timestamp 1607194113
transform 1 0 30360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_323
timestamp 1607194113
transform 1 0 30820 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_331
timestamp 1607194113
transform 1 0 31556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:196.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 32752 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_336
timestamp 1607194113
transform 1 0 32016 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_347
timestamp 1607194113
transform 1 0 33028 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:175.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:181.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33764 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607194113
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_358
timestamp 1607194113
transform 1 0 34040 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_367
timestamp 1607194113
transform 1 0 34868 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:179.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36616 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_378
timestamp 1607194113
transform 1 0 35880 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_389
timestamp 1607194113
transform 1 0 36892 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:184.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37628 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_400
timestamp 1607194113
transform 1 0 37904 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_412
timestamp 1607194113
transform 1 0 39008 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607194113
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_424
timestamp 1607194113
transform 1 0 40112 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_428
timestamp 1607194113
transform 1 0 40480 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_440
timestamp 1607194113
transform 1 0 41584 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_452
timestamp 1607194113
transform 1 0 42688 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_464
timestamp 1607194113
transform 1 0 43792 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_476
timestamp 1607194113
transform 1 0 44896 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607194113
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_489
timestamp 1607194113
transform 1 0 46092 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_501
timestamp 1607194113
transform 1 0 47196 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_513
timestamp 1607194113
transform 1 0 48300 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_525
timestamp 1607194113
transform 1 0 49404 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_537
timestamp 1607194113
transform 1 0 50508 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607194113
transform 1 0 51612 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_550
timestamp 1607194113
transform 1 0 51704 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_562
timestamp 1607194113
transform 1 0 52808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607194113
transform -1 0 54832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_574
timestamp 1607194113
transform 1 0 53912 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_580
timestamp 1607194113
transform 1 0 54464 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:4.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607194113
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607194113
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1607194113
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1607194113
transform 1 0 2852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:8.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4784 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607194113
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1607194113
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1607194113
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:18.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_43
timestamp 1607194113
transform 1 0 5060 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_55
timestamp 1607194113
transform 1 0 6164 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_61
timestamp 1607194113
transform 1 0 6716 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:13.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:16.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8464 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_72
timestamp 1607194113
transform 1 0 7728 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1607194113
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:35.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607194113
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1607194113
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1607194113
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_104
timestamp 1607194113
transform 1 0 10672 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:36.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:38.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 12420 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_115
timestamp 1607194113
transform 1 0 11684 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:45.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_126
timestamp 1607194113
transform 1 0 12696 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_137
timestamp 1607194113
transform 1 0 13708 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:103.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607194113
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1607194113
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_154
timestamp 1607194113
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_165
timestamp 1607194113
transform 1 0 16284 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:7.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17020 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:81.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18032 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_delay_line.g_taps:7.g_subtaps:7.inst_tap.g_clkbuf_1.dly_A
timestamp 1607194113
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_176
timestamp 1607194113
transform 1 0 17296 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1607194113
transform 1 0 18308 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:86.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19044 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:90.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20056 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_198
timestamp 1607194113
transform 1 0 19320 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:21.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607194113
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1607194113
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1607194113
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1607194113
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_226
timestamp 1607194113
transform 1 0 21896 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:233.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:237.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23092 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_238
timestamp 1607194113
transform 1 0 23000 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_242
timestamp 1607194113
transform 1 0 23368 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:225.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25116 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1607194113
transform 1 0 24380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_264
timestamp 1607194113
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:213.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27692 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:219.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607194113
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1607194113
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_288
timestamp 1607194113
transform 1 0 27600 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:203.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:207.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_292
timestamp 1607194113
transform 1 0 27968 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_303
timestamp 1607194113
transform 1 0 28980 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:195.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:201.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_314
timestamp 1607194113
transform 1 0 29992 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_325
timestamp 1607194113
transform 1 0 31004 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:192.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33120 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607194113
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_337
timestamp 1607194113
transform 1 0 32108 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_345
timestamp 1607194113
transform 1 0 32844 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_351
timestamp 1607194113
transform 1 0 33396 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:177.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:182.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 34132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_362
timestamp 1607194113
transform 1 0 34408 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_373
timestamp 1607194113
transform 1 0 35420 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:183.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_384
timestamp 1607194113
transform 1 0 36432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:189.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 38456 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607194113
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_396
timestamp 1607194113
transform 1 0 37536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1607194113
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_409
timestamp 1607194113
transform 1 0 38732 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1607194113
transform 1 0 39836 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1607194113
transform 1 0 40940 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607194113
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1607194113
transform 1 0 42044 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_457
timestamp 1607194113
transform 1 0 43148 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_459
timestamp 1607194113
transform 1 0 43332 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_471
timestamp 1607194113
transform 1 0 44436 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_483
timestamp 1607194113
transform 1 0 45540 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_495
timestamp 1607194113
transform 1 0 46644 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607194113
transform 1 0 48852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_507
timestamp 1607194113
transform 1 0 47748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_520
timestamp 1607194113
transform 1 0 48944 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_532
timestamp 1607194113
transform 1 0 50048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_544
timestamp 1607194113
transform 1 0 51152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_556
timestamp 1607194113
transform 1 0 52256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607194113
transform -1 0 54832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607194113
transform 1 0 54464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_568
timestamp 1607194113
transform 1 0 53360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1607194113
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1607194113
transform 1 0 1380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607194113
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607194113
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_15
timestamp 1607194113
transform 1 0 2484 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1607194113
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_17
timestamp 1607194113
transform 1 0 2668 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_11
timestamp 1607194113
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:13.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2392 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:11.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2208 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1607194113
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_28
timestamp 1607194113
transform 1 0 3680 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:7.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:15.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3404 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1607194113
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1607194113
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607194113
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:18.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 1607194113
transform 1 0 4692 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:16.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4784 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:17.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:6.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607194113
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 1607194113
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1607194113
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1607194113
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_43
timestamp 1607194113
transform 1 0 5060 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_54
timestamp 1607194113
transform 1 0 6072 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1607194113
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:10.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:11.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8004 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:12.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:14.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_73
timestamp 1607194113
transform 1 0 7820 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_67
timestamp 1607194113
transform 1 0 7268 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1607194113
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:37.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10488 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:40.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:41.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607194113
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_84
timestamp 1607194113
transform 1 0 8832 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_96
timestamp 1607194113
transform 1 0 9936 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_86
timestamp 1607194113
transform 1 0 9016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1607194113
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_101
timestamp 1607194113
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:43.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11500 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:48.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 12512 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607194113
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_105
timestamp 1607194113
transform 1 0 10764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1607194113
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1607194113
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_123
timestamp 1607194113
transform 1 0 12420 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_105
timestamp 1607194113
transform 1 0 10764 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_116
timestamp 1607194113
transform 1 0 11776 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:44.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:49.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:53.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_134
timestamp 1607194113
transform 1 0 13432 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_145
timestamp 1607194113
transform 1 0 14444 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_127
timestamp 1607194113
transform 1 0 12788 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_138
timestamp 1607194113
transform 1 0 13800 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:102.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15180 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:104.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16192 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:106.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607194113
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_156
timestamp 1607194113
transform 1 0 15456 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1607194113
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1607194113
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1607194113
transform 1 0 16284 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_167
timestamp 1607194113
transform 1 0 16468 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:109.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17020 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:107.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17204 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_176
timestamp 1607194113
transform 1 0 17296 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_184
timestamp 1607194113
transform 1 0 18032 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1607194113
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1607194113
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607194113
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:114.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18032 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1607194113
transform 1 0 18308 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:87.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:89.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:91.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19780 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:12.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20056 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_195
timestamp 1607194113
transform 1 0 19044 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_206
timestamp 1607194113
transform 1 0 20056 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_198
timestamp 1607194113
transform 1 0 19320 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1607194113
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1607194113
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1607194113
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_217
timestamp 1607194113
transform 1 0 21068 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607194113
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:93.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20792 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_226
timestamp 1607194113
transform 1 0 21896 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:19.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21804 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:15.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_228
timestamp 1607194113
transform 1 0 22080 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:18.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22632 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:22.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22816 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607194113
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1607194113
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1607194113
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_245
timestamp 1607194113
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1607194113
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_249
timestamp 1607194113
transform 1 0 24012 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:228.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25392 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:230.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 25392 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:231.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:232.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_256
timestamp 1607194113
transform 1 0 24656 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_267
timestamp 1607194113
transform 1 0 25668 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_256
timestamp 1607194113
transform 1 0 24656 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_267
timestamp 1607194113
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:220.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 26404 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:222.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27232 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:223.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607194113
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_278
timestamp 1607194113
transform 1 0 26680 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_289
timestamp 1607194113
transform 1 0 27692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_276
timestamp 1607194113
transform 1 0 26496 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_287
timestamp 1607194113
transform 1 0 27508 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:206.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:224.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 28244 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:227.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607194113
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_301
timestamp 1607194113
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_306
timestamp 1607194113
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1607194113
transform 1 0 28520 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1607194113
transform 1 0 29532 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:199.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31740 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:202.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30728 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:205.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 30268 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_318
timestamp 1607194113
transform 1 0 30360 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_325
timestamp 1607194113
transform 1 0 31004 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_320
timestamp 1607194113
transform 1 0 30544 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_332
timestamp 1607194113
transform 1 0 31648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:194.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 32752 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:197.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33028 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607194113
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_336
timestamp 1607194113
transform 1 0 32016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_347
timestamp 1607194113
transform 1 0 33028 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_337
timestamp 1607194113
transform 1 0 32108 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_345
timestamp 1607194113
transform 1 0 32844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_350
timestamp 1607194113
transform 1 0 33304 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:180.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:185.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35052 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:191.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 33764 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:193.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 34040 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607194113
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_358
timestamp 1607194113
transform 1 0 34040 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_367
timestamp 1607194113
transform 1 0 34868 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_361
timestamp 1607194113
transform 1 0 34316 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_372
timestamp 1607194113
transform 1 0 35328 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:186.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36616 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:187.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 36064 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_378
timestamp 1607194113
transform 1 0 35880 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_389
timestamp 1607194113
transform 1 0 36892 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_383
timestamp 1607194113
transform 1 0 36340 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_395
timestamp 1607194113
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:188.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 37628 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607194113
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_400
timestamp 1607194113
transform 1 0 37904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_412
timestamp 1607194113
transform 1 0 39008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_398
timestamp 1607194113
transform 1 0 37720 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_410
timestamp 1607194113
transform 1 0 38824 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607194113
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_424
timestamp 1607194113
transform 1 0 40112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_428
timestamp 1607194113
transform 1 0 40480 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_422
timestamp 1607194113
transform 1 0 39928 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_434
timestamp 1607194113
transform 1 0 41032 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607194113
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_440
timestamp 1607194113
transform 1 0 41584 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_452
timestamp 1607194113
transform 1 0 42688 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_446
timestamp 1607194113
transform 1 0 42136 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_464
timestamp 1607194113
transform 1 0 43792 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_476
timestamp 1607194113
transform 1 0 44896 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_459
timestamp 1607194113
transform 1 0 43332 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_471
timestamp 1607194113
transform 1 0 44436 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607194113
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_489
timestamp 1607194113
transform 1 0 46092 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_483
timestamp 1607194113
transform 1 0 45540 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_495
timestamp 1607194113
transform 1 0 46644 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607194113
transform 1 0 48852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_501
timestamp 1607194113
transform 1 0 47196 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_513
timestamp 1607194113
transform 1 0 48300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_507
timestamp 1607194113
transform 1 0 47748 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_520
timestamp 1607194113
transform 1 0 48944 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_525
timestamp 1607194113
transform 1 0 49404 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_537
timestamp 1607194113
transform 1 0 50508 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_532
timestamp 1607194113
transform 1 0 50048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607194113
transform 1 0 51612 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_550
timestamp 1607194113
transform 1 0 51704 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_562
timestamp 1607194113
transform 1 0 52808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_544
timestamp 1607194113
transform 1 0 51152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_556
timestamp 1607194113
transform 1 0 52256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607194113
transform -1 0 54832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607194113
transform -1 0 54832 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607194113
transform 1 0 54464 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_574
timestamp 1607194113
transform 1 0 53912 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_580
timestamp 1607194113
transform 1 0 54464 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_568
timestamp 1607194113
transform 1 0 53360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:9.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607194113
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1607194113
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_14
timestamp 1607194113
transform 1 0 2392 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:10.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3128 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:12.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4140 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_25
timestamp 1607194113
transform 1 0 3404 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_36
timestamp 1607194113
transform 1 0 4416 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:14.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5152 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:20.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6164 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607194113
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1607194113
transform 1 0 5428 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1607194113
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1607194113
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:9.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:4.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_73
timestamp 1607194113
transform 1 0 7820 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:42.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_84
timestamp 1607194113
transform 1 0 8832 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1607194113
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 1607194113
transform 1 0 10304 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1607194113
transform 1 0 10672 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:47.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11408 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607194113
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1607194113
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1607194113
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_123
timestamp 1607194113
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:52.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:55.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_134
timestamp 1607194113
transform 1 0 13432 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_145
timestamp 1607194113
transform 1 0 14444 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:105.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:108.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_156
timestamp 1607194113
transform 1 0 15456 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:112.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17204 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607194113
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_167
timestamp 1607194113
transform 1 0 16468 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1607194113
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1607194113
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_184
timestamp 1607194113
transform 1 0 18032 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:117.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:10.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19780 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_195
timestamp 1607194113
transform 1 0 19044 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_206
timestamp 1607194113
transform 1 0 20056 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:13.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20792 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:14.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21804 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_217
timestamp 1607194113
transform 1 0 21068 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_228
timestamp 1607194113
transform 1 0 22080 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:16.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607194113
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_239
timestamp 1607194113
transform 1 0 23092 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1607194113
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_245
timestamp 1607194113
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 25576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:234.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24564 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_253
timestamp 1607194113
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_258
timestamp 1607194113
transform 1 0 24840 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1607194113
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:226.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27232 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_281
timestamp 1607194113
transform 1 0 26956 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_287
timestamp 1607194113
transform 1 0 27508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607194113
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_299
timestamp 1607194113
transform 1 0 28612 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_306
timestamp 1607194113
transform 1 0 29256 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 30728 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:251.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_317
timestamp 1607194113
transform 1 0 30268 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_321
timestamp 1607194113
transform 1 0 30636 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__848__CLK
timestamp 1607194113
transform 1 0 32476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_343
timestamp 1607194113
transform 1 0 32660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:190.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 35604 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607194113
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_355
timestamp 1607194113
transform 1 0 33764 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_363
timestamp 1607194113
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_367
timestamp 1607194113
transform 1 0 34868 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_378
timestamp 1607194113
transform 1 0 35880 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_390
timestamp 1607194113
transform 1 0 36984 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_402
timestamp 1607194113
transform 1 0 38088 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_414
timestamp 1607194113
transform 1 0 39192 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607194113
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_426
timestamp 1607194113
transform 1 0 40296 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_428
timestamp 1607194113
transform 1 0 40480 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_440
timestamp 1607194113
transform 1 0 41584 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_452
timestamp 1607194113
transform 1 0 42688 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_464
timestamp 1607194113
transform 1 0 43792 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_476
timestamp 1607194113
transform 1 0 44896 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607194113
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_489
timestamp 1607194113
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_501
timestamp 1607194113
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_513
timestamp 1607194113
transform 1 0 48300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_525
timestamp 1607194113
transform 1 0 49404 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_537
timestamp 1607194113
transform 1 0 50508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607194113
transform 1 0 51612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_550
timestamp 1607194113
transform 1 0 51704 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_562
timestamp 1607194113
transform 1 0 52808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607194113
transform -1 0 54832 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_574
timestamp 1607194113
transform 1 0 53912 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_580
timestamp 1607194113
transform 1 0 54464 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:7.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607194113
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1607194113
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_14
timestamp 1607194113
transform 1 0 2392 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:19.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4784 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607194113
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1607194113
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1607194113
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_32
timestamp 1607194113
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:21.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:23.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6808 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_43
timestamp 1607194113
transform 1 0 5060 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_54
timestamp 1607194113
transform 1 0 6072 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:26.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7820 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1607194113
transform 1 0 7084 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1607194113
transform 1 0 8096 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8832 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:46.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607194113
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1607194113
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1607194113
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1607194113
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_104
timestamp 1607194113
transform 1 0 10672 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:51.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11408 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:54.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 12420 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_115
timestamp 1607194113
transform 1 0 11684 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:57.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13432 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_126
timestamp 1607194113
transform 1 0 12696 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_137
timestamp 1607194113
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:111.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607194113
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1607194113
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_154
timestamp 1607194113
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_165
timestamp 1607194113
transform 1 0 16284 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:113.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 17020 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:118.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18032 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_176
timestamp 1607194113
transform 1 0 17296 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1607194113
transform 1 0 18308 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:121.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 19044 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:11.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 20056 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_198
timestamp 1607194113
transform 1 0 19320 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1607194113
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:17.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607194113
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1607194113
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1607194113
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_218
timestamp 1607194113
transform 1 0 21160 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_229
timestamp 1607194113
transform 1 0 22172 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:23.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22908 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:235.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 23920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_240
timestamp 1607194113
transform 1 0 23184 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 24656 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A
timestamp 1607194113
transform 1 0 25484 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_251
timestamp 1607194113
transform 1 0 24196 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_255
timestamp 1607194113
transform 1 0 24564 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1607194113
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:229.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 27232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607194113
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_276
timestamp 1607194113
transform 1 0 26496 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_287
timestamp 1607194113
transform 1 0 27508 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_291
timestamp 1607194113
transform 1 0 27876 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 29532 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _523_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 27968 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_301
timestamp 1607194113
transform 1 0 28796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_316
timestamp 1607194113
transform 1 0 30176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_328
timestamp 1607194113
transform 1 0 31280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1607194113
transform 1 0 32108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _511_
timestamp 1607194113
transform 1 0 33120 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607194113
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_340
timestamp 1607194113
transform 1 0 32384 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _517_
timestamp 1607194113
transform 1 0 34500 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 1607194113
transform 1 0 33764 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_370
timestamp 1607194113
transform 1 0 35144 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_382
timestamp 1607194113
transform 1 0 36248 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_394
timestamp 1607194113
transform 1 0 37352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607194113
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_398
timestamp 1607194113
transform 1 0 37720 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_410
timestamp 1607194113
transform 1 0 38824 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_422
timestamp 1607194113
transform 1 0 39928 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_434
timestamp 1607194113
transform 1 0 41032 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607194113
transform 1 0 43240 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_446
timestamp 1607194113
transform 1 0 42136 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_459
timestamp 1607194113
transform 1 0 43332 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_471
timestamp 1607194113
transform 1 0 44436 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_483
timestamp 1607194113
transform 1 0 45540 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_495
timestamp 1607194113
transform 1 0 46644 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607194113
transform 1 0 48852 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_507
timestamp 1607194113
transform 1 0 47748 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_520
timestamp 1607194113
transform 1 0 48944 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_532
timestamp 1607194113
transform 1 0 50048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_544
timestamp 1607194113
transform 1 0 51152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_556
timestamp 1607194113
transform 1 0 52256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607194113
transform -1 0 54832 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607194113
transform 1 0 54464 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_568
timestamp 1607194113
transform 1 0 53360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:6.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607194113
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1607194113
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_14
timestamp 1607194113
transform 1 0 2392 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:22.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4324 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:27.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3312 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_22
timestamp 1607194113
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_27
timestamp 1607194113
transform 1 0 3588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1607194113
transform 1 0 4600 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:24.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607194113
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_49
timestamp 1607194113
transform 1 0 5612 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1607194113
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:29.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:31.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_73
timestamp 1607194113
transform 1 0 7820 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:3.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 9568 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:5.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10580 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_84
timestamp 1607194113
transform 1 0 8832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_95
timestamp 1607194113
transform 1 0 9844 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:50.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11592 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607194113
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1607194113
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1607194113
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1607194113
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1607194113
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:56.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:60.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_134
timestamp 1607194113
transform 1 0 13432 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_145
timestamp 1607194113
transform 1 0 14444 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 16008 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:62.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15180 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_156
timestamp 1607194113
transform 1 0 15456 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607194113
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_174
timestamp 1607194113
transform 1 0 17112 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1607194113
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_184
timestamp 1607194113
transform 1 0 18032 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _841_
timestamp 1607194113
transform 1 0 19228 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:124.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__841__CLK
timestamp 1607194113
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:20.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21712 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1607194113
transform 1 0 20976 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_227
timestamp 1607194113
transform 1 0 21988 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607194113
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1607194113
transform 1 0 23092 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1607194113
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_245
timestamp 1607194113
transform 1 0 23644 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _845_
timestamp 1607194113
transform 1 0 24472 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__845__CLK
timestamp 1607194113
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_251
timestamp 1607194113
transform 1 0 24196 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _515_
timestamp 1607194113
transform 1 0 26956 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_273
timestamp 1607194113
transform 1 0 26220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_288
timestamp 1607194113
transform 1 0 27600 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607194113
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1607194113
transform 1 0 28704 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_304
timestamp 1607194113
transform 1 0 29072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_306
timestamp 1607194113
transform 1 0 29256 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 31556 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:254.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 29992 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:255.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 31004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_317
timestamp 1607194113
transform 1 0 30268 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_328
timestamp 1607194113
transform 1 0 31280 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _509_
timestamp 1607194113
transform 1 0 33488 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__B1
timestamp 1607194113
transform 1 0 32752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_346
timestamp 1607194113
transform 1 0 32936 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _521_
timestamp 1607194113
transform 1 0 34868 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607194113
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_355
timestamp 1607194113
transform 1 0 33764 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_363
timestamp 1607194113
transform 1 0 34500 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _847_
timestamp 1607194113
transform 1 0 36984 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__847__CLK
timestamp 1607194113
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_376
timestamp 1607194113
transform 1 0 35696 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_409
timestamp 1607194113
transform 1 0 38732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607194113
transform 1 0 40388 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_421
timestamp 1607194113
transform 1 0 39836 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_428
timestamp 1607194113
transform 1 0 40480 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_440
timestamp 1607194113
transform 1 0 41584 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_452
timestamp 1607194113
transform 1 0 42688 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_464
timestamp 1607194113
transform 1 0 43792 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_476
timestamp 1607194113
transform 1 0 44896 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607194113
transform 1 0 46000 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_489
timestamp 1607194113
transform 1 0 46092 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_501
timestamp 1607194113
transform 1 0 47196 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_513
timestamp 1607194113
transform 1 0 48300 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_525
timestamp 1607194113
transform 1 0 49404 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_537
timestamp 1607194113
transform 1 0 50508 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607194113
transform 1 0 51612 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_550
timestamp 1607194113
transform 1 0 51704 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_562
timestamp 1607194113
transform 1 0 52808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607194113
transform -1 0 54832 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_574
timestamp 1607194113
transform 1 0 53912 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_580
timestamp 1607194113
transform 1 0 54464 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:14.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2852 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607194113
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607194113
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1607194113
transform 1 0 2484 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4784 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607194113
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1607194113
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1607194113
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1607194113
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:25.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:28.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_43
timestamp 1607194113
transform 1 0 5060 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_54
timestamp 1607194113
transform 1 0 6072 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:3.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7820 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_65
timestamp 1607194113
transform 1 0 7084 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 1607194113
transform 1 0 8096 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 9660 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:30.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8832 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607194113
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1607194113
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1607194113
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _752_
timestamp 1607194113
transform 1 0 12420 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_18_107
timestamp 1607194113
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1607194113
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__752__B2
timestamp 1607194113
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_139
timestamp 1607194113
transform 1 0 13892 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:116.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607194113
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1607194113
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_154
timestamp 1607194113
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1607194113
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _534_
timestamp 1607194113
transform 1 0 16468 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__B1
timestamp 1607194113
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_182
timestamp 1607194113
transform 1 0 17848 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _536_
timestamp 1607194113
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_194
timestamp 1607194113
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1607194113
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _533_
timestamp 1607194113
transform 1 0 20884 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607194113
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__844__CLK
timestamp 1607194113
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_222
timestamp 1607194113
transform 1 0 21528 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _844_
timestamp 1607194113
transform 1 0 22264 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_18_249
timestamp 1607194113
transform 1 0 24012 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _525_
timestamp 1607194113
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1607194113
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1607194113
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _528_
timestamp 1607194113
transform 1 0 26496 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607194113
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_283
timestamp 1607194113
transform 1 0 27140 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_291
timestamp 1607194113
transform 1 0 27876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _524_
timestamp 1607194113
transform 1 0 28152 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1607194113
transform 1 0 28980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_305
timestamp 1607194113
transform 1 0 29164 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 30452 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_317
timestamp 1607194113
transform 1 0 30268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_328
timestamp 1607194113
transform 1 0 31280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _519_
timestamp 1607194113
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607194113
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_349
timestamp 1607194113
transform 1 0 33212 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1607194113
transform 1 0 34132 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _522_
timestamp 1607194113
transform 1 0 35144 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1607194113
transform 1 0 34408 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_357
timestamp 1607194113
transform 1 0 33948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_364
timestamp 1607194113
transform 1 0 34592 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1607194113
transform 1 0 35972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_381
timestamp 1607194113
transform 1 0 36156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_393
timestamp 1607194113
transform 1 0 37260 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _837_
timestamp 1607194113
transform 1 0 39376 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607194113
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_398
timestamp 1607194113
transform 1 0 37720 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_410
timestamp 1607194113
transform 1 0 38824 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__837__CLK
timestamp 1607194113
transform 1 0 41124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_437
timestamp 1607194113
transform 1 0 41308 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607194113
transform 1 0 43240 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__864__CLK
timestamp 1607194113
transform 1 0 43056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_449
timestamp 1607194113
transform 1 0 42412 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_455
timestamp 1607194113
transform 1 0 42964 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _864_
timestamp 1607194113
transform 1 0 43332 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_478
timestamp 1607194113
transform 1 0 45080 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_490
timestamp 1607194113
transform 1 0 46184 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607194113
transform 1 0 48852 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_502
timestamp 1607194113
transform 1 0 47288 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_514
timestamp 1607194113
transform 1 0 48392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_518
timestamp 1607194113
transform 1 0 48760 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_520
timestamp 1607194113
transform 1 0 48944 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_532
timestamp 1607194113
transform 1 0 50048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_544
timestamp 1607194113
transform 1 0 51152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_556
timestamp 1607194113
transform 1 0 52256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607194113
transform -1 0 54832 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607194113
transform 1 0 54464 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_568
timestamp 1607194113
transform 1 0 53360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:10.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:12.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2208 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607194113
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607194113
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1607194113
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1607194113
transform 1 0 2116 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1607194113
transform 1 0 2484 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1607194113
transform 1 0 1380 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_14
timestamp 1607194113
transform 1 0 2392 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _755_
timestamp 1607194113
transform 1 0 4324 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:13.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:8.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607194113
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_26
timestamp 1607194113
transform 1 0 3496 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_37
timestamp 1607194113
transform 1 0 4508 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1607194113
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1607194113
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1607194113
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _754_
timestamp 1607194113
transform 1 0 6808 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5244 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607194113
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_48
timestamp 1607194113
transform 1 0 5520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1607194113
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_49
timestamp 1607194113
transform 1 0 5612 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1607194113
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _775_
timestamp 1607194113
transform 1 0 6900 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__775__CLK
timestamp 1607194113
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_76
timestamp 1607194113
transform 1 0 8096 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1607194113
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _776_
timestamp 1607194113
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607194113
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_87
timestamp 1607194113
transform 1 0 9108 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_99
timestamp 1607194113
transform 1 0 10212 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1607194113
transform 1 0 10580 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1607194113
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _777_
timestamp 1607194113
transform 1 0 12144 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:58.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607194113
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__776__CLK
timestamp 1607194113
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1607194113
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1607194113
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_114
timestamp 1607194113
transform 1 0 11592 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1607194113
transform 1 0 12972 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__777__CLK
timestamp 1607194113
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_132
timestamp 1607194113
transform 1 0 13248 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_143
timestamp 1607194113
transform 1 0 14260 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1607194113
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _842_
timestamp 1607194113
transform 1 0 15088 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:123.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607194113
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__842__CLK
timestamp 1607194113
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1607194113
transform 1 0 14812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1607194113
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1607194113
transform 1 0 16284 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1607194113
transform 1 0 16652 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _532_
timestamp 1607194113
transform 1 0 17848 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607194113
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1607194113
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_184
timestamp 1607194113
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_172
timestamp 1607194113
transform 1 0 16928 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1607194113
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _432_
timestamp 1607194113
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _537_
timestamp 1607194113
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:128.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__A
timestamp 1607194113
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_195
timestamp 1607194113
transform 1 0 19044 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_189
timestamp 1607194113
transform 1 0 18492 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1607194113
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _840_
timestamp 1607194113
transform 1 0 20976 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:249.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607194113
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__840__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_209
timestamp 1607194113
transform 1 0 20332 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1607194113
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_223
timestamp 1607194113
transform 1 0 21620 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1607194113
transform 1 0 20884 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _434_
timestamp 1607194113
transform 1 0 23828 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:244.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22356 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607194113
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_234
timestamp 1607194113
transform 1 0 22632 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1607194113
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1607194113
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_235
timestamp 1607194113
transform 1 0 22724 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_247
timestamp 1607194113
transform 1 0 23828 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _529_
timestamp 1607194113
transform 1 0 25208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 24380 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__B1
timestamp 1607194113
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_254
timestamp 1607194113
transform 1 0 24472 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_269
timestamp 1607194113
transform 1 0 25852 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _422_
timestamp 1607194113
transform 1 0 27784 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1607194113
transform 1 0 26772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _433_
timestamp 1607194113
transform 1 0 26496 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607194113
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__A
timestamp 1607194113
transform 1 0 26036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1607194113
transform 1 0 26220 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_282
timestamp 1607194113
transform 1 0 27048 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_283
timestamp 1607194113
transform 1 0 27140 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_291
timestamp 1607194113
transform 1 0 27876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _513_
timestamp 1607194113
transform 1 0 29532 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__dfxtp_4  _846_
timestamp 1607194113
transform 1 0 28152 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607194113
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_297
timestamp 1607194113
transform 1 0 28428 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_306
timestamp 1607194113
transform 1 0 29256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1607194113
transform 1 0 31004 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _508_
timestamp 1607194113
transform 1 0 31740 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__B1
timestamp 1607194113
transform 1 0 30820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__846__CLK
timestamp 1607194113
transform 1 0 29900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1607194113
transform 1 0 31004 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_315
timestamp 1607194113
transform 1 0 30084 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_323
timestamp 1607194113
transform 1 0 30820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_328
timestamp 1607194113
transform 1 0 31280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _436_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 32108 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _510_
timestamp 1607194113
transform 1 0 33396 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607194113
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_340
timestamp 1607194113
transform 1 0 32384 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_348
timestamp 1607194113
transform 1 0 33120 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_346
timestamp 1607194113
transform 1 0 32936 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _512_
timestamp 1607194113
transform 1 0 34224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _850_
timestamp 1607194113
transform 1 0 35052 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607194113
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_358
timestamp 1607194113
transform 1 0 34040 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_367
timestamp 1607194113
transform 1 0 34868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_358
timestamp 1607194113
transform 1 0 34040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_369
timestamp 1607194113
transform 1 0 35052 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _504_
timestamp 1607194113
transform 1 0 35972 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__850__CLK
timestamp 1607194113
transform 1 0 36800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_390
timestamp 1607194113
transform 1 0 36984 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_377
timestamp 1607194113
transform 1 0 35788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_386
timestamp 1607194113
transform 1 0 36616 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_394
timestamp 1607194113
transform 1 0 37352 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 1607194113
transform 1 0 37536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 38824 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _852_
timestamp 1607194113
transform 1 0 37904 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607194113
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_399
timestamp 1607194113
transform 1 0 37812 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_407
timestamp 1607194113
transform 1 0 38548 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_398
timestamp 1607194113
transform 1 0 37720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_421
timestamp 1607194113
transform 1 0 39836 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_423
timestamp 1607194113
transform 1 0 40020 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__852__CLK
timestamp 1607194113
transform 1 0 39652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__B
timestamp 1607194113
transform 1 0 39836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1607194113
transform 1 0 39652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_429
timestamp 1607194113
transform 1 0 40572 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_428
timestamp 1607194113
transform 1 0 40480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__A
timestamp 1607194113
transform 1 0 41032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607194113
transform 1 0 40388 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 40664 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _463_
timestamp 1607194113
transform 1 0 40848 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_436
timestamp 1607194113
transform 1 0 41216 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_436
timestamp 1607194113
transform 1 0 41216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _481_
timestamp 1607194113
transform 1 0 41952 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _520_
timestamp 1607194113
transform 1 0 41768 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607194113
transform 1 0 43240 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__A
timestamp 1607194113
transform 1 0 41584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__A
timestamp 1607194113
transform 1 0 42320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_446
timestamp 1607194113
transform 1 0 42136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_458
timestamp 1607194113
transform 1 0 43240 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_450
timestamp 1607194113
transform 1 0 42504 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _465_
timestamp 1607194113
transform 1 0 43792 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_4  _466_
timestamp 1607194113
transform 1 0 43608 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__B1
timestamp 1607194113
transform 1 0 43608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_477
timestamp 1607194113
transform 1 0 44988 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_459
timestamp 1607194113
transform 1 0 43332 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_474
timestamp 1607194113
transform 1 0 44712 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_487
timestamp 1607194113
transform 1 0 45908 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_489
timestamp 1607194113
transform 1 0 46092 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_485
timestamp 1607194113
transform 1 0 45724 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1607194113
transform 1 0 45724 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607194113
transform 1 0 46000 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1607194113
transform 1 0 45448 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_495
timestamp 1607194113
transform 1 0 46644 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_493
timestamp 1607194113
transform 1 0 46460 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _467_
timestamp 1607194113
transform 1 0 46920 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _462_
timestamp 1607194113
transform 1 0 46552 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _863_
timestamp 1607194113
transform 1 0 47932 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607194113
transform 1 0 48852 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__863__CLK
timestamp 1607194113
transform 1 0 47748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_501
timestamp 1607194113
transform 1 0 47196 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_507
timestamp 1607194113
transform 1 0 47748 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_520
timestamp 1607194113
transform 1 0 48944 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _861_
timestamp 1607194113
transform 1 0 50048 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__861__CLK
timestamp 1607194113
transform 1 0 49864 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_528
timestamp 1607194113
transform 1 0 49680 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_540
timestamp 1607194113
transform 1 0 50784 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_528
timestamp 1607194113
transform 1 0 49680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607194113
transform 1 0 51612 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_548
timestamp 1607194113
transform 1 0 51520 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_550
timestamp 1607194113
transform 1 0 51704 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_562
timestamp 1607194113
transform 1 0 52808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_551
timestamp 1607194113
transform 1 0 51796 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607194113
transform -1 0 54832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607194113
transform -1 0 54832 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607194113
transform 1 0 54464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_574
timestamp 1607194113
transform 1 0 53912 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_580
timestamp 1607194113
transform 1 0 54464 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_563
timestamp 1607194113
transform 1 0 52900 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_575
timestamp 1607194113
transform 1 0 54004 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_579
timestamp 1607194113
transform 1 0 54372 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:11.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607194113
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1607194113
transform 1 0 1380 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_14
timestamp 1607194113
transform 1 0 2392 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:15.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:16.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4232 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_22
timestamp 1607194113
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_26
timestamp 1607194113
transform 1 0 3496 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_37
timestamp 1607194113
transform 1 0 4508 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _592_
timestamp 1607194113
transform 1 0 5336 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607194113
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_45
timestamp 1607194113
transform 1 0 5244 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_49
timestamp 1607194113
transform 1 0 5612 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1607194113
transform 1 0 6808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _588_
timestamp 1607194113
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:5.g_subtaps:32.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1607194113
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1607194113
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:59.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 9752 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_90
timestamp 1607194113
transform 1 0 9384 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_97
timestamp 1607194113
transform 1 0 10028 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:61.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10764 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607194113
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_108
timestamp 1607194113
transform 1 0 11040 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1607194113
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1607194113
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _783_
timestamp 1607194113
transform 1 0 13248 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1607194113
transform 1 0 13156 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15732 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__783__CLK
timestamp 1607194113
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_153
timestamp 1607194113
transform 1 0 15180 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607194113
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1607194113
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_184
timestamp 1607194113
transform 1 0 18032 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _538_
timestamp 1607194113
transform 1 0 19228 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_195
timestamp 1607194113
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_206
timestamp 1607194113
transform 1 0 20056 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _539_
timestamp 1607194113
transform 1 0 20792 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A
timestamp 1607194113
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1607194113
transform 1 0 21804 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:248.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607194113
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_236
timestamp 1607194113
transform 1 0 22816 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_245
timestamp 1607194113
transform 1 0 23644 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _531_
timestamp 1607194113
transform 1 0 24196 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _648_
timestamp 1607194113
transform 1 0 25208 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__A1_N
timestamp 1607194113
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_254
timestamp 1607194113
transform 1 0 24472 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_278
timestamp 1607194113
transform 1 0 26680 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_290
timestamp 1607194113
transform 1 0 27784 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _500_
timestamp 1607194113
transform 1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _514_
timestamp 1607194113
transform 1 0 28152 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607194113
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_297
timestamp 1607194113
transform 1 0 28428 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_309
timestamp 1607194113
transform 1 0 29532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _851_
timestamp 1607194113
transform 1 0 31188 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_21_321
timestamp 1607194113
transform 1 0 30636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__851__CLK
timestamp 1607194113
transform 1 0 32936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_348
timestamp 1607194113
transform 1 0 33120 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_354
timestamp 1607194113
transform 1 0 33672 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1607194113
transform 1 0 33764 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _501_
timestamp 1607194113
transform 1 0 35236 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607194113
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1607194113
transform 1 0 34040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_360
timestamp 1607194113
transform 1 0 34224 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_367
timestamp 1607194113
transform 1 0 34868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _505_
timestamp 1607194113
transform 1 0 37352 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_378
timestamp 1607194113
transform 1 0 35880 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_390
timestamp 1607194113
transform 1 0 36984 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1607194113
transform 1 0 39376 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__A
timestamp 1607194113
transform 1 0 39192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_403
timestamp 1607194113
transform 1 0 38180 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_411
timestamp 1607194113
transform 1 0 38916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _450_
timestamp 1607194113
transform 1 0 41216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607194113
transform 1 0 40388 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_419
timestamp 1607194113
transform 1 0 39652 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_428
timestamp 1607194113
transform 1 0 40480 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _857_
timestamp 1607194113
transform 1 0 42320 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__857__CLK
timestamp 1607194113
transform 1 0 42136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_440
timestamp 1607194113
transform 1 0 41584 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _395_
timestamp 1607194113
transform 1 0 44804 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1607194113
transform 1 0 44620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_467
timestamp 1607194113
transform 1 0 44068 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_479
timestamp 1607194113
transform 1 0 45172 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _396_
timestamp 1607194113
transform 1 0 46092 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607194113
transform 1 0 46000 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1607194113
transform 1 0 46460 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_487
timestamp 1607194113
transform 1 0 45908 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_495
timestamp 1607194113
transform 1 0 46644 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _468_
timestamp 1607194113
transform 1 0 47196 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_510
timestamp 1607194113
transform 1 0 48024 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1607194113
transform 1 0 50600 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 1607194113
transform 1 0 49588 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_522
timestamp 1607194113
transform 1 0 49128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_526
timestamp 1607194113
transform 1 0 49496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_530
timestamp 1607194113
transform 1 0 49864 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_541
timestamp 1607194113
transform 1 0 50876 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _470_
timestamp 1607194113
transform 1 0 51704 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607194113
transform 1 0 51612 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__A
timestamp 1607194113
transform 1 0 52348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_559
timestamp 1607194113
transform 1 0 52532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607194113
transform -1 0 54832 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_571
timestamp 1607194113
transform 1 0 53636 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_579
timestamp 1607194113
transform 1 0 54372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2208 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607194113
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1607194113
transform 1 0 1380 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1607194113
transform 1 0 2116 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp 1607194113
transform 1 0 2484 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _774_
timestamp 1607194113
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:3.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3220 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607194113
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_26
timestamp 1607194113
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1607194113
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:5.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__774__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_53
timestamp 1607194113
transform 1 0 5980 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_62
timestamp 1607194113
transform 1 0 6808 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:63.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:9.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7544 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1607194113
transform 1 0 7820 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _740_
timestamp 1607194113
transform 1 0 10580 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607194113
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__740__B1
timestamp 1607194113
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1607194113
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1607194113
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_119
timestamp 1607194113
transform 1 0 12052 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:119.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 12788 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:122.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 13800 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1607194113
transform 1 0 13064 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1607194113
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _591_
timestamp 1607194113
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607194113
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_157
timestamp 1607194113
transform 1 0 15548 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1607194113
transform 1 0 16284 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _839_
timestamp 1607194113
transform 1 0 16560 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__839__CLK
timestamp 1607194113
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _541_
timestamp 1607194113
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1607194113
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_189
timestamp 1607194113
transform 1 0 18492 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1607194113
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _543_
timestamp 1607194113
transform 1 0 21804 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607194113
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1607194113
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_223
timestamp 1607194113
transform 1 0 21620 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _542_
timestamp 1607194113
transform 1 0 23368 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1607194113
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1607194113
transform 1 0 24012 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_236
timestamp 1607194113
transform 1 0 22816 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _527_
timestamp 1607194113
transform 1 0 25116 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_251
timestamp 1607194113
transform 1 0 24196 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_259
timestamp 1607194113
transform 1 0 24932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_264
timestamp 1607194113
transform 1 0 25392 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1607194113
transform 1 0 26496 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _849_
timestamp 1607194113
transform 1 0 27784 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607194113
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_272
timestamp 1607194113
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_279
timestamp 1607194113
transform 1 0 26772 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_287
timestamp 1607194113
transform 1 0 27508 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__849__CLK
timestamp 1607194113
transform 1 0 29532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_311
timestamp 1607194113
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _496_
timestamp 1607194113
transform 1 0 31004 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_323
timestamp 1607194113
transform 1 0 30820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_328
timestamp 1607194113
transform 1 0 31280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _506_
timestamp 1607194113
transform 1 0 33028 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607194113
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_337
timestamp 1607194113
transform 1 0 32108 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_345
timestamp 1607194113
transform 1 0 32844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _437_
timestamp 1607194113
transform 1 0 35236 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__B1
timestamp 1607194113
transform 1 0 34316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_363
timestamp 1607194113
transform 1 0 34500 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_380
timestamp 1607194113
transform 1 0 36064 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_392
timestamp 1607194113
transform 1 0 37168 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _503_
timestamp 1607194113
transform 1 0 37720 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607194113
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__A
timestamp 1607194113
transform 1 0 38364 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_396
timestamp 1607194113
transform 1 0 37536 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_407
timestamp 1607194113
transform 1 0 38548 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _482_
timestamp 1607194113
transform 1 0 41124 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1607194113
transform 1 0 40112 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_419
timestamp 1607194113
transform 1 0 39652 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_423
timestamp 1607194113
transform 1 0 40020 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_427
timestamp 1607194113
transform 1 0 40388 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607194113
transform 1 0 43240 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_442
timestamp 1607194113
transform 1 0 41768 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_454
timestamp 1607194113
transform 1 0 42872 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1607194113
transform 1 0 43976 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1607194113
transform 1 0 44252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_459
timestamp 1607194113
transform 1 0 43332 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_465
timestamp 1607194113
transform 1 0 43884 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_471
timestamp 1607194113
transform 1 0 44436 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _460_
timestamp 1607194113
transform 1 0 47012 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _461_
timestamp 1607194113
transform 1 0 45632 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_22_483
timestamp 1607194113
transform 1 0 45540 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_491
timestamp 1607194113
transform 1 0 46276 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607194113
transform 1 0 48852 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_506
timestamp 1607194113
transform 1 0 47656 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_518
timestamp 1607194113
transform 1 0 48760 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_520
timestamp 1607194113
transform 1 0 48944 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _472_
timestamp 1607194113
transform 1 0 49036 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_22_535
timestamp 1607194113
transform 1 0 50324 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _862_
timestamp 1607194113
transform 1 0 51980 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__862__CLK
timestamp 1607194113
transform 1 0 51796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_547
timestamp 1607194113
transform 1 0 51428 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607194113
transform -1 0 54832 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607194113
transform 1 0 54464 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_572
timestamp 1607194113
transform 1 0 53728 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607194113
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1607194113
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_14
timestamp 1607194113
transform 1 0 2392 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_4  _756_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3128 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_23_39
timestamp 1607194113
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _743_
timestamp 1607194113
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:4.g_subtaps:4.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607194113
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__743__B1
timestamp 1607194113
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_50
timestamp 1607194113
transform 1 0 5704 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_58
timestamp 1607194113
transform 1 0 6440 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_78
timestamp 1607194113
transform 1 0 8280 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _741_
timestamp 1607194113
transform 1 0 9016 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__741__B1
timestamp 1607194113
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1607194113
transform 1 0 10488 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _730_
timestamp 1607194113
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:125.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607194113
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__730__B1
timestamp 1607194113
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_110
timestamp 1607194113
transform 1 0 11224 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_114
timestamp 1607194113
transform 1 0 11592 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_139
timestamp 1607194113
transform 1 0 13892 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:127.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14628 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 15640 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_150
timestamp 1607194113
transform 1 0 14904 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_161
timestamp 1607194113
transform 1 0 15916 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:3.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 16652 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607194113
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1607194113
transform 1 0 16928 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1607194113
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1607194113
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _429_
timestamp 1607194113
transform 1 0 19504 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:30.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1607194113
transform 1 0 19044 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1607194113
transform 1 0 19412 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_207
timestamp 1607194113
transform 1 0 20148 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 22172 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1607194113
transform 1 0 20884 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_218
timestamp 1607194113
transform 1 0 21160 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_226
timestamp 1607194113
transform 1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607194113
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1607194113
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_238
timestamp 1607194113
transform 1 0 23000 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_245
timestamp 1607194113
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _843_
timestamp 1607194113
transform 1 0 24840 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:253.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__843__CLK
timestamp 1607194113
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1607194113
transform 1 0 27508 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1607194113
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_285
timestamp 1607194113
transform 1 0 27324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_290
timestamp 1607194113
transform 1 0 27784 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607194113
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_302
timestamp 1607194113
transform 1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_306
timestamp 1607194113
transform 1 0 29256 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _499_
timestamp 1607194113
transform 1 0 30084 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__B1
timestamp 1607194113
transform 1 0 31372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_314
timestamp 1607194113
transform 1 0 29992 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_331
timestamp 1607194113
transform 1 0 31556 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1607194113
transform 1 0 33488 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _489_
timestamp 1607194113
transform 1 0 32108 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1607194113
transform 1 0 33304 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_344
timestamp 1607194113
transform 1 0 32752 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _491_
timestamp 1607194113
transform 1 0 34960 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607194113
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_355
timestamp 1607194113
transform 1 0 33764 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_363
timestamp 1607194113
transform 1 0 34500 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_367
timestamp 1607194113
transform 1 0 34868 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_375
timestamp 1607194113
transform 1 0 35604 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _438_
timestamp 1607194113
transform 1 0 36340 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_392
timestamp 1607194113
transform 1 0 37168 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _492_
timestamp 1607194113
transform 1 0 38272 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1607194113
transform 1 0 40480 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607194113
transform 1 0 40388 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__B1
timestamp 1607194113
transform 1 0 39468 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_419
timestamp 1607194113
transform 1 0 39652 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_431
timestamp 1607194113
transform 1 0 40756 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _487_
timestamp 1607194113
transform 1 0 41492 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_23_453
timestamp 1607194113
transform 1 0 42780 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1607194113
transform 1 0 44988 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1607194113
transform 1 0 43700 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_461
timestamp 1607194113
transform 1 0 43516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_466
timestamp 1607194113
transform 1 0 43976 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_474
timestamp 1607194113
transform 1 0 44712 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _441_
timestamp 1607194113
transform 1 0 46920 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607194113
transform 1 0 46000 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1607194113
transform 1 0 45264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_482
timestamp 1607194113
transform 1 0 45448 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_489
timestamp 1607194113
transform 1 0 46092 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_497
timestamp 1607194113
transform 1 0 46828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_507
timestamp 1607194113
transform 1 0 47748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_519
timestamp 1607194113
transform 1 0 48852 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1607194113
transform 1 0 49220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475_
timestamp 1607194113
transform 1 0 50508 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_526
timestamp 1607194113
transform 1 0 49496 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_534
timestamp 1607194113
transform 1 0 50232 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_540
timestamp 1607194113
transform 1 0 50784 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _471_
timestamp 1607194113
transform 1 0 51704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607194113
transform 1 0 51612 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_548
timestamp 1607194113
transform 1 0 51520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_559
timestamp 1607194113
transform 1 0 52532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607194113
transform -1 0 54832 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_571
timestamp 1607194113
transform 1 0 53636 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_579
timestamp 1607194113
transform 1 0 54372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:3.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607194113
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1607194113
transform 1 0 1380 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_14
timestamp 1607194113
transform 1 0 2392 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:5.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:6.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4784 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607194113
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_25
timestamp 1607194113
transform 1 0 3404 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_32
timestamp 1607194113
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _744_
timestamp 1607194113
transform 1 0 5336 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__744__B1
timestamp 1607194113
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_43
timestamp 1607194113
transform 1 0 5060 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_62
timestamp 1607194113
transform 1 0 6808 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _593_
timestamp 1607194113
transform 1 0 7544 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:6.g_subtaps:64.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10396 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607194113
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_84
timestamp 1607194113
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_93
timestamp 1607194113
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_104
timestamp 1607194113
transform 1 0 10672 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _729_
timestamp 1607194113
transform 1 0 11868 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 11408 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__729__B1
timestamp 1607194113
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:126.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14076 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__729__A1_N
timestamp 1607194113
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_135
timestamp 1607194113
transform 1 0 13524 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1607194113
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1607194113
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607194113
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1607194113
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_157
timestamp 1607194113
transform 1 0 15548 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _786_
timestamp 1607194113
transform 1 0 16744 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_169
timestamp 1607194113
transform 1 0 16652 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _540_
timestamp 1607194113
transform 1 0 19320 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__786__CLK
timestamp 1607194113
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_191
timestamp 1607194113
transform 1 0 18676 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1607194113
transform 1 0 19228 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_205
timestamp 1607194113
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1607194113
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _838_
timestamp 1607194113
transform 1 0 21896 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607194113
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__838__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1607194113
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_218
timestamp 1607194113
transform 1 0 21160 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1607194113
transform 1 0 23644 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:256.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 24380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_delay_line.g_taps:8.g_subtaps:256.inst_tap.g_clkbuf_1.dly_A
timestamp 1607194113
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_256
timestamp 1607194113
transform 1 0 24656 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_268
timestamp 1607194113
transform 1 0 25760 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _853_
timestamp 1607194113
transform 1 0 27876 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607194113
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1607194113
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1607194113
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_288
timestamp 1607194113
transform 1 0 27600 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__853__CLK
timestamp 1607194113
transform 1 0 29624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_312
timestamp 1607194113
transform 1 0 29808 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1607194113
transform 1 0 30360 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1607194113
transform 1 0 30636 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_333
timestamp 1607194113
transform 1 0 31740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _413_
timestamp 1607194113
transform 1 0 32292 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _490_
timestamp 1607194113
transform 1 0 33672 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607194113
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_337
timestamp 1607194113
transform 1 0 32108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_346
timestamp 1607194113
transform 1 0 32936 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _494_
timestamp 1607194113
transform 1 0 35420 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_361
timestamp 1607194113
transform 1 0 34316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_382
timestamp 1607194113
transform 1 0 36248 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_394
timestamp 1607194113
transform 1 0 37352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _493_
timestamp 1607194113
transform 1 0 38180 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607194113
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_398
timestamp 1607194113
transform 1 0 37720 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_402
timestamp 1607194113
transform 1 0 38088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_415
timestamp 1607194113
transform 1 0 39284 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _485_
timestamp 1607194113
transform 1 0 40296 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_24_423
timestamp 1607194113
transform 1 0 40020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_433
timestamp 1607194113
transform 1 0 40940 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _486_
timestamp 1607194113
transform 1 0 41676 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607194113
transform 1 0 43240 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_450
timestamp 1607194113
transform 1 0 42504 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _858_
timestamp 1607194113
transform 1 0 44068 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__858__CLK
timestamp 1607194113
transform 1 0 43884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_459
timestamp 1607194113
transform 1 0 43332 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _404_
timestamp 1607194113
transform 1 0 46736 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_24_486
timestamp 1607194113
transform 1 0 45816 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_494
timestamp 1607194113
transform 1 0 46552 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _440_
timestamp 1607194113
transform 1 0 48944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607194113
transform 1 0 48852 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_503
timestamp 1607194113
transform 1 0 47380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_515
timestamp 1607194113
transform 1 0 48484 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_529
timestamp 1607194113
transform 1 0 49772 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_541
timestamp 1607194113
transform 1 0 50876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _476_
timestamp 1607194113
transform 1 0 51152 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__A
timestamp 1607194113
transform 1 0 51796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_553
timestamp 1607194113
transform 1 0 51980 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607194113
transform -1 0 54832 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607194113
transform 1 0 54464 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_565
timestamp 1607194113
transform 1 0 53084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_577
timestamp 1607194113
transform 1 0 54188 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _773_
timestamp 1607194113
transform 1 0 2116 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607194113
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1607194113
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _596_
timestamp 1607194113
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__773__CLK
timestamp 1607194113
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_32
timestamp 1607194113
transform 1 0 4048 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_41
timestamp 1607194113
transform 1 0 4876 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:7.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5612 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607194113
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_52
timestamp 1607194113
transform 1 0 5888 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1607194113
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1607194113
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _589_
timestamp 1607194113
transform 1 0 8556 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _739_
timestamp 1607194113
transform 1 0 7084 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1607194113
transform 1 0 7452 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:7.g_subtaps:4.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 10580 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__A1
timestamp 1607194113
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_delay_line.g_taps:7.g_subtaps:4.inst_tap.g_clkbuf_1.dly_A
timestamp 1607194113
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1607194113
transform 1 0 10028 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607194113
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_106
timestamp 1607194113
transform 1 0 10856 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1607194113
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1607194113
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _784_
timestamp 1607194113
transform 1 0 13248 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1607194113
transform 1 0 13156 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _726_
timestamp 1607194113
transform 1 0 15732 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__726__B1
timestamp 1607194113
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__784__CLK
timestamp 1607194113
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1607194113
transform 1 0 15180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607194113
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1607194113
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_184
timestamp 1607194113
transform 1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _649_
timestamp 1607194113
transform 1 0 19136 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:4.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_delay_line.g_taps:8.g_subtaps:4.inst_tap.g_clkbuf_1.dly_A
timestamp 1607194113
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_195
timestamp 1607194113
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _676_
timestamp 1607194113
transform 1 0 21344 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_212
timestamp 1607194113
transform 1 0 20608 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607194113
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_236
timestamp 1607194113
transform 1 0 22816 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1607194113
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _647_
timestamp 1607194113
transform 1 0 24472 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_253
timestamp 1607194113
transform 1 0 24380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1607194113
transform 1 0 25944 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _650_
timestamp 1607194113
transform 1 0 26680 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_287
timestamp 1607194113
transform 1 0 27508 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1607194113
transform 1 0 29256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607194113
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_299
timestamp 1607194113
transform 1 0 28612 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_309
timestamp 1607194113
transform 1 0 29532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _497_
timestamp 1607194113
transform 1 0 31004 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_321
timestamp 1607194113
transform 1 0 30636 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_332
timestamp 1607194113
transform 1 0 31648 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _498_
timestamp 1607194113
transform 1 0 32384 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1607194113
transform 1 0 33212 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _495_
timestamp 1607194113
transform 1 0 35420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607194113
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_361
timestamp 1607194113
transform 1 0 34316 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_365
timestamp 1607194113
transform 1 0 34684 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_367
timestamp 1607194113
transform 1 0 34868 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_382
timestamp 1607194113
transform 1 0 36248 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_394
timestamp 1607194113
transform 1 0 37352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1607194113
transform 1 0 39100 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_406
timestamp 1607194113
transform 1 0 38456 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_412
timestamp 1607194113
transform 1 0 39008 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_416
timestamp 1607194113
transform 1 0 39376 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607194113
transform 1 0 40388 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_424
timestamp 1607194113
transform 1 0 40112 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_428
timestamp 1607194113
transform 1 0 40480 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _439_
timestamp 1607194113
transform 1 0 43240 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _484_
timestamp 1607194113
transform 1 0 41860 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_25_440
timestamp 1607194113
transform 1 0 41584 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_450
timestamp 1607194113
transform 1 0 42504 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_467
timestamp 1607194113
transform 1 0 44068 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_479
timestamp 1607194113
transform 1 0 45172 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607194113
transform 1 0 46000 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_487
timestamp 1607194113
transform 1 0 45908 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_489
timestamp 1607194113
transform 1 0 46092 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _479_
timestamp 1607194113
transform 1 0 47564 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_25_501
timestamp 1607194113
transform 1 0 47196 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_519
timestamp 1607194113
transform 1 0 48852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _474_
timestamp 1607194113
transform 1 0 49588 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_534
timestamp 1607194113
transform 1 0 50232 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _860_
timestamp 1607194113
transform 1 0 52072 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607194113
transform 1 0 51612 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__860__CLK
timestamp 1607194113
transform 1 0 51888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_546
timestamp 1607194113
transform 1 0 51336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_550
timestamp 1607194113
transform 1 0 51704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607194113
transform -1 0 54832 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_573
timestamp 1607194113
transform 1 0 53820 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:2.g_subtaps:4.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607194113
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607194113
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607194113
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1607194113
transform 1 0 2484 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1607194113
transform 1 0 2852 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1607194113
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_14
timestamp 1607194113
transform 1 0 2392 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _757_
timestamp 1607194113
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _758_
timestamp 1607194113
transform 1 0 3588 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3128 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:4.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3588 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607194113
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1607194113
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_35
timestamp 1607194113
transform 1 0 4324 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_25
timestamp 1607194113
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _745_
timestamp 1607194113
transform 1 0 5612 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607194113
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__745__B1
timestamp 1607194113
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_43
timestamp 1607194113
transform 1 0 5060 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_55
timestamp 1607194113
transform 1 0 6164 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_62
timestamp 1607194113
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _597_
timestamp 1607194113
transform 1 0 7084 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:3.g_subtaps:8.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 7820 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_65
timestamp 1607194113
transform 1 0 7084 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_76
timestamp 1607194113
transform 1 0 8096 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_79
timestamp 1607194113
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _581_
timestamp 1607194113
transform 1 0 10488 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _585_
timestamp 1607194113
transform 1 0 9752 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607194113
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1607194113
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_93
timestamp 1607194113
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_101
timestamp 1607194113
transform 1 0 10396 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_91
timestamp 1607194113
transform 1 0 9476 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607194113
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_116
timestamp 1607194113
transform 1 0 11776 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_108
timestamp 1607194113
transform 1 0 11040 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1607194113
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_123
timestamp 1607194113
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _595_
timestamp 1607194113
transform 1 0 13340 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _782_
timestamp 1607194113
transform 1 0 12696 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk_i
timestamp 1607194113
transform 1 0 14352 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__782__CLK
timestamp 1607194113
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_128
timestamp 1607194113
transform 1 0 12880 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_132
timestamp 1607194113
transform 1 0 13248 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_136
timestamp 1607194113
transform 1 0 13616 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _727_
timestamp 1607194113
transform 1 0 15272 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _785_
timestamp 1607194113
transform 1 0 16192 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607194113
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__727__B1
timestamp 1607194113
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__785__CLK
timestamp 1607194113
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_147
timestamp 1607194113
transform 1 0 14628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1607194113
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1607194113
transform 1 0 14628 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 1607194113
transform 1 0 14996 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607194113
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_183
timestamp 1607194113
transform 1 0 17940 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_170
timestamp 1607194113
transform 1 0 16744 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1607194113
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_184
timestamp 1607194113
transform 1 0 18032 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1607194113
transform 1 0 19320 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _667_
timestamp 1607194113
transform 1 0 18860 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk_i
timestamp 1607194113
transform 1 0 18676 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_194
timestamp 1607194113
transform 1 0 18952 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1607194113
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_192
timestamp 1607194113
transform 1 0 18768 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1607194113
transform 1 0 21068 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _655_
timestamp 1607194113
transform 1 0 21988 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607194113
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__655__B1
timestamp 1607194113
transform 1 0 21804 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__655__A1_N
timestamp 1607194113
transform 1 0 21620 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1607194113
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1607194113
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_209
timestamp 1607194113
transform 1 0 20332 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1607194113
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607194113
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1607194113
transform 1 0 23460 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1607194113
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_245
timestamp 1607194113
transform 1 0 23644 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _671_
timestamp 1607194113
transform 1 0 24196 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _673_
timestamp 1607194113
transform 1 0 24196 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__B1
timestamp 1607194113
transform 1 0 25668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__B2
timestamp 1607194113
transform 1 0 25852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_260
timestamp 1607194113
transform 1 0 25024 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _646_
timestamp 1607194113
transform 1 0 26496 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _657_
timestamp 1607194113
transform 1 0 27600 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607194113
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1607194113
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_272
timestamp 1607194113
transform 1 0 26128 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_284
timestamp 1607194113
transform 1 0 27232 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _620_
timestamp 1607194113
transform 1 0 29440 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _653_
timestamp 1607194113
transform 1 0 28888 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607194113
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__B1
timestamp 1607194113
transform 1 0 27968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__A1
timestamp 1607194113
transform 1 0 29256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__A1_N
timestamp 1607194113
transform 1 0 28704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__657__B
timestamp 1607194113
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_294
timestamp 1607194113
transform 1 0 28152 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_299
timestamp 1607194113
transform 1 0 28612 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1607194113
transform 1 0 31740 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__B1
timestamp 1607194113
transform 1 0 30728 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__B1
timestamp 1607194113
transform 1 0 30360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__B2
timestamp 1607194113
transform 1 0 30544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_322
timestamp 1607194113
transform 1 0 30728 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_324
timestamp 1607194113
transform 1 0 30912 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_332
timestamp 1607194113
transform 1 0 31648 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _854_
timestamp 1607194113
transform 1 0 32200 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607194113
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_334
timestamp 1607194113
transform 1 0 31832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1607194113
transform 1 0 32108 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_336
timestamp 1607194113
transform 1 0 32016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_348
timestamp 1607194113
transform 1 0 33120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _669_
timestamp 1607194113
transform 1 0 34868 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _855_
timestamp 1607194113
transform 1 0 35144 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607194113
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__B1
timestamp 1607194113
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__854__CLK
timestamp 1607194113
transform 1 0 33948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_359
timestamp 1607194113
transform 1 0 34132 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_367
timestamp 1607194113
transform 1 0 34868 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1607194113
transform 1 0 34224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__B1
timestamp 1607194113
transform 1 0 37444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__B2
timestamp 1607194113
transform 1 0 36340 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__855__CLK
timestamp 1607194113
transform 1 0 36892 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_391
timestamp 1607194113
transform 1 0 37076 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_385
timestamp 1607194113
transform 1 0 36524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1607194113
transform 1 0 37260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _679_
timestamp 1607194113
transform 1 0 37628 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _856_
timestamp 1607194113
transform 1 0 38088 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607194113
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__A2_N
timestamp 1607194113
transform 1 0 39100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_398
timestamp 1607194113
transform 1 0 37720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_415
timestamp 1607194113
transform 1 0 39284 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _680_
timestamp 1607194113
transform 1 0 40572 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607194113
transform 1 0 40388 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk_i
timestamp 1607194113
transform 1 0 39836 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__B
timestamp 1607194113
transform 1 0 40388 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__856__CLK
timestamp 1607194113
transform 1 0 39836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_423
timestamp 1607194113
transform 1 0 40020 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_424
timestamp 1607194113
transform 1 0 40112 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_428
timestamp 1607194113
transform 1 0 40480 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_436
timestamp 1607194113
transform 1 0 41216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _652_
timestamp 1607194113
transform 1 0 42136 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _654_
timestamp 1607194113
transform 1 0 41584 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607194113
transform 1 0 43240 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__A1_N
timestamp 1607194113
transform 1 0 41400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_438
timestamp 1607194113
transform 1 0 41400 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_449
timestamp 1607194113
transform 1 0 42412 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_457
timestamp 1607194113
transform 1 0 43148 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_456
timestamp 1607194113
transform 1 0 43056 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1607194113
transform 1 0 44988 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1607194113
transform 1 0 43332 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1607194113
transform 1 0 43976 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_462
timestamp 1607194113
transform 1 0 43608 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_474
timestamp 1607194113
transform 1 0 44712 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_464
timestamp 1607194113
transform 1 0 43792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_469
timestamp 1607194113
transform 1 0 44252 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _859_
timestamp 1607194113
transform 1 0 46920 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607194113
transform 1 0 46000 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__859__CLK
timestamp 1607194113
transform 1 0 46736 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_486
timestamp 1607194113
transform 1 0 45816 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_498
timestamp 1607194113
transform 1 0 46920 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_480
timestamp 1607194113
transform 1 0 45264 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_489
timestamp 1607194113
transform 1 0 46092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_495
timestamp 1607194113
transform 1 0 46644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1607194113
transform 1 0 48944 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _480_
timestamp 1607194113
transform 1 0 47380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607194113
transform 1 0 48852 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_502
timestamp 1607194113
transform 1 0 47288 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_506
timestamp 1607194113
transform 1 0 47656 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_518
timestamp 1607194113
transform 1 0 48760 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1607194113
transform 1 0 48668 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _455_
timestamp 1607194113
transform 1 0 50232 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _477_
timestamp 1607194113
transform 1 0 50232 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__A
timestamp 1607194113
transform 1 0 50876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_523
timestamp 1607194113
transform 1 0 49220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_531
timestamp 1607194113
transform 1 0 49956 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_541
timestamp 1607194113
transform 1 0 50876 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_529
timestamp 1607194113
transform 1 0 49772 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_533
timestamp 1607194113
transform 1 0 50140 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _478_
timestamp 1607194113
transform 1 0 51612 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _866_
timestamp 1607194113
transform 1 0 52072 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607194113
transform 1 0 51612 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__866__CLK
timestamp 1607194113
transform 1 0 51888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_558
timestamp 1607194113
transform 1 0 52440 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_543
timestamp 1607194113
transform 1 0 51060 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_550
timestamp 1607194113
transform 1 0 51704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1607194113
transform 1 0 53176 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607194113
transform -1 0 54832 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607194113
transform -1 0 54832 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607194113
transform 1 0 54464 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1607194113
transform 1 0 53452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_571
timestamp 1607194113
transform 1 0 53636 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_579
timestamp 1607194113
transform 1 0 54372 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_573
timestamp 1607194113
transform 1 0 53820 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:2.g_subtaps:3.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607194113
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607194113
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1607194113
transform 1 0 2484 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp 1607194113
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:2.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 4784 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607194113
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1607194113
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1607194113
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _738_
timestamp 1607194113
transform 1 0 6624 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:2.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5796 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_43
timestamp 1607194113
transform 1 0 5060 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_54
timestamp 1607194113
transform 1 0 6072 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _580_
timestamp 1607194113
transform 1 0 7820 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_64
timestamp 1607194113
transform 1 0 6992 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_72
timestamp 1607194113
transform 1 0 7728 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_77
timestamp 1607194113
transform 1 0 8188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _576_
timestamp 1607194113
transform 1 0 10488 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607194113
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_89
timestamp 1607194113
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_93
timestamp 1607194113
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_101
timestamp 1607194113
transform 1 0 10396 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _732_
timestamp 1607194113
transform 1 0 11776 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__732__B1
timestamp 1607194113
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_106
timestamp 1607194113
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:8.g_subtaps:6.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_delay_line.g_taps:8.g_subtaps:6.inst_tap.g_clkbuf_1.dly_A
timestamp 1607194113
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1607194113
transform 1 0 13248 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_140
timestamp 1607194113
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _599_
timestamp 1607194113
transform 1 0 16008 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607194113
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_147
timestamp 1607194113
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_154
timestamp 1607194113
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_165
timestamp 1607194113
transform 1 0 16284 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1607194113
transform 1 0 17020 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk_i
timestamp 1607194113
transform 1 0 18032 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_176
timestamp 1607194113
transform 1 0 17296 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1607194113
transform 1 0 18308 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _603_
timestamp 1607194113
transform 1 0 19136 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1607194113
transform 1 0 19044 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_199
timestamp 1607194113
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _651_
timestamp 1607194113
transform 1 0 21068 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _672_
timestamp 1607194113
transform 1 0 22080 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607194113
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__A1_N
timestamp 1607194113
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1607194113
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1607194113
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_220
timestamp 1607194113
transform 1 0 21344 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__A2_N
timestamp 1607194113
transform 1 0 23552 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_246
timestamp 1607194113
transform 1 0 23736 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _681_
timestamp 1607194113
transform 1 0 24840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__D
timestamp 1607194113
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_269
timestamp 1607194113
transform 1 0 25852 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607194113
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1607194113
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1607194113
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 28612 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A2
timestamp 1607194113
transform 1 0 29808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1607194113
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_314
timestamp 1607194113
transform 1 0 29992 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_326
timestamp 1607194113
transform 1 0 31096 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _633_
timestamp 1607194113
transform 1 0 32108 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607194113
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__B1
timestamp 1607194113
transform 1 0 31832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_353
timestamp 1607194113
transform 1 0 33580 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1607194113
transform 1 0 34316 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_364
timestamp 1607194113
transform 1 0 34592 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1607194113
transform 1 0 36156 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk_i
timestamp 1607194113
transform 1 0 37352 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk_i
timestamp 1607194113
transform 1 0 35880 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_376
timestamp 1607194113
transform 1 0 35696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_384
timestamp 1607194113
transform 1 0 36432 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_392
timestamp 1607194113
transform 1 0 37168 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _644_
timestamp 1607194113
transform 1 0 37720 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607194113
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__A1_N
timestamp 1607194113
transform 1 0 39192 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_416
timestamp 1607194113
transform 1 0 39376 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _677_
timestamp 1607194113
transform 1 0 40112 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__677__A1_N
timestamp 1607194113
transform 1 0 39928 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607194113
transform 1 0 43240 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__677__A2_N
timestamp 1607194113
transform 1 0 41584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_442
timestamp 1607194113
transform 1 0 41768 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_454
timestamp 1607194113
transform 1 0 42872 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _865_
timestamp 1607194113
transform 1 0 43792 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__865__CLK
timestamp 1607194113
transform 1 0 43608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_459
timestamp 1607194113
transform 1 0 43332 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _458_
timestamp 1607194113
transform 1 0 46368 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_28_483
timestamp 1607194113
transform 1 0 45540 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_491
timestamp 1607194113
transform 1 0 46276 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _453_
timestamp 1607194113
transform 1 0 48944 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607194113
transform 1 0 48852 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_506
timestamp 1607194113
transform 1 0 47656 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_518
timestamp 1607194113
transform 1 0 48760 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1607194113
transform 1 0 50324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_527
timestamp 1607194113
transform 1 0 49588 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_538
timestamp 1607194113
transform 1 0 50600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _457_
timestamp 1607194113
transform 1 0 51336 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_555
timestamp 1607194113
transform 1 0 52164 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1607194113
transform 1 0 52900 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607194113
transform -1 0 54832 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607194113
transform 1 0 54464 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_566
timestamp 1607194113
transform 1 0 53176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_578
timestamp 1607194113
transform 1 0 54280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _771_
timestamp 1607194113
transform 1 0 1564 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607194113
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1607194113
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a22oi_4  _759_
timestamp 1607194113
transform 1 0 4048 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__771__CLK
timestamp 1607194113
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_26
timestamp 1607194113
transform 1 0 3496 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _742_
timestamp 1607194113
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607194113
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_49
timestamp 1607194113
transform 1 0 5612 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _772_
timestamp 1607194113
transform 1 0 8372 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_29_66
timestamp 1607194113
transform 1 0 7176 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_78
timestamp 1607194113
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__772__CLK
timestamp 1607194113
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_100
timestamp 1607194113
transform 1 0 10304 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _600_
timestamp 1607194113
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _734_
timestamp 1607194113
transform 1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607194113
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__734__B1
timestamp 1607194113
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_109
timestamp 1607194113
transform 1 0 11132 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_117
timestamp 1607194113
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_139
timestamp 1607194113
transform 1 0 13892 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_145
timestamp 1607194113
transform 1 0 14444 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _781_
timestamp 1607194113
transform 1 0 14720 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__781__CLK
timestamp 1607194113
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _780_
timestamp 1607194113
transform 1 0 18032 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607194113
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_167
timestamp 1607194113
transform 1 0 16468 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1607194113
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__780__CLK
timestamp 1607194113
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_205
timestamp 1607194113
transform 1 0 19964 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _811_
timestamp 1607194113
transform 1 0 21068 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__811__CLK
timestamp 1607194113
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp 1607194113
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607194113
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_236
timestamp 1607194113
transform 1 0 22816 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1607194113
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _660_
timestamp 1607194113
transform 1 0 24748 0 1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 26772 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1607194113
transform 1 0 26588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_271
timestamp 1607194113
transform 1 0 26036 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _682_
timestamp 1607194113
transform 1 0 29256 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607194113
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_299
timestamp 1607194113
transform 1 0 28612 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _624_
timestamp 1607194113
transform 1 0 31004 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_315
timestamp 1607194113
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_323
timestamp 1607194113
transform 1 0 30820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _629_
timestamp 1607194113
transform 1 0 33212 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A1_N
timestamp 1607194113
transform 1 0 32476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__B2
timestamp 1607194113
transform 1 0 32660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A2_N
timestamp 1607194113
transform 1 0 32844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_347
timestamp 1607194113
transform 1 0 33028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _628_
timestamp 1607194113
transform 1 0 34960 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607194113
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_358
timestamp 1607194113
transform 1 0 34040 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_367
timestamp 1607194113
transform 1 0 34868 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__B1
timestamp 1607194113
transform 1 0 36432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__B2
timestamp 1607194113
transform 1 0 36616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_388
timestamp 1607194113
transform 1 0 36800 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _645_
timestamp 1607194113
transform 1 0 38824 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_400
timestamp 1607194113
transform 1 0 37904 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_408
timestamp 1607194113
transform 1 0 38640 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _670_
timestamp 1607194113
transform 1 0 40756 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607194113
transform 1 0 40388 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__B
timestamp 1607194113
transform 1 0 39652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_421
timestamp 1607194113
transform 1 0 39836 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_428
timestamp 1607194113
transform 1 0 40480 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_434
timestamp 1607194113
transform 1 0 41032 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _631_
timestamp 1607194113
transform 1 0 41768 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__A1_N
timestamp 1607194113
transform 1 0 43240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _637_
timestamp 1607194113
transform 1 0 43976 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_460
timestamp 1607194113
transform 1 0 43424 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_475
timestamp 1607194113
transform 1 0 44804 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _675_
timestamp 1607194113
transform 1 0 46092 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607194113
transform 1 0 46000 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__A1_N
timestamp 1607194113
transform 1 0 45816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_483
timestamp 1607194113
transform 1 0 45540 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _442_
timestamp 1607194113
transform 1 0 48300 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__B
timestamp 1607194113
transform 1 0 48116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_505
timestamp 1607194113
transform 1 0 47564 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _456_
timestamp 1607194113
transform 1 0 49864 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__A
timestamp 1607194113
transform 1 0 49680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_522
timestamp 1607194113
transform 1 0 49128 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_537
timestamp 1607194113
transform 1 0 50508 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _448_
timestamp 1607194113
transform 1 0 52348 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607194113
transform 1 0 51612 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_550
timestamp 1607194113
transform 1 0 51704 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_556
timestamp 1607194113
transform 1 0 52256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607194113
transform -1 0 54832 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_566
timestamp 1607194113
transform 1 0 53176 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_578
timestamp 1607194113
transform 1 0 54280 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:1.g_subtaps:2.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607194113
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607194113
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1607194113
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_19
timestamp 1607194113
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _604_
timestamp 1607194113
transform 1 0 4232 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607194113
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1607194113
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1607194113
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_37
timestamp 1607194113
transform 1 0 4508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _748_
timestamp 1607194113
transform 1 0 6164 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__748__B1
timestamp 1607194113
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_49
timestamp 1607194113
transform 1 0 5612 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_71
timestamp 1607194113
transform 1 0 7636 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_83
timestamp 1607194113
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _601_
timestamp 1607194113
transform 1 0 9660 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607194113
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1607194113
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_107
timestamp 1607194113
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_119
timestamp 1607194113
transform 1 0 12052 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1607194113
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _733_
timestamp 1607194113
transform 1 0 12696 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_142
timestamp 1607194113
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _728_
timestamp 1607194113
transform 1 0 15824 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607194113
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__728__A
timestamp 1607194113
transform 1 0 15640 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1607194113
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1607194113
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_164
timestamp 1607194113
transform 1 0 16192 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _724_
timestamp 1607194113
transform 1 0 17020 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__724__A
timestamp 1607194113
transform 1 0 17388 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_172
timestamp 1607194113
transform 1 0 16928 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_179
timestamp 1607194113
transform 1 0 17572 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_191
timestamp 1607194113
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_203
timestamp 1607194113
transform 1 0 19780 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _683_
timestamp 1607194113
transform 1 0 21712 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607194113
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1607194113
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1607194113
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_223
timestamp 1607194113
transform 1 0 21620 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1607194113
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _790_
timestamp 1607194113
transform 1 0 23920 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__790__CLK
timestamp 1607194113
transform 1 0 23736 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_239
timestamp 1607194113
transform 1 0 23092 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_245
timestamp 1607194113
transform 1 0 23644 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_267
timestamp 1607194113
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _659_
timestamp 1607194113
transform 1 0 26496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607194113
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_279
timestamp 1607194113
transform 1 0 26772 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1607194113
transform 1 0 27876 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _658_
timestamp 1607194113
transform 1 0 28336 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__A
timestamp 1607194113
transform 1 0 29164 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__A
timestamp 1607194113
transform 1 0 29716 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_295
timestamp 1607194113
transform 1 0 28244 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_307
timestamp 1607194113
transform 1 0 29348 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1607194113
transform 1 0 29900 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_316
timestamp 1607194113
transform 1 0 30176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_328
timestamp 1607194113
transform 1 0 31280 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _623_
timestamp 1607194113
transform 1 0 32108 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607194113
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__B1
timestamp 1607194113
transform 1 0 33580 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__A1_N
timestamp 1607194113
transform 1 0 31832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__B2
timestamp 1607194113
transform 1 0 33764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_357
timestamp 1607194113
transform 1 0 33948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_369
timestamp 1607194113
transform 1 0 35052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk_i
timestamp 1607194113
transform 1 0 36340 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_i_A
timestamp 1607194113
transform 1 0 36156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_386
timestamp 1607194113
transform 1 0 36616 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_394
timestamp 1607194113
transform 1 0 37352 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _643_
timestamp 1607194113
transform 1 0 38548 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607194113
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__B1
timestamp 1607194113
transform 1 0 38364 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__B2
timestamp 1607194113
transform 1 0 38180 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_398
timestamp 1607194113
transform 1 0 37720 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_402
timestamp 1607194113
transform 1 0 38088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_423
timestamp 1607194113
transform 1 0 40020 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_435
timestamp 1607194113
transform 1 0 41124 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _634_
timestamp 1607194113
transform 1 0 41860 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607194113
transform 1 0 43240 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__A
timestamp 1607194113
transform 1 0 41676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_446
timestamp 1607194113
transform 1 0 42136 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _635_
timestamp 1607194113
transform 1 0 43884 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_459
timestamp 1607194113
transform 1 0 43332 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_481
timestamp 1607194113
transform 1 0 45356 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_493
timestamp 1607194113
transform 1 0 46460 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1607194113
transform 1 0 47840 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607194113
transform 1 0 48852 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1607194113
transform 1 0 48116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_505
timestamp 1607194113
transform 1 0 47564 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_513
timestamp 1607194113
transform 1 0 48300 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_520
timestamp 1607194113
transform 1 0 48944 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _443_
timestamp 1607194113
transform 1 0 49036 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _636_
timestamp 1607194113
transform 1 0 50692 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__B1
timestamp 1607194113
transform 1 0 50508 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_528
timestamp 1607194113
transform 1 0 49680 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_536
timestamp 1607194113
transform 1 0 50416 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_555
timestamp 1607194113
transform 1 0 52164 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _445_
timestamp 1607194113
transform 1 0 52900 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607194113
transform -1 0 54832 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607194113
transform 1 0 54464 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_570
timestamp 1607194113
transform 1 0 53544 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_578
timestamp 1607194113
transform 1 0 54280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607194113
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607194113
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_15
timestamp 1607194113
transform 1 0 2484 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _760_
timestamp 1607194113
transform 1 0 4048 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:1.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 3036 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_24
timestamp 1607194113
transform 1 0 3312 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_35
timestamp 1607194113
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _746_
timestamp 1607194113
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  inst_delay_line.g_taps:0.g_subtaps:1.inst_tap.g_clkbuf_1.dly
timestamp 1607194113
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607194113
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_47
timestamp 1607194113
transform 1 0 5428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1607194113
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _747_
timestamp 1607194113
transform 1 0 8004 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_66
timestamp 1607194113
transform 1 0 7176 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_74
timestamp 1607194113
transform 1 0 7912 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _605_
timestamp 1607194113
transform 1 0 10212 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_31_91
timestamp 1607194113
transform 1 0 9476 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607194113
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1607194113
transform 1 0 11500 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1607194113
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1607194113
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1607194113
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _688_
timestamp 1607194113
transform 1 0 16284 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _731_
timestamp 1607194113
transform 1 0 15180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_147
timestamp 1607194113
transform 1 0 14628 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_157
timestamp 1607194113
transform 1 0 15548 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _721_
timestamp 1607194113
transform 1 0 18308 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607194113
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk_i
timestamp 1607194113
transform 1 0 17388 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__721__A
timestamp 1607194113
transform 1 0 18124 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_i_A
timestamp 1607194113
transform 1 0 17664 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1607194113
transform 1 0 16652 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1607194113
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1607194113
transform 1 0 18032 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _787_
timestamp 1607194113
transform 1 0 19412 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__787__CLK
timestamp 1607194113
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_191
timestamp 1607194113
transform 1 0 18676 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_218
timestamp 1607194113
transform 1 0 21160 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _720_
timestamp 1607194113
transform 1 0 23644 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607194113
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_230
timestamp 1607194113
transform 1 0 22264 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_242
timestamp 1607194113
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1607194113
transform 1 0 25116 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _719_
timestamp 1607194113
transform 1 0 26404 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_273
timestamp 1607194113
transform 1 0 26220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_291
timestamp 1607194113
transform 1 0 27876 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607194113
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_303
timestamp 1607194113
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_306
timestamp 1607194113
transform 1 0 29256 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _665_
timestamp 1607194113
transform 1 0 30176 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_31_314
timestamp 1607194113
transform 1 0 29992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_330
timestamp 1607194113
transform 1 0 31464 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1607194113
transform 1 0 32292 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_338
timestamp 1607194113
transform 1 0 32200 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_342
timestamp 1607194113
transform 1 0 32568 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_354
timestamp 1607194113
transform 1 0 33672 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607194113
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1607194113
transform 1 0 34868 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _625_
timestamp 1607194113
transform 1 0 36064 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_379
timestamp 1607194113
transform 1 0 35972 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _563_
timestamp 1607194113
transform 1 0 38272 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _678_
timestamp 1607194113
transform 1 0 39284 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__B2
timestamp 1607194113
transform 1 0 37536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__B1
timestamp 1607194113
transform 1 0 37720 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_400
timestamp 1607194113
transform 1 0 37904 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_407
timestamp 1607194113
transform 1 0 38548 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607194113
transform 1 0 40388 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__A
timestamp 1607194113
transform 1 0 39560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_420
timestamp 1607194113
transform 1 0 39744 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_426
timestamp 1607194113
transform 1 0 40296 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_428
timestamp 1607194113
transform 1 0 40480 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _696_
timestamp 1607194113
transform 1 0 41676 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__696__A1_N
timestamp 1607194113
transform 1 0 43148 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_440
timestamp 1607194113
transform 1 0 41584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _674_
timestamp 1607194113
transform 1 0 44988 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_459
timestamp 1607194113
transform 1 0 43332 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_471
timestamp 1607194113
transform 1 0 44436 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _627_
timestamp 1607194113
transform 1 0 46092 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607194113
transform 1 0 46000 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__A
timestamp 1607194113
transform 1 0 46368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_480
timestamp 1607194113
transform 1 0 45264 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_494
timestamp 1607194113
transform 1 0 46552 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _451_
timestamp 1607194113
transform 1 0 47932 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_31_506
timestamp 1607194113
transform 1 0 47656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1607194113
transform 1 0 49956 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_523
timestamp 1607194113
transform 1 0 49220 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_534
timestamp 1607194113
transform 1 0 50232 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _447_
timestamp 1607194113
transform 1 0 51888 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607194113
transform 1 0 51612 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_546
timestamp 1607194113
transform 1 0 51336 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_550
timestamp 1607194113
transform 1 0 51704 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_559
timestamp 1607194113
transform 1 0 52532 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1607194113
transform 1 0 53268 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607194113
transform -1 0 54832 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_570
timestamp 1607194113
transform 1 0 53544 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_578
timestamp 1607194113
transform 1 0 54280 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _770_
timestamp 1607194113
transform 1 0 1472 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607194113
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1607194113
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1607194113
transform 1 0 4508 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607194113
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__770__CLK
timestamp 1607194113
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_25
timestamp 1607194113
transform 1 0 3404 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1607194113
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1607194113
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_40
timestamp 1607194113
transform 1 0 4784 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _749_
timestamp 1607194113
transform 1 0 6072 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_52
timestamp 1607194113
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _762_
timestamp 1607194113
transform 1 0 8280 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_70
timestamp 1607194113
transform 1 0 7544 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_81
timestamp 1607194113
transform 1 0 8556 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _609_
timestamp 1607194113
transform 1 0 9660 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607194113
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1607194113
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _735_
timestamp 1607194113
transform 1 0 11960 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__A1
timestamp 1607194113
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1607194113
transform 1 0 11132 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_117
timestamp 1607194113
transform 1 0 11868 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _607_
timestamp 1607194113
transform 1 0 14168 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__735__A1_N
timestamp 1607194113
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__735__B2
timestamp 1607194113
transform 1 0 13616 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__735__A2_N
timestamp 1607194113
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_140
timestamp 1607194113
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_145
timestamp 1607194113
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _697_
timestamp 1607194113
transform 1 0 15548 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607194113
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_154
timestamp 1607194113
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_161
timestamp 1607194113
transform 1 0 15916 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _687_
timestamp 1607194113
transform 1 0 16652 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _725_
timestamp 1607194113
transform 1 0 17848 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_32_173
timestamp 1607194113
transform 1 0 17020 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_181
timestamp 1607194113
transform 1 0 17756 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__725__A1_N
timestamp 1607194113
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_200
timestamp 1607194113
transform 1 0 19504 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _788_
timestamp 1607194113
transform 1 0 20884 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607194113
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__788__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _717_
timestamp 1607194113
transform 1 0 23460 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__717__A
timestamp 1607194113
transform 1 0 23276 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_234
timestamp 1607194113
transform 1 0 22632 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1607194113
transform 1 0 23184 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_247
timestamp 1607194113
transform 1 0 23828 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _663_
timestamp 1607194113
transform 1 0 25024 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__663__B
timestamp 1607194113
transform 1 0 25668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_259
timestamp 1607194113
transform 1 0 24932 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_269
timestamp 1607194113
transform 1 0 25852 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _662_
timestamp 1607194113
transform 1 0 26496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _791_
timestamp 1607194113
transform 1 0 27784 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607194113
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__A
timestamp 1607194113
transform 1 0 26772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_281
timestamp 1607194113
transform 1 0 26956 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_289
timestamp 1607194113
transform 1 0 27692 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__791__CLK
timestamp 1607194113
transform 1 0 29532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_311
timestamp 1607194113
transform 1 0 29716 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1607194113
transform 1 0 30912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_323
timestamp 1607194113
transform 1 0 30820 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_327
timestamp 1607194113
transform 1 0 31188 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _796_
timestamp 1607194113
transform 1 0 32936 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607194113
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_335
timestamp 1607194113
transform 1 0 31924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_337
timestamp 1607194113
transform 1 0 32108 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_345
timestamp 1607194113
transform 1 0 32844 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__796__CLK
timestamp 1607194113
transform 1 0 34684 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_367
timestamp 1607194113
transform 1 0 34868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_379
timestamp 1607194113
transform 1 0 35972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_391
timestamp 1607194113
transform 1 0 37076 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _638_
timestamp 1607194113
transform 1 0 39008 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607194113
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk_i
timestamp 1607194113
transform 1 0 38456 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_398
timestamp 1607194113
transform 1 0 37720 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_409
timestamp 1607194113
transform 1 0 38732 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _693_
timestamp 1607194113
transform 1 0 41216 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A
timestamp 1607194113
transform 1 0 41032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__B1
timestamp 1607194113
transform 1 0 40480 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_430
timestamp 1607194113
transform 1 0 40664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607194113
transform 1 0 43240 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_440
timestamp 1607194113
transform 1 0 41584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_452
timestamp 1607194113
transform 1 0 42688 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_459
timestamp 1607194113
transform 1 0 43332 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_471
timestamp 1607194113
transform 1 0 44436 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _806_
timestamp 1607194113
transform 1 0 46000 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__806__CLK
timestamp 1607194113
transform 1 0 45816 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_483
timestamp 1607194113
transform 1 0 45540 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _867_
timestamp 1607194113
transform 1 0 48944 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607194113
transform 1 0 48852 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__867__CLK
timestamp 1607194113
transform 1 0 48668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_507
timestamp 1607194113
transform 1 0 47748 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_515
timestamp 1607194113
transform 1 0 48484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_539
timestamp 1607194113
transform 1 0 50692 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _868_
timestamp 1607194113
transform 1 0 51980 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__868__CLK
timestamp 1607194113
transform 1 0 51796 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607194113
transform -1 0 54832 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607194113
transform 1 0 54464 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_572
timestamp 1607194113
transform 1 0 53728 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607194113
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607194113
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607194113
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1607194113
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607194113
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607194113
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _751_
timestamp 1607194113
transform 1 0 4416 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _761_
timestamp 1607194113
transform 1 0 3496 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607194113
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_23
timestamp 1607194113
transform 1 0 3220 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1607194113
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1607194113
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _750_
timestamp 1607194113
transform 1 0 5704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607194113
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_42
timestamp 1607194113
transform 1 0 4968 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_53
timestamp 1607194113
transform 1 0 5980 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_62
timestamp 1607194113
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_52
timestamp 1607194113
transform 1 0 5888 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _612_
timestamp 1607194113
transform 1 0 7176 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_4  _763_
timestamp 1607194113
transform 1 0 7268 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__A
timestamp 1607194113
transform 1 0 8004 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_66
timestamp 1607194113
transform 1 0 7176 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_83
timestamp 1607194113
transform 1 0 8740 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_64
timestamp 1607194113
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_77
timestamp 1607194113
transform 1 0 8188 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _615_
timestamp 1607194113
transform 1 0 9660 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _736_
timestamp 1607194113
transform 1 0 10120 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607194113
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_95
timestamp 1607194113
transform 1 0 9844 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_89
timestamp 1607194113
transform 1 0 9292 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_100
timestamp 1607194113
transform 1 0 10304 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_112
timestamp 1607194113
transform 1 0 11408 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__736__A1_N
timestamp 1607194113
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _564_
timestamp 1607194113
transform 1 0 11040 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_120
timestamp 1607194113
transform 1 0 12144 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1607194113
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1607194113
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__736__A2_N
timestamp 1607194113
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__736__B2
timestamp 1607194113
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607194113
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _778_
timestamp 1607194113
transform 1 0 12328 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _779_
timestamp 1607194113
transform 1 0 13248 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__778__CLK
timestamp 1607194113
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_131
timestamp 1607194113
transform 1 0 13156 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_143
timestamp 1607194113
transform 1 0 14260 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _565_
timestamp 1607194113
transform 1 0 15824 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _572_
timestamp 1607194113
transform 1 0 15732 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607194113
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk_i
timestamp 1607194113
transform 1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1607194113
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__779__CLK
timestamp 1607194113
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_153
timestamp 1607194113
transform 1 0 15180 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1607194113
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_154
timestamp 1607194113
transform 1 0 15272 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_169
timestamp 1607194113
transform 1 0 16652 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_168
timestamp 1607194113
transform 1 0 16560 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1607194113
transform 1 0 16468 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__686__A
timestamp 1607194113
transform 1 0 17020 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk_i
timestamp 1607194113
transform 1 0 17112 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1607194113
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__686__B
timestamp 1607194113
transform 1 0 17848 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _686_
timestamp 1607194113
transform 1 0 17204 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_34_184
timestamp 1607194113
transform 1 0 18032 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607194113
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _692_
timestamp 1607194113
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _722_
timestamp 1607194113
transform 1 0 18584 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _723_
timestamp 1607194113
transform 1 0 19136 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__722__A1_N
timestamp 1607194113
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_188
timestamp 1607194113
transform 1 0 18400 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_208
timestamp 1607194113
transform 1 0 20240 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _619_
timestamp 1607194113
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _642_
timestamp 1607194113
transform 1 0 21712 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607194113
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__723__A1_N
timestamp 1607194113
transform 1 0 20608 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1607194113
transform 1 0 20792 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1607194113
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_227
timestamp 1607194113
transform 1 0 21988 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_218
timestamp 1607194113
transform 1 0 21160 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _666_
timestamp 1607194113
transform 1 0 24104 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _876_
timestamp 1607194113
transform 1 0 22448 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607194113
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__876__CLK
timestamp 1607194113
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_239
timestamp 1607194113
transform 1 0 23092 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1607194113
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_245
timestamp 1607194113
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_249
timestamp 1607194113
transform 1 0 24012 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _611_
timestamp 1607194113
transform 1 0 24932 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _718_
timestamp 1607194113
transform 1 0 25668 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__A
timestamp 1607194113
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A
timestamp 1607194113
transform 1 0 24748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_261
timestamp 1607194113
transform 1 0 25116 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_251
timestamp 1607194113
transform 1 0 24196 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_262
timestamp 1607194113
transform 1 0 25208 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _792_
timestamp 1607194113
transform 1 0 27048 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607194113
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_283
timestamp 1607194113
transform 1 0 27140 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1607194113
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_276
timestamp 1607194113
transform 1 0 26496 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _713_
timestamp 1607194113
transform 1 0 29808 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607194113
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__710__A
timestamp 1607194113
transform 1 0 29808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__792__CLK
timestamp 1607194113
transform 1 0 28796 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_295
timestamp 1607194113
transform 1 0 28244 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_303
timestamp 1607194113
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_306
timestamp 1607194113
transform 1 0 29256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_303
timestamp 1607194113
transform 1 0 28980 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_311
timestamp 1607194113
transform 1 0 29716 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _710_
timestamp 1607194113
transform 1 0 29992 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _712_
timestamp 1607194113
transform 1 0 31464 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_33_318
timestamp 1607194113
transform 1 0 30360 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_328
timestamp 1607194113
transform 1 0 31280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _711_
timestamp 1607194113
transform 1 0 33212 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607194113
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_346
timestamp 1607194113
transform 1 0 32936 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_337
timestamp 1607194113
transform 1 0 32108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _797_
timestamp 1607194113
transform 1 0 35604 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607194113
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__711__A1_N
timestamp 1607194113
transform 1 0 34684 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_358
timestamp 1607194113
transform 1 0 34040 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_367
timestamp 1607194113
transform 1 0 34868 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_367
timestamp 1607194113
transform 1 0 34868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _706_
timestamp 1607194113
transform 1 0 36248 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk_i
timestamp 1607194113
transform 1 0 35972 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__706__A
timestamp 1607194113
transform 1 0 36616 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__797__CLK
timestamp 1607194113
transform 1 0 37352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_388
timestamp 1607194113
transform 1 0 36800 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _707_
timestamp 1607194113
transform 1 0 38088 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _799_
timestamp 1607194113
transform 1 0 38640 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607194113
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_396
timestamp 1607194113
transform 1 0 37536 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_396
timestamp 1607194113
transform 1 0 37536 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_398
timestamp 1607194113
transform 1 0 37720 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_406
timestamp 1607194113
transform 1 0 38456 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607194113
transform 1 0 40388 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk_i
timestamp 1607194113
transform 1 0 41216 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__799__CLK
timestamp 1607194113
transform 1 0 40388 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_418
timestamp 1607194113
transform 1 0 39560 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_426
timestamp 1607194113
transform 1 0 40296 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_428
timestamp 1607194113
transform 1 0 40480 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_429
timestamp 1607194113
transform 1 0 40572 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_437
timestamp 1607194113
transform 1 0 41308 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _698_
timestamp 1607194113
transform 1 0 41676 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _805_
timestamp 1607194113
transform 1 0 42228 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607194113
transform 1 0 43240 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__698__A
timestamp 1607194113
transform 1 0 41492 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__805__CLK
timestamp 1607194113
transform 1 0 42044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_439
timestamp 1607194113
transform 1 0 41492 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1607194113
transform 1 0 42044 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_457
timestamp 1607194113
transform 1 0 43148 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _689_
timestamp 1607194113
transform 1 0 44620 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__689__A
timestamp 1607194113
transform 1 0 44436 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_466
timestamp 1607194113
transform 1 0 43976 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_478
timestamp 1607194113
transform 1 0 45080 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_459
timestamp 1607194113
transform 1 0 43332 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_477
timestamp 1607194113
transform 1 0 44988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _694_
timestamp 1607194113
transform 1 0 45724 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _695_
timestamp 1607194113
transform 1 0 46092 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607194113
transform 1 0 46000 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_486
timestamp 1607194113
transform 1 0 45816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1607194113
transform 1 0 48392 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607194113
transform 1 0 48852 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__694__A1_N
timestamp 1607194113
transform 1 0 47196 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1607194113
transform 1 0 47564 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_513
timestamp 1607194113
transform 1 0 48300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1607194113
transform 1 0 48668 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_503
timestamp 1607194113
transform 1 0 47380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_515
timestamp 1607194113
transform 1 0 48484 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_520
timestamp 1607194113
transform 1 0 48944 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1607194113
transform 1 0 50600 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1607194113
transform 1 0 49588 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _691_
timestamp 1607194113
transform 1 0 49496 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__A
timestamp 1607194113
transform 1 0 49864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1607194113
transform 1 0 49404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_532
timestamp 1607194113
transform 1 0 50048 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_541
timestamp 1607194113
transform 1 0 50876 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _641_
timestamp 1607194113
transform 1 0 51704 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _808_
timestamp 1607194113
transform 1 0 51980 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607194113
transform 1 0 51612 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__808__CLK
timestamp 1607194113
transform 1 0 51796 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_542
timestamp 1607194113
transform 1 0 50968 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_550
timestamp 1607194113
transform 1 0 51704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607194113
transform -1 0 54832 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607194113
transform -1 0 54832 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607194113
transform 1 0 54464 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_566
timestamp 1607194113
transform 1 0 53176 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_578
timestamp 1607194113
transform 1 0 54280 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_572
timestamp 1607194113
transform 1 0 53728 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _769_
timestamp 1607194113
transform 1 0 2116 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607194113
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1607194113
transform 1 0 1380 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__769__CLK
timestamp 1607194113
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1607194113
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1607194113
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607194113
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_44
timestamp 1607194113
transform 1 0 5152 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_53
timestamp 1607194113
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1607194113
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _381_
timestamp 1607194113
transform 1 0 6992 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_35_73
timestamp 1607194113
transform 1 0 7820 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _737_
timestamp 1607194113
transform 1 0 9384 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__737__B
timestamp 1607194113
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp 1607194113
transform 1 0 8924 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_89
timestamp 1607194113
transform 1 0 9292 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_99
timestamp 1607194113
transform 1 0 10212 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1607194113
transform 1 0 11040 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _616_
timestamp 1607194113
transform 1 0 12420 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607194113
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_107
timestamp 1607194113
transform 1 0 10948 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_111
timestamp 1607194113
transform 1 0 11316 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_119
timestamp 1607194113
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _668_
timestamp 1607194113
transform 1 0 13800 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__B
timestamp 1607194113
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_132
timestamp 1607194113
transform 1 0 13248 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_141
timestamp 1607194113
transform 1 0 14076 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _568_
timestamp 1607194113
transform 1 0 14996 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__B1
timestamp 1607194113
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_164
timestamp 1607194113
transform 1 0 16192 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607194113
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk_i
timestamp 1607194113
transform 1 0 17664 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1607194113
transform 1 0 17296 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1607194113
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _789_
timestamp 1607194113
transform 1 0 19412 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__789__CLK
timestamp 1607194113
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_196
timestamp 1607194113
transform 1 0 19136 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1607194113
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _661_
timestamp 1607194113
transform 1 0 22540 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _765_
timestamp 1607194113
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607194113
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__661__A
timestamp 1607194113
transform 1 0 22356 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__765__B
timestamp 1607194113
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_230
timestamp 1607194113
transform 1 0 22264 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_236
timestamp 1607194113
transform 1 0 22816 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _685_
timestamp 1607194113
transform 1 0 25208 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_254
timestamp 1607194113
transform 1 0 24472 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_266
timestamp 1607194113
transform 1 0 25576 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _716_
timestamp 1607194113
transform 1 0 26588 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_35_274
timestamp 1607194113
transform 1 0 26312 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _571_
timestamp 1607194113
transform 1 0 29716 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607194113
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1607194113
transform 1 0 28060 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_306
timestamp 1607194113
transform 1 0 29256 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_310
timestamp 1607194113
transform 1 0 29624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _795_
timestamp 1607194113
transform 1 0 31004 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_35_314
timestamp 1607194113
transform 1 0 29992 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_322
timestamp 1607194113
transform 1 0 30728 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__795__CLK
timestamp 1607194113
transform 1 0 32752 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_346
timestamp 1607194113
transform 1 0 32936 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_354
timestamp 1607194113
transform 1 0 33672 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _708_
timestamp 1607194113
transform 1 0 33764 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _798_
timestamp 1607194113
transform 1 0 35328 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607194113
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_358
timestamp 1607194113
transform 1 0 34040 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_367
timestamp 1607194113
transform 1 0 34868 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_371
timestamp 1607194113
transform 1 0 35236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__798__CLK
timestamp 1607194113
transform 1 0 37076 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1607194113
transform 1 0 37260 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _704_
timestamp 1607194113
transform 1 0 38180 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_35_401
timestamp 1607194113
transform 1 0 37996 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _702_
timestamp 1607194113
transform 1 0 40848 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607194113
transform 1 0 40388 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__702__A
timestamp 1607194113
transform 1 0 40664 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_419
timestamp 1607194113
transform 1 0 39652 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_428
timestamp 1607194113
transform 1 0 40480 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_436
timestamp 1607194113
transform 1 0 41216 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _804_
timestamp 1607194113
transform 1 0 43240 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__804__CLK
timestamp 1607194113
transform 1 0 43056 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_448
timestamp 1607194113
transform 1 0 42320 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_477
timestamp 1607194113
transform 1 0 44988 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _807_
timestamp 1607194113
transform 1 0 46736 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607194113
transform 1 0 46000 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__807__CLK
timestamp 1607194113
transform 1 0 46552 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_485
timestamp 1607194113
transform 1 0 45724 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_489
timestamp 1607194113
transform 1 0 46092 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_493
timestamp 1607194113
transform 1 0 46460 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_515
timestamp 1607194113
transform 1 0 48484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_527
timestamp 1607194113
transform 1 0 49588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_539
timestamp 1607194113
transform 1 0 50692 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _809_
timestamp 1607194113
transform 1 0 51704 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607194113
transform 1 0 51612 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__809__CLK
timestamp 1607194113
transform 1 0 51428 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607194113
transform -1 0 54832 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_569
timestamp 1607194113
transform 1 0 53452 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _610_
timestamp 1607194113
transform 1 0 1932 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607194113
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__A
timestamp 1607194113
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1607194113
transform 1 0 1380 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1607194113
transform 1 0 2944 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _602_
timestamp 1607194113
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607194113
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__A
timestamp 1607194113
transform 1 0 4876 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_28
timestamp 1607194113
transform 1 0 3680 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1607194113
transform 1 0 5888 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_43
timestamp 1607194113
transform 1 0 5060 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_51
timestamp 1607194113
transform 1 0 5796 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_55
timestamp 1607194113
transform 1 0 6164 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _579_
timestamp 1607194113
transform 1 0 6900 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1607194113
transform 1 0 8556 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_72
timestamp 1607194113
transform 1 0 7728 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_80
timestamp 1607194113
transform 1 0 8464 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_4  _617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 9844 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607194113
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_84
timestamp 1607194113
transform 1 0 8832 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1607194113
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _574_
timestamp 1607194113
transform 1 0 12512 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__B1
timestamp 1607194113
transform 1 0 11408 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_114
timestamp 1607194113
transform 1 0 11592 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_122
timestamp 1607194113
transform 1 0 12328 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1607194113
transform 1 0 13616 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_128
timestamp 1607194113
transform 1 0 12880 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_139
timestamp 1607194113
transform 1 0 13892 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607194113
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1607194113
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1607194113
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_166
timestamp 1607194113
transform 1 0 16376 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _824_
timestamp 1607194113
transform 1 0 17112 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__824__CLK
timestamp 1607194113
transform 1 0 18860 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_195
timestamp 1607194113
transform 1 0 19044 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_207
timestamp 1607194113
transform 1 0 20148 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _394_
timestamp 1607194113
transform 1 0 20884 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607194113
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1607194113
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__B
timestamp 1607194113
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1607194113
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_228
timestamp 1607194113
transform 1 0 22080 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _764_
timestamp 1607194113
transform 1 0 23552 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _766_
timestamp 1607194113
transform 1 0 22540 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__764__A1
timestamp 1607194113
transform 1 0 23368 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__764__A2
timestamp 1607194113
transform 1 0 23184 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_232
timestamp 1607194113
transform 1 0 22448 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1607194113
transform 1 0 22816 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__764__B1
timestamp 1607194113
transform 1 0 24748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_259
timestamp 1607194113
transform 1 0 24932 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _714_
timestamp 1607194113
transform 1 0 26956 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607194113
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__714__A
timestamp 1607194113
transform 1 0 26772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1607194113
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_276
timestamp 1607194113
transform 1 0 26496 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_285
timestamp 1607194113
transform 1 0 27324 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _794_
timestamp 1607194113
transform 1 0 28336 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_36_293
timestamp 1607194113
transform 1 0 28060 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__794__CLK
timestamp 1607194113
transform 1 0 30084 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_317
timestamp 1607194113
transform 1 0 30268 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_329
timestamp 1607194113
transform 1 0 31372 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607194113
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_335
timestamp 1607194113
transform 1 0 31924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_337
timestamp 1607194113
transform 1 0 32108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_349
timestamp 1607194113
transform 1 0 33212 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _709_
timestamp 1607194113
transform 1 0 33948 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_36_373
timestamp 1607194113
transform 1 0 35420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_385
timestamp 1607194113
transform 1 0 36524 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607194113
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__801__CLK
timestamp 1607194113
transform 1 0 39376 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_398
timestamp 1607194113
transform 1 0 37720 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_410
timestamp 1607194113
transform 1 0 38824 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _801_
timestamp 1607194113
transform 1 0 39560 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_36_437
timestamp 1607194113
transform 1 0 41308 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _701_
timestamp 1607194113
transform 1 0 42228 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607194113
transform 1 0 43240 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__701__A
timestamp 1607194113
transform 1 0 42504 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_445
timestamp 1607194113
transform 1 0 42044 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_452
timestamp 1607194113
transform 1 0 42688 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _700_
timestamp 1607194113
transform 1 0 43332 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__700__A1_N
timestamp 1607194113
transform 1 0 44804 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_477
timestamp 1607194113
transform 1 0 44988 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _767_
timestamp 1607194113
transform 1 0 46276 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__767__D
timestamp 1607194113
transform 1 0 46092 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__767__CLK
timestamp 1607194113
transform 1 0 45908 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_485
timestamp 1607194113
transform 1 0 45724 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607194113
transform 1 0 48852 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_510
timestamp 1607194113
transform 1 0 48024 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_518
timestamp 1607194113
transform 1 0 48760 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_520
timestamp 1607194113
transform 1 0 48944 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _690_
timestamp 1607194113
transform 1 0 49864 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_36_528
timestamp 1607194113
transform 1 0 49680 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _546_
timestamp 1607194113
transform 1 0 52072 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1607194113
transform 1 0 51888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__B
timestamp 1607194113
transform 1 0 51704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_546
timestamp 1607194113
transform 1 0 51336 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607194113
transform -1 0 54832 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607194113
transform 1 0 54464 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__C
timestamp 1607194113
transform 1 0 52900 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_565
timestamp 1607194113
transform 1 0 53084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_577
timestamp 1607194113
transform 1 0 54188 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _813_
timestamp 1607194113
transform 1 0 1472 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607194113
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1607194113
transform 1 0 1380 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _606_
timestamp 1607194113
transform 1 0 3956 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__A
timestamp 1607194113
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__813__CLK
timestamp 1607194113
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_25
timestamp 1607194113
transform 1 0 3404 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607194113
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1607194113
transform 1 0 4968 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_54
timestamp 1607194113
transform 1 0 6072 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_60
timestamp 1607194113
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_62
timestamp 1607194113
transform 1 0 6808 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _561_
timestamp 1607194113
transform 1 0 6900 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_37_72
timestamp 1607194113
transform 1 0 7728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _586_
timestamp 1607194113
transform 1 0 9476 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_37_84
timestamp 1607194113
transform 1 0 8832 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_90
timestamp 1607194113
transform 1 0 9384 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_100
timestamp 1607194113
transform 1 0 10304 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _613_
timestamp 1607194113
transform 1 0 11040 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607194113
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_111
timestamp 1607194113
transform 1 0 11316 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_119
timestamp 1607194113
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1607194113
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _567_
timestamp 1607194113
transform 1 0 12880 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_127
timestamp 1607194113
transform 1 0 12788 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_132
timestamp 1607194113
transform 1 0 13248 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_144
timestamp 1607194113
transform 1 0 14352 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _821_
timestamp 1607194113
transform 1 0 15088 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__821__CLK
timestamp 1607194113
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607194113
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1607194113
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_184
timestamp 1607194113
transform 1 0 18032 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _387_
timestamp 1607194113
transform 1 0 19136 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1607194113
transform 1 0 18952 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__C
timestamp 1607194113
transform 1 0 19964 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_192
timestamp 1607194113
transform 1 0 18768 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_207
timestamp 1607194113
transform 1 0 20148 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _391_
timestamp 1607194113
transform 1 0 20700 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1607194113
transform 1 0 21528 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_224
timestamp 1607194113
transform 1 0 21712 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607194113
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__684__B
timestamp 1607194113
transform 1 0 24012 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__684__A
timestamp 1607194113
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_236
timestamp 1607194113
transform 1 0 22816 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_245
timestamp 1607194113
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _384_
timestamp 1607194113
transform 1 0 25576 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _684_
timestamp 1607194113
transform 1 0 24196 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_37_258
timestamp 1607194113
transform 1 0 24840 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1607194113
transform 1 0 25944 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _715_
timestamp 1607194113
transform 1 0 26864 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1607194113
transform 1 0 26680 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1607194113
transform 1 0 29256 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607194113
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__715__A1_N
timestamp 1607194113
transform 1 0 28336 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_298
timestamp 1607194113
transform 1 0 28520 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_304
timestamp 1607194113
transform 1 0 29072 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_309
timestamp 1607194113
transform 1 0 29532 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _569_
timestamp 1607194113
transform 1 0 31372 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_321
timestamp 1607194113
transform 1 0 30636 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _558_
timestamp 1607194113
transform 1 0 33212 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_338
timestamp 1607194113
transform 1 0 32200 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_346
timestamp 1607194113
transform 1 0 32936 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _557_
timestamp 1607194113
transform 1 0 34868 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607194113
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_358
timestamp 1607194113
transform 1 0 34040 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _549_
timestamp 1607194113
transform 1 0 36432 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__C
timestamp 1607194113
transform 1 0 35696 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_378
timestamp 1607194113
transform 1 0 35880 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_388
timestamp 1607194113
transform 1 0 36800 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _705_
timestamp 1607194113
transform 1 0 37536 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_37_412
timestamp 1607194113
transform 1 0 39008 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _390_
timestamp 1607194113
transform 1 0 40480 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607194113
transform 1 0 40388 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_424
timestamp 1607194113
transform 1 0 40112 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_432
timestamp 1607194113
transform 1 0 40848 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _699_
timestamp 1607194113
transform 1 0 42228 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__699__A1_N
timestamp 1607194113
transform 1 0 42044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_444
timestamp 1607194113
transform 1 0 41952 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_463
timestamp 1607194113
transform 1 0 43700 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_475
timestamp 1607194113
transform 1 0 44804 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _622_
timestamp 1607194113
transform 1 0 46092 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607194113
transform 1 0 46000 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_487
timestamp 1607194113
transform 1 0 45908 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_492
timestamp 1607194113
transform 1 0 46368 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _802_
timestamp 1607194113
transform 1 0 48576 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__802__CLK
timestamp 1607194113
transform 1 0 48392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_504
timestamp 1607194113
transform 1 0 47472 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_512
timestamp 1607194113
transform 1 0 48208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_535
timestamp 1607194113
transform 1 0 50324 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _835_
timestamp 1607194113
transform 1 0 52072 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607194113
transform 1 0 51612 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__835__CLK
timestamp 1607194113
transform 1 0 51888 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_547
timestamp 1607194113
transform 1 0 51428 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_550
timestamp 1607194113
transform 1 0 51704 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607194113
transform -1 0 54832 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_573
timestamp 1607194113
transform 1 0 53820 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607194113
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1607194113
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1607194113
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _814_
timestamp 1607194113
transform 1 0 4048 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607194113
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1607194113
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__814__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1607194113
transform 1 0 5980 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _590_
timestamp 1607194113
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_38_65
timestamp 1607194113
transform 1 0 7084 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_73
timestamp 1607194113
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607194113
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_84
timestamp 1607194113
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1607194113
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _582_
timestamp 1607194113
transform 1 0 10948 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_38_105
timestamp 1607194113
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_116
timestamp 1607194113
transform 1 0 11776 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _379_
timestamp 1607194113
transform 1 0 13340 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1607194113
transform 1 0 13156 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_128
timestamp 1607194113
transform 1 0 12880 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_137
timestamp 1607194113
transform 1 0 13708 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _573_
timestamp 1607194113
transform 1 0 15272 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607194113
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__B1
timestamp 1607194113
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1607194113
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1607194113
transform 1 0 18308 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_167
timestamp 1607194113
transform 1 0 16468 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_179
timestamp 1607194113
transform 1 0 17572 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _388_
timestamp 1607194113
transform 1 0 18492 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_38_198
timestamp 1607194113
transform 1 0 19320 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _393_
timestamp 1607194113
transform 1 0 20976 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607194113
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1607194113
transform 1 0 21804 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__B
timestamp 1607194113
transform 1 0 21988 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1607194113
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_215
timestamp 1607194113
transform 1 0 20884 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_229
timestamp 1607194113
transform 1 0 22172 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _385_
timestamp 1607194113
transform 1 0 23092 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1607194113
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_248
timestamp 1607194113
transform 1 0 23920 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _383_
timestamp 1607194113
transform 1 0 24656 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1607194113
transform 1 0 24472 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_260
timestamp 1607194113
transform 1 0 25024 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _392_
timestamp 1607194113
transform 1 0 26496 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _793_
timestamp 1607194113
transform 1 0 27692 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607194113
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_272
timestamp 1607194113
transform 1 0 26128 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_280
timestamp 1607194113
transform 1 0 26864 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_288
timestamp 1607194113
transform 1 0 27600 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__793__CLK
timestamp 1607194113
transform 1 0 29440 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_310
timestamp 1607194113
transform 1 0 29624 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _570_
timestamp 1607194113
transform 1 0 30452 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_38_318
timestamp 1607194113
transform 1 0 30360 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_328
timestamp 1607194113
transform 1 0 31280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _556_
timestamp 1607194113
transform 1 0 32108 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607194113
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_341
timestamp 1607194113
transform 1 0 32476 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_353
timestamp 1607194113
transform 1 0 33580 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _559_
timestamp 1607194113
transform 1 0 33764 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__C
timestamp 1607194113
transform 1 0 34592 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_366
timestamp 1607194113
transform 1 0 34776 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _555_
timestamp 1607194113
transform 1 0 36064 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__C
timestamp 1607194113
transform 1 0 36892 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_378
timestamp 1607194113
transform 1 0 35880 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_391
timestamp 1607194113
transform 1 0 37076 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _800_
timestamp 1607194113
transform 1 0 38548 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607194113
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__800__CLK
timestamp 1607194113
transform 1 0 38364 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_398
timestamp 1607194113
transform 1 0 37720 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_404
timestamp 1607194113
transform 1 0 38272 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _703_
timestamp 1607194113
transform 1 0 41032 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_38_426
timestamp 1607194113
transform 1 0 40296 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607194113
transform 1 0 43240 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_450
timestamp 1607194113
transform 1 0 42504 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _803_
timestamp 1607194113
transform 1 0 44620 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__803__CLK
timestamp 1607194113
transform 1 0 44436 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_459
timestamp 1607194113
transform 1 0 43332 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__B
timestamp 1607194113
transform 1 0 47104 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_492
timestamp 1607194113
transform 1 0 46368 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _548_
timestamp 1607194113
transform 1 0 47288 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607194113
transform 1 0 48852 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__C
timestamp 1607194113
transform 1 0 48116 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_513
timestamp 1607194113
transform 1 0 48300 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_520
timestamp 1607194113
transform 1 0 48944 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_532
timestamp 1607194113
transform 1 0 50048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _545_
timestamp 1607194113
transform 1 0 51612 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A
timestamp 1607194113
transform 1 0 51428 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__B
timestamp 1607194113
transform 1 0 51244 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_544
timestamp 1607194113
transform 1 0 51152 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_558
timestamp 1607194113
transform 1 0 52440 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607194113
transform -1 0 54832 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607194113
transform 1 0 54464 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_570
timestamp 1607194113
transform 1 0 53544 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_578
timestamp 1607194113
transform 1 0 54280 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _812_
timestamp 1607194113
transform 1 0 1380 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607194113
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607194113
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1607194113
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1607194113
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _815_
timestamp 1607194113
transform 1 0 4048 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607194113
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__812__CLK
timestamp 1607194113
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1607194113
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1607194113
transform 1 0 4692 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_24
timestamp 1607194113
transform 1 0 3312 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_30
timestamp 1607194113
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _594_
timestamp 1607194113
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _598_
timestamp 1607194113
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _816_
timestamp 1607194113
transform 1 0 6532 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607194113
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__815__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_43
timestamp 1607194113
transform 1 0 5060 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_53
timestamp 1607194113
transform 1 0 5980 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_53
timestamp 1607194113
transform 1 0 5980 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _818_
timestamp 1607194113
transform 1 0 8464 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__816__CLK
timestamp 1607194113
transform 1 0 8280 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_71
timestamp 1607194113
transform 1 0 7636 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_79
timestamp 1607194113
transform 1 0 8372 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1607194113
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _819_
timestamp 1607194113
transform 1 0 9936 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607194113
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__818__CLK
timestamp 1607194113
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_101
timestamp 1607194113
transform 1 0 10396 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1607194113
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1607194113
transform 1 0 12604 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _820_
timestamp 1607194113
transform 1 0 12420 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607194113
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1607194113
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__819__CLK
timestamp 1607194113
transform 1 0 11684 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1607194113
transform 1 0 11500 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1607194113
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_117
timestamp 1607194113
transform 1 0 11868 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _869_
timestamp 1607194113
transform 1 0 13616 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__820__CLK
timestamp 1607194113
transform 1 0 14168 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_128
timestamp 1607194113
transform 1 0 12880 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_144
timestamp 1607194113
transform 1 0 14352 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _870_
timestamp 1607194113
transform 1 0 15272 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607194113
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__869__CLK
timestamp 1607194113
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__870__CLK
timestamp 1607194113
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_157
timestamp 1607194113
transform 1 0 15548 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_150
timestamp 1607194113
transform 1 0 14904 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _871_
timestamp 1607194113
transform 1 0 17756 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _872_
timestamp 1607194113
transform 1 0 18032 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607194113
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__871__CLK
timestamp 1607194113
transform 1 0 17572 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__872__CLK
timestamp 1607194113
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1607194113
transform 1 0 16652 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_173
timestamp 1607194113
transform 1 0 17020 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_203
timestamp 1607194113
transform 1 0 19780 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_200
timestamp 1607194113
transform 1 0 19504 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _386_
timestamp 1607194113
transform 1 0 21988 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _873_
timestamp 1607194113
transform 1 0 20884 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607194113
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1607194113
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__873__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1607194113
transform 1 0 20884 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_223
timestamp 1607194113
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _875_
timestamp 1607194113
transform 1 0 23368 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607194113
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__C
timestamp 1607194113
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__875__CLK
timestamp 1607194113
transform 1 0 23184 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_238
timestamp 1607194113
transform 1 0 23000 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1607194113
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_234
timestamp 1607194113
transform 1 0 22632 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _822_
timestamp 1607194113
transform 1 0 25392 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__822__CLK
timestamp 1607194113
transform 1 0 25208 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_257
timestamp 1607194113
transform 1 0 24748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_261
timestamp 1607194113
transform 1 0 25116 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_261
timestamp 1607194113
transform 1 0 25116 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _823_
timestamp 1607194113
transform 1 0 26496 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607194113
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__823__CLK
timestamp 1607194113
transform 1 0 26220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_283
timestamp 1607194113
transform 1 0 27140 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _825_
timestamp 1607194113
transform 1 0 28980 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607194113
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_295
timestamp 1607194113
transform 1 0 28244 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_303
timestamp 1607194113
transform 1 0 28980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_306
timestamp 1607194113
transform 1 0 29256 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_295
timestamp 1607194113
transform 1 0 28244 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _826_
timestamp 1607194113
transform 1 0 30544 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__825__CLK
timestamp 1607194113
transform 1 0 30728 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_318
timestamp 1607194113
transform 1 0 30360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_324
timestamp 1607194113
transform 1 0 30912 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _560_
timestamp 1607194113
transform 1 0 33212 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _827_
timestamp 1607194113
transform 1 0 32292 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607194113
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__826__CLK
timestamp 1607194113
transform 1 0 32292 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_341
timestamp 1607194113
transform 1 0 32476 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1607194113
transform 1 0 32108 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _554_
timestamp 1607194113
transform 1 0 34960 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _828_
timestamp 1607194113
transform 1 0 34776 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607194113
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__827__CLK
timestamp 1607194113
transform 1 0 34040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_358
timestamp 1607194113
transform 1 0 34040 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_367
timestamp 1607194113
transform 1 0 34868 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_372
timestamp 1607194113
transform 1 0 35328 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_360
timestamp 1607194113
transform 1 0 34224 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _829_
timestamp 1607194113
transform 1 0 36064 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__828__CLK
timestamp 1607194113
transform 1 0 36524 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__829__CLK
timestamp 1607194113
transform 1 0 35880 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_387
timestamp 1607194113
transform 1 0 36708 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_395
timestamp 1607194113
transform 1 0 37444 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _552_
timestamp 1607194113
transform 1 0 38824 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _831_
timestamp 1607194113
transform 1 0 38456 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607194113
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_399
timestamp 1607194113
transform 1 0 37812 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_407
timestamp 1607194113
transform 1 0 38548 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_398
timestamp 1607194113
transform 1 0 37720 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1607194113
transform 1 0 40480 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607194113
transform 1 0 40388 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__831__CLK
timestamp 1607194113
transform 1 0 40204 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_419
timestamp 1607194113
transform 1 0 39652 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_431
timestamp 1607194113
transform 1 0 40756 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_427
timestamp 1607194113
transform 1 0 40388 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _551_
timestamp 1607194113
transform 1 0 41492 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607194113
transform 1 0 43240 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_448
timestamp 1607194113
transform 1 0 42320 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_439
timestamp 1607194113
transform 1 0 41492 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_451
timestamp 1607194113
transform 1 0 42596 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_457
timestamp 1607194113
transform 1 0 43148 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _550_
timestamp 1607194113
transform 1 0 43792 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_39_460
timestamp 1607194113
transform 1 0 43424 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1607194113
transform 1 0 44620 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_459
timestamp 1607194113
transform 1 0 43332 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_471
timestamp 1607194113
transform 1 0 44436 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _553_
timestamp 1607194113
transform 1 0 46092 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _830_
timestamp 1607194113
transform 1 0 45908 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607194113
transform 1 0 46000 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__830__CLK
timestamp 1607194113
transform 1 0 45724 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_485
timestamp 1607194113
transform 1 0 45724 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_498
timestamp 1607194113
transform 1 0 46920 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_483
timestamp 1607194113
transform 1 0 45540 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _810_
timestamp 1607194113
transform 1 0 48116 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607194113
transform 1 0 48852 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__810__D
timestamp 1607194113
transform 1 0 47932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__810__CLK
timestamp 1607194113
transform 1 0 47748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_506
timestamp 1607194113
transform 1 0 47656 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_506
timestamp 1607194113
transform 1 0 47656 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_518
timestamp 1607194113
transform 1 0 48760 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_520
timestamp 1607194113
transform 1 0 48944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__768__D
timestamp 1607194113
transform 1 0 50784 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__768__CLK
timestamp 1607194113
transform 1 0 50600 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_530
timestamp 1607194113
transform 1 0 49864 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_532
timestamp 1607194113
transform 1 0 50048 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _768_
timestamp 1607194113
transform 1 0 50968 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _836_
timestamp 1607194113
transform 1 0 52072 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607194113
transform 1 0 51612 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__836__CLK
timestamp 1607194113
transform 1 0 51888 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_542
timestamp 1607194113
transform 1 0 50968 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_548
timestamp 1607194113
transform 1 0 51520 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_550
timestamp 1607194113
transform 1 0 51704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_561
timestamp 1607194113
transform 1 0 52716 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607194113
transform -1 0 54832 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607194113
transform -1 0 54832 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607194113
transform 1 0 54464 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_573
timestamp 1607194113
transform 1 0 53820 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_573
timestamp 1607194113
transform 1 0 53820 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_579
timestamp 1607194113
transform 1 0 54372 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607194113
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1607194113
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1607194113
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607194113
transform 1 0 3956 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1607194113
transform 1 0 3588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_32
timestamp 1607194113
transform 1 0 4048 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607194113
transform 1 0 6808 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_44
timestamp 1607194113
transform 1 0 5152 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_56
timestamp 1607194113
transform 1 0 6256 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _817_
timestamp 1607194113
transform 1 0 6900 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__817__CLK
timestamp 1607194113
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607194113
transform 1 0 9660 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_84
timestamp 1607194113
transform 1 0 8832 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_92
timestamp 1607194113
transform 1 0 9568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1607194113
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607194113
transform 1 0 12512 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_106
timestamp 1607194113
transform 1 0 10856 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_118
timestamp 1607194113
transform 1 0 11960 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1607194113
transform 1 0 12604 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1607194113
transform 1 0 13708 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607194113
transform 1 0 15364 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_149
timestamp 1607194113
transform 1 0 14812 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_156
timestamp 1607194113
transform 1 0 15456 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607194113
transform 1 0 18216 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_168
timestamp 1607194113
transform 1 0 16560 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_180
timestamp 1607194113
transform 1 0 17664 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_187
timestamp 1607194113
transform 1 0 18308 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_199
timestamp 1607194113
transform 1 0 19412 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _874_
timestamp 1607194113
transform 1 0 21436 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607194113
transform 1 0 21068 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__874__CLK
timestamp 1607194113
transform 1 0 21252 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_211
timestamp 1607194113
transform 1 0 20516 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_218
timestamp 1607194113
transform 1 0 21160 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607194113
transform 1 0 23920 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_240
timestamp 1607194113
transform 1 0 23184 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1607194113
transform 1 0 24012 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1607194113
transform 1 0 25116 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607194113
transform 1 0 26772 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1607194113
transform 1 0 26220 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_280
timestamp 1607194113
transform 1 0 26864 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607194113
transform 1 0 29624 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_292
timestamp 1607194113
transform 1 0 27968 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_304
timestamp 1607194113
transform 1 0 29072 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_311
timestamp 1607194113
transform 1 0 29716 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_323
timestamp 1607194113
transform 1 0 30820 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607194113
transform 1 0 32476 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_335
timestamp 1607194113
transform 1 0 31924 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_342
timestamp 1607194113
transform 1 0 32568 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_354
timestamp 1607194113
transform 1 0 33672 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607194113
transform 1 0 35328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_366
timestamp 1607194113
transform 1 0 34776 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1607194113
transform 1 0 35420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_385
timestamp 1607194113
transform 1 0 36524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _389_
timestamp 1607194113
transform 1 0 38640 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607194113
transform 1 0 38180 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1607194113
transform 1 0 38456 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_397
timestamp 1607194113
transform 1 0 37628 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_404
timestamp 1607194113
transform 1 0 38272 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_412
timestamp 1607194113
transform 1 0 39008 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _547_
timestamp 1607194113
transform 1 0 39744 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _832_
timestamp 1607194113
transform 1 0 41216 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607194113
transform 1 0 41032 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_424
timestamp 1607194113
transform 1 0 40112 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_432
timestamp 1607194113
transform 1 0 40848 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_435
timestamp 1607194113
transform 1 0 41124 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__832__CLK
timestamp 1607194113
transform 1 0 42964 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_457
timestamp 1607194113
transform 1 0 43148 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _833_
timestamp 1607194113
transform 1 0 43976 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607194113
transform 1 0 43884 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__833__CLK
timestamp 1607194113
transform 1 0 43700 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607194113
transform 1 0 46736 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_485
timestamp 1607194113
transform 1 0 45724 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_493
timestamp 1607194113
transform 1 0 46460 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_497
timestamp 1607194113
transform 1 0 46828 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_509
timestamp 1607194113
transform 1 0 47932 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _834_
timestamp 1607194113
transform 1 0 49680 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607194113
transform 1 0 49588 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__834__CLK
timestamp 1607194113
transform 1 0 49404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_521
timestamp 1607194113
transform 1 0 49036 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607194113
transform 1 0 52440 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_547
timestamp 1607194113
transform 1 0 51428 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_555
timestamp 1607194113
transform 1 0 52164 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_559
timestamp 1607194113
transform 1 0 52532 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607194113
transform -1 0 54832 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_571
timestamp 1607194113
transform 1 0 53636 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_579
timestamp 1607194113
transform 1 0 54372 0 1 24480
box -38 -48 222 592
<< labels >>
rlabel metal2 s 938 26400 994 27200 6 bus_in[0]
port 0 nsew default input
rlabel metal2 s 15290 26400 15346 27200 6 bus_in[10]
port 1 nsew default input
rlabel metal2 s 16762 26400 16818 27200 6 bus_in[11]
port 2 nsew default input
rlabel metal2 s 18234 26400 18290 27200 6 bus_in[12]
port 3 nsew default input
rlabel metal2 s 19614 26400 19670 27200 6 bus_in[13]
port 4 nsew default input
rlabel metal2 s 21086 26400 21142 27200 6 bus_in[14]
port 5 nsew default input
rlabel metal2 s 22558 26400 22614 27200 6 bus_in[15]
port 6 nsew default input
rlabel metal2 s 23938 26400 23994 27200 6 bus_in[16]
port 7 nsew default input
rlabel metal2 s 25410 26400 25466 27200 6 bus_in[17]
port 8 nsew default input
rlabel metal2 s 26790 26400 26846 27200 6 bus_in[18]
port 9 nsew default input
rlabel metal2 s 28262 26400 28318 27200 6 bus_in[19]
port 10 nsew default input
rlabel metal2 s 2410 26400 2466 27200 6 bus_in[1]
port 11 nsew default input
rlabel metal2 s 29734 26400 29790 27200 6 bus_in[20]
port 12 nsew default input
rlabel metal2 s 31114 26400 31170 27200 6 bus_in[21]
port 13 nsew default input
rlabel metal2 s 32586 26400 32642 27200 6 bus_in[22]
port 14 nsew default input
rlabel metal2 s 33966 26400 34022 27200 6 bus_in[23]
port 15 nsew default input
rlabel metal2 s 35438 26400 35494 27200 6 bus_in[24]
port 16 nsew default input
rlabel metal2 s 36910 26400 36966 27200 6 bus_in[25]
port 17 nsew default input
rlabel metal2 s 38290 26400 38346 27200 6 bus_in[26]
port 18 nsew default input
rlabel metal2 s 39762 26400 39818 27200 6 bus_in[27]
port 19 nsew default input
rlabel metal2 s 41234 26400 41290 27200 6 bus_in[28]
port 20 nsew default input
rlabel metal2 s 42614 26400 42670 27200 6 bus_in[29]
port 21 nsew default input
rlabel metal2 s 3882 26400 3938 27200 6 bus_in[2]
port 22 nsew default input
rlabel metal2 s 44086 26400 44142 27200 6 bus_in[30]
port 23 nsew default input
rlabel metal2 s 45466 26400 45522 27200 6 bus_in[31]
port 24 nsew default input
rlabel metal2 s 46938 26400 46994 27200 6 bus_in[32]
port 25 nsew default input
rlabel metal2 s 48410 26400 48466 27200 6 bus_in[33]
port 26 nsew default input
rlabel metal2 s 49790 26400 49846 27200 6 bus_in[34]
port 27 nsew default input
rlabel metal2 s 51262 26400 51318 27200 6 bus_in[35]
port 28 nsew default input
rlabel metal2 s 51998 26400 52054 27200 6 bus_in[36]
port 29 nsew default input
rlabel metal2 s 52642 26400 52698 27200 6 bus_in[37]
port 30 nsew default input
rlabel metal2 s 53378 26400 53434 27200 6 bus_in[38]
port 31 nsew default input
rlabel metal2 s 54114 26400 54170 27200 6 bus_in[39]
port 32 nsew default input
rlabel metal2 s 5262 26400 5318 27200 6 bus_in[3]
port 33 nsew default input
rlabel metal2 s 54850 26400 54906 27200 6 bus_in[40]
port 34 nsew default input
rlabel metal2 s 55586 26400 55642 27200 6 bus_in[41]
port 35 nsew default input
rlabel metal2 s 6734 26400 6790 27200 6 bus_in[4]
port 36 nsew default input
rlabel metal2 s 8114 26400 8170 27200 6 bus_in[5]
port 37 nsew default input
rlabel metal2 s 9586 26400 9642 27200 6 bus_in[6]
port 38 nsew default input
rlabel metal2 s 11058 26400 11114 27200 6 bus_in[7]
port 39 nsew default input
rlabel metal2 s 12438 26400 12494 27200 6 bus_in[8]
port 40 nsew default input
rlabel metal2 s 13910 26400 13966 27200 6 bus_in[9]
port 41 nsew default input
rlabel metal2 s 1674 26400 1730 27200 6 bus_out[0]
port 42 nsew default tristate
rlabel metal2 s 16026 26400 16082 27200 6 bus_out[10]
port 43 nsew default tristate
rlabel metal2 s 17498 26400 17554 27200 6 bus_out[11]
port 44 nsew default tristate
rlabel metal2 s 18970 26400 19026 27200 6 bus_out[12]
port 45 nsew default tristate
rlabel metal2 s 20350 26400 20406 27200 6 bus_out[13]
port 46 nsew default tristate
rlabel metal2 s 21822 26400 21878 27200 6 bus_out[14]
port 47 nsew default tristate
rlabel metal2 s 23202 26400 23258 27200 6 bus_out[15]
port 48 nsew default tristate
rlabel metal2 s 24674 26400 24730 27200 6 bus_out[16]
port 49 nsew default tristate
rlabel metal2 s 26146 26400 26202 27200 6 bus_out[17]
port 50 nsew default tristate
rlabel metal2 s 27526 26400 27582 27200 6 bus_out[18]
port 51 nsew default tristate
rlabel metal2 s 28998 26400 29054 27200 6 bus_out[19]
port 52 nsew default tristate
rlabel metal2 s 3146 26400 3202 27200 6 bus_out[1]
port 53 nsew default tristate
rlabel metal2 s 30378 26400 30434 27200 6 bus_out[20]
port 54 nsew default tristate
rlabel metal2 s 31850 26400 31906 27200 6 bus_out[21]
port 55 nsew default tristate
rlabel metal2 s 33322 26400 33378 27200 6 bus_out[22]
port 56 nsew default tristate
rlabel metal2 s 34702 26400 34758 27200 6 bus_out[23]
port 57 nsew default tristate
rlabel metal2 s 36174 26400 36230 27200 6 bus_out[24]
port 58 nsew default tristate
rlabel metal2 s 37646 26400 37702 27200 6 bus_out[25]
port 59 nsew default tristate
rlabel metal2 s 39026 26400 39082 27200 6 bus_out[26]
port 60 nsew default tristate
rlabel metal2 s 40498 26400 40554 27200 6 bus_out[27]
port 61 nsew default tristate
rlabel metal2 s 41878 26400 41934 27200 6 bus_out[28]
port 62 nsew default tristate
rlabel metal2 s 43350 26400 43406 27200 6 bus_out[29]
port 63 nsew default tristate
rlabel metal2 s 4526 26400 4582 27200 6 bus_out[2]
port 64 nsew default tristate
rlabel metal2 s 44822 26400 44878 27200 6 bus_out[30]
port 65 nsew default tristate
rlabel metal2 s 46202 26400 46258 27200 6 bus_out[31]
port 66 nsew default tristate
rlabel metal2 s 47674 26400 47730 27200 6 bus_out[32]
port 67 nsew default tristate
rlabel metal2 s 49054 26400 49110 27200 6 bus_out[33]
port 68 nsew default tristate
rlabel metal2 s 50526 26400 50582 27200 6 bus_out[34]
port 69 nsew default tristate
rlabel metal2 s 5998 26400 6054 27200 6 bus_out[3]
port 70 nsew default tristate
rlabel metal2 s 7470 26400 7526 27200 6 bus_out[4]
port 71 nsew default tristate
rlabel metal2 s 8850 26400 8906 27200 6 bus_out[5]
port 72 nsew default tristate
rlabel metal2 s 10322 26400 10378 27200 6 bus_out[6]
port 73 nsew default tristate
rlabel metal2 s 11702 26400 11758 27200 6 bus_out[7]
port 74 nsew default tristate
rlabel metal2 s 13174 26400 13230 27200 6 bus_out[8]
port 75 nsew default tristate
rlabel metal2 s 14646 26400 14702 27200 6 bus_out[9]
port 76 nsew default tristate
rlabel metal3 s 55200 6808 56000 6928 6 clk_i
port 77 nsew default input
rlabel metal3 s 55200 20408 56000 20528 6 out_o
port 78 nsew default tristate
rlabel metal2 s 294 26400 350 27200 6 rst_n_i
port 79 nsew default input
rlabel metal4 s 9909 2128 10229 25072 6 VPWR
port 80 nsew default input
rlabel metal4 s 18875 2128 19195 25072 6 VGND
port 81 nsew default input
<< properties >>
string FIXED_BBOX 0 0 56000 27200
<< end >>
