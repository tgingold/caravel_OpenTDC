VERSION 5.7 ;
NOWIREEXTENSIONATPIN ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
MACRO rescue_top
  CLASS BLOCK ;
  FOREIGN rescue_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 736.000 BY 223.040 ;
  PIN clk_i
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 732.000 111.560 736.000 112.160 ;
    END
  END clk_i
  PIN fd_oen_o
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 0.000 167.320 4.000 167.920 ;
    END
  END fd_oen_o
  PIN fd_out_o
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 0.000 55.800 4.000 56.400 ;
    END
  END fd_out_o
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 1.010 0.000 1.290 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 576.010 0.000 576.290 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 581.530 0.000 581.810 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 587.510 0.000 587.790 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 593.030 0.000 593.310 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 604.530 0.000 604.810 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 616.030 0.000 616.310 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 622.010 0.000 622.290 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 627.530 0.000 627.810 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 58.510 0.000 58.790 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 633.510 0.000 633.790 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 639.030 0.000 639.310 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 645.010 0.000 645.290 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 662.030 0.000 662.310 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 668.010 0.000 668.290 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 679.510 0.000 679.790 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 685.030 0.000 685.310 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 64.030 0.000 64.310 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 691.010 0.000 691.290 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 696.530 0.000 696.810 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 708.030 0.000 708.310 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 714.010 0.000 714.290 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 719.530 0.000 719.810 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 731.030 0.000 731.310 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 70.010 0.000 70.290 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 75.530 0.000 75.810 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 81.510 0.000 81.790 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 87.030 0.000 87.310 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 93.010 0.000 93.290 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 98.530 0.000 98.810 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 104.510 0.000 104.790 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 110.030 0.000 110.310 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 6.530 0.000 6.810 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 116.010 0.000 116.290 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 121.530 0.000 121.810 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 127.510 0.000 127.790 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 133.030 0.000 133.310 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 139.010 0.000 139.290 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 144.530 0.000 144.810 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 150.510 0.000 150.790 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 156.030 0.000 156.310 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 162.010 0.000 162.290 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 167.530 0.000 167.810 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 12.510 0.000 12.790 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 173.510 0.000 173.790 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 179.030 0.000 179.310 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 185.010 0.000 185.290 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 190.530 0.000 190.810 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 196.510 0.000 196.790 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 202.030 0.000 202.310 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 208.010 0.000 208.290 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 213.530 0.000 213.810 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 219.510 0.000 219.790 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 225.030 0.000 225.310 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 18.030 0.000 18.310 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 231.010 0.000 231.290 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 242.510 0.000 242.790 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 248.030 0.000 248.310 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 254.010 0.000 254.290 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 259.530 0.000 259.810 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 265.510 0.000 265.790 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 271.030 0.000 271.310 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 277.010 0.000 277.290 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 282.530 0.000 282.810 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 24.010 0.000 24.290 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 288.510 0.000 288.790 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 294.030 0.000 294.310 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 300.010 0.000 300.290 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 305.530 0.000 305.810 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 311.510 0.000 311.790 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 317.030 0.000 317.310 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 323.010 0.000 323.290 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 334.510 0.000 334.790 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 29.530 0.000 29.810 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 346.010 0.000 346.290 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 351.530 0.000 351.810 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 363.030 0.000 363.310 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 369.010 0.000 369.290 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 374.530 0.000 374.810 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 380.510 0.000 380.790 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 392.010 0.000 392.290 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 397.530 0.000 397.810 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 35.510 0.000 35.790 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 403.510 0.000 403.790 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 409.030 0.000 409.310 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 415.010 0.000 415.290 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 420.530 0.000 420.810 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 426.510 0.000 426.790 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 432.030 0.000 432.310 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 443.530 0.000 443.810 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 455.030 0.000 455.310 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 41.030 0.000 41.310 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 466.530 0.000 466.810 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 472.510 0.000 472.790 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 484.010 0.000 484.290 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 489.530 0.000 489.810 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 495.510 0.000 495.790 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 501.030 0.000 501.310 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 507.010 0.000 507.290 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 512.530 0.000 512.810 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 47.010 0.000 47.290 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 524.030 0.000 524.310 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 530.010 0.000 530.290 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 541.510 0.000 541.790 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 547.030 0.000 547.310 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 553.010 0.000 553.290 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 558.530 0.000 558.810 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 564.510 0.000 564.790 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 52.530 0.000 52.810 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 577.850 0.000 578.130 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 583.370 0.000 583.650 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 600.850 0.000 601.130 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 606.370 0.000 606.650 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 612.350 0.000 612.630 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 617.870 0.000 618.150 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 623.850 0.000 624.130 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 629.370 0.000 629.650 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 60.350 0.000 60.630 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 635.350 0.000 635.630 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 640.870 0.000 641.150 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 646.850 0.000 647.130 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 652.370 0.000 652.650 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 658.350 0.000 658.630 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 675.370 0.000 675.650 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 681.350 0.000 681.630 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 686.870 0.000 687.150 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 65.870 0.000 66.150 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 704.350 0.000 704.630 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 709.870 0.000 710.150 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 715.850 0.000 716.130 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 721.370 0.000 721.650 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 71.850 0.000 72.130 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 83.350 0.000 83.630 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 88.870 0.000 89.150 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 94.850 0.000 95.130 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 100.370 0.000 100.650 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 106.350 0.000 106.630 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 111.870 0.000 112.150 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 8.370 0.000 8.650 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 117.850 0.000 118.130 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 123.370 0.000 123.650 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 129.350 0.000 129.630 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 134.870 0.000 135.150 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 140.850 0.000 141.130 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 146.370 0.000 146.650 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 152.350 0.000 152.630 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 163.850 0.000 164.130 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 169.370 0.000 169.650 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 14.350 0.000 14.630 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 180.870 0.000 181.150 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 186.850 0.000 187.130 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 192.370 0.000 192.650 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 198.350 0.000 198.630 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 209.850 0.000 210.130 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 215.370 0.000 215.650 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 221.350 0.000 221.630 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 226.870 0.000 227.150 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 19.870 0.000 20.150 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 232.850 0.000 233.130 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 238.370 0.000 238.650 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 244.350 0.000 244.630 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 249.870 0.000 250.150 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 255.850 0.000 256.130 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 261.370 0.000 261.650 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 267.350 0.000 267.630 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 272.870 0.000 273.150 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 284.370 0.000 284.650 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 290.350 0.000 290.630 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 295.870 0.000 296.150 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 301.850 0.000 302.130 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 307.370 0.000 307.650 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 313.350 0.000 313.630 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 318.870 0.000 319.150 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 324.850 0.000 325.130 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 330.370 0.000 330.650 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 336.350 0.000 336.630 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 341.870 0.000 342.150 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 31.370 0.000 31.650 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 353.370 0.000 353.650 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 359.350 0.000 359.630 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 364.870 0.000 365.150 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 370.850 0.000 371.130 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 376.370 0.000 376.650 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 387.870 0.000 388.150 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 393.850 0.000 394.130 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 37.350 0.000 37.630 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 405.350 0.000 405.630 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 410.870 0.000 411.150 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 416.850 0.000 417.130 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 422.370 0.000 422.650 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 428.350 0.000 428.630 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 433.870 0.000 434.150 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 439.850 0.000 440.130 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 445.370 0.000 445.650 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 456.870 0.000 457.150 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 42.870 0.000 43.150 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 462.850 0.000 463.130 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 468.370 0.000 468.650 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 474.350 0.000 474.630 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 479.870 0.000 480.150 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 491.370 0.000 491.650 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 497.350 0.000 497.630 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 502.870 0.000 503.150 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 514.370 0.000 514.650 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 48.850 0.000 49.130 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 520.350 0.000 520.630 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 525.870 0.000 526.150 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 531.850 0.000 532.130 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 537.370 0.000 537.650 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 543.350 0.000 543.630 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 548.870 0.000 549.150 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 554.850 0.000 555.130 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 566.350 0.000 566.630 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 571.870 0.000 572.150 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met2 ;
      RECT 54.370 0.000 54.650 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 4.690 0.000 4.970 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 579.690 0.000 579.970 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 585.210 0.000 585.490 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 591.190 0.000 591.470 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 596.710 0.000 596.990 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 602.690 0.000 602.970 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 608.210 0.000 608.490 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 631.210 0.000 631.490 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 62.190 0.000 62.470 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 637.190 0.000 637.470 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 648.690 0.000 648.970 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 654.210 0.000 654.490 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 665.710 0.000 665.990 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 671.690 0.000 671.970 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 677.210 0.000 677.490 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 683.190 0.000 683.470 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 688.710 0.000 688.990 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 694.690 0.000 694.970 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 706.190 0.000 706.470 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 717.690 0.000 717.970 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 723.210 0.000 723.490 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 734.710 0.000 734.990 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 73.690 0.000 73.970 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 79.210 0.000 79.490 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 85.190 0.000 85.470 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 90.710 0.000 90.990 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 102.210 0.000 102.490 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 108.190 0.000 108.470 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 113.710 0.000 113.990 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 10.210 0.000 10.490 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 119.690 0.000 119.970 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 125.210 0.000 125.490 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 131.190 0.000 131.470 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 136.710 0.000 136.990 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 142.690 0.000 142.970 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 148.210 0.000 148.490 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 154.190 0.000 154.470 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 159.710 0.000 159.990 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 165.690 0.000 165.970 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 171.210 0.000 171.490 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 177.190 0.000 177.470 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 182.710 0.000 182.990 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 188.690 0.000 188.970 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 194.210 0.000 194.490 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 200.190 0.000 200.470 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 205.710 0.000 205.990 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 211.690 0.000 211.970 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 217.210 0.000 217.490 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 223.190 0.000 223.470 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 21.710 0.000 21.990 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 234.690 0.000 234.970 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 240.210 0.000 240.490 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 246.190 0.000 246.470 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 251.710 0.000 251.990 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 257.690 0.000 257.970 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 263.210 0.000 263.490 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 274.710 0.000 274.990 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 280.690 0.000 280.970 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 286.210 0.000 286.490 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 27.690 0.000 27.970 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 292.190 0.000 292.470 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 297.710 0.000 297.990 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 303.690 0.000 303.970 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 309.210 0.000 309.490 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 320.710 0.000 320.990 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 326.690 0.000 326.970 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 332.210 0.000 332.490 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 343.710 0.000 343.990 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 33.210 0.000 33.490 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 349.690 0.000 349.970 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 355.210 0.000 355.490 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 361.190 0.000 361.470 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 366.710 0.000 366.990 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 372.690 0.000 372.970 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 401.210 0.000 401.490 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 39.190 0.000 39.470 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 407.190 0.000 407.470 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 412.710 0.000 412.990 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 424.210 0.000 424.490 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 430.190 0.000 430.470 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 435.710 0.000 435.990 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 441.690 0.000 441.970 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 458.710 0.000 458.990 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 44.710 0.000 44.990 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 464.690 0.000 464.970 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 470.210 0.000 470.490 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 476.190 0.000 476.470 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 487.690 0.000 487.970 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 493.210 0.000 493.490 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 499.190 0.000 499.470 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 504.710 0.000 504.990 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 510.690 0.000 510.970 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 516.210 0.000 516.490 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 50.690 0.000 50.970 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 527.710 0.000 527.990 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 533.690 0.000 533.970 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 545.190 0.000 545.470 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 550.710 0.000 550.990 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 562.210 0.000 562.490 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 568.190 0.000 568.470 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 573.710 0.000 573.990 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 56.210 0.000 56.490 4.000 ;
    END
  END la_oen[9]
  PIN tdc_inp_i
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 368.090 219.040 368.370 223.040 ;
    END
  END tdc_inp_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT 
      LAYER met4 ;
      RECT 174.64 10.64 176.24 212.4 ;
      RECT 328.24 10.64 329.84 212.4 ;
      RECT 481.84 10.64 483.44 212.4 ;
      RECT 635.44 10.64 637.04 212.4 ;
      RECT 21.040 10.640 22.640 212.400 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT 
      LAYER met4 ;
      RECT 251.44 10.64 253.04 212.4 ;
      RECT 405.04 10.64 406.64 212.4 ;
      RECT 558.64 10.64 560.24 212.4 ;
      RECT 712.24 10.64 713.84 212.4 ;
      RECT 97.840 10.640 99.440 212.400 ;
    END
  END VGND
  OBS 
    LAYER li1 ;
    RECT 5.520 10.795 730.480 212.245 ;
    LAYER met1 ;
    RECT 2.830 7.180 733.170 212.400 ;
    LAYER met2 ;
    RECT 2.860 218.760 367.810 219.040 ;
    RECT 368.650 218.760 733.140 219.040 ;
    RECT 2.860 4.280 733.140 218.760 ;
    RECT 3.410 4.000 4.410 4.280 ;
    RECT 5.250 4.000 6.250 4.280 ;
    RECT 7.090 4.000 8.090 4.280 ;
    RECT 8.930 4.000 9.930 4.280 ;
    RECT 10.770 4.000 12.230 4.280 ;
    RECT 13.070 4.000 14.070 4.280 ;
    RECT 14.910 4.000 15.910 4.280 ;
    RECT 16.750 4.000 17.750 4.280 ;
    RECT 18.590 4.000 19.590 4.280 ;
    RECT 20.430 4.000 21.430 4.280 ;
    RECT 22.270 4.000 23.730 4.280 ;
    RECT 24.570 4.000 25.570 4.280 ;
    RECT 26.410 4.000 27.410 4.280 ;
    RECT 28.250 4.000 29.250 4.280 ;
    RECT 30.090 4.000 31.090 4.280 ;
    RECT 31.930 4.000 32.930 4.280 ;
    RECT 33.770 4.000 35.230 4.280 ;
    RECT 36.070 4.000 37.070 4.280 ;
    RECT 37.910 4.000 38.910 4.280 ;
    RECT 39.750 4.000 40.750 4.280 ;
    RECT 41.590 4.000 42.590 4.280 ;
    RECT 43.430 4.000 44.430 4.280 ;
    RECT 45.270 4.000 46.730 4.280 ;
    RECT 47.570 4.000 48.570 4.280 ;
    RECT 49.410 4.000 50.410 4.280 ;
    RECT 51.250 4.000 52.250 4.280 ;
    RECT 53.090 4.000 54.090 4.280 ;
    RECT 54.930 4.000 55.930 4.280 ;
    RECT 56.770 4.000 58.230 4.280 ;
    RECT 59.070 4.000 60.070 4.280 ;
    RECT 60.910 4.000 61.910 4.280 ;
    RECT 62.750 4.000 63.750 4.280 ;
    RECT 64.590 4.000 65.590 4.280 ;
    RECT 66.430 4.000 67.430 4.280 ;
    RECT 68.270 4.000 69.730 4.280 ;
    RECT 70.570 4.000 71.570 4.280 ;
    RECT 72.410 4.000 73.410 4.280 ;
    RECT 74.250 4.000 75.250 4.280 ;
    RECT 76.090 4.000 77.090 4.280 ;
    RECT 77.930 4.000 78.930 4.280 ;
    RECT 79.770 4.000 81.230 4.280 ;
    RECT 82.070 4.000 83.070 4.280 ;
    RECT 83.910 4.000 84.910 4.280 ;
    RECT 85.750 4.000 86.750 4.280 ;
    RECT 87.590 4.000 88.590 4.280 ;
    RECT 89.430 4.000 90.430 4.280 ;
    RECT 91.270 4.000 92.730 4.280 ;
    RECT 93.570 4.000 94.570 4.280 ;
    RECT 95.410 4.000 96.410 4.280 ;
    RECT 97.250 4.000 98.250 4.280 ;
    RECT 99.090 4.000 100.090 4.280 ;
    RECT 100.930 4.000 101.930 4.280 ;
    RECT 102.770 4.000 104.230 4.280 ;
    RECT 105.070 4.000 106.070 4.280 ;
    RECT 106.910 4.000 107.910 4.280 ;
    RECT 108.750 4.000 109.750 4.280 ;
    RECT 110.590 4.000 111.590 4.280 ;
    RECT 112.430 4.000 113.430 4.280 ;
    RECT 114.270 4.000 115.730 4.280 ;
    RECT 116.570 4.000 117.570 4.280 ;
    RECT 118.410 4.000 119.410 4.280 ;
    RECT 120.250 4.000 121.250 4.280 ;
    RECT 122.090 4.000 123.090 4.280 ;
    RECT 123.930 4.000 124.930 4.280 ;
    RECT 125.770 4.000 127.230 4.280 ;
    RECT 128.070 4.000 129.070 4.280 ;
    RECT 129.910 4.000 130.910 4.280 ;
    RECT 131.750 4.000 132.750 4.280 ;
    RECT 133.590 4.000 134.590 4.280 ;
    RECT 135.430 4.000 136.430 4.280 ;
    RECT 137.270 4.000 138.730 4.280 ;
    RECT 139.570 4.000 140.570 4.280 ;
    RECT 141.410 4.000 142.410 4.280 ;
    RECT 143.250 4.000 144.250 4.280 ;
    RECT 145.090 4.000 146.090 4.280 ;
    RECT 146.930 4.000 147.930 4.280 ;
    RECT 148.770 4.000 150.230 4.280 ;
    RECT 151.070 4.000 152.070 4.280 ;
    RECT 152.910 4.000 153.910 4.280 ;
    RECT 154.750 4.000 155.750 4.280 ;
    RECT 156.590 4.000 157.590 4.280 ;
    RECT 158.430 4.000 159.430 4.280 ;
    RECT 160.270 4.000 161.730 4.280 ;
    RECT 162.570 4.000 163.570 4.280 ;
    RECT 164.410 4.000 165.410 4.280 ;
    RECT 166.250 4.000 167.250 4.280 ;
    RECT 168.090 4.000 169.090 4.280 ;
    RECT 169.930 4.000 170.930 4.280 ;
    RECT 171.770 4.000 173.230 4.280 ;
    RECT 174.070 4.000 175.070 4.280 ;
    RECT 175.910 4.000 176.910 4.280 ;
    RECT 177.750 4.000 178.750 4.280 ;
    RECT 179.590 4.000 180.590 4.280 ;
    RECT 181.430 4.000 182.430 4.280 ;
    RECT 183.270 4.000 184.730 4.280 ;
    RECT 185.570 4.000 186.570 4.280 ;
    RECT 187.410 4.000 188.410 4.280 ;
    RECT 189.250 4.000 190.250 4.280 ;
    RECT 191.090 4.000 192.090 4.280 ;
    RECT 192.930 4.000 193.930 4.280 ;
    RECT 194.770 4.000 196.230 4.280 ;
    RECT 197.070 4.000 198.070 4.280 ;
    RECT 198.910 4.000 199.910 4.280 ;
    RECT 200.750 4.000 201.750 4.280 ;
    RECT 202.590 4.000 203.590 4.280 ;
    RECT 204.430 4.000 205.430 4.280 ;
    RECT 206.270 4.000 207.730 4.280 ;
    RECT 208.570 4.000 209.570 4.280 ;
    RECT 210.410 4.000 211.410 4.280 ;
    RECT 212.250 4.000 213.250 4.280 ;
    RECT 214.090 4.000 215.090 4.280 ;
    RECT 215.930 4.000 216.930 4.280 ;
    RECT 217.770 4.000 219.230 4.280 ;
    RECT 220.070 4.000 221.070 4.280 ;
    RECT 221.910 4.000 222.910 4.280 ;
    RECT 223.750 4.000 224.750 4.280 ;
    RECT 225.590 4.000 226.590 4.280 ;
    RECT 227.430 4.000 228.430 4.280 ;
    RECT 229.270 4.000 230.730 4.280 ;
    RECT 231.570 4.000 232.570 4.280 ;
    RECT 233.410 4.000 234.410 4.280 ;
    RECT 235.250 4.000 236.250 4.280 ;
    RECT 237.090 4.000 238.090 4.280 ;
    RECT 238.930 4.000 239.930 4.280 ;
    RECT 240.770 4.000 242.230 4.280 ;
    RECT 243.070 4.000 244.070 4.280 ;
    RECT 244.910 4.000 245.910 4.280 ;
    RECT 246.750 4.000 247.750 4.280 ;
    RECT 248.590 4.000 249.590 4.280 ;
    RECT 250.430 4.000 251.430 4.280 ;
    RECT 252.270 4.000 253.730 4.280 ;
    RECT 254.570 4.000 255.570 4.280 ;
    RECT 256.410 4.000 257.410 4.280 ;
    RECT 258.250 4.000 259.250 4.280 ;
    RECT 260.090 4.000 261.090 4.280 ;
    RECT 261.930 4.000 262.930 4.280 ;
    RECT 263.770 4.000 265.230 4.280 ;
    RECT 266.070 4.000 267.070 4.280 ;
    RECT 267.910 4.000 268.910 4.280 ;
    RECT 269.750 4.000 270.750 4.280 ;
    RECT 271.590 4.000 272.590 4.280 ;
    RECT 273.430 4.000 274.430 4.280 ;
    RECT 275.270 4.000 276.730 4.280 ;
    RECT 277.570 4.000 278.570 4.280 ;
    RECT 279.410 4.000 280.410 4.280 ;
    RECT 281.250 4.000 282.250 4.280 ;
    RECT 283.090 4.000 284.090 4.280 ;
    RECT 284.930 4.000 285.930 4.280 ;
    RECT 286.770 4.000 288.230 4.280 ;
    RECT 289.070 4.000 290.070 4.280 ;
    RECT 290.910 4.000 291.910 4.280 ;
    RECT 292.750 4.000 293.750 4.280 ;
    RECT 294.590 4.000 295.590 4.280 ;
    RECT 296.430 4.000 297.430 4.280 ;
    RECT 298.270 4.000 299.730 4.280 ;
    RECT 300.570 4.000 301.570 4.280 ;
    RECT 302.410 4.000 303.410 4.280 ;
    RECT 304.250 4.000 305.250 4.280 ;
    RECT 306.090 4.000 307.090 4.280 ;
    RECT 307.930 4.000 308.930 4.280 ;
    RECT 309.770 4.000 311.230 4.280 ;
    RECT 312.070 4.000 313.070 4.280 ;
    RECT 313.910 4.000 314.910 4.280 ;
    RECT 315.750 4.000 316.750 4.280 ;
    RECT 317.590 4.000 318.590 4.280 ;
    RECT 319.430 4.000 320.430 4.280 ;
    RECT 321.270 4.000 322.730 4.280 ;
    RECT 323.570 4.000 324.570 4.280 ;
    RECT 325.410 4.000 326.410 4.280 ;
    RECT 327.250 4.000 328.250 4.280 ;
    RECT 329.090 4.000 330.090 4.280 ;
    RECT 330.930 4.000 331.930 4.280 ;
    RECT 332.770 4.000 334.230 4.280 ;
    RECT 335.070 4.000 336.070 4.280 ;
    RECT 336.910 4.000 337.910 4.280 ;
    RECT 338.750 4.000 339.750 4.280 ;
    RECT 340.590 4.000 341.590 4.280 ;
    RECT 342.430 4.000 343.430 4.280 ;
    RECT 344.270 4.000 345.730 4.280 ;
    RECT 346.570 4.000 347.570 4.280 ;
    RECT 348.410 4.000 349.410 4.280 ;
    RECT 350.250 4.000 351.250 4.280 ;
    RECT 352.090 4.000 353.090 4.280 ;
    RECT 353.930 4.000 354.930 4.280 ;
    RECT 355.770 4.000 357.230 4.280 ;
    RECT 358.070 4.000 359.070 4.280 ;
    RECT 359.910 4.000 360.910 4.280 ;
    RECT 361.750 4.000 362.750 4.280 ;
    RECT 363.590 4.000 364.590 4.280 ;
    RECT 365.430 4.000 366.430 4.280 ;
    RECT 367.270 4.000 368.730 4.280 ;
    RECT 369.570 4.000 370.570 4.280 ;
    RECT 371.410 4.000 372.410 4.280 ;
    RECT 373.250 4.000 374.250 4.280 ;
    RECT 375.090 4.000 376.090 4.280 ;
    RECT 376.930 4.000 377.930 4.280 ;
    RECT 378.770 4.000 380.230 4.280 ;
    RECT 381.070 4.000 382.070 4.280 ;
    RECT 382.910 4.000 383.910 4.280 ;
    RECT 384.750 4.000 385.750 4.280 ;
    RECT 386.590 4.000 387.590 4.280 ;
    RECT 388.430 4.000 389.430 4.280 ;
    RECT 390.270 4.000 391.730 4.280 ;
    RECT 392.570 4.000 393.570 4.280 ;
    RECT 394.410 4.000 395.410 4.280 ;
    RECT 396.250 4.000 397.250 4.280 ;
    RECT 398.090 4.000 399.090 4.280 ;
    RECT 399.930 4.000 400.930 4.280 ;
    RECT 401.770 4.000 403.230 4.280 ;
    RECT 404.070 4.000 405.070 4.280 ;
    RECT 405.910 4.000 406.910 4.280 ;
    RECT 407.750 4.000 408.750 4.280 ;
    RECT 409.590 4.000 410.590 4.280 ;
    RECT 411.430 4.000 412.430 4.280 ;
    RECT 413.270 4.000 414.730 4.280 ;
    RECT 415.570 4.000 416.570 4.280 ;
    RECT 417.410 4.000 418.410 4.280 ;
    RECT 419.250 4.000 420.250 4.280 ;
    RECT 421.090 4.000 422.090 4.280 ;
    RECT 422.930 4.000 423.930 4.280 ;
    RECT 424.770 4.000 426.230 4.280 ;
    RECT 427.070 4.000 428.070 4.280 ;
    RECT 428.910 4.000 429.910 4.280 ;
    RECT 430.750 4.000 431.750 4.280 ;
    RECT 432.590 4.000 433.590 4.280 ;
    RECT 434.430 4.000 435.430 4.280 ;
    RECT 436.270 4.000 437.730 4.280 ;
    RECT 438.570 4.000 439.570 4.280 ;
    RECT 440.410 4.000 441.410 4.280 ;
    RECT 442.250 4.000 443.250 4.280 ;
    RECT 444.090 4.000 445.090 4.280 ;
    RECT 445.930 4.000 446.930 4.280 ;
    RECT 447.770 4.000 449.230 4.280 ;
    RECT 450.070 4.000 451.070 4.280 ;
    RECT 451.910 4.000 452.910 4.280 ;
    RECT 453.750 4.000 454.750 4.280 ;
    RECT 455.590 4.000 456.590 4.280 ;
    RECT 457.430 4.000 458.430 4.280 ;
    RECT 459.270 4.000 460.730 4.280 ;
    RECT 461.570 4.000 462.570 4.280 ;
    RECT 463.410 4.000 464.410 4.280 ;
    RECT 465.250 4.000 466.250 4.280 ;
    RECT 467.090 4.000 468.090 4.280 ;
    RECT 468.930 4.000 469.930 4.280 ;
    RECT 470.770 4.000 472.230 4.280 ;
    RECT 473.070 4.000 474.070 4.280 ;
    RECT 474.910 4.000 475.910 4.280 ;
    RECT 476.750 4.000 477.750 4.280 ;
    RECT 478.590 4.000 479.590 4.280 ;
    RECT 480.430 4.000 481.430 4.280 ;
    RECT 482.270 4.000 483.730 4.280 ;
    RECT 484.570 4.000 485.570 4.280 ;
    RECT 486.410 4.000 487.410 4.280 ;
    RECT 488.250 4.000 489.250 4.280 ;
    RECT 490.090 4.000 491.090 4.280 ;
    RECT 491.930 4.000 492.930 4.280 ;
    RECT 493.770 4.000 495.230 4.280 ;
    RECT 496.070 4.000 497.070 4.280 ;
    RECT 497.910 4.000 498.910 4.280 ;
    RECT 499.750 4.000 500.750 4.280 ;
    RECT 501.590 4.000 502.590 4.280 ;
    RECT 503.430 4.000 504.430 4.280 ;
    RECT 505.270 4.000 506.730 4.280 ;
    RECT 507.570 4.000 508.570 4.280 ;
    RECT 509.410 4.000 510.410 4.280 ;
    RECT 511.250 4.000 512.250 4.280 ;
    RECT 513.090 4.000 514.090 4.280 ;
    RECT 514.930 4.000 515.930 4.280 ;
    RECT 516.770 4.000 518.230 4.280 ;
    RECT 519.070 4.000 520.070 4.280 ;
    RECT 520.910 4.000 521.910 4.280 ;
    RECT 522.750 4.000 523.750 4.280 ;
    RECT 524.590 4.000 525.590 4.280 ;
    RECT 526.430 4.000 527.430 4.280 ;
    RECT 528.270 4.000 529.730 4.280 ;
    RECT 530.570 4.000 531.570 4.280 ;
    RECT 532.410 4.000 533.410 4.280 ;
    RECT 534.250 4.000 535.250 4.280 ;
    RECT 536.090 4.000 537.090 4.280 ;
    RECT 537.930 4.000 538.930 4.280 ;
    RECT 539.770 4.000 541.230 4.280 ;
    RECT 542.070 4.000 543.070 4.280 ;
    RECT 543.910 4.000 544.910 4.280 ;
    RECT 545.750 4.000 546.750 4.280 ;
    RECT 547.590 4.000 548.590 4.280 ;
    RECT 549.430 4.000 550.430 4.280 ;
    RECT 551.270 4.000 552.730 4.280 ;
    RECT 553.570 4.000 554.570 4.280 ;
    RECT 555.410 4.000 556.410 4.280 ;
    RECT 557.250 4.000 558.250 4.280 ;
    RECT 559.090 4.000 560.090 4.280 ;
    RECT 560.930 4.000 561.930 4.280 ;
    RECT 562.770 4.000 564.230 4.280 ;
    RECT 565.070 4.000 566.070 4.280 ;
    RECT 566.910 4.000 567.910 4.280 ;
    RECT 568.750 4.000 569.750 4.280 ;
    RECT 570.590 4.000 571.590 4.280 ;
    RECT 572.430 4.000 573.430 4.280 ;
    RECT 574.270 4.000 575.730 4.280 ;
    RECT 576.570 4.000 577.570 4.280 ;
    RECT 578.410 4.000 579.410 4.280 ;
    RECT 580.250 4.000 581.250 4.280 ;
    RECT 582.090 4.000 583.090 4.280 ;
    RECT 583.930 4.000 584.930 4.280 ;
    RECT 585.770 4.000 587.230 4.280 ;
    RECT 588.070 4.000 589.070 4.280 ;
    RECT 589.910 4.000 590.910 4.280 ;
    RECT 591.750 4.000 592.750 4.280 ;
    RECT 593.590 4.000 594.590 4.280 ;
    RECT 595.430 4.000 596.430 4.280 ;
    RECT 597.270 4.000 598.730 4.280 ;
    RECT 599.570 4.000 600.570 4.280 ;
    RECT 601.410 4.000 602.410 4.280 ;
    RECT 603.250 4.000 604.250 4.280 ;
    RECT 605.090 4.000 606.090 4.280 ;
    RECT 606.930 4.000 607.930 4.280 ;
    RECT 608.770 4.000 610.230 4.280 ;
    RECT 611.070 4.000 612.070 4.280 ;
    RECT 612.910 4.000 613.910 4.280 ;
    RECT 614.750 4.000 615.750 4.280 ;
    RECT 616.590 4.000 617.590 4.280 ;
    RECT 618.430 4.000 619.430 4.280 ;
    RECT 620.270 4.000 621.730 4.280 ;
    RECT 622.570 4.000 623.570 4.280 ;
    RECT 624.410 4.000 625.410 4.280 ;
    RECT 626.250 4.000 627.250 4.280 ;
    RECT 628.090 4.000 629.090 4.280 ;
    RECT 629.930 4.000 630.930 4.280 ;
    RECT 631.770 4.000 633.230 4.280 ;
    RECT 634.070 4.000 635.070 4.280 ;
    RECT 635.910 4.000 636.910 4.280 ;
    RECT 637.750 4.000 638.750 4.280 ;
    RECT 639.590 4.000 640.590 4.280 ;
    RECT 641.430 4.000 642.430 4.280 ;
    RECT 643.270 4.000 644.730 4.280 ;
    RECT 645.570 4.000 646.570 4.280 ;
    RECT 647.410 4.000 648.410 4.280 ;
    RECT 649.250 4.000 650.250 4.280 ;
    RECT 651.090 4.000 652.090 4.280 ;
    RECT 652.930 4.000 653.930 4.280 ;
    RECT 654.770 4.000 656.230 4.280 ;
    RECT 657.070 4.000 658.070 4.280 ;
    RECT 658.910 4.000 659.910 4.280 ;
    RECT 660.750 4.000 661.750 4.280 ;
    RECT 662.590 4.000 663.590 4.280 ;
    RECT 664.430 4.000 665.430 4.280 ;
    RECT 666.270 4.000 667.730 4.280 ;
    RECT 668.570 4.000 669.570 4.280 ;
    RECT 670.410 4.000 671.410 4.280 ;
    RECT 672.250 4.000 673.250 4.280 ;
    RECT 674.090 4.000 675.090 4.280 ;
    RECT 675.930 4.000 676.930 4.280 ;
    RECT 677.770 4.000 679.230 4.280 ;
    RECT 680.070 4.000 681.070 4.280 ;
    RECT 681.910 4.000 682.910 4.280 ;
    RECT 683.750 4.000 684.750 4.280 ;
    RECT 685.590 4.000 686.590 4.280 ;
    RECT 687.430 4.000 688.430 4.280 ;
    RECT 689.270 4.000 690.730 4.280 ;
    RECT 691.570 4.000 692.570 4.280 ;
    RECT 693.410 4.000 694.410 4.280 ;
    RECT 695.250 4.000 696.250 4.280 ;
    RECT 697.090 4.000 698.090 4.280 ;
    RECT 698.930 4.000 699.930 4.280 ;
    RECT 700.770 4.000 702.230 4.280 ;
    RECT 703.070 4.000 704.070 4.280 ;
    RECT 704.910 4.000 705.910 4.280 ;
    RECT 706.750 4.000 707.750 4.280 ;
    RECT 708.590 4.000 709.590 4.280 ;
    RECT 710.430 4.000 711.430 4.280 ;
    RECT 712.270 4.000 713.730 4.280 ;
    RECT 714.570 4.000 715.570 4.280 ;
    RECT 716.410 4.000 717.410 4.280 ;
    RECT 718.250 4.000 719.250 4.280 ;
    RECT 720.090 4.000 721.090 4.280 ;
    RECT 721.930 4.000 722.930 4.280 ;
    RECT 723.770 4.000 725.230 4.280 ;
    RECT 726.070 4.000 727.070 4.280 ;
    RECT 727.910 4.000 728.910 4.280 ;
    RECT 729.750 4.000 730.750 4.280 ;
    RECT 731.590 4.000 732.590 4.280 ;
    LAYER met3 ;
    RECT 4.000 168.320 732.000 212.325 ;
    RECT 4.400 166.920 732.000 168.320 ;
    RECT 4.000 112.560 732.000 166.920 ;
    RECT 4.000 111.160 731.600 112.560 ;
    RECT 4.000 56.800 732.000 111.160 ;
    RECT 4.400 55.400 732.000 56.800 ;
    RECT 4.000 4.255 732.000 55.400 ;
    LAYER met4 ;
    RECT 174.640 10.640 713.840 212.400 ;
  END
END rescue_top
END LIBRARY
