magic
tech sky130A
magscale 1 2
timestamp 1607274956
<< metal1 >>
rect 1064 52846 9556 52868
rect 1064 52794 3606 52846
rect 3658 52794 3670 52846
rect 3722 52794 3734 52846
rect 3786 52794 3798 52846
rect 3850 52794 8934 52846
rect 8986 52794 8998 52846
rect 9050 52794 9062 52846
rect 9114 52794 9126 52846
rect 9178 52794 9556 52846
rect 1064 52772 9556 52794
rect 1350 52513 1402 52519
rect 1350 52455 1402 52461
rect 1446 52276 1452 52328
rect 1504 52276 1510 52328
rect 2022 52291 2074 52297
rect 1302 52254 1354 52260
rect 2022 52233 2074 52239
rect 1302 52196 1354 52202
rect 1104 52128 1110 52180
rect 1162 52128 1168 52180
rect 1872 52128 1878 52180
rect 1930 52128 1936 52180
rect 1296 52017 1302 52069
rect 1354 52057 1360 52069
rect 1872 52057 1878 52069
rect 1354 52029 1878 52057
rect 1354 52017 1360 52029
rect 1872 52017 1878 52029
rect 1930 52017 1936 52069
rect 1064 51514 9556 51536
rect 1064 51462 6270 51514
rect 6322 51462 6334 51514
rect 6386 51462 6398 51514
rect 6450 51462 6462 51514
rect 6514 51462 9556 51514
rect 1064 51440 9556 51462
rect 1926 50848 1978 50854
rect 1104 50796 1110 50848
rect 1162 50796 1168 50848
rect 1302 50774 1354 50780
rect 1392 50759 1398 50811
rect 1450 50799 1456 50811
rect 1450 50771 1822 50799
rect 1926 50790 1978 50796
rect 1450 50759 1456 50771
rect 1302 50716 1354 50722
rect 1446 50648 1452 50700
rect 1504 50648 1510 50700
rect 1350 50626 1402 50632
rect 1794 50589 1822 50771
rect 2022 50663 2074 50669
rect 2022 50605 2074 50611
rect 1350 50568 1402 50574
rect 1776 50537 1782 50589
rect 1834 50537 1840 50589
rect 1064 50182 9556 50204
rect 1064 50130 3606 50182
rect 3658 50130 3670 50182
rect 3722 50130 3734 50182
rect 3786 50130 3798 50182
rect 3850 50130 8934 50182
rect 8986 50130 8998 50182
rect 9050 50130 9062 50182
rect 9114 50130 9126 50182
rect 9178 50130 9556 50182
rect 1064 50108 9556 50130
rect 2022 49849 2074 49855
rect 2022 49791 2074 49797
rect 1872 49464 1878 49516
rect 1930 49464 1936 49516
rect 1064 48850 9556 48872
rect 1064 48798 6270 48850
rect 6322 48798 6334 48850
rect 6386 48798 6398 48850
rect 6450 48798 6462 48850
rect 6514 48798 9556 48850
rect 1064 48776 9556 48798
rect 1872 48243 1878 48295
rect 1930 48283 1936 48295
rect 2496 48283 2502 48295
rect 1930 48255 2502 48283
rect 1930 48243 1936 48255
rect 2496 48243 2502 48255
rect 2554 48243 2560 48295
rect 1104 48132 1110 48184
rect 1162 48132 1168 48184
rect 1302 48110 1354 48116
rect 1776 48095 1782 48147
rect 1834 48095 1840 48147
rect 1872 48132 1878 48184
rect 1930 48132 1936 48184
rect 2352 48132 2358 48184
rect 2410 48132 2416 48184
rect 1302 48052 1354 48058
rect 1446 47984 1452 48036
rect 1504 47984 1510 48036
rect 1488 47873 1494 47925
rect 1546 47913 1552 47925
rect 1794 47913 1822 48095
rect 2502 48073 2554 48079
rect 2502 48015 2554 48021
rect 2022 47999 2074 48005
rect 2022 47941 2074 47947
rect 1546 47885 1822 47913
rect 1546 47873 1552 47885
rect 1350 47851 1402 47857
rect 1350 47793 1402 47799
rect 1064 47518 9556 47540
rect 1064 47466 3606 47518
rect 3658 47466 3670 47518
rect 3722 47466 3734 47518
rect 3786 47466 3798 47518
rect 3850 47466 8934 47518
rect 8986 47466 8998 47518
rect 9050 47466 9062 47518
rect 9114 47466 9126 47518
rect 9178 47466 9556 47518
rect 1064 47444 9556 47466
rect 2502 47185 2554 47191
rect 2502 47127 2554 47133
rect 2022 46963 2074 46969
rect 2022 46905 2074 46911
rect 1200 46763 1206 46815
rect 1258 46803 1264 46815
rect 1776 46803 1782 46815
rect 1258 46775 1782 46803
rect 1258 46763 1264 46775
rect 1776 46763 1782 46775
rect 1834 46763 1840 46815
rect 1872 46800 1878 46852
rect 1930 46800 1936 46852
rect 2352 46800 2358 46852
rect 2410 46800 2416 46852
rect 1064 46186 9556 46208
rect 1064 46134 6270 46186
rect 6322 46134 6334 46186
rect 6386 46134 6398 46186
rect 6450 46134 6462 46186
rect 6514 46134 9556 46186
rect 1064 46112 9556 46134
rect 1926 45520 1978 45526
rect 1104 45468 1110 45520
rect 1162 45468 1168 45520
rect 1302 45446 1354 45452
rect 1392 45431 1398 45483
rect 1450 45471 1456 45483
rect 1450 45443 1822 45471
rect 1926 45462 1978 45468
rect 2406 45520 2458 45526
rect 2406 45462 2458 45468
rect 2838 45520 2890 45526
rect 2838 45462 2890 45468
rect 3318 45520 3370 45526
rect 3318 45462 3370 45468
rect 1450 45431 1456 45443
rect 1302 45388 1354 45394
rect 1446 45320 1452 45372
rect 1504 45320 1510 45372
rect 1350 45298 1402 45304
rect 1794 45261 1822 45443
rect 3462 45409 3514 45415
rect 3462 45351 3514 45357
rect 2022 45335 2074 45341
rect 2022 45277 2074 45283
rect 2502 45335 2554 45341
rect 2502 45277 2554 45283
rect 2982 45335 3034 45341
rect 2982 45277 3034 45283
rect 1350 45240 1402 45246
rect 1776 45209 1782 45261
rect 1834 45209 1840 45261
rect 1064 44854 9556 44876
rect 1064 44802 3606 44854
rect 3658 44802 3670 44854
rect 3722 44802 3734 44854
rect 3786 44802 3798 44854
rect 3850 44802 8934 44854
rect 8986 44802 8998 44854
rect 9050 44802 9062 44854
rect 9114 44802 9126 44854
rect 9178 44802 9556 44854
rect 1064 44780 9556 44802
rect 3462 44521 3514 44527
rect 3462 44463 3514 44469
rect 2982 44447 3034 44453
rect 2982 44389 3034 44395
rect 2022 44299 2074 44305
rect 2022 44241 2074 44247
rect 2502 44299 2554 44305
rect 2502 44241 2554 44247
rect 2838 44188 2890 44194
rect 1872 44136 1878 44188
rect 1930 44136 1936 44188
rect 2352 44136 2358 44188
rect 2410 44136 2416 44188
rect 2838 44130 2890 44136
rect 3318 44188 3370 44194
rect 3318 44130 3370 44136
rect 1064 43522 9556 43544
rect 1064 43470 6270 43522
rect 6322 43470 6334 43522
rect 6386 43470 6398 43522
rect 6450 43470 6462 43522
rect 6514 43470 9556 43522
rect 1064 43448 9556 43470
rect 4752 42915 4758 42967
rect 4810 42955 4816 42967
rect 5376 42955 5382 42967
rect 4810 42927 5382 42955
rect 4810 42915 4816 42927
rect 5376 42915 5382 42927
rect 5434 42915 5440 42967
rect 1926 42856 1978 42862
rect 1104 42804 1110 42856
rect 1162 42804 1168 42856
rect 1302 42782 1354 42788
rect 1776 42767 1782 42819
rect 1834 42767 1840 42819
rect 1926 42798 1978 42804
rect 2406 42856 2458 42862
rect 2880 42804 2886 42856
rect 2938 42804 2944 42856
rect 3360 42804 3366 42856
rect 3418 42804 3424 42856
rect 3843 42804 3849 42856
rect 3901 42804 3907 42856
rect 4327 42804 4333 42856
rect 4385 42804 4391 42856
rect 4752 42804 4758 42856
rect 4810 42804 4816 42856
rect 5295 42804 5301 42856
rect 5353 42804 5359 42856
rect 2406 42798 2458 42804
rect 1302 42724 1354 42730
rect 1446 42656 1452 42708
rect 1504 42656 1510 42708
rect 1488 42545 1494 42597
rect 1546 42585 1552 42597
rect 1794 42585 1822 42767
rect 5382 42745 5434 42751
rect 5382 42687 5434 42693
rect 2022 42671 2074 42677
rect 2022 42613 2074 42619
rect 2502 42671 2554 42677
rect 2502 42613 2554 42619
rect 2982 42671 3034 42677
rect 2982 42613 3034 42619
rect 3462 42671 3514 42677
rect 3462 42613 3514 42619
rect 3942 42671 3994 42677
rect 3942 42613 3994 42619
rect 4422 42671 4474 42677
rect 4422 42613 4474 42619
rect 4902 42671 4954 42677
rect 4902 42613 4954 42619
rect 1546 42557 1822 42585
rect 1546 42545 1552 42557
rect 1350 42523 1402 42529
rect 1350 42465 1402 42471
rect 1200 42323 1206 42375
rect 1258 42363 1264 42375
rect 1776 42363 1782 42375
rect 1258 42335 1782 42363
rect 1258 42323 1264 42335
rect 1776 42323 1782 42335
rect 1834 42323 1840 42375
rect 1064 42190 9556 42212
rect 1064 42138 3606 42190
rect 3658 42138 3670 42190
rect 3722 42138 3734 42190
rect 3786 42138 3798 42190
rect 3850 42138 8934 42190
rect 8986 42138 8998 42190
rect 9050 42138 9062 42190
rect 9114 42138 9126 42190
rect 9178 42138 9556 42190
rect 1064 42116 9556 42138
rect 5382 41857 5434 41863
rect 5382 41799 5434 41805
rect 2022 41635 2074 41641
rect 2022 41577 2074 41583
rect 2502 41635 2554 41641
rect 2502 41577 2554 41583
rect 2982 41635 3034 41641
rect 2982 41577 3034 41583
rect 3462 41635 3514 41641
rect 3462 41577 3514 41583
rect 3942 41635 3994 41641
rect 3942 41577 3994 41583
rect 4422 41635 4474 41641
rect 4422 41577 4474 41583
rect 4902 41635 4954 41641
rect 4902 41577 4954 41583
rect 2838 41524 2890 41530
rect 1872 41472 1878 41524
rect 1930 41472 1936 41524
rect 2352 41472 2358 41524
rect 2410 41472 2416 41524
rect 2838 41466 2890 41472
rect 3318 41524 3370 41530
rect 3318 41466 3370 41472
rect 3798 41524 3850 41530
rect 3798 41466 3850 41472
rect 4278 41524 4330 41530
rect 4752 41472 4758 41524
rect 4810 41472 4816 41524
rect 5278 41472 5284 41524
rect 5336 41472 5342 41524
rect 4278 41466 4330 41472
rect 1064 40858 9556 40880
rect 1064 40806 6270 40858
rect 6322 40806 6334 40858
rect 6386 40806 6398 40858
rect 6450 40806 6462 40858
rect 6514 40806 9556 40858
rect 1064 40784 9556 40806
rect 5280 40325 5286 40377
rect 5338 40365 5344 40377
rect 5904 40365 5910 40377
rect 5338 40337 5910 40365
rect 5338 40325 5344 40337
rect 5904 40325 5910 40337
rect 5962 40325 5968 40377
rect 6263 40325 6269 40377
rect 6321 40365 6327 40377
rect 6864 40365 6870 40377
rect 6321 40337 6870 40365
rect 6321 40325 6327 40337
rect 6864 40325 6870 40337
rect 6922 40325 6928 40377
rect 4752 40251 4758 40303
rect 4810 40291 4816 40303
rect 5376 40291 5382 40303
rect 4810 40263 5382 40291
rect 4810 40251 4816 40263
rect 5376 40251 5382 40263
rect 5434 40251 5440 40303
rect 5779 40251 5785 40303
rect 5837 40291 5843 40303
rect 6384 40291 6390 40303
rect 5837 40263 6390 40291
rect 5837 40251 5843 40263
rect 6384 40251 6390 40263
rect 6442 40251 6448 40303
rect 6768 40251 6774 40303
rect 6826 40291 6832 40303
rect 7344 40291 7350 40303
rect 6826 40263 7350 40291
rect 6826 40251 6832 40263
rect 7344 40251 7350 40263
rect 7402 40251 7408 40303
rect 8688 40251 8694 40303
rect 8746 40291 8752 40303
rect 9264 40291 9270 40303
rect 8746 40263 9270 40291
rect 8746 40251 8752 40263
rect 9264 40251 9270 40263
rect 9322 40251 9328 40303
rect 1926 40192 1978 40198
rect 1104 40140 1110 40192
rect 1162 40140 1168 40192
rect 1926 40134 1978 40140
rect 2406 40192 2458 40198
rect 6774 40192 6826 40198
rect 2880 40140 2886 40192
rect 2938 40140 2944 40192
rect 3360 40140 3366 40192
rect 3418 40140 3424 40192
rect 3843 40140 3849 40192
rect 3901 40140 3907 40192
rect 4327 40140 4333 40192
rect 4385 40140 4391 40192
rect 4752 40140 4758 40192
rect 4810 40140 4816 40192
rect 5280 40140 5286 40192
rect 5338 40140 5344 40192
rect 5779 40140 5785 40192
rect 5837 40140 5843 40192
rect 6263 40140 6269 40192
rect 6321 40140 6327 40192
rect 2406 40134 2458 40140
rect 6774 40134 6826 40140
rect 7254 40192 7306 40198
rect 7254 40134 7306 40140
rect 7734 40192 7786 40198
rect 7734 40134 7786 40140
rect 8214 40192 8266 40198
rect 8688 40140 8694 40192
rect 8746 40140 8752 40192
rect 9168 40140 9174 40192
rect 9226 40140 9232 40192
rect 8214 40134 8266 40140
rect 5910 40118 5962 40124
rect 1268 40066 1274 40118
rect 1326 40066 1332 40118
rect 2502 40081 2554 40087
rect 1446 39992 1452 40044
rect 1504 39992 1510 40044
rect 2502 40023 2554 40029
rect 2982 40081 3034 40087
rect 2982 40023 3034 40029
rect 3462 40081 3514 40087
rect 3462 40023 3514 40029
rect 3942 40081 3994 40087
rect 3942 40023 3994 40029
rect 4422 40081 4474 40087
rect 4422 40023 4474 40029
rect 4902 40081 4954 40087
rect 4902 40023 4954 40029
rect 5382 40081 5434 40087
rect 5910 40060 5962 40066
rect 6390 40118 6442 40124
rect 6390 40060 6442 40066
rect 6870 40118 6922 40124
rect 6870 40060 6922 40066
rect 7350 40081 7402 40087
rect 5382 40023 5434 40029
rect 7350 40023 7402 40029
rect 8310 40081 8362 40087
rect 8310 40023 8362 40029
rect 8790 40081 8842 40087
rect 8790 40023 8842 40029
rect 9270 40081 9322 40087
rect 9270 40023 9322 40029
rect 2022 40007 2074 40013
rect 1350 39970 1402 39976
rect 2022 39949 2074 39955
rect 1350 39912 1402 39918
rect 7830 39933 7882 39939
rect 7830 39875 7882 39881
rect 1064 39526 9556 39548
rect 1064 39474 3606 39526
rect 3658 39474 3670 39526
rect 3722 39474 3734 39526
rect 3786 39474 3798 39526
rect 3850 39474 8934 39526
rect 8986 39474 8998 39526
rect 9050 39474 9062 39526
rect 9114 39474 9126 39526
rect 9178 39474 9556 39526
rect 1064 39452 9556 39474
rect 9270 39193 9322 39199
rect 9270 39135 9322 39141
rect 2022 38971 2074 38977
rect 2022 38913 2074 38919
rect 2502 38971 2554 38977
rect 2502 38913 2554 38919
rect 2982 38971 3034 38977
rect 2982 38913 3034 38919
rect 3462 38971 3514 38977
rect 3462 38913 3514 38919
rect 3942 38971 3994 38977
rect 3942 38913 3994 38919
rect 4422 38971 4474 38977
rect 4422 38913 4474 38919
rect 4902 38971 4954 38977
rect 4902 38913 4954 38919
rect 5382 38971 5434 38977
rect 7350 38971 7402 38977
rect 5382 38913 5434 38919
rect 5910 38934 5962 38940
rect 5910 38876 5962 38882
rect 6390 38934 6442 38940
rect 6390 38876 6442 38882
rect 6870 38934 6922 38940
rect 7350 38913 7402 38919
rect 7830 38971 7882 38977
rect 7830 38913 7882 38919
rect 8310 38971 8362 38977
rect 8310 38913 8362 38919
rect 8790 38971 8842 38977
rect 8790 38913 8842 38919
rect 6870 38876 6922 38882
rect 2838 38860 2890 38866
rect 1872 38808 1878 38860
rect 1930 38808 1936 38860
rect 2352 38808 2358 38860
rect 2410 38808 2416 38860
rect 2838 38802 2890 38808
rect 3318 38860 3370 38866
rect 3318 38802 3370 38808
rect 3798 38860 3850 38866
rect 3798 38802 3850 38808
rect 4278 38860 4330 38866
rect 7254 38860 7306 38866
rect 4752 38808 4758 38860
rect 4810 38808 4816 38860
rect 5278 38808 5284 38860
rect 5336 38808 5342 38860
rect 5760 38808 5766 38860
rect 5818 38808 5824 38860
rect 6240 38808 6246 38860
rect 6298 38808 6304 38860
rect 6720 38808 6726 38860
rect 6778 38808 6784 38860
rect 4278 38802 4330 38808
rect 7254 38802 7306 38808
rect 7734 38860 7786 38866
rect 7734 38802 7786 38808
rect 8214 38860 8266 38866
rect 8688 38808 8694 38860
rect 8746 38808 8752 38860
rect 9168 38808 9174 38860
rect 9226 38808 9232 38860
rect 8214 38802 8266 38808
rect 1200 38697 1206 38749
rect 1258 38737 1264 38749
rect 1872 38737 1878 38749
rect 1258 38709 1878 38737
rect 1258 38697 1264 38709
rect 1872 38697 1878 38709
rect 1930 38697 1936 38749
rect 1064 38194 9556 38216
rect 1064 38142 6270 38194
rect 6322 38142 6334 38194
rect 6386 38142 6398 38194
rect 6450 38142 6462 38194
rect 6514 38142 9556 38194
rect 1064 38120 9556 38142
rect 5779 37661 5785 37713
rect 5837 37701 5843 37713
rect 5837 37673 6046 37701
rect 5837 37661 5843 37673
rect 5295 37587 5301 37639
rect 5353 37627 5359 37639
rect 5904 37627 5910 37639
rect 5353 37599 5910 37627
rect 5353 37587 5359 37599
rect 5904 37587 5910 37599
rect 5962 37587 5968 37639
rect 6018 37627 6046 37673
rect 6263 37661 6269 37713
rect 6321 37701 6327 37713
rect 6864 37701 6870 37713
rect 6321 37673 6870 37701
rect 6321 37661 6327 37673
rect 6864 37661 6870 37673
rect 6922 37661 6928 37713
rect 6384 37627 6390 37639
rect 6018 37599 6390 37627
rect 6384 37587 6390 37599
rect 6442 37587 6448 37639
rect 6768 37587 6774 37639
rect 6826 37627 6832 37639
rect 7344 37627 7350 37639
rect 6826 37599 7350 37627
rect 6826 37587 6832 37599
rect 7344 37587 7350 37599
rect 7402 37587 7408 37639
rect 8688 37587 8694 37639
rect 8746 37627 8752 37639
rect 9264 37627 9270 37639
rect 8746 37599 9270 37627
rect 8746 37587 8752 37599
rect 9264 37587 9270 37599
rect 9322 37587 9328 37639
rect 1926 37528 1978 37534
rect 1104 37476 1110 37528
rect 1162 37476 1168 37528
rect 1302 37454 1354 37460
rect 1392 37439 1398 37491
rect 1450 37479 1456 37491
rect 1450 37451 1822 37479
rect 1926 37470 1978 37476
rect 2406 37528 2458 37534
rect 6774 37528 6826 37534
rect 2880 37476 2886 37528
rect 2938 37476 2944 37528
rect 3360 37476 3366 37528
rect 3418 37476 3424 37528
rect 3843 37476 3849 37528
rect 3901 37476 3907 37528
rect 4327 37476 4333 37528
rect 4385 37476 4391 37528
rect 4811 37476 4817 37528
rect 4869 37476 4875 37528
rect 5295 37476 5301 37528
rect 5353 37476 5359 37528
rect 5779 37476 5785 37528
rect 5837 37476 5843 37528
rect 6263 37476 6269 37528
rect 6321 37476 6327 37528
rect 2406 37470 2458 37476
rect 6774 37470 6826 37476
rect 7254 37528 7306 37534
rect 7254 37470 7306 37476
rect 7734 37528 7786 37534
rect 7734 37470 7786 37476
rect 8214 37528 8266 37534
rect 8688 37476 8694 37528
rect 8746 37476 8752 37528
rect 9168 37476 9174 37528
rect 9226 37476 9232 37528
rect 8214 37470 8266 37476
rect 1450 37439 1456 37451
rect 1302 37396 1354 37402
rect 1446 37328 1452 37380
rect 1504 37328 1510 37380
rect 1350 37306 1402 37312
rect 1794 37269 1822 37451
rect 5910 37454 5962 37460
rect 2502 37417 2554 37423
rect 2502 37359 2554 37365
rect 2982 37417 3034 37423
rect 2982 37359 3034 37365
rect 3462 37417 3514 37423
rect 3462 37359 3514 37365
rect 3942 37417 3994 37423
rect 3942 37359 3994 37365
rect 4422 37417 4474 37423
rect 4422 37359 4474 37365
rect 4902 37417 4954 37423
rect 4902 37359 4954 37365
rect 5382 37417 5434 37423
rect 5910 37396 5962 37402
rect 6390 37454 6442 37460
rect 6390 37396 6442 37402
rect 6870 37454 6922 37460
rect 6870 37396 6922 37402
rect 7350 37417 7402 37423
rect 5382 37359 5434 37365
rect 7350 37359 7402 37365
rect 8310 37417 8362 37423
rect 8310 37359 8362 37365
rect 8790 37417 8842 37423
rect 8790 37359 8842 37365
rect 9270 37417 9322 37423
rect 9270 37359 9322 37365
rect 2022 37343 2074 37349
rect 2022 37285 2074 37291
rect 7830 37343 7882 37349
rect 7830 37285 7882 37291
rect 1350 37248 1402 37254
rect 1776 37217 1782 37269
rect 1834 37217 1840 37269
rect 1064 36862 9556 36884
rect 1064 36810 3606 36862
rect 3658 36810 3670 36862
rect 3722 36810 3734 36862
rect 3786 36810 3798 36862
rect 3850 36810 8934 36862
rect 8986 36810 8998 36862
rect 9050 36810 9062 36862
rect 9114 36810 9126 36862
rect 9178 36810 9556 36862
rect 1064 36788 9556 36810
rect 9270 36529 9322 36535
rect 9270 36471 9322 36477
rect 2022 36307 2074 36313
rect 2022 36249 2074 36255
rect 2502 36307 2554 36313
rect 2502 36249 2554 36255
rect 2982 36307 3034 36313
rect 2982 36249 3034 36255
rect 3462 36307 3514 36313
rect 3462 36249 3514 36255
rect 3942 36307 3994 36313
rect 3942 36249 3994 36255
rect 4422 36307 4474 36313
rect 4422 36249 4474 36255
rect 4902 36307 4954 36313
rect 4902 36249 4954 36255
rect 5382 36307 5434 36313
rect 7350 36307 7402 36313
rect 5382 36249 5434 36255
rect 5910 36270 5962 36276
rect 5910 36212 5962 36218
rect 6390 36270 6442 36276
rect 6390 36212 6442 36218
rect 6870 36270 6922 36276
rect 7350 36249 7402 36255
rect 7830 36307 7882 36313
rect 7830 36249 7882 36255
rect 8310 36307 8362 36313
rect 8310 36249 8362 36255
rect 8790 36307 8842 36313
rect 8790 36249 8842 36255
rect 6870 36212 6922 36218
rect 1926 36196 1978 36202
rect 2838 36196 2890 36202
rect 2352 36144 2358 36196
rect 2410 36144 2416 36196
rect 1926 36138 1978 36144
rect 2838 36138 2890 36144
rect 3318 36196 3370 36202
rect 3318 36138 3370 36144
rect 3798 36196 3850 36202
rect 3798 36138 3850 36144
rect 4278 36196 4330 36202
rect 8646 36196 8698 36202
rect 4752 36144 4758 36196
rect 4810 36144 4816 36196
rect 5278 36144 5284 36196
rect 5336 36144 5342 36196
rect 5760 36144 5766 36196
rect 5818 36144 5824 36196
rect 6240 36144 6246 36196
rect 6298 36144 6304 36196
rect 6720 36144 6726 36196
rect 6778 36144 6784 36196
rect 7200 36144 7206 36196
rect 7258 36144 7264 36196
rect 7680 36144 7686 36196
rect 7738 36144 7744 36196
rect 8160 36144 8166 36196
rect 8218 36144 8224 36196
rect 4278 36138 4330 36144
rect 8646 36138 8698 36144
rect 9126 36196 9178 36202
rect 9126 36138 9178 36144
rect 1064 35530 9556 35552
rect 1064 35478 6270 35530
rect 6322 35478 6334 35530
rect 6386 35478 6398 35530
rect 6450 35478 6462 35530
rect 6514 35478 9556 35530
rect 1064 35456 9556 35478
rect 5779 34923 5785 34975
rect 5837 34963 5843 34975
rect 5837 34935 6430 34963
rect 5837 34923 5843 34935
rect 6402 34901 6430 34935
rect 2406 34864 2458 34870
rect 1872 34812 1878 34864
rect 1930 34812 1936 34864
rect 2880 34812 2886 34864
rect 2938 34812 2944 34864
rect 3360 34812 3366 34864
rect 3418 34812 3424 34864
rect 3843 34812 3849 34864
rect 3901 34812 3907 34864
rect 4327 34812 4333 34864
rect 4385 34812 4391 34864
rect 4811 34812 4817 34864
rect 4869 34812 4875 34864
rect 5295 34812 5301 34864
rect 5353 34812 5359 34864
rect 5779 34812 5785 34864
rect 5837 34812 5843 34864
rect 6263 34812 6269 34864
rect 6321 34812 6327 34864
rect 6384 34849 6390 34901
rect 6442 34849 6448 34901
rect 6774 34864 6826 34870
rect 2406 34806 2458 34812
rect 6774 34806 6826 34812
rect 7254 34864 7306 34870
rect 7254 34806 7306 34812
rect 7734 34864 7786 34870
rect 7734 34806 7786 34812
rect 8214 34864 8266 34870
rect 8688 34812 8694 34864
rect 8746 34812 8752 34864
rect 9168 34812 9174 34864
rect 9226 34812 9232 34864
rect 8214 34806 8266 34812
rect 6390 34790 6442 34796
rect 2022 34753 2074 34759
rect 6390 34732 6442 34738
rect 9270 34753 9322 34759
rect 2022 34695 2074 34701
rect 9270 34695 9322 34701
rect 2502 34679 2554 34685
rect 2502 34621 2554 34627
rect 2982 34679 3034 34685
rect 2982 34621 3034 34627
rect 3462 34679 3514 34685
rect 3462 34621 3514 34627
rect 3942 34679 3994 34685
rect 3942 34621 3994 34627
rect 4422 34679 4474 34685
rect 4422 34621 4474 34627
rect 4902 34679 4954 34685
rect 4902 34621 4954 34627
rect 5382 34679 5434 34685
rect 5382 34621 5434 34627
rect 7350 34679 7402 34685
rect 7350 34621 7402 34627
rect 7830 34679 7882 34685
rect 7830 34621 7882 34627
rect 8310 34679 8362 34685
rect 8310 34621 8362 34627
rect 8790 34679 8842 34685
rect 8790 34621 8842 34627
rect 5910 34494 5962 34500
rect 5910 34436 5962 34442
rect 6870 34494 6922 34500
rect 6870 34436 6922 34442
rect 6288 34331 6294 34383
rect 6346 34371 6352 34383
rect 6864 34371 6870 34383
rect 6346 34343 6870 34371
rect 6346 34331 6352 34343
rect 6864 34331 6870 34343
rect 6922 34331 6928 34383
rect 1064 34198 9556 34220
rect 1064 34146 3606 34198
rect 3658 34146 3670 34198
rect 3722 34146 3734 34198
rect 3786 34146 3798 34198
rect 3850 34146 8934 34198
rect 8986 34146 8998 34198
rect 9050 34146 9062 34198
rect 9114 34146 9126 34198
rect 9178 34146 9556 34198
rect 1064 34124 9556 34146
rect 6390 33902 6442 33908
rect 6390 33844 6442 33850
rect 9270 33865 9322 33871
rect 9270 33807 9322 33813
rect 2982 33791 3034 33797
rect 2982 33733 3034 33739
rect 3942 33791 3994 33797
rect 3942 33733 3994 33739
rect 5382 33791 5434 33797
rect 5382 33733 5434 33739
rect 2022 33643 2074 33649
rect 2022 33585 2074 33591
rect 2502 33643 2554 33649
rect 2502 33585 2554 33591
rect 3462 33643 3514 33649
rect 3462 33585 3514 33591
rect 4422 33643 4474 33649
rect 4422 33585 4474 33591
rect 4902 33643 4954 33649
rect 7350 33643 7402 33649
rect 4902 33585 4954 33591
rect 5910 33606 5962 33612
rect 5910 33548 5962 33554
rect 6870 33606 6922 33612
rect 7350 33585 7402 33591
rect 7830 33643 7882 33649
rect 7830 33585 7882 33591
rect 8310 33643 8362 33649
rect 8310 33585 8362 33591
rect 8790 33643 8842 33649
rect 8790 33585 8842 33591
rect 6870 33548 6922 33554
rect 2838 33532 2890 33538
rect 1872 33480 1878 33532
rect 1930 33480 1936 33532
rect 2352 33480 2358 33532
rect 2410 33480 2416 33532
rect 2838 33474 2890 33480
rect 3318 33532 3370 33538
rect 3318 33474 3370 33480
rect 3798 33532 3850 33538
rect 3798 33474 3850 33480
rect 4278 33532 4330 33538
rect 6774 33532 6826 33538
rect 7734 33532 7786 33538
rect 4752 33480 4758 33532
rect 4810 33480 4816 33532
rect 5278 33480 5284 33532
rect 5336 33480 5342 33532
rect 5760 33480 5766 33532
rect 5818 33480 5824 33532
rect 6240 33480 6246 33532
rect 6298 33480 6304 33532
rect 7200 33480 7206 33532
rect 7258 33480 7264 33532
rect 4278 33474 4330 33480
rect 6774 33474 6826 33480
rect 7734 33474 7786 33480
rect 8214 33532 8266 33538
rect 8688 33480 8694 33532
rect 8746 33480 8752 33532
rect 9168 33480 9174 33532
rect 9226 33480 9232 33532
rect 8214 33474 8266 33480
rect 1064 32866 9556 32888
rect 1064 32814 6270 32866
rect 6322 32814 6334 32866
rect 6386 32814 6398 32866
rect 6450 32814 6462 32866
rect 6514 32814 9556 32866
rect 1064 32792 9556 32814
rect 5280 32333 5286 32385
rect 5338 32373 5344 32385
rect 5904 32373 5910 32385
rect 5338 32345 5910 32373
rect 5338 32333 5344 32345
rect 5904 32333 5910 32345
rect 5962 32333 5968 32385
rect 6263 32333 6269 32385
rect 6321 32373 6327 32385
rect 6864 32373 6870 32385
rect 6321 32345 6870 32373
rect 6321 32333 6327 32345
rect 6864 32333 6870 32345
rect 6922 32333 6928 32385
rect 4752 32259 4758 32311
rect 4810 32299 4816 32311
rect 5376 32299 5382 32311
rect 4810 32271 5382 32299
rect 4810 32259 4816 32271
rect 5376 32259 5382 32271
rect 5434 32259 5440 32311
rect 5779 32259 5785 32311
rect 5837 32299 5843 32311
rect 6384 32299 6390 32311
rect 5837 32271 6390 32299
rect 5837 32259 5843 32271
rect 6384 32259 6390 32271
rect 6442 32259 6448 32311
rect 6768 32259 6774 32311
rect 6826 32299 6832 32311
rect 7344 32299 7350 32311
rect 6826 32271 7350 32299
rect 6826 32259 6832 32271
rect 7344 32259 7350 32271
rect 7402 32259 7408 32311
rect 8688 32259 8694 32311
rect 8746 32299 8752 32311
rect 9264 32299 9270 32311
rect 8746 32271 9270 32299
rect 8746 32259 8752 32271
rect 9264 32259 9270 32271
rect 9322 32259 9328 32311
rect 1926 32200 1978 32206
rect 1104 32148 1110 32200
rect 1162 32148 1168 32200
rect 1926 32142 1978 32148
rect 2406 32200 2458 32206
rect 6774 32200 6826 32206
rect 2880 32148 2886 32200
rect 2938 32148 2944 32200
rect 3360 32148 3366 32200
rect 3418 32148 3424 32200
rect 3843 32148 3849 32200
rect 3901 32148 3907 32200
rect 4327 32148 4333 32200
rect 4385 32148 4391 32200
rect 4752 32148 4758 32200
rect 4810 32148 4816 32200
rect 5280 32148 5286 32200
rect 5338 32148 5344 32200
rect 5779 32148 5785 32200
rect 5837 32148 5843 32200
rect 6263 32148 6269 32200
rect 6321 32148 6327 32200
rect 2406 32142 2458 32148
rect 6774 32142 6826 32148
rect 7254 32200 7306 32206
rect 7254 32142 7306 32148
rect 7734 32200 7786 32206
rect 7734 32142 7786 32148
rect 8214 32200 8266 32206
rect 8688 32148 8694 32200
rect 8746 32148 8752 32200
rect 9168 32148 9174 32200
rect 9226 32148 9232 32200
rect 8214 32142 8266 32148
rect 5910 32126 5962 32132
rect 1268 32074 1274 32126
rect 1326 32074 1332 32126
rect 2502 32089 2554 32095
rect 1446 32000 1452 32052
rect 1504 32000 1510 32052
rect 2502 32031 2554 32037
rect 2982 32089 3034 32095
rect 2982 32031 3034 32037
rect 3462 32089 3514 32095
rect 3462 32031 3514 32037
rect 3942 32089 3994 32095
rect 3942 32031 3994 32037
rect 4422 32089 4474 32095
rect 4422 32031 4474 32037
rect 4902 32089 4954 32095
rect 4902 32031 4954 32037
rect 5382 32089 5434 32095
rect 5910 32068 5962 32074
rect 6390 32126 6442 32132
rect 6390 32068 6442 32074
rect 6870 32126 6922 32132
rect 6870 32068 6922 32074
rect 7350 32089 7402 32095
rect 5382 32031 5434 32037
rect 7350 32031 7402 32037
rect 8310 32089 8362 32095
rect 8310 32031 8362 32037
rect 8790 32089 8842 32095
rect 8790 32031 8842 32037
rect 9270 32089 9322 32095
rect 9270 32031 9322 32037
rect 2022 32015 2074 32021
rect 1350 31978 1402 31984
rect 2022 31957 2074 31963
rect 1350 31920 1402 31926
rect 7830 31941 7882 31947
rect 7830 31883 7882 31889
rect 1296 31667 1302 31719
rect 1354 31707 1360 31719
rect 1776 31707 1782 31719
rect 1354 31679 1782 31707
rect 1354 31667 1360 31679
rect 1776 31667 1782 31679
rect 1834 31667 1840 31719
rect 1064 31534 9556 31556
rect 1064 31482 3606 31534
rect 3658 31482 3670 31534
rect 3722 31482 3734 31534
rect 3786 31482 3798 31534
rect 3850 31482 8934 31534
rect 8986 31482 8998 31534
rect 9050 31482 9062 31534
rect 9114 31482 9126 31534
rect 9178 31482 9556 31534
rect 1064 31460 9556 31482
rect 9270 31201 9322 31207
rect 9270 31143 9322 31149
rect 2022 30979 2074 30985
rect 2022 30921 2074 30927
rect 2502 30979 2554 30985
rect 2502 30921 2554 30927
rect 2982 30979 3034 30985
rect 2982 30921 3034 30927
rect 3462 30979 3514 30985
rect 3462 30921 3514 30927
rect 3942 30979 3994 30985
rect 3942 30921 3994 30927
rect 4422 30979 4474 30985
rect 4422 30921 4474 30927
rect 4902 30979 4954 30985
rect 4902 30921 4954 30927
rect 5382 30979 5434 30985
rect 7350 30979 7402 30985
rect 5382 30921 5434 30927
rect 5910 30942 5962 30948
rect 5910 30884 5962 30890
rect 6390 30942 6442 30948
rect 6390 30884 6442 30890
rect 6870 30942 6922 30948
rect 7350 30921 7402 30927
rect 7830 30979 7882 30985
rect 7830 30921 7882 30927
rect 8310 30979 8362 30985
rect 8310 30921 8362 30927
rect 8790 30979 8842 30985
rect 8790 30921 8842 30927
rect 6870 30884 6922 30890
rect 2838 30868 2890 30874
rect 1872 30816 1878 30868
rect 1930 30816 1936 30868
rect 2352 30816 2358 30868
rect 2410 30816 2416 30868
rect 2838 30810 2890 30816
rect 3318 30868 3370 30874
rect 3318 30810 3370 30816
rect 3798 30868 3850 30874
rect 3798 30810 3850 30816
rect 4278 30868 4330 30874
rect 6774 30868 6826 30874
rect 4752 30816 4758 30868
rect 4810 30816 4816 30868
rect 5278 30816 5284 30868
rect 5336 30816 5342 30868
rect 5760 30816 5766 30868
rect 5818 30816 5824 30868
rect 6240 30816 6246 30868
rect 6298 30816 6304 30868
rect 4278 30810 4330 30816
rect 6774 30810 6826 30816
rect 7254 30868 7306 30874
rect 7254 30810 7306 30816
rect 7734 30868 7786 30874
rect 7734 30810 7786 30816
rect 8214 30868 8266 30874
rect 8688 30816 8694 30868
rect 8746 30816 8752 30868
rect 9168 30816 9174 30868
rect 9226 30816 9232 30868
rect 8214 30810 8266 30816
rect 1064 30202 9556 30224
rect 1064 30150 6270 30202
rect 6322 30150 6334 30202
rect 6386 30150 6398 30202
rect 6450 30150 6462 30202
rect 6514 30150 9556 30202
rect 1064 30128 9556 30150
rect 5280 29669 5286 29721
rect 5338 29709 5344 29721
rect 5904 29709 5910 29721
rect 5338 29681 5910 29709
rect 5338 29669 5344 29681
rect 5904 29669 5910 29681
rect 5962 29669 5968 29721
rect 6263 29669 6269 29721
rect 6321 29709 6327 29721
rect 6864 29709 6870 29721
rect 6321 29681 6870 29709
rect 6321 29669 6327 29681
rect 6864 29669 6870 29681
rect 6922 29669 6928 29721
rect 4752 29595 4758 29647
rect 4810 29635 4816 29647
rect 5376 29635 5382 29647
rect 4810 29607 5382 29635
rect 4810 29595 4816 29607
rect 5376 29595 5382 29607
rect 5434 29595 5440 29647
rect 5779 29595 5785 29647
rect 5837 29635 5843 29647
rect 6384 29635 6390 29647
rect 5837 29607 6390 29635
rect 5837 29595 5843 29607
rect 6384 29595 6390 29607
rect 6442 29595 6448 29647
rect 6768 29595 6774 29647
rect 6826 29635 6832 29647
rect 7344 29635 7350 29647
rect 6826 29607 7350 29635
rect 6826 29595 6832 29607
rect 7344 29595 7350 29607
rect 7402 29595 7408 29647
rect 8688 29595 8694 29647
rect 8746 29635 8752 29647
rect 9264 29635 9270 29647
rect 8746 29607 9270 29635
rect 8746 29595 8752 29607
rect 9264 29595 9270 29607
rect 9322 29595 9328 29647
rect 2406 29536 2458 29542
rect 6774 29536 6826 29542
rect 1872 29484 1878 29536
rect 1930 29484 1936 29536
rect 2880 29484 2886 29536
rect 2938 29484 2944 29536
rect 3360 29484 3366 29536
rect 3418 29484 3424 29536
rect 3843 29484 3849 29536
rect 3901 29484 3907 29536
rect 4327 29484 4333 29536
rect 4385 29484 4391 29536
rect 4752 29484 4758 29536
rect 4810 29484 4816 29536
rect 5280 29484 5286 29536
rect 5338 29484 5344 29536
rect 5779 29484 5785 29536
rect 5837 29484 5843 29536
rect 6263 29484 6269 29536
rect 6321 29484 6327 29536
rect 2406 29478 2458 29484
rect 6774 29478 6826 29484
rect 7254 29536 7306 29542
rect 7254 29478 7306 29484
rect 7734 29536 7786 29542
rect 7734 29478 7786 29484
rect 8214 29536 8266 29542
rect 8688 29484 8694 29536
rect 8746 29484 8752 29536
rect 9168 29484 9174 29536
rect 9226 29484 9232 29536
rect 8214 29478 8266 29484
rect 5910 29462 5962 29468
rect 2022 29425 2074 29431
rect 2022 29367 2074 29373
rect 2982 29425 3034 29431
rect 2982 29367 3034 29373
rect 3462 29425 3514 29431
rect 3462 29367 3514 29373
rect 3942 29425 3994 29431
rect 3942 29367 3994 29373
rect 4422 29425 4474 29431
rect 4422 29367 4474 29373
rect 4902 29425 4954 29431
rect 4902 29367 4954 29373
rect 5382 29425 5434 29431
rect 5910 29404 5962 29410
rect 6390 29462 6442 29468
rect 6390 29404 6442 29410
rect 6870 29462 6922 29468
rect 6870 29404 6922 29410
rect 7350 29425 7402 29431
rect 5382 29367 5434 29373
rect 7350 29367 7402 29373
rect 8310 29425 8362 29431
rect 8310 29367 8362 29373
rect 8790 29425 8842 29431
rect 8790 29367 8842 29373
rect 9270 29425 9322 29431
rect 9270 29367 9322 29373
rect 2502 29351 2554 29357
rect 2502 29293 2554 29299
rect 7830 29277 7882 29283
rect 7830 29219 7882 29225
rect 1064 28870 9556 28892
rect 1064 28818 3606 28870
rect 3658 28818 3670 28870
rect 3722 28818 3734 28870
rect 3786 28818 3798 28870
rect 3850 28818 8934 28870
rect 8986 28818 8998 28870
rect 9050 28818 9062 28870
rect 9114 28818 9126 28870
rect 9178 28818 9556 28870
rect 1064 28796 9556 28818
rect 9270 28537 9322 28543
rect 9270 28479 9322 28485
rect 2022 28315 2074 28321
rect 2022 28257 2074 28263
rect 2502 28315 2554 28321
rect 2502 28257 2554 28263
rect 2982 28315 3034 28321
rect 2982 28257 3034 28263
rect 3462 28315 3514 28321
rect 3462 28257 3514 28263
rect 3942 28315 3994 28321
rect 3942 28257 3994 28263
rect 4422 28315 4474 28321
rect 4422 28257 4474 28263
rect 4902 28315 4954 28321
rect 4902 28257 4954 28263
rect 5382 28315 5434 28321
rect 7350 28315 7402 28321
rect 5382 28257 5434 28263
rect 5910 28278 5962 28284
rect 5910 28220 5962 28226
rect 6390 28278 6442 28284
rect 6390 28220 6442 28226
rect 6870 28278 6922 28284
rect 7350 28257 7402 28263
rect 7830 28315 7882 28321
rect 7830 28257 7882 28263
rect 8310 28315 8362 28321
rect 8310 28257 8362 28263
rect 8790 28315 8842 28321
rect 8790 28257 8842 28263
rect 6870 28220 6922 28226
rect 2838 28204 2890 28210
rect 1872 28152 1878 28204
rect 1930 28152 1936 28204
rect 2352 28152 2358 28204
rect 2410 28152 2416 28204
rect 2838 28146 2890 28152
rect 3318 28204 3370 28210
rect 3318 28146 3370 28152
rect 3798 28204 3850 28210
rect 3798 28146 3850 28152
rect 4278 28204 4330 28210
rect 6774 28204 6826 28210
rect 4752 28152 4758 28204
rect 4810 28152 4816 28204
rect 5278 28152 5284 28204
rect 5336 28152 5342 28204
rect 5760 28152 5766 28204
rect 5818 28152 5824 28204
rect 6240 28152 6246 28204
rect 6298 28152 6304 28204
rect 4278 28146 4330 28152
rect 6774 28146 6826 28152
rect 7254 28204 7306 28210
rect 7254 28146 7306 28152
rect 7734 28204 7786 28210
rect 7734 28146 7786 28152
rect 8214 28204 8266 28210
rect 8688 28152 8694 28204
rect 8746 28152 8752 28204
rect 9168 28152 9174 28204
rect 9226 28152 9232 28204
rect 8214 28146 8266 28152
rect 1064 27538 9556 27560
rect 1064 27486 6270 27538
rect 6322 27486 6334 27538
rect 6386 27486 6398 27538
rect 6450 27486 6462 27538
rect 6514 27486 9556 27538
rect 1064 27464 9556 27486
rect 5280 27005 5286 27057
rect 5338 27045 5344 27057
rect 5904 27045 5910 27057
rect 5338 27017 5910 27045
rect 5338 27005 5344 27017
rect 5904 27005 5910 27017
rect 5962 27005 5968 27057
rect 6263 27005 6269 27057
rect 6321 27045 6327 27057
rect 6864 27045 6870 27057
rect 6321 27017 6870 27045
rect 6321 27005 6327 27017
rect 6864 27005 6870 27017
rect 6922 27005 6928 27057
rect 4752 26931 4758 26983
rect 4810 26971 4816 26983
rect 5376 26971 5382 26983
rect 4810 26943 5382 26971
rect 4810 26931 4816 26943
rect 5376 26931 5382 26943
rect 5434 26931 5440 26983
rect 5779 26931 5785 26983
rect 5837 26971 5843 26983
rect 6384 26971 6390 26983
rect 5837 26943 6390 26971
rect 5837 26931 5843 26943
rect 6384 26931 6390 26943
rect 6442 26931 6448 26983
rect 6768 26931 6774 26983
rect 6826 26971 6832 26983
rect 7344 26971 7350 26983
rect 6826 26943 7350 26971
rect 6826 26931 6832 26943
rect 7344 26931 7350 26943
rect 7402 26931 7408 26983
rect 8688 26931 8694 26983
rect 8746 26971 8752 26983
rect 9264 26971 9270 26983
rect 8746 26943 9270 26971
rect 8746 26931 8752 26943
rect 9264 26931 9270 26943
rect 9322 26931 9328 26983
rect 2406 26872 2458 26878
rect 6774 26872 6826 26878
rect 1872 26820 1878 26872
rect 1930 26820 1936 26872
rect 2880 26820 2886 26872
rect 2938 26820 2944 26872
rect 3360 26820 3366 26872
rect 3418 26820 3424 26872
rect 3843 26820 3849 26872
rect 3901 26820 3907 26872
rect 4327 26820 4333 26872
rect 4385 26820 4391 26872
rect 4752 26820 4758 26872
rect 4810 26820 4816 26872
rect 5280 26820 5286 26872
rect 5338 26820 5344 26872
rect 5779 26820 5785 26872
rect 5837 26820 5843 26872
rect 6263 26820 6269 26872
rect 6321 26820 6327 26872
rect 2406 26814 2458 26820
rect 6774 26814 6826 26820
rect 7254 26872 7306 26878
rect 7254 26814 7306 26820
rect 7734 26872 7786 26878
rect 7734 26814 7786 26820
rect 8214 26872 8266 26878
rect 8688 26820 8694 26872
rect 8746 26820 8752 26872
rect 9168 26820 9174 26872
rect 9226 26820 9232 26872
rect 8214 26814 8266 26820
rect 5910 26798 5962 26804
rect 2022 26761 2074 26767
rect 2022 26703 2074 26709
rect 2982 26761 3034 26767
rect 2982 26703 3034 26709
rect 3462 26761 3514 26767
rect 3462 26703 3514 26709
rect 3942 26761 3994 26767
rect 3942 26703 3994 26709
rect 4422 26761 4474 26767
rect 4422 26703 4474 26709
rect 4902 26761 4954 26767
rect 4902 26703 4954 26709
rect 5382 26761 5434 26767
rect 5910 26740 5962 26746
rect 6390 26798 6442 26804
rect 6390 26740 6442 26746
rect 6870 26798 6922 26804
rect 6870 26740 6922 26746
rect 7350 26761 7402 26767
rect 5382 26703 5434 26709
rect 7350 26703 7402 26709
rect 8310 26761 8362 26767
rect 8310 26703 8362 26709
rect 8790 26761 8842 26767
rect 8790 26703 8842 26709
rect 9270 26761 9322 26767
rect 9270 26703 9322 26709
rect 2502 26687 2554 26693
rect 2502 26629 2554 26635
rect 7830 26687 7882 26693
rect 7830 26629 7882 26635
rect 1064 26206 9556 26228
rect 1064 26154 3606 26206
rect 3658 26154 3670 26206
rect 3722 26154 3734 26206
rect 3786 26154 3798 26206
rect 3850 26154 8934 26206
rect 8986 26154 8998 26206
rect 9050 26154 9062 26206
rect 9114 26154 9126 26206
rect 9178 26154 9556 26206
rect 1064 26132 9556 26154
rect 9270 25873 9322 25879
rect 9270 25815 9322 25821
rect 2022 25651 2074 25657
rect 2022 25593 2074 25599
rect 2502 25651 2554 25657
rect 2502 25593 2554 25599
rect 2982 25651 3034 25657
rect 2982 25593 3034 25599
rect 3462 25651 3514 25657
rect 3462 25593 3514 25599
rect 3942 25651 3994 25657
rect 3942 25593 3994 25599
rect 4422 25651 4474 25657
rect 4422 25593 4474 25599
rect 4902 25651 4954 25657
rect 4902 25593 4954 25599
rect 5382 25651 5434 25657
rect 7350 25651 7402 25657
rect 5382 25593 5434 25599
rect 5910 25614 5962 25620
rect 5910 25556 5962 25562
rect 6390 25614 6442 25620
rect 6390 25556 6442 25562
rect 6870 25614 6922 25620
rect 7350 25593 7402 25599
rect 7830 25651 7882 25657
rect 7830 25593 7882 25599
rect 8310 25651 8362 25657
rect 8310 25593 8362 25599
rect 8790 25651 8842 25657
rect 8790 25593 8842 25599
rect 6870 25556 6922 25562
rect 1926 25540 1978 25546
rect 2838 25540 2890 25546
rect 2352 25488 2358 25540
rect 2410 25488 2416 25540
rect 1926 25482 1978 25488
rect 2838 25482 2890 25488
rect 3318 25540 3370 25546
rect 3318 25482 3370 25488
rect 3798 25540 3850 25546
rect 3798 25482 3850 25488
rect 4278 25540 4330 25546
rect 6774 25540 6826 25546
rect 4752 25488 4758 25540
rect 4810 25488 4816 25540
rect 5278 25488 5284 25540
rect 5336 25488 5342 25540
rect 5760 25488 5766 25540
rect 5818 25488 5824 25540
rect 6240 25488 6246 25540
rect 6298 25488 6304 25540
rect 4278 25482 4330 25488
rect 6774 25482 6826 25488
rect 7254 25540 7306 25546
rect 7254 25482 7306 25488
rect 7734 25540 7786 25546
rect 7734 25482 7786 25488
rect 8214 25540 8266 25546
rect 8688 25488 8694 25540
rect 8746 25488 8752 25540
rect 9168 25488 9174 25540
rect 9226 25488 9232 25540
rect 8214 25482 8266 25488
rect 1064 24874 9556 24896
rect 1064 24822 6270 24874
rect 6322 24822 6334 24874
rect 6386 24822 6398 24874
rect 6450 24822 6462 24874
rect 6514 24822 9556 24874
rect 1064 24800 9556 24822
rect 5779 24267 5785 24319
rect 5837 24307 5843 24319
rect 5837 24279 6430 24307
rect 5837 24267 5843 24279
rect 6402 24245 6430 24279
rect 2406 24208 2458 24214
rect 1872 24156 1878 24208
rect 1930 24156 1936 24208
rect 2880 24156 2886 24208
rect 2938 24156 2944 24208
rect 3360 24156 3366 24208
rect 3418 24156 3424 24208
rect 3843 24156 3849 24208
rect 3901 24156 3907 24208
rect 4327 24156 4333 24208
rect 4385 24156 4391 24208
rect 4811 24156 4817 24208
rect 4869 24156 4875 24208
rect 5295 24156 5301 24208
rect 5353 24156 5359 24208
rect 5779 24156 5785 24208
rect 5837 24156 5843 24208
rect 6263 24156 6269 24208
rect 6321 24156 6327 24208
rect 6384 24193 6390 24245
rect 6442 24193 6448 24245
rect 6774 24208 6826 24214
rect 2406 24150 2458 24156
rect 6774 24150 6826 24156
rect 7254 24208 7306 24214
rect 7254 24150 7306 24156
rect 7734 24208 7786 24214
rect 7734 24150 7786 24156
rect 8214 24208 8266 24214
rect 8688 24156 8694 24208
rect 8746 24156 8752 24208
rect 9168 24156 9174 24208
rect 9226 24156 9232 24208
rect 8214 24150 8266 24156
rect 6390 24134 6442 24140
rect 2022 24097 2074 24103
rect 6390 24076 6442 24082
rect 8310 24097 8362 24103
rect 2022 24039 2074 24045
rect 8310 24039 8362 24045
rect 9270 24097 9322 24103
rect 9270 24039 9322 24045
rect 2502 24023 2554 24029
rect 2502 23965 2554 23971
rect 2982 24023 3034 24029
rect 2982 23965 3034 23971
rect 3462 24023 3514 24029
rect 3462 23965 3514 23971
rect 3942 24023 3994 24029
rect 3942 23965 3994 23971
rect 4422 24023 4474 24029
rect 4422 23965 4474 23971
rect 4902 24023 4954 24029
rect 4902 23965 4954 23971
rect 5382 24023 5434 24029
rect 5382 23965 5434 23971
rect 7350 24023 7402 24029
rect 7350 23965 7402 23971
rect 7830 24023 7882 24029
rect 7830 23965 7882 23971
rect 8790 24023 8842 24029
rect 8790 23965 8842 23971
rect 5910 23838 5962 23844
rect 5910 23780 5962 23786
rect 6870 23838 6922 23844
rect 6870 23780 6922 23786
rect 6288 23675 6294 23727
rect 6346 23715 6352 23727
rect 6864 23715 6870 23727
rect 6346 23687 6870 23715
rect 6346 23675 6352 23687
rect 6864 23675 6870 23687
rect 6922 23675 6928 23727
rect 1064 23542 9556 23564
rect 1064 23490 3606 23542
rect 3658 23490 3670 23542
rect 3722 23490 3734 23542
rect 3786 23490 3798 23542
rect 3850 23490 8934 23542
rect 8986 23490 8998 23542
rect 9050 23490 9062 23542
rect 9114 23490 9126 23542
rect 9178 23490 9556 23542
rect 1064 23468 9556 23490
rect 6390 23246 6442 23252
rect 6390 23188 6442 23194
rect 9270 23209 9322 23215
rect 9270 23151 9322 23157
rect 3942 23135 3994 23141
rect 3942 23077 3994 23083
rect 5382 23135 5434 23141
rect 5382 23077 5434 23083
rect 7830 23135 7882 23141
rect 7830 23077 7882 23083
rect 2022 22987 2074 22993
rect 2022 22929 2074 22935
rect 2502 22987 2554 22993
rect 2502 22929 2554 22935
rect 2982 22987 3034 22993
rect 2982 22929 3034 22935
rect 3462 22987 3514 22993
rect 3462 22929 3514 22935
rect 4422 22987 4474 22993
rect 4422 22929 4474 22935
rect 4902 22987 4954 22993
rect 7350 22987 7402 22993
rect 4902 22929 4954 22935
rect 5910 22950 5962 22956
rect 5910 22892 5962 22898
rect 6870 22950 6922 22956
rect 7350 22929 7402 22935
rect 8310 22987 8362 22993
rect 8310 22929 8362 22935
rect 8790 22987 8842 22993
rect 8790 22929 8842 22935
rect 6870 22892 6922 22898
rect 2838 22876 2890 22882
rect 1872 22824 1878 22876
rect 1930 22824 1936 22876
rect 2352 22824 2358 22876
rect 2410 22824 2416 22876
rect 2838 22818 2890 22824
rect 3318 22876 3370 22882
rect 3318 22818 3370 22824
rect 3798 22876 3850 22882
rect 6774 22876 6826 22882
rect 4310 22824 4316 22876
rect 4368 22824 4374 22876
rect 4752 22824 4758 22876
rect 4810 22824 4816 22876
rect 5278 22824 5284 22876
rect 5336 22824 5342 22876
rect 5760 22824 5766 22876
rect 5818 22824 5824 22876
rect 6240 22824 6246 22876
rect 6298 22824 6304 22876
rect 3798 22818 3850 22824
rect 6774 22818 6826 22824
rect 7254 22876 7306 22882
rect 7254 22818 7306 22824
rect 7734 22876 7786 22882
rect 8160 22824 8166 22876
rect 8218 22824 8224 22876
rect 8688 22824 8694 22876
rect 8746 22824 8752 22876
rect 9168 22824 9174 22876
rect 9226 22824 9232 22876
rect 7734 22818 7786 22824
rect 1064 22210 9556 22232
rect 1064 22158 6270 22210
rect 6322 22158 6334 22210
rect 6386 22158 6398 22210
rect 6450 22158 6462 22210
rect 6514 22158 9556 22210
rect 1064 22136 9556 22158
rect 5280 21677 5286 21729
rect 5338 21717 5344 21729
rect 5904 21717 5910 21729
rect 5338 21689 5910 21717
rect 5338 21677 5344 21689
rect 5904 21677 5910 21689
rect 5962 21677 5968 21729
rect 6263 21677 6269 21729
rect 6321 21717 6327 21729
rect 6864 21717 6870 21729
rect 6321 21689 6870 21717
rect 6321 21677 6327 21689
rect 6864 21677 6870 21689
rect 6922 21677 6928 21729
rect 4752 21603 4758 21655
rect 4810 21643 4816 21655
rect 5376 21643 5382 21655
rect 4810 21615 5382 21643
rect 4810 21603 4816 21615
rect 5376 21603 5382 21615
rect 5434 21603 5440 21655
rect 5779 21603 5785 21655
rect 5837 21643 5843 21655
rect 6384 21643 6390 21655
rect 5837 21615 6390 21643
rect 5837 21603 5843 21615
rect 6384 21603 6390 21615
rect 6442 21603 6448 21655
rect 6768 21603 6774 21655
rect 6826 21643 6832 21655
rect 7344 21643 7350 21655
rect 6826 21615 7350 21643
rect 6826 21603 6832 21615
rect 7344 21603 7350 21615
rect 7402 21603 7408 21655
rect 8688 21603 8694 21655
rect 8746 21643 8752 21655
rect 9264 21643 9270 21655
rect 8746 21615 9270 21643
rect 8746 21603 8752 21615
rect 9264 21603 9270 21615
rect 9322 21603 9328 21655
rect 1926 21544 1978 21550
rect 1104 21492 1110 21544
rect 1162 21492 1168 21544
rect 1926 21486 1978 21492
rect 2406 21544 2458 21550
rect 6774 21544 6826 21550
rect 2880 21492 2886 21544
rect 2938 21492 2944 21544
rect 3360 21492 3366 21544
rect 3418 21492 3424 21544
rect 3843 21492 3849 21544
rect 3901 21492 3907 21544
rect 4327 21492 4333 21544
rect 4385 21492 4391 21544
rect 4752 21492 4758 21544
rect 4810 21492 4816 21544
rect 5280 21492 5286 21544
rect 5338 21492 5344 21544
rect 5779 21492 5785 21544
rect 5837 21492 5843 21544
rect 6263 21492 6269 21544
rect 6321 21492 6327 21544
rect 2406 21486 2458 21492
rect 6774 21486 6826 21492
rect 7254 21544 7306 21550
rect 7254 21486 7306 21492
rect 7734 21544 7786 21550
rect 7734 21486 7786 21492
rect 8214 21544 8266 21550
rect 8688 21492 8694 21544
rect 8746 21492 8752 21544
rect 9168 21492 9174 21544
rect 9226 21492 9232 21544
rect 8214 21486 8266 21492
rect 5910 21470 5962 21476
rect 1268 21418 1274 21470
rect 1326 21418 1332 21470
rect 2502 21433 2554 21439
rect 1446 21344 1452 21396
rect 1504 21344 1510 21396
rect 2502 21375 2554 21381
rect 2982 21433 3034 21439
rect 2982 21375 3034 21381
rect 3462 21433 3514 21439
rect 3462 21375 3514 21381
rect 3942 21433 3994 21439
rect 3942 21375 3994 21381
rect 4422 21433 4474 21439
rect 4422 21375 4474 21381
rect 4902 21433 4954 21439
rect 4902 21375 4954 21381
rect 5382 21433 5434 21439
rect 5910 21412 5962 21418
rect 6390 21470 6442 21476
rect 6390 21412 6442 21418
rect 6870 21470 6922 21476
rect 6870 21412 6922 21418
rect 7350 21433 7402 21439
rect 5382 21375 5434 21381
rect 7350 21375 7402 21381
rect 8310 21433 8362 21439
rect 8310 21375 8362 21381
rect 8790 21433 8842 21439
rect 8790 21375 8842 21381
rect 9270 21433 9322 21439
rect 9270 21375 9322 21381
rect 2022 21359 2074 21365
rect 1350 21322 1402 21328
rect 2022 21301 2074 21307
rect 1350 21264 1402 21270
rect 7830 21285 7882 21291
rect 7830 21227 7882 21233
rect 1296 21011 1302 21063
rect 1354 21051 1360 21063
rect 1776 21051 1782 21063
rect 1354 21023 1782 21051
rect 1354 21011 1360 21023
rect 1776 21011 1782 21023
rect 1834 21011 1840 21063
rect 1064 20878 9556 20900
rect 1064 20826 3606 20878
rect 3658 20826 3670 20878
rect 3722 20826 3734 20878
rect 3786 20826 3798 20878
rect 3850 20826 8934 20878
rect 8986 20826 8998 20878
rect 9050 20826 9062 20878
rect 9114 20826 9126 20878
rect 9178 20826 9556 20878
rect 1064 20804 9556 20826
rect 9270 20545 9322 20551
rect 9270 20487 9322 20493
rect 2022 20323 2074 20329
rect 2022 20265 2074 20271
rect 2502 20323 2554 20329
rect 2502 20265 2554 20271
rect 2982 20323 3034 20329
rect 2982 20265 3034 20271
rect 3462 20323 3514 20329
rect 3462 20265 3514 20271
rect 3942 20323 3994 20329
rect 3942 20265 3994 20271
rect 4422 20323 4474 20329
rect 4422 20265 4474 20271
rect 4902 20323 4954 20329
rect 4902 20265 4954 20271
rect 5382 20323 5434 20329
rect 7350 20323 7402 20329
rect 5382 20265 5434 20271
rect 5910 20286 5962 20292
rect 5910 20228 5962 20234
rect 6390 20286 6442 20292
rect 6390 20228 6442 20234
rect 6870 20286 6922 20292
rect 7350 20265 7402 20271
rect 7830 20323 7882 20329
rect 7830 20265 7882 20271
rect 8310 20323 8362 20329
rect 8310 20265 8362 20271
rect 8790 20323 8842 20329
rect 8790 20265 8842 20271
rect 6870 20228 6922 20234
rect 2838 20212 2890 20218
rect 1872 20160 1878 20212
rect 1930 20160 1936 20212
rect 2352 20160 2358 20212
rect 2410 20160 2416 20212
rect 2838 20154 2890 20160
rect 3318 20212 3370 20218
rect 3318 20154 3370 20160
rect 3798 20212 3850 20218
rect 3798 20154 3850 20160
rect 4278 20212 4330 20218
rect 6774 20212 6826 20218
rect 4752 20160 4758 20212
rect 4810 20160 4816 20212
rect 5278 20160 5284 20212
rect 5336 20160 5342 20212
rect 5760 20160 5766 20212
rect 5818 20160 5824 20212
rect 6240 20160 6246 20212
rect 6298 20160 6304 20212
rect 4278 20154 4330 20160
rect 6774 20154 6826 20160
rect 7254 20212 7306 20218
rect 7254 20154 7306 20160
rect 7734 20212 7786 20218
rect 7734 20154 7786 20160
rect 8214 20212 8266 20218
rect 8688 20160 8694 20212
rect 8746 20160 8752 20212
rect 9168 20160 9174 20212
rect 9226 20160 9232 20212
rect 8214 20154 8266 20160
rect 1064 19546 9556 19568
rect 1064 19494 6270 19546
rect 6322 19494 6334 19546
rect 6386 19494 6398 19546
rect 6450 19494 6462 19546
rect 6514 19494 9556 19546
rect 1064 19472 9556 19494
rect 5280 19013 5286 19065
rect 5338 19053 5344 19065
rect 5904 19053 5910 19065
rect 5338 19025 5910 19053
rect 5338 19013 5344 19025
rect 5904 19013 5910 19025
rect 5962 19013 5968 19065
rect 6263 19013 6269 19065
rect 6321 19053 6327 19065
rect 6864 19053 6870 19065
rect 6321 19025 6870 19053
rect 6321 19013 6327 19025
rect 6864 19013 6870 19025
rect 6922 19013 6928 19065
rect 4752 18939 4758 18991
rect 4810 18979 4816 18991
rect 5376 18979 5382 18991
rect 4810 18951 5382 18979
rect 4810 18939 4816 18951
rect 5376 18939 5382 18951
rect 5434 18939 5440 18991
rect 5779 18939 5785 18991
rect 5837 18979 5843 18991
rect 6384 18979 6390 18991
rect 5837 18951 6390 18979
rect 5837 18939 5843 18951
rect 6384 18939 6390 18951
rect 6442 18939 6448 18991
rect 6768 18939 6774 18991
rect 6826 18979 6832 18991
rect 7344 18979 7350 18991
rect 6826 18951 7350 18979
rect 6826 18939 6832 18951
rect 7344 18939 7350 18951
rect 7402 18939 7408 18991
rect 8688 18939 8694 18991
rect 8746 18979 8752 18991
rect 9264 18979 9270 18991
rect 8746 18951 9270 18979
rect 8746 18939 8752 18951
rect 9264 18939 9270 18951
rect 9322 18939 9328 18991
rect 2406 18880 2458 18886
rect 6774 18880 6826 18886
rect 1872 18828 1878 18880
rect 1930 18828 1936 18880
rect 2880 18828 2886 18880
rect 2938 18828 2944 18880
rect 3360 18828 3366 18880
rect 3418 18828 3424 18880
rect 3843 18828 3849 18880
rect 3901 18828 3907 18880
rect 4327 18828 4333 18880
rect 4385 18828 4391 18880
rect 4752 18828 4758 18880
rect 4810 18828 4816 18880
rect 5280 18828 5286 18880
rect 5338 18828 5344 18880
rect 5779 18828 5785 18880
rect 5837 18828 5843 18880
rect 6263 18828 6269 18880
rect 6321 18828 6327 18880
rect 2406 18822 2458 18828
rect 6774 18822 6826 18828
rect 7254 18880 7306 18886
rect 7254 18822 7306 18828
rect 7734 18880 7786 18886
rect 7734 18822 7786 18828
rect 8214 18880 8266 18886
rect 8688 18828 8694 18880
rect 8746 18828 8752 18880
rect 9168 18828 9174 18880
rect 9226 18828 9232 18880
rect 8214 18822 8266 18828
rect 5910 18806 5962 18812
rect 2022 18769 2074 18775
rect 2022 18711 2074 18717
rect 2982 18769 3034 18775
rect 2982 18711 3034 18717
rect 3462 18769 3514 18775
rect 3462 18711 3514 18717
rect 3942 18769 3994 18775
rect 3942 18711 3994 18717
rect 4422 18769 4474 18775
rect 4422 18711 4474 18717
rect 4902 18769 4954 18775
rect 4902 18711 4954 18717
rect 5382 18769 5434 18775
rect 5910 18748 5962 18754
rect 6390 18806 6442 18812
rect 6390 18748 6442 18754
rect 6870 18806 6922 18812
rect 6870 18748 6922 18754
rect 7350 18769 7402 18775
rect 5382 18711 5434 18717
rect 7350 18711 7402 18717
rect 8310 18769 8362 18775
rect 8310 18711 8362 18717
rect 8790 18769 8842 18775
rect 8790 18711 8842 18717
rect 9270 18769 9322 18775
rect 9270 18711 9322 18717
rect 2502 18695 2554 18701
rect 2502 18637 2554 18643
rect 7830 18621 7882 18627
rect 7830 18563 7882 18569
rect 1064 18214 9556 18236
rect 1064 18162 3606 18214
rect 3658 18162 3670 18214
rect 3722 18162 3734 18214
rect 3786 18162 3798 18214
rect 3850 18162 8934 18214
rect 8986 18162 8998 18214
rect 9050 18162 9062 18214
rect 9114 18162 9126 18214
rect 9178 18162 9556 18214
rect 1064 18140 9556 18162
rect 9270 17881 9322 17887
rect 9270 17823 9322 17829
rect 2022 17659 2074 17665
rect 2022 17601 2074 17607
rect 2502 17659 2554 17665
rect 2502 17601 2554 17607
rect 2982 17659 3034 17665
rect 2982 17601 3034 17607
rect 3462 17659 3514 17665
rect 3462 17601 3514 17607
rect 3942 17659 3994 17665
rect 3942 17601 3994 17607
rect 4422 17659 4474 17665
rect 4422 17601 4474 17607
rect 4902 17659 4954 17665
rect 4902 17601 4954 17607
rect 5382 17659 5434 17665
rect 7350 17659 7402 17665
rect 5382 17601 5434 17607
rect 5910 17622 5962 17628
rect 5910 17564 5962 17570
rect 6390 17622 6442 17628
rect 6390 17564 6442 17570
rect 6870 17622 6922 17628
rect 7350 17601 7402 17607
rect 7830 17659 7882 17665
rect 7830 17601 7882 17607
rect 8310 17659 8362 17665
rect 8310 17601 8362 17607
rect 8790 17659 8842 17665
rect 8790 17601 8842 17607
rect 6870 17564 6922 17570
rect 2838 17548 2890 17554
rect 1872 17496 1878 17548
rect 1930 17496 1936 17548
rect 2352 17496 2358 17548
rect 2410 17496 2416 17548
rect 2838 17490 2890 17496
rect 3318 17548 3370 17554
rect 3318 17490 3370 17496
rect 3798 17548 3850 17554
rect 3798 17490 3850 17496
rect 4278 17548 4330 17554
rect 6774 17548 6826 17554
rect 4752 17496 4758 17548
rect 4810 17496 4816 17548
rect 5278 17496 5284 17548
rect 5336 17496 5342 17548
rect 5760 17496 5766 17548
rect 5818 17496 5824 17548
rect 6240 17496 6246 17548
rect 6298 17496 6304 17548
rect 4278 17490 4330 17496
rect 6774 17490 6826 17496
rect 7254 17548 7306 17554
rect 7254 17490 7306 17496
rect 7734 17548 7786 17554
rect 7734 17490 7786 17496
rect 8214 17548 8266 17554
rect 8688 17496 8694 17548
rect 8746 17496 8752 17548
rect 9168 17496 9174 17548
rect 9226 17496 9232 17548
rect 8214 17490 8266 17496
rect 1064 16882 9556 16904
rect 1064 16830 6270 16882
rect 6322 16830 6334 16882
rect 6386 16830 6398 16882
rect 6450 16830 6462 16882
rect 6514 16830 9556 16882
rect 1064 16808 9556 16830
rect 5280 16349 5286 16401
rect 5338 16389 5344 16401
rect 5904 16389 5910 16401
rect 5338 16361 5910 16389
rect 5338 16349 5344 16361
rect 5904 16349 5910 16361
rect 5962 16349 5968 16401
rect 6263 16349 6269 16401
rect 6321 16389 6327 16401
rect 6864 16389 6870 16401
rect 6321 16361 6870 16389
rect 6321 16349 6327 16361
rect 6864 16349 6870 16361
rect 6922 16349 6928 16401
rect 4752 16275 4758 16327
rect 4810 16315 4816 16327
rect 5376 16315 5382 16327
rect 4810 16287 5382 16315
rect 4810 16275 4816 16287
rect 5376 16275 5382 16287
rect 5434 16275 5440 16327
rect 5779 16275 5785 16327
rect 5837 16315 5843 16327
rect 6384 16315 6390 16327
rect 5837 16287 6390 16315
rect 5837 16275 5843 16287
rect 6384 16275 6390 16287
rect 6442 16275 6448 16327
rect 6768 16275 6774 16327
rect 6826 16315 6832 16327
rect 7344 16315 7350 16327
rect 6826 16287 7350 16315
rect 6826 16275 6832 16287
rect 7344 16275 7350 16287
rect 7402 16275 7408 16327
rect 8688 16275 8694 16327
rect 8746 16315 8752 16327
rect 9264 16315 9270 16327
rect 8746 16287 9270 16315
rect 8746 16275 8752 16287
rect 9264 16275 9270 16287
rect 9322 16275 9328 16327
rect 2406 16216 2458 16222
rect 6774 16216 6826 16222
rect 1872 16164 1878 16216
rect 1930 16164 1936 16216
rect 2880 16164 2886 16216
rect 2938 16164 2944 16216
rect 3360 16164 3366 16216
rect 3418 16164 3424 16216
rect 3843 16164 3849 16216
rect 3901 16164 3907 16216
rect 4327 16164 4333 16216
rect 4385 16164 4391 16216
rect 4752 16164 4758 16216
rect 4810 16164 4816 16216
rect 5280 16164 5286 16216
rect 5338 16164 5344 16216
rect 5779 16164 5785 16216
rect 5837 16164 5843 16216
rect 6263 16164 6269 16216
rect 6321 16164 6327 16216
rect 2406 16158 2458 16164
rect 6774 16158 6826 16164
rect 7254 16216 7306 16222
rect 7254 16158 7306 16164
rect 7734 16216 7786 16222
rect 7734 16158 7786 16164
rect 8214 16216 8266 16222
rect 8688 16164 8694 16216
rect 8746 16164 8752 16216
rect 9168 16164 9174 16216
rect 9226 16164 9232 16216
rect 8214 16158 8266 16164
rect 5910 16142 5962 16148
rect 2022 16105 2074 16111
rect 2022 16047 2074 16053
rect 2982 16105 3034 16111
rect 2982 16047 3034 16053
rect 3462 16105 3514 16111
rect 3462 16047 3514 16053
rect 3942 16105 3994 16111
rect 3942 16047 3994 16053
rect 4422 16105 4474 16111
rect 4422 16047 4474 16053
rect 4902 16105 4954 16111
rect 4902 16047 4954 16053
rect 5382 16105 5434 16111
rect 5910 16084 5962 16090
rect 6390 16142 6442 16148
rect 6390 16084 6442 16090
rect 6870 16142 6922 16148
rect 6870 16084 6922 16090
rect 7350 16105 7402 16111
rect 5382 16047 5434 16053
rect 7350 16047 7402 16053
rect 9270 16105 9322 16111
rect 9270 16047 9322 16053
rect 2502 16031 2554 16037
rect 2502 15973 2554 15979
rect 7830 16031 7882 16037
rect 7830 15973 7882 15979
rect 8310 16031 8362 16037
rect 8310 15973 8362 15979
rect 8790 16031 8842 16037
rect 8790 15973 8842 15979
rect 1064 15550 9556 15572
rect 1064 15498 3606 15550
rect 3658 15498 3670 15550
rect 3722 15498 3734 15550
rect 3786 15498 3798 15550
rect 3850 15498 8934 15550
rect 8986 15498 8998 15550
rect 9050 15498 9062 15550
rect 9114 15498 9126 15550
rect 9178 15498 9556 15550
rect 1064 15476 9556 15498
rect 9270 15217 9322 15223
rect 9270 15159 9322 15165
rect 2022 14995 2074 15001
rect 2022 14937 2074 14943
rect 2502 14995 2554 15001
rect 2502 14937 2554 14943
rect 2982 14995 3034 15001
rect 2982 14937 3034 14943
rect 3462 14995 3514 15001
rect 3462 14937 3514 14943
rect 3942 14995 3994 15001
rect 3942 14937 3994 14943
rect 4422 14995 4474 15001
rect 4422 14937 4474 14943
rect 4902 14995 4954 15001
rect 4902 14937 4954 14943
rect 5382 14995 5434 15001
rect 7350 14995 7402 15001
rect 5382 14937 5434 14943
rect 5910 14958 5962 14964
rect 5910 14900 5962 14906
rect 6390 14958 6442 14964
rect 6390 14900 6442 14906
rect 6870 14958 6922 14964
rect 7350 14937 7402 14943
rect 7830 14995 7882 15001
rect 7830 14937 7882 14943
rect 8310 14995 8362 15001
rect 8310 14937 8362 14943
rect 8790 14995 8842 15001
rect 8790 14937 8842 14943
rect 6870 14900 6922 14906
rect 1926 14884 1978 14890
rect 2838 14884 2890 14890
rect 2352 14832 2358 14884
rect 2410 14832 2416 14884
rect 1926 14826 1978 14832
rect 2838 14826 2890 14832
rect 3318 14884 3370 14890
rect 3318 14826 3370 14832
rect 3798 14884 3850 14890
rect 3798 14826 3850 14832
rect 4278 14884 4330 14890
rect 8646 14884 8698 14890
rect 4752 14832 4758 14884
rect 4810 14832 4816 14884
rect 5278 14832 5284 14884
rect 5336 14832 5342 14884
rect 5760 14832 5766 14884
rect 5818 14832 5824 14884
rect 6240 14832 6246 14884
rect 6298 14832 6304 14884
rect 6720 14832 6726 14884
rect 6778 14832 6784 14884
rect 7200 14832 7206 14884
rect 7258 14832 7264 14884
rect 7680 14832 7686 14884
rect 7738 14832 7744 14884
rect 8160 14832 8166 14884
rect 8218 14832 8224 14884
rect 4278 14826 4330 14832
rect 8646 14826 8698 14832
rect 9126 14884 9178 14890
rect 9126 14826 9178 14832
rect 1064 14218 9556 14240
rect 1064 14166 6270 14218
rect 6322 14166 6334 14218
rect 6386 14166 6398 14218
rect 6450 14166 6462 14218
rect 6514 14166 9556 14218
rect 1064 14144 9556 14166
rect 5779 13611 5785 13663
rect 5837 13651 5843 13663
rect 5837 13623 6430 13651
rect 5837 13611 5843 13623
rect 6402 13589 6430 13623
rect 2406 13552 2458 13558
rect 1872 13500 1878 13552
rect 1930 13500 1936 13552
rect 2880 13500 2886 13552
rect 2938 13500 2944 13552
rect 3360 13500 3366 13552
rect 3418 13500 3424 13552
rect 3843 13500 3849 13552
rect 3901 13500 3907 13552
rect 4327 13500 4333 13552
rect 4385 13500 4391 13552
rect 4811 13500 4817 13552
rect 4869 13500 4875 13552
rect 5295 13500 5301 13552
rect 5353 13500 5359 13552
rect 5779 13500 5785 13552
rect 5837 13500 5843 13552
rect 6263 13500 6269 13552
rect 6321 13500 6327 13552
rect 6384 13537 6390 13589
rect 6442 13537 6448 13589
rect 6774 13552 6826 13558
rect 2406 13494 2458 13500
rect 6774 13494 6826 13500
rect 7254 13552 7306 13558
rect 7254 13494 7306 13500
rect 7734 13552 7786 13558
rect 7734 13494 7786 13500
rect 8214 13552 8266 13558
rect 8688 13500 8694 13552
rect 8746 13500 8752 13552
rect 9168 13500 9174 13552
rect 9226 13500 9232 13552
rect 8214 13494 8266 13500
rect 6390 13478 6442 13484
rect 2022 13441 2074 13447
rect 6390 13420 6442 13426
rect 9270 13441 9322 13447
rect 2022 13383 2074 13389
rect 9270 13383 9322 13389
rect 2502 13367 2554 13373
rect 2502 13309 2554 13315
rect 2982 13367 3034 13373
rect 2982 13309 3034 13315
rect 3462 13367 3514 13373
rect 3462 13309 3514 13315
rect 3942 13367 3994 13373
rect 3942 13309 3994 13315
rect 4422 13367 4474 13373
rect 4422 13309 4474 13315
rect 4902 13367 4954 13373
rect 4902 13309 4954 13315
rect 5382 13367 5434 13373
rect 5382 13309 5434 13315
rect 7350 13367 7402 13373
rect 7350 13309 7402 13315
rect 7830 13367 7882 13373
rect 7830 13309 7882 13315
rect 8310 13367 8362 13373
rect 8310 13309 8362 13315
rect 8790 13367 8842 13373
rect 8790 13309 8842 13315
rect 5910 13182 5962 13188
rect 5910 13124 5962 13130
rect 6870 13182 6922 13188
rect 6870 13124 6922 13130
rect 6288 13019 6294 13071
rect 6346 13059 6352 13071
rect 6864 13059 6870 13071
rect 6346 13031 6870 13059
rect 6346 13019 6352 13031
rect 6864 13019 6870 13031
rect 6922 13019 6928 13071
rect 1064 12886 9556 12908
rect 1064 12834 3606 12886
rect 3658 12834 3670 12886
rect 3722 12834 3734 12886
rect 3786 12834 3798 12886
rect 3850 12834 8934 12886
rect 8986 12834 8998 12886
rect 9050 12834 9062 12886
rect 9114 12834 9126 12886
rect 9178 12834 9556 12886
rect 1064 12812 9556 12834
rect 6390 12590 6442 12596
rect 3942 12553 3994 12559
rect 3942 12495 3994 12501
rect 5382 12553 5434 12559
rect 6390 12532 6442 12538
rect 9270 12553 9322 12559
rect 5382 12495 5434 12501
rect 9270 12495 9322 12501
rect 2022 12331 2074 12337
rect 2022 12273 2074 12279
rect 2502 12331 2554 12337
rect 2502 12273 2554 12279
rect 2982 12331 3034 12337
rect 2982 12273 3034 12279
rect 3462 12331 3514 12337
rect 3462 12273 3514 12279
rect 4422 12331 4474 12337
rect 4422 12273 4474 12279
rect 4902 12331 4954 12337
rect 7350 12331 7402 12337
rect 4902 12273 4954 12279
rect 5910 12294 5962 12300
rect 5910 12236 5962 12242
rect 6870 12294 6922 12300
rect 7350 12273 7402 12279
rect 7830 12331 7882 12337
rect 7830 12273 7882 12279
rect 8310 12331 8362 12337
rect 8310 12273 8362 12279
rect 8790 12331 8842 12337
rect 8790 12273 8842 12279
rect 6870 12236 6922 12242
rect 2838 12220 2890 12226
rect 1872 12168 1878 12220
rect 1930 12168 1936 12220
rect 2352 12168 2358 12220
rect 2410 12168 2416 12220
rect 2838 12162 2890 12168
rect 3318 12220 3370 12226
rect 3318 12162 3370 12168
rect 3798 12220 3850 12226
rect 3798 12162 3850 12168
rect 4278 12220 4330 12226
rect 6774 12220 6826 12226
rect 8646 12220 8698 12226
rect 4752 12168 4758 12220
rect 4810 12168 4816 12220
rect 5278 12168 5284 12220
rect 5336 12168 5342 12220
rect 5762 12168 5768 12220
rect 5820 12168 5826 12220
rect 6240 12168 6246 12220
rect 6298 12168 6304 12220
rect 7200 12168 7206 12220
rect 7258 12168 7264 12220
rect 7680 12168 7686 12220
rect 7738 12168 7744 12220
rect 8160 12168 8166 12220
rect 8218 12168 8224 12220
rect 4278 12162 4330 12168
rect 6774 12162 6826 12168
rect 8646 12162 8698 12168
rect 9126 12220 9178 12226
rect 9126 12162 9178 12168
rect 1064 11554 9556 11576
rect 1064 11502 6270 11554
rect 6322 11502 6334 11554
rect 6386 11502 6398 11554
rect 6450 11502 6462 11554
rect 6514 11502 9556 11554
rect 1064 11480 9556 11502
rect 5280 11021 5286 11073
rect 5338 11061 5344 11073
rect 5904 11061 5910 11073
rect 5338 11033 5910 11061
rect 5338 11021 5344 11033
rect 5904 11021 5910 11033
rect 5962 11021 5968 11073
rect 6263 11021 6269 11073
rect 6321 11061 6327 11073
rect 6864 11061 6870 11073
rect 6321 11033 6870 11061
rect 6321 11021 6327 11033
rect 6864 11021 6870 11033
rect 6922 11021 6928 11073
rect 4752 10947 4758 10999
rect 4810 10987 4816 10999
rect 5376 10987 5382 10999
rect 4810 10959 5382 10987
rect 4810 10947 4816 10959
rect 5376 10947 5382 10959
rect 5434 10947 5440 10999
rect 5779 10947 5785 10999
rect 5837 10987 5843 10999
rect 6384 10987 6390 10999
rect 5837 10959 6390 10987
rect 5837 10947 5843 10959
rect 6384 10947 6390 10959
rect 6442 10947 6448 10999
rect 6768 10947 6774 10999
rect 6826 10987 6832 10999
rect 7344 10987 7350 10999
rect 6826 10959 7350 10987
rect 6826 10947 6832 10959
rect 7344 10947 7350 10959
rect 7402 10947 7408 10999
rect 8688 10947 8694 10999
rect 8746 10987 8752 10999
rect 9264 10987 9270 10999
rect 8746 10959 9270 10987
rect 8746 10947 8752 10959
rect 9264 10947 9270 10959
rect 9322 10947 9328 10999
rect 2406 10888 2458 10894
rect 6774 10888 6826 10894
rect 1872 10836 1878 10888
rect 1930 10836 1936 10888
rect 2880 10836 2886 10888
rect 2938 10836 2944 10888
rect 3360 10836 3366 10888
rect 3418 10836 3424 10888
rect 3843 10836 3849 10888
rect 3901 10836 3907 10888
rect 4327 10836 4333 10888
rect 4385 10836 4391 10888
rect 4752 10836 4758 10888
rect 4810 10836 4816 10888
rect 5280 10836 5286 10888
rect 5338 10836 5344 10888
rect 5779 10836 5785 10888
rect 5837 10836 5843 10888
rect 6263 10836 6269 10888
rect 6321 10836 6327 10888
rect 2406 10830 2458 10836
rect 6774 10830 6826 10836
rect 7254 10888 7306 10894
rect 7254 10830 7306 10836
rect 7734 10888 7786 10894
rect 7734 10830 7786 10836
rect 8214 10888 8266 10894
rect 8688 10836 8694 10888
rect 8746 10836 8752 10888
rect 9168 10836 9174 10888
rect 9226 10836 9232 10888
rect 8214 10830 8266 10836
rect 5910 10814 5962 10820
rect 2022 10777 2074 10783
rect 2022 10719 2074 10725
rect 2982 10777 3034 10783
rect 2982 10719 3034 10725
rect 3462 10777 3514 10783
rect 3462 10719 3514 10725
rect 3942 10777 3994 10783
rect 3942 10719 3994 10725
rect 4422 10777 4474 10783
rect 4422 10719 4474 10725
rect 4902 10777 4954 10783
rect 4902 10719 4954 10725
rect 5382 10777 5434 10783
rect 5910 10756 5962 10762
rect 6390 10814 6442 10820
rect 6390 10756 6442 10762
rect 6870 10814 6922 10820
rect 6870 10756 6922 10762
rect 7350 10777 7402 10783
rect 5382 10719 5434 10725
rect 7350 10719 7402 10725
rect 9270 10777 9322 10783
rect 9270 10719 9322 10725
rect 2502 10703 2554 10709
rect 2502 10645 2554 10651
rect 8310 10703 8362 10709
rect 8310 10645 8362 10651
rect 8790 10703 8842 10709
rect 8790 10645 8842 10651
rect 7830 10629 7882 10635
rect 7830 10571 7882 10577
rect 1064 10222 9556 10244
rect 1064 10170 3606 10222
rect 3658 10170 3670 10222
rect 3722 10170 3734 10222
rect 3786 10170 3798 10222
rect 3850 10170 8934 10222
rect 8986 10170 8998 10222
rect 9050 10170 9062 10222
rect 9114 10170 9126 10222
rect 9178 10170 9556 10222
rect 1064 10148 9556 10170
rect 9270 9889 9322 9895
rect 9270 9831 9322 9837
rect 2022 9667 2074 9673
rect 2022 9609 2074 9615
rect 2502 9667 2554 9673
rect 2502 9609 2554 9615
rect 2982 9667 3034 9673
rect 2982 9609 3034 9615
rect 3462 9667 3514 9673
rect 3462 9609 3514 9615
rect 3942 9667 3994 9673
rect 3942 9609 3994 9615
rect 4422 9667 4474 9673
rect 4422 9609 4474 9615
rect 4902 9667 4954 9673
rect 4902 9609 4954 9615
rect 5382 9667 5434 9673
rect 7350 9667 7402 9673
rect 5382 9609 5434 9615
rect 5910 9630 5962 9636
rect 5910 9572 5962 9578
rect 6390 9630 6442 9636
rect 6390 9572 6442 9578
rect 6870 9630 6922 9636
rect 7350 9609 7402 9615
rect 7830 9667 7882 9673
rect 7830 9609 7882 9615
rect 8310 9667 8362 9673
rect 8310 9609 8362 9615
rect 8790 9667 8842 9673
rect 8790 9609 8842 9615
rect 6870 9572 6922 9578
rect 2838 9556 2890 9562
rect 1872 9504 1878 9556
rect 1930 9504 1936 9556
rect 2352 9504 2358 9556
rect 2410 9504 2416 9556
rect 2838 9498 2890 9504
rect 3318 9556 3370 9562
rect 3318 9498 3370 9504
rect 3798 9556 3850 9562
rect 3798 9498 3850 9504
rect 4278 9556 4330 9562
rect 8646 9556 8698 9562
rect 4752 9504 4758 9556
rect 4810 9504 4816 9556
rect 5278 9504 5284 9556
rect 5336 9504 5342 9556
rect 5760 9504 5766 9556
rect 5818 9504 5824 9556
rect 6240 9504 6246 9556
rect 6298 9504 6304 9556
rect 6720 9504 6726 9556
rect 6778 9504 6784 9556
rect 7200 9504 7206 9556
rect 7258 9504 7264 9556
rect 7680 9504 7686 9556
rect 7738 9504 7744 9556
rect 8160 9504 8166 9556
rect 8218 9504 8224 9556
rect 4278 9498 4330 9504
rect 8646 9498 8698 9504
rect 9126 9556 9178 9562
rect 9126 9498 9178 9504
rect 1064 8890 9556 8912
rect 1064 8838 6270 8890
rect 6322 8838 6334 8890
rect 6386 8838 6398 8890
rect 6450 8838 6462 8890
rect 6514 8838 9556 8890
rect 1064 8816 9556 8838
rect 5280 8357 5286 8409
rect 5338 8397 5344 8409
rect 5904 8397 5910 8409
rect 5338 8369 5910 8397
rect 5338 8357 5344 8369
rect 5904 8357 5910 8369
rect 5962 8357 5968 8409
rect 6263 8357 6269 8409
rect 6321 8397 6327 8409
rect 6864 8397 6870 8409
rect 6321 8369 6870 8397
rect 6321 8357 6327 8369
rect 6864 8357 6870 8369
rect 6922 8357 6928 8409
rect 4752 8283 4758 8335
rect 4810 8323 4816 8335
rect 5376 8323 5382 8335
rect 4810 8295 5382 8323
rect 4810 8283 4816 8295
rect 5376 8283 5382 8295
rect 5434 8283 5440 8335
rect 5779 8283 5785 8335
rect 5837 8323 5843 8335
rect 6384 8323 6390 8335
rect 5837 8295 6390 8323
rect 5837 8283 5843 8295
rect 6384 8283 6390 8295
rect 6442 8283 6448 8335
rect 6768 8283 6774 8335
rect 6826 8323 6832 8335
rect 7344 8323 7350 8335
rect 6826 8295 7350 8323
rect 6826 8283 6832 8295
rect 7344 8283 7350 8295
rect 7402 8283 7408 8335
rect 8688 8283 8694 8335
rect 8746 8323 8752 8335
rect 9264 8323 9270 8335
rect 8746 8295 9270 8323
rect 8746 8283 8752 8295
rect 9264 8283 9270 8295
rect 9322 8283 9328 8335
rect 2406 8224 2458 8230
rect 6774 8224 6826 8230
rect 1872 8172 1878 8224
rect 1930 8172 1936 8224
rect 2880 8172 2886 8224
rect 2938 8172 2944 8224
rect 3360 8172 3366 8224
rect 3418 8172 3424 8224
rect 3843 8172 3849 8224
rect 3901 8172 3907 8224
rect 4327 8172 4333 8224
rect 4385 8172 4391 8224
rect 4752 8172 4758 8224
rect 4810 8172 4816 8224
rect 5280 8172 5286 8224
rect 5338 8172 5344 8224
rect 5779 8172 5785 8224
rect 5837 8172 5843 8224
rect 6263 8172 6269 8224
rect 6321 8172 6327 8224
rect 2406 8166 2458 8172
rect 6774 8166 6826 8172
rect 7254 8224 7306 8230
rect 7254 8166 7306 8172
rect 7734 8224 7786 8230
rect 7734 8166 7786 8172
rect 8214 8224 8266 8230
rect 8688 8172 8694 8224
rect 8746 8172 8752 8224
rect 9168 8172 9174 8224
rect 9226 8172 9232 8224
rect 8214 8166 8266 8172
rect 5910 8150 5962 8156
rect 2022 8113 2074 8119
rect 2022 8055 2074 8061
rect 2982 8113 3034 8119
rect 2982 8055 3034 8061
rect 3462 8113 3514 8119
rect 3462 8055 3514 8061
rect 3942 8113 3994 8119
rect 3942 8055 3994 8061
rect 4422 8113 4474 8119
rect 4422 8055 4474 8061
rect 4902 8113 4954 8119
rect 4902 8055 4954 8061
rect 5382 8113 5434 8119
rect 5910 8092 5962 8098
rect 6390 8150 6442 8156
rect 6390 8092 6442 8098
rect 6870 8150 6922 8156
rect 6870 8092 6922 8098
rect 7350 8113 7402 8119
rect 5382 8055 5434 8061
rect 7350 8055 7402 8061
rect 9270 8113 9322 8119
rect 9270 8055 9322 8061
rect 2502 8039 2554 8045
rect 2502 7981 2554 7987
rect 8310 8039 8362 8045
rect 8310 7981 8362 7987
rect 8790 8039 8842 8045
rect 8790 7981 8842 7987
rect 7830 7965 7882 7971
rect 7830 7907 7882 7913
rect 1064 7558 9556 7580
rect 1064 7506 3606 7558
rect 3658 7506 3670 7558
rect 3722 7506 3734 7558
rect 3786 7506 3798 7558
rect 3850 7506 8934 7558
rect 8986 7506 8998 7558
rect 9050 7506 9062 7558
rect 9114 7506 9126 7558
rect 9178 7506 9556 7558
rect 1064 7484 9556 7506
rect 9270 7225 9322 7231
rect 9270 7167 9322 7173
rect 2022 7003 2074 7009
rect 2022 6945 2074 6951
rect 2502 7003 2554 7009
rect 2502 6945 2554 6951
rect 2982 7003 3034 7009
rect 2982 6945 3034 6951
rect 3462 7003 3514 7009
rect 3462 6945 3514 6951
rect 3942 7003 3994 7009
rect 3942 6945 3994 6951
rect 4422 7003 4474 7009
rect 4422 6945 4474 6951
rect 4902 7003 4954 7009
rect 4902 6945 4954 6951
rect 5382 7003 5434 7009
rect 7350 7003 7402 7009
rect 5382 6945 5434 6951
rect 5910 6966 5962 6972
rect 5910 6908 5962 6914
rect 6390 6966 6442 6972
rect 6390 6908 6442 6914
rect 6870 6966 6922 6972
rect 7350 6945 7402 6951
rect 7830 7003 7882 7009
rect 7830 6945 7882 6951
rect 8310 7003 8362 7009
rect 8310 6945 8362 6951
rect 8790 7003 8842 7009
rect 8790 6945 8842 6951
rect 6870 6908 6922 6914
rect 2838 6892 2890 6898
rect 1872 6840 1878 6892
rect 1930 6840 1936 6892
rect 2352 6840 2358 6892
rect 2410 6840 2416 6892
rect 2838 6834 2890 6840
rect 3318 6892 3370 6898
rect 3318 6834 3370 6840
rect 3798 6892 3850 6898
rect 3798 6834 3850 6840
rect 4278 6892 4330 6898
rect 8646 6892 8698 6898
rect 4752 6840 4758 6892
rect 4810 6840 4816 6892
rect 5278 6840 5284 6892
rect 5336 6840 5342 6892
rect 5760 6840 5766 6892
rect 5818 6840 5824 6892
rect 6240 6840 6246 6892
rect 6298 6840 6304 6892
rect 6720 6840 6726 6892
rect 6778 6840 6784 6892
rect 7200 6840 7206 6892
rect 7258 6840 7264 6892
rect 7680 6840 7686 6892
rect 7738 6840 7744 6892
rect 8160 6840 8166 6892
rect 8218 6840 8224 6892
rect 4278 6834 4330 6840
rect 8646 6834 8698 6840
rect 9126 6892 9178 6898
rect 9126 6834 9178 6840
rect 1064 6226 9556 6248
rect 1064 6174 6270 6226
rect 6322 6174 6334 6226
rect 6386 6174 6398 6226
rect 6450 6174 6462 6226
rect 6514 6174 9556 6226
rect 1064 6152 9556 6174
rect 5280 5693 5286 5745
rect 5338 5733 5344 5745
rect 5904 5733 5910 5745
rect 5338 5705 5910 5733
rect 5338 5693 5344 5705
rect 5904 5693 5910 5705
rect 5962 5693 5968 5745
rect 6263 5693 6269 5745
rect 6321 5733 6327 5745
rect 6864 5733 6870 5745
rect 6321 5705 6870 5733
rect 6321 5693 6327 5705
rect 6864 5693 6870 5705
rect 6922 5693 6928 5745
rect 4752 5619 4758 5671
rect 4810 5659 4816 5671
rect 5376 5659 5382 5671
rect 4810 5631 5382 5659
rect 4810 5619 4816 5631
rect 5376 5619 5382 5631
rect 5434 5619 5440 5671
rect 5779 5619 5785 5671
rect 5837 5659 5843 5671
rect 6384 5659 6390 5671
rect 5837 5631 6390 5659
rect 5837 5619 5843 5631
rect 6384 5619 6390 5631
rect 6442 5619 6448 5671
rect 6768 5619 6774 5671
rect 6826 5659 6832 5671
rect 7344 5659 7350 5671
rect 6826 5631 7350 5659
rect 6826 5619 6832 5631
rect 7344 5619 7350 5631
rect 7402 5619 7408 5671
rect 8688 5619 8694 5671
rect 8746 5659 8752 5671
rect 9264 5659 9270 5671
rect 8746 5631 9270 5659
rect 8746 5619 8752 5631
rect 9264 5619 9270 5631
rect 9322 5619 9328 5671
rect 2406 5560 2458 5566
rect 6774 5560 6826 5566
rect 1872 5508 1878 5560
rect 1930 5508 1936 5560
rect 2880 5508 2886 5560
rect 2938 5508 2944 5560
rect 3360 5508 3366 5560
rect 3418 5508 3424 5560
rect 3843 5508 3849 5560
rect 3901 5508 3907 5560
rect 4327 5508 4333 5560
rect 4385 5508 4391 5560
rect 4752 5508 4758 5560
rect 4810 5508 4816 5560
rect 5280 5508 5286 5560
rect 5338 5508 5344 5560
rect 5779 5508 5785 5560
rect 5837 5508 5843 5560
rect 6263 5508 6269 5560
rect 6321 5508 6327 5560
rect 2406 5502 2458 5508
rect 6774 5502 6826 5508
rect 7254 5560 7306 5566
rect 7254 5502 7306 5508
rect 7734 5560 7786 5566
rect 7734 5502 7786 5508
rect 8214 5560 8266 5566
rect 8688 5508 8694 5560
rect 8746 5508 8752 5560
rect 9168 5508 9174 5560
rect 9226 5508 9232 5560
rect 8214 5502 8266 5508
rect 5910 5486 5962 5492
rect 2022 5449 2074 5455
rect 2022 5391 2074 5397
rect 2982 5449 3034 5455
rect 2982 5391 3034 5397
rect 3462 5449 3514 5455
rect 3462 5391 3514 5397
rect 3942 5449 3994 5455
rect 3942 5391 3994 5397
rect 4422 5449 4474 5455
rect 4422 5391 4474 5397
rect 4902 5449 4954 5455
rect 4902 5391 4954 5397
rect 5382 5449 5434 5455
rect 5910 5428 5962 5434
rect 6390 5486 6442 5492
rect 6390 5428 6442 5434
rect 6870 5486 6922 5492
rect 6870 5428 6922 5434
rect 7350 5449 7402 5455
rect 5382 5391 5434 5397
rect 7350 5391 7402 5397
rect 9270 5449 9322 5455
rect 9270 5391 9322 5397
rect 2502 5375 2554 5381
rect 2502 5317 2554 5323
rect 7830 5375 7882 5381
rect 7830 5317 7882 5323
rect 8310 5375 8362 5381
rect 8310 5317 8362 5323
rect 8790 5375 8842 5381
rect 8790 5317 8842 5323
rect 1064 4894 9556 4916
rect 1064 4842 3606 4894
rect 3658 4842 3670 4894
rect 3722 4842 3734 4894
rect 3786 4842 3798 4894
rect 3850 4842 8934 4894
rect 8986 4842 8998 4894
rect 9050 4842 9062 4894
rect 9114 4842 9126 4894
rect 9178 4842 9556 4894
rect 1064 4820 9556 4842
rect 9270 4561 9322 4567
rect 9270 4503 9322 4509
rect 2022 4339 2074 4345
rect 2022 4281 2074 4287
rect 2502 4339 2554 4345
rect 2502 4281 2554 4287
rect 2982 4339 3034 4345
rect 2982 4281 3034 4287
rect 3462 4339 3514 4345
rect 3462 4281 3514 4287
rect 3942 4339 3994 4345
rect 3942 4281 3994 4287
rect 4422 4339 4474 4345
rect 4422 4281 4474 4287
rect 4902 4339 4954 4345
rect 4902 4281 4954 4287
rect 5382 4339 5434 4345
rect 7350 4339 7402 4345
rect 5382 4281 5434 4287
rect 5910 4302 5962 4308
rect 5910 4244 5962 4250
rect 6390 4302 6442 4308
rect 6390 4244 6442 4250
rect 6870 4302 6922 4308
rect 7350 4281 7402 4287
rect 7830 4339 7882 4345
rect 7830 4281 7882 4287
rect 8310 4339 8362 4345
rect 8310 4281 8362 4287
rect 8790 4339 8842 4345
rect 8790 4281 8842 4287
rect 6870 4244 6922 4250
rect 2838 4228 2890 4234
rect 1872 4176 1878 4228
rect 1930 4176 1936 4228
rect 2352 4176 2358 4228
rect 2410 4176 2416 4228
rect 2838 4170 2890 4176
rect 3318 4228 3370 4234
rect 3318 4170 3370 4176
rect 3798 4228 3850 4234
rect 3798 4170 3850 4176
rect 4278 4228 4330 4234
rect 8646 4228 8698 4234
rect 4752 4176 4758 4228
rect 4810 4176 4816 4228
rect 5278 4176 5284 4228
rect 5336 4176 5342 4228
rect 5760 4176 5766 4228
rect 5818 4176 5824 4228
rect 6240 4176 6246 4228
rect 6298 4176 6304 4228
rect 6720 4176 6726 4228
rect 6778 4176 6784 4228
rect 7200 4176 7206 4228
rect 7258 4176 7264 4228
rect 7680 4176 7686 4228
rect 7738 4176 7744 4228
rect 8160 4176 8166 4228
rect 8218 4176 8224 4228
rect 4278 4170 4330 4176
rect 8646 4170 8698 4176
rect 9126 4228 9178 4234
rect 9126 4170 9178 4176
rect 1064 3562 9556 3584
rect 1064 3510 6270 3562
rect 6322 3510 6334 3562
rect 6386 3510 6398 3562
rect 6450 3510 6462 3562
rect 6514 3510 9556 3562
rect 1064 3488 9556 3510
rect 5779 2955 5785 3007
rect 5837 2995 5843 3007
rect 5837 2967 6430 2995
rect 5837 2955 5843 2967
rect 6402 2933 6430 2967
rect 2406 2896 2458 2902
rect 1872 2844 1878 2896
rect 1930 2844 1936 2896
rect 2880 2844 2886 2896
rect 2938 2844 2944 2896
rect 3360 2844 3366 2896
rect 3418 2844 3424 2896
rect 3843 2844 3849 2896
rect 3901 2844 3907 2896
rect 4327 2844 4333 2896
rect 4385 2844 4391 2896
rect 4811 2844 4817 2896
rect 4869 2844 4875 2896
rect 5295 2844 5301 2896
rect 5353 2844 5359 2896
rect 5779 2844 5785 2896
rect 5837 2844 5843 2896
rect 6263 2844 6269 2896
rect 6321 2844 6327 2896
rect 6384 2881 6390 2933
rect 6442 2881 6448 2933
rect 6774 2896 6826 2902
rect 2406 2838 2458 2844
rect 6774 2838 6826 2844
rect 7254 2896 7306 2902
rect 7254 2838 7306 2844
rect 7734 2896 7786 2902
rect 7734 2838 7786 2844
rect 8214 2896 8266 2902
rect 8688 2844 8694 2896
rect 8746 2844 8752 2896
rect 9168 2844 9174 2896
rect 9226 2844 9232 2896
rect 8214 2838 8266 2844
rect 6390 2822 6442 2828
rect 2022 2785 2074 2791
rect 6390 2764 6442 2770
rect 7350 2785 7402 2791
rect 2022 2727 2074 2733
rect 7350 2727 7402 2733
rect 7830 2785 7882 2791
rect 7830 2727 7882 2733
rect 8310 2785 8362 2791
rect 8310 2727 8362 2733
rect 8790 2785 8842 2791
rect 8790 2727 8842 2733
rect 9270 2785 9322 2791
rect 9270 2727 9322 2733
rect 2502 2711 2554 2717
rect 2502 2653 2554 2659
rect 2982 2711 3034 2717
rect 2982 2653 3034 2659
rect 3462 2711 3514 2717
rect 3462 2653 3514 2659
rect 3942 2711 3994 2717
rect 3942 2653 3994 2659
rect 4422 2711 4474 2717
rect 4422 2653 4474 2659
rect 4902 2711 4954 2717
rect 4902 2653 4954 2659
rect 5382 2711 5434 2717
rect 5382 2653 5434 2659
rect 5910 2526 5962 2532
rect 5910 2468 5962 2474
rect 6870 2526 6922 2532
rect 6870 2468 6922 2474
rect 6288 2363 6294 2415
rect 6346 2403 6352 2415
rect 6864 2403 6870 2415
rect 6346 2375 6870 2403
rect 6346 2363 6352 2375
rect 6864 2363 6870 2375
rect 6922 2363 6928 2415
rect 1064 2230 9556 2252
rect 1064 2178 3606 2230
rect 3658 2178 3670 2230
rect 3722 2178 3734 2230
rect 3786 2178 3798 2230
rect 3850 2178 8934 2230
rect 8986 2178 8998 2230
rect 9050 2178 9062 2230
rect 9114 2178 9126 2230
rect 9178 2178 9556 2230
rect 1064 2156 9556 2178
rect 6390 1934 6442 1940
rect 6390 1876 6442 1882
rect 9270 1897 9322 1903
rect 9270 1839 9322 1845
rect 3942 1823 3994 1829
rect 3942 1765 3994 1771
rect 5382 1823 5434 1829
rect 5382 1765 5434 1771
rect 2022 1675 2074 1681
rect 2022 1617 2074 1623
rect 2502 1675 2554 1681
rect 2502 1617 2554 1623
rect 2982 1675 3034 1681
rect 2982 1617 3034 1623
rect 3462 1675 3514 1681
rect 3462 1617 3514 1623
rect 4422 1675 4474 1681
rect 4422 1617 4474 1623
rect 4902 1675 4954 1681
rect 7350 1675 7402 1681
rect 4902 1617 4954 1623
rect 5910 1638 5962 1644
rect 5910 1580 5962 1586
rect 6870 1638 6922 1644
rect 7350 1617 7402 1623
rect 7830 1675 7882 1681
rect 7830 1617 7882 1623
rect 8310 1675 8362 1681
rect 8310 1617 8362 1623
rect 8790 1675 8842 1681
rect 8790 1617 8842 1623
rect 6870 1580 6922 1586
rect 2838 1564 2890 1570
rect 1872 1512 1878 1564
rect 1930 1512 1936 1564
rect 2352 1512 2358 1564
rect 2410 1512 2416 1564
rect 2838 1506 2890 1512
rect 3318 1564 3370 1570
rect 3318 1506 3370 1512
rect 3798 1564 3850 1570
rect 6774 1564 6826 1570
rect 8646 1564 8698 1570
rect 4327 1512 4333 1564
rect 4385 1512 4391 1564
rect 4752 1512 4758 1564
rect 4810 1512 4816 1564
rect 5278 1512 5284 1564
rect 5336 1512 5342 1564
rect 5760 1512 5766 1564
rect 5818 1512 5824 1564
rect 6240 1512 6246 1564
rect 6298 1512 6304 1564
rect 7200 1512 7206 1564
rect 7258 1512 7264 1564
rect 7680 1512 7686 1564
rect 7738 1512 7744 1564
rect 8160 1512 8166 1564
rect 8218 1512 8224 1564
rect 3798 1506 3850 1512
rect 6774 1506 6826 1512
rect 8646 1506 8698 1512
rect 9126 1564 9178 1570
rect 9126 1506 9178 1512
rect 1064 898 9556 920
rect 1064 846 6270 898
rect 6322 846 6334 898
rect 6386 846 6398 898
rect 6450 846 6462 898
rect 6514 846 9556 898
rect 1064 824 9556 846
<< via1 >>
rect 3606 52794 3658 52846
rect 3670 52794 3722 52846
rect 3734 52794 3786 52846
rect 3798 52794 3850 52846
rect 8934 52794 8986 52846
rect 8998 52794 9050 52846
rect 9062 52794 9114 52846
rect 9126 52794 9178 52846
rect 1350 52461 1402 52513
rect 1452 52276 1504 52328
rect 1302 52202 1354 52254
rect 2022 52239 2074 52291
rect 1110 52128 1162 52180
rect 1878 52128 1930 52180
rect 1302 52017 1354 52069
rect 1878 52017 1930 52069
rect 6270 51462 6322 51514
rect 6334 51462 6386 51514
rect 6398 51462 6450 51514
rect 6462 51462 6514 51514
rect 1110 50796 1162 50848
rect 1302 50722 1354 50774
rect 1398 50759 1450 50811
rect 1926 50796 1978 50848
rect 1452 50648 1504 50700
rect 1350 50574 1402 50626
rect 2022 50611 2074 50663
rect 1782 50537 1834 50589
rect 3606 50130 3658 50182
rect 3670 50130 3722 50182
rect 3734 50130 3786 50182
rect 3798 50130 3850 50182
rect 8934 50130 8986 50182
rect 8998 50130 9050 50182
rect 9062 50130 9114 50182
rect 9126 50130 9178 50182
rect 2022 49797 2074 49849
rect 1878 49464 1930 49516
rect 6270 48798 6322 48850
rect 6334 48798 6386 48850
rect 6398 48798 6450 48850
rect 6462 48798 6514 48850
rect 1878 48243 1930 48295
rect 2502 48243 2554 48295
rect 1110 48132 1162 48184
rect 1302 48058 1354 48110
rect 1782 48095 1834 48147
rect 1878 48132 1930 48184
rect 2358 48132 2410 48184
rect 1452 47984 1504 48036
rect 1494 47873 1546 47925
rect 2502 48021 2554 48073
rect 2022 47947 2074 47999
rect 1350 47799 1402 47851
rect 3606 47466 3658 47518
rect 3670 47466 3722 47518
rect 3734 47466 3786 47518
rect 3798 47466 3850 47518
rect 8934 47466 8986 47518
rect 8998 47466 9050 47518
rect 9062 47466 9114 47518
rect 9126 47466 9178 47518
rect 2502 47133 2554 47185
rect 2022 46911 2074 46963
rect 1206 46763 1258 46815
rect 1782 46763 1834 46815
rect 1878 46800 1930 46852
rect 2358 46800 2410 46852
rect 6270 46134 6322 46186
rect 6334 46134 6386 46186
rect 6398 46134 6450 46186
rect 6462 46134 6514 46186
rect 1110 45468 1162 45520
rect 1302 45394 1354 45446
rect 1398 45431 1450 45483
rect 1926 45468 1978 45520
rect 2406 45468 2458 45520
rect 2838 45468 2890 45520
rect 3318 45468 3370 45520
rect 1452 45320 1504 45372
rect 1350 45246 1402 45298
rect 3462 45357 3514 45409
rect 2022 45283 2074 45335
rect 2502 45283 2554 45335
rect 2982 45283 3034 45335
rect 1782 45209 1834 45261
rect 3606 44802 3658 44854
rect 3670 44802 3722 44854
rect 3734 44802 3786 44854
rect 3798 44802 3850 44854
rect 8934 44802 8986 44854
rect 8998 44802 9050 44854
rect 9062 44802 9114 44854
rect 9126 44802 9178 44854
rect 3462 44469 3514 44521
rect 2982 44395 3034 44447
rect 2022 44247 2074 44299
rect 2502 44247 2554 44299
rect 1878 44136 1930 44188
rect 2358 44136 2410 44188
rect 2838 44136 2890 44188
rect 3318 44136 3370 44188
rect 6270 43470 6322 43522
rect 6334 43470 6386 43522
rect 6398 43470 6450 43522
rect 6462 43470 6514 43522
rect 4758 42915 4810 42967
rect 5382 42915 5434 42967
rect 1110 42804 1162 42856
rect 1302 42730 1354 42782
rect 1782 42767 1834 42819
rect 1926 42804 1978 42856
rect 2406 42804 2458 42856
rect 2886 42804 2938 42856
rect 3366 42804 3418 42856
rect 3849 42804 3901 42856
rect 4333 42804 4385 42856
rect 4758 42804 4810 42856
rect 5301 42804 5353 42856
rect 1452 42656 1504 42708
rect 1494 42545 1546 42597
rect 5382 42693 5434 42745
rect 2022 42619 2074 42671
rect 2502 42619 2554 42671
rect 2982 42619 3034 42671
rect 3462 42619 3514 42671
rect 3942 42619 3994 42671
rect 4422 42619 4474 42671
rect 4902 42619 4954 42671
rect 1350 42471 1402 42523
rect 1206 42323 1258 42375
rect 1782 42323 1834 42375
rect 3606 42138 3658 42190
rect 3670 42138 3722 42190
rect 3734 42138 3786 42190
rect 3798 42138 3850 42190
rect 8934 42138 8986 42190
rect 8998 42138 9050 42190
rect 9062 42138 9114 42190
rect 9126 42138 9178 42190
rect 5382 41805 5434 41857
rect 2022 41583 2074 41635
rect 2502 41583 2554 41635
rect 2982 41583 3034 41635
rect 3462 41583 3514 41635
rect 3942 41583 3994 41635
rect 4422 41583 4474 41635
rect 4902 41583 4954 41635
rect 1878 41472 1930 41524
rect 2358 41472 2410 41524
rect 2838 41472 2890 41524
rect 3318 41472 3370 41524
rect 3798 41472 3850 41524
rect 4278 41472 4330 41524
rect 4758 41472 4810 41524
rect 5284 41472 5336 41524
rect 6270 40806 6322 40858
rect 6334 40806 6386 40858
rect 6398 40806 6450 40858
rect 6462 40806 6514 40858
rect 5286 40325 5338 40377
rect 5910 40325 5962 40377
rect 6269 40325 6321 40377
rect 6870 40325 6922 40377
rect 4758 40251 4810 40303
rect 5382 40251 5434 40303
rect 5785 40251 5837 40303
rect 6390 40251 6442 40303
rect 6774 40251 6826 40303
rect 7350 40251 7402 40303
rect 8694 40251 8746 40303
rect 9270 40251 9322 40303
rect 1110 40140 1162 40192
rect 1926 40140 1978 40192
rect 2406 40140 2458 40192
rect 2886 40140 2938 40192
rect 3366 40140 3418 40192
rect 3849 40140 3901 40192
rect 4333 40140 4385 40192
rect 4758 40140 4810 40192
rect 5286 40140 5338 40192
rect 5785 40140 5837 40192
rect 6269 40140 6321 40192
rect 6774 40140 6826 40192
rect 7254 40140 7306 40192
rect 7734 40140 7786 40192
rect 8214 40140 8266 40192
rect 8694 40140 8746 40192
rect 9174 40140 9226 40192
rect 1274 40066 1326 40118
rect 1452 39992 1504 40044
rect 2502 40029 2554 40081
rect 2982 40029 3034 40081
rect 3462 40029 3514 40081
rect 3942 40029 3994 40081
rect 4422 40029 4474 40081
rect 4902 40029 4954 40081
rect 5382 40029 5434 40081
rect 5910 40066 5962 40118
rect 6390 40066 6442 40118
rect 6870 40066 6922 40118
rect 7350 40029 7402 40081
rect 8310 40029 8362 40081
rect 8790 40029 8842 40081
rect 9270 40029 9322 40081
rect 1350 39918 1402 39970
rect 2022 39955 2074 40007
rect 7830 39881 7882 39933
rect 3606 39474 3658 39526
rect 3670 39474 3722 39526
rect 3734 39474 3786 39526
rect 3798 39474 3850 39526
rect 8934 39474 8986 39526
rect 8998 39474 9050 39526
rect 9062 39474 9114 39526
rect 9126 39474 9178 39526
rect 9270 39141 9322 39193
rect 2022 38919 2074 38971
rect 2502 38919 2554 38971
rect 2982 38919 3034 38971
rect 3462 38919 3514 38971
rect 3942 38919 3994 38971
rect 4422 38919 4474 38971
rect 4902 38919 4954 38971
rect 5382 38919 5434 38971
rect 5910 38882 5962 38934
rect 6390 38882 6442 38934
rect 6870 38882 6922 38934
rect 7350 38919 7402 38971
rect 7830 38919 7882 38971
rect 8310 38919 8362 38971
rect 8790 38919 8842 38971
rect 1878 38808 1930 38860
rect 2358 38808 2410 38860
rect 2838 38808 2890 38860
rect 3318 38808 3370 38860
rect 3798 38808 3850 38860
rect 4278 38808 4330 38860
rect 4758 38808 4810 38860
rect 5284 38808 5336 38860
rect 5766 38808 5818 38860
rect 6246 38808 6298 38860
rect 6726 38808 6778 38860
rect 7254 38808 7306 38860
rect 7734 38808 7786 38860
rect 8214 38808 8266 38860
rect 8694 38808 8746 38860
rect 9174 38808 9226 38860
rect 1206 38697 1258 38749
rect 1878 38697 1930 38749
rect 6270 38142 6322 38194
rect 6334 38142 6386 38194
rect 6398 38142 6450 38194
rect 6462 38142 6514 38194
rect 5785 37661 5837 37713
rect 5301 37587 5353 37639
rect 5910 37587 5962 37639
rect 6269 37661 6321 37713
rect 6870 37661 6922 37713
rect 6390 37587 6442 37639
rect 6774 37587 6826 37639
rect 7350 37587 7402 37639
rect 8694 37587 8746 37639
rect 9270 37587 9322 37639
rect 1110 37476 1162 37528
rect 1302 37402 1354 37454
rect 1398 37439 1450 37491
rect 1926 37476 1978 37528
rect 2406 37476 2458 37528
rect 2886 37476 2938 37528
rect 3366 37476 3418 37528
rect 3849 37476 3901 37528
rect 4333 37476 4385 37528
rect 4817 37476 4869 37528
rect 5301 37476 5353 37528
rect 5785 37476 5837 37528
rect 6269 37476 6321 37528
rect 6774 37476 6826 37528
rect 7254 37476 7306 37528
rect 7734 37476 7786 37528
rect 8214 37476 8266 37528
rect 8694 37476 8746 37528
rect 9174 37476 9226 37528
rect 1452 37328 1504 37380
rect 1350 37254 1402 37306
rect 2502 37365 2554 37417
rect 2982 37365 3034 37417
rect 3462 37365 3514 37417
rect 3942 37365 3994 37417
rect 4422 37365 4474 37417
rect 4902 37365 4954 37417
rect 5382 37365 5434 37417
rect 5910 37402 5962 37454
rect 6390 37402 6442 37454
rect 6870 37402 6922 37454
rect 7350 37365 7402 37417
rect 8310 37365 8362 37417
rect 8790 37365 8842 37417
rect 9270 37365 9322 37417
rect 2022 37291 2074 37343
rect 7830 37291 7882 37343
rect 1782 37217 1834 37269
rect 3606 36810 3658 36862
rect 3670 36810 3722 36862
rect 3734 36810 3786 36862
rect 3798 36810 3850 36862
rect 8934 36810 8986 36862
rect 8998 36810 9050 36862
rect 9062 36810 9114 36862
rect 9126 36810 9178 36862
rect 9270 36477 9322 36529
rect 2022 36255 2074 36307
rect 2502 36255 2554 36307
rect 2982 36255 3034 36307
rect 3462 36255 3514 36307
rect 3942 36255 3994 36307
rect 4422 36255 4474 36307
rect 4902 36255 4954 36307
rect 5382 36255 5434 36307
rect 5910 36218 5962 36270
rect 6390 36218 6442 36270
rect 6870 36218 6922 36270
rect 7350 36255 7402 36307
rect 7830 36255 7882 36307
rect 8310 36255 8362 36307
rect 8790 36255 8842 36307
rect 1926 36144 1978 36196
rect 2358 36144 2410 36196
rect 2838 36144 2890 36196
rect 3318 36144 3370 36196
rect 3798 36144 3850 36196
rect 4278 36144 4330 36196
rect 4758 36144 4810 36196
rect 5284 36144 5336 36196
rect 5766 36144 5818 36196
rect 6246 36144 6298 36196
rect 6726 36144 6778 36196
rect 7206 36144 7258 36196
rect 7686 36144 7738 36196
rect 8166 36144 8218 36196
rect 8646 36144 8698 36196
rect 9126 36144 9178 36196
rect 6270 35478 6322 35530
rect 6334 35478 6386 35530
rect 6398 35478 6450 35530
rect 6462 35478 6514 35530
rect 5785 34923 5837 34975
rect 1878 34812 1930 34864
rect 2406 34812 2458 34864
rect 2886 34812 2938 34864
rect 3366 34812 3418 34864
rect 3849 34812 3901 34864
rect 4333 34812 4385 34864
rect 4817 34812 4869 34864
rect 5301 34812 5353 34864
rect 5785 34812 5837 34864
rect 6269 34812 6321 34864
rect 6390 34849 6442 34901
rect 6774 34812 6826 34864
rect 7254 34812 7306 34864
rect 7734 34812 7786 34864
rect 8214 34812 8266 34864
rect 8694 34812 8746 34864
rect 9174 34812 9226 34864
rect 2022 34701 2074 34753
rect 6390 34738 6442 34790
rect 9270 34701 9322 34753
rect 2502 34627 2554 34679
rect 2982 34627 3034 34679
rect 3462 34627 3514 34679
rect 3942 34627 3994 34679
rect 4422 34627 4474 34679
rect 4902 34627 4954 34679
rect 5382 34627 5434 34679
rect 7350 34627 7402 34679
rect 7830 34627 7882 34679
rect 8310 34627 8362 34679
rect 8790 34627 8842 34679
rect 5910 34442 5962 34494
rect 6870 34442 6922 34494
rect 6294 34331 6346 34383
rect 6870 34331 6922 34383
rect 3606 34146 3658 34198
rect 3670 34146 3722 34198
rect 3734 34146 3786 34198
rect 3798 34146 3850 34198
rect 8934 34146 8986 34198
rect 8998 34146 9050 34198
rect 9062 34146 9114 34198
rect 9126 34146 9178 34198
rect 6390 33850 6442 33902
rect 9270 33813 9322 33865
rect 2982 33739 3034 33791
rect 3942 33739 3994 33791
rect 5382 33739 5434 33791
rect 2022 33591 2074 33643
rect 2502 33591 2554 33643
rect 3462 33591 3514 33643
rect 4422 33591 4474 33643
rect 4902 33591 4954 33643
rect 5910 33554 5962 33606
rect 6870 33554 6922 33606
rect 7350 33591 7402 33643
rect 7830 33591 7882 33643
rect 8310 33591 8362 33643
rect 8790 33591 8842 33643
rect 1878 33480 1930 33532
rect 2358 33480 2410 33532
rect 2838 33480 2890 33532
rect 3318 33480 3370 33532
rect 3798 33480 3850 33532
rect 4278 33480 4330 33532
rect 4758 33480 4810 33532
rect 5284 33480 5336 33532
rect 5766 33480 5818 33532
rect 6246 33480 6298 33532
rect 6774 33480 6826 33532
rect 7206 33480 7258 33532
rect 7734 33480 7786 33532
rect 8214 33480 8266 33532
rect 8694 33480 8746 33532
rect 9174 33480 9226 33532
rect 6270 32814 6322 32866
rect 6334 32814 6386 32866
rect 6398 32814 6450 32866
rect 6462 32814 6514 32866
rect 5286 32333 5338 32385
rect 5910 32333 5962 32385
rect 6269 32333 6321 32385
rect 6870 32333 6922 32385
rect 4758 32259 4810 32311
rect 5382 32259 5434 32311
rect 5785 32259 5837 32311
rect 6390 32259 6442 32311
rect 6774 32259 6826 32311
rect 7350 32259 7402 32311
rect 8694 32259 8746 32311
rect 9270 32259 9322 32311
rect 1110 32148 1162 32200
rect 1926 32148 1978 32200
rect 2406 32148 2458 32200
rect 2886 32148 2938 32200
rect 3366 32148 3418 32200
rect 3849 32148 3901 32200
rect 4333 32148 4385 32200
rect 4758 32148 4810 32200
rect 5286 32148 5338 32200
rect 5785 32148 5837 32200
rect 6269 32148 6321 32200
rect 6774 32148 6826 32200
rect 7254 32148 7306 32200
rect 7734 32148 7786 32200
rect 8214 32148 8266 32200
rect 8694 32148 8746 32200
rect 9174 32148 9226 32200
rect 1274 32074 1326 32126
rect 1452 32000 1504 32052
rect 2502 32037 2554 32089
rect 2982 32037 3034 32089
rect 3462 32037 3514 32089
rect 3942 32037 3994 32089
rect 4422 32037 4474 32089
rect 4902 32037 4954 32089
rect 5382 32037 5434 32089
rect 5910 32074 5962 32126
rect 6390 32074 6442 32126
rect 6870 32074 6922 32126
rect 7350 32037 7402 32089
rect 8310 32037 8362 32089
rect 8790 32037 8842 32089
rect 9270 32037 9322 32089
rect 1350 31926 1402 31978
rect 2022 31963 2074 32015
rect 7830 31889 7882 31941
rect 1302 31667 1354 31719
rect 1782 31667 1834 31719
rect 3606 31482 3658 31534
rect 3670 31482 3722 31534
rect 3734 31482 3786 31534
rect 3798 31482 3850 31534
rect 8934 31482 8986 31534
rect 8998 31482 9050 31534
rect 9062 31482 9114 31534
rect 9126 31482 9178 31534
rect 9270 31149 9322 31201
rect 2022 30927 2074 30979
rect 2502 30927 2554 30979
rect 2982 30927 3034 30979
rect 3462 30927 3514 30979
rect 3942 30927 3994 30979
rect 4422 30927 4474 30979
rect 4902 30927 4954 30979
rect 5382 30927 5434 30979
rect 5910 30890 5962 30942
rect 6390 30890 6442 30942
rect 6870 30890 6922 30942
rect 7350 30927 7402 30979
rect 7830 30927 7882 30979
rect 8310 30927 8362 30979
rect 8790 30927 8842 30979
rect 1878 30816 1930 30868
rect 2358 30816 2410 30868
rect 2838 30816 2890 30868
rect 3318 30816 3370 30868
rect 3798 30816 3850 30868
rect 4278 30816 4330 30868
rect 4758 30816 4810 30868
rect 5284 30816 5336 30868
rect 5766 30816 5818 30868
rect 6246 30816 6298 30868
rect 6774 30816 6826 30868
rect 7254 30816 7306 30868
rect 7734 30816 7786 30868
rect 8214 30816 8266 30868
rect 8694 30816 8746 30868
rect 9174 30816 9226 30868
rect 6270 30150 6322 30202
rect 6334 30150 6386 30202
rect 6398 30150 6450 30202
rect 6462 30150 6514 30202
rect 5286 29669 5338 29721
rect 5910 29669 5962 29721
rect 6269 29669 6321 29721
rect 6870 29669 6922 29721
rect 4758 29595 4810 29647
rect 5382 29595 5434 29647
rect 5785 29595 5837 29647
rect 6390 29595 6442 29647
rect 6774 29595 6826 29647
rect 7350 29595 7402 29647
rect 8694 29595 8746 29647
rect 9270 29595 9322 29647
rect 1878 29484 1930 29536
rect 2406 29484 2458 29536
rect 2886 29484 2938 29536
rect 3366 29484 3418 29536
rect 3849 29484 3901 29536
rect 4333 29484 4385 29536
rect 4758 29484 4810 29536
rect 5286 29484 5338 29536
rect 5785 29484 5837 29536
rect 6269 29484 6321 29536
rect 6774 29484 6826 29536
rect 7254 29484 7306 29536
rect 7734 29484 7786 29536
rect 8214 29484 8266 29536
rect 8694 29484 8746 29536
rect 9174 29484 9226 29536
rect 2022 29373 2074 29425
rect 2982 29373 3034 29425
rect 3462 29373 3514 29425
rect 3942 29373 3994 29425
rect 4422 29373 4474 29425
rect 4902 29373 4954 29425
rect 5382 29373 5434 29425
rect 5910 29410 5962 29462
rect 6390 29410 6442 29462
rect 6870 29410 6922 29462
rect 7350 29373 7402 29425
rect 8310 29373 8362 29425
rect 8790 29373 8842 29425
rect 9270 29373 9322 29425
rect 2502 29299 2554 29351
rect 7830 29225 7882 29277
rect 3606 28818 3658 28870
rect 3670 28818 3722 28870
rect 3734 28818 3786 28870
rect 3798 28818 3850 28870
rect 8934 28818 8986 28870
rect 8998 28818 9050 28870
rect 9062 28818 9114 28870
rect 9126 28818 9178 28870
rect 9270 28485 9322 28537
rect 2022 28263 2074 28315
rect 2502 28263 2554 28315
rect 2982 28263 3034 28315
rect 3462 28263 3514 28315
rect 3942 28263 3994 28315
rect 4422 28263 4474 28315
rect 4902 28263 4954 28315
rect 5382 28263 5434 28315
rect 5910 28226 5962 28278
rect 6390 28226 6442 28278
rect 6870 28226 6922 28278
rect 7350 28263 7402 28315
rect 7830 28263 7882 28315
rect 8310 28263 8362 28315
rect 8790 28263 8842 28315
rect 1878 28152 1930 28204
rect 2358 28152 2410 28204
rect 2838 28152 2890 28204
rect 3318 28152 3370 28204
rect 3798 28152 3850 28204
rect 4278 28152 4330 28204
rect 4758 28152 4810 28204
rect 5284 28152 5336 28204
rect 5766 28152 5818 28204
rect 6246 28152 6298 28204
rect 6774 28152 6826 28204
rect 7254 28152 7306 28204
rect 7734 28152 7786 28204
rect 8214 28152 8266 28204
rect 8694 28152 8746 28204
rect 9174 28152 9226 28204
rect 6270 27486 6322 27538
rect 6334 27486 6386 27538
rect 6398 27486 6450 27538
rect 6462 27486 6514 27538
rect 5286 27005 5338 27057
rect 5910 27005 5962 27057
rect 6269 27005 6321 27057
rect 6870 27005 6922 27057
rect 4758 26931 4810 26983
rect 5382 26931 5434 26983
rect 5785 26931 5837 26983
rect 6390 26931 6442 26983
rect 6774 26931 6826 26983
rect 7350 26931 7402 26983
rect 8694 26931 8746 26983
rect 9270 26931 9322 26983
rect 1878 26820 1930 26872
rect 2406 26820 2458 26872
rect 2886 26820 2938 26872
rect 3366 26820 3418 26872
rect 3849 26820 3901 26872
rect 4333 26820 4385 26872
rect 4758 26820 4810 26872
rect 5286 26820 5338 26872
rect 5785 26820 5837 26872
rect 6269 26820 6321 26872
rect 6774 26820 6826 26872
rect 7254 26820 7306 26872
rect 7734 26820 7786 26872
rect 8214 26820 8266 26872
rect 8694 26820 8746 26872
rect 9174 26820 9226 26872
rect 2022 26709 2074 26761
rect 2982 26709 3034 26761
rect 3462 26709 3514 26761
rect 3942 26709 3994 26761
rect 4422 26709 4474 26761
rect 4902 26709 4954 26761
rect 5382 26709 5434 26761
rect 5910 26746 5962 26798
rect 6390 26746 6442 26798
rect 6870 26746 6922 26798
rect 7350 26709 7402 26761
rect 8310 26709 8362 26761
rect 8790 26709 8842 26761
rect 9270 26709 9322 26761
rect 2502 26635 2554 26687
rect 7830 26635 7882 26687
rect 3606 26154 3658 26206
rect 3670 26154 3722 26206
rect 3734 26154 3786 26206
rect 3798 26154 3850 26206
rect 8934 26154 8986 26206
rect 8998 26154 9050 26206
rect 9062 26154 9114 26206
rect 9126 26154 9178 26206
rect 9270 25821 9322 25873
rect 2022 25599 2074 25651
rect 2502 25599 2554 25651
rect 2982 25599 3034 25651
rect 3462 25599 3514 25651
rect 3942 25599 3994 25651
rect 4422 25599 4474 25651
rect 4902 25599 4954 25651
rect 5382 25599 5434 25651
rect 5910 25562 5962 25614
rect 6390 25562 6442 25614
rect 6870 25562 6922 25614
rect 7350 25599 7402 25651
rect 7830 25599 7882 25651
rect 8310 25599 8362 25651
rect 8790 25599 8842 25651
rect 1926 25488 1978 25540
rect 2358 25488 2410 25540
rect 2838 25488 2890 25540
rect 3318 25488 3370 25540
rect 3798 25488 3850 25540
rect 4278 25488 4330 25540
rect 4758 25488 4810 25540
rect 5284 25488 5336 25540
rect 5766 25488 5818 25540
rect 6246 25488 6298 25540
rect 6774 25488 6826 25540
rect 7254 25488 7306 25540
rect 7734 25488 7786 25540
rect 8214 25488 8266 25540
rect 8694 25488 8746 25540
rect 9174 25488 9226 25540
rect 6270 24822 6322 24874
rect 6334 24822 6386 24874
rect 6398 24822 6450 24874
rect 6462 24822 6514 24874
rect 5785 24267 5837 24319
rect 1878 24156 1930 24208
rect 2406 24156 2458 24208
rect 2886 24156 2938 24208
rect 3366 24156 3418 24208
rect 3849 24156 3901 24208
rect 4333 24156 4385 24208
rect 4817 24156 4869 24208
rect 5301 24156 5353 24208
rect 5785 24156 5837 24208
rect 6269 24156 6321 24208
rect 6390 24193 6442 24245
rect 6774 24156 6826 24208
rect 7254 24156 7306 24208
rect 7734 24156 7786 24208
rect 8214 24156 8266 24208
rect 8694 24156 8746 24208
rect 9174 24156 9226 24208
rect 2022 24045 2074 24097
rect 6390 24082 6442 24134
rect 8310 24045 8362 24097
rect 9270 24045 9322 24097
rect 2502 23971 2554 24023
rect 2982 23971 3034 24023
rect 3462 23971 3514 24023
rect 3942 23971 3994 24023
rect 4422 23971 4474 24023
rect 4902 23971 4954 24023
rect 5382 23971 5434 24023
rect 7350 23971 7402 24023
rect 7830 23971 7882 24023
rect 8790 23971 8842 24023
rect 5910 23786 5962 23838
rect 6870 23786 6922 23838
rect 6294 23675 6346 23727
rect 6870 23675 6922 23727
rect 3606 23490 3658 23542
rect 3670 23490 3722 23542
rect 3734 23490 3786 23542
rect 3798 23490 3850 23542
rect 8934 23490 8986 23542
rect 8998 23490 9050 23542
rect 9062 23490 9114 23542
rect 9126 23490 9178 23542
rect 6390 23194 6442 23246
rect 9270 23157 9322 23209
rect 3942 23083 3994 23135
rect 5382 23083 5434 23135
rect 7830 23083 7882 23135
rect 2022 22935 2074 22987
rect 2502 22935 2554 22987
rect 2982 22935 3034 22987
rect 3462 22935 3514 22987
rect 4422 22935 4474 22987
rect 4902 22935 4954 22987
rect 5910 22898 5962 22950
rect 6870 22898 6922 22950
rect 7350 22935 7402 22987
rect 8310 22935 8362 22987
rect 8790 22935 8842 22987
rect 1878 22824 1930 22876
rect 2358 22824 2410 22876
rect 2838 22824 2890 22876
rect 3318 22824 3370 22876
rect 3798 22824 3850 22876
rect 4316 22824 4368 22876
rect 4758 22824 4810 22876
rect 5284 22824 5336 22876
rect 5766 22824 5818 22876
rect 6246 22824 6298 22876
rect 6774 22824 6826 22876
rect 7254 22824 7306 22876
rect 7734 22824 7786 22876
rect 8166 22824 8218 22876
rect 8694 22824 8746 22876
rect 9174 22824 9226 22876
rect 6270 22158 6322 22210
rect 6334 22158 6386 22210
rect 6398 22158 6450 22210
rect 6462 22158 6514 22210
rect 5286 21677 5338 21729
rect 5910 21677 5962 21729
rect 6269 21677 6321 21729
rect 6870 21677 6922 21729
rect 4758 21603 4810 21655
rect 5382 21603 5434 21655
rect 5785 21603 5837 21655
rect 6390 21603 6442 21655
rect 6774 21603 6826 21655
rect 7350 21603 7402 21655
rect 8694 21603 8746 21655
rect 9270 21603 9322 21655
rect 1110 21492 1162 21544
rect 1926 21492 1978 21544
rect 2406 21492 2458 21544
rect 2886 21492 2938 21544
rect 3366 21492 3418 21544
rect 3849 21492 3901 21544
rect 4333 21492 4385 21544
rect 4758 21492 4810 21544
rect 5286 21492 5338 21544
rect 5785 21492 5837 21544
rect 6269 21492 6321 21544
rect 6774 21492 6826 21544
rect 7254 21492 7306 21544
rect 7734 21492 7786 21544
rect 8214 21492 8266 21544
rect 8694 21492 8746 21544
rect 9174 21492 9226 21544
rect 1274 21418 1326 21470
rect 1452 21344 1504 21396
rect 2502 21381 2554 21433
rect 2982 21381 3034 21433
rect 3462 21381 3514 21433
rect 3942 21381 3994 21433
rect 4422 21381 4474 21433
rect 4902 21381 4954 21433
rect 5382 21381 5434 21433
rect 5910 21418 5962 21470
rect 6390 21418 6442 21470
rect 6870 21418 6922 21470
rect 7350 21381 7402 21433
rect 8310 21381 8362 21433
rect 8790 21381 8842 21433
rect 9270 21381 9322 21433
rect 1350 21270 1402 21322
rect 2022 21307 2074 21359
rect 7830 21233 7882 21285
rect 1302 21011 1354 21063
rect 1782 21011 1834 21063
rect 3606 20826 3658 20878
rect 3670 20826 3722 20878
rect 3734 20826 3786 20878
rect 3798 20826 3850 20878
rect 8934 20826 8986 20878
rect 8998 20826 9050 20878
rect 9062 20826 9114 20878
rect 9126 20826 9178 20878
rect 9270 20493 9322 20545
rect 2022 20271 2074 20323
rect 2502 20271 2554 20323
rect 2982 20271 3034 20323
rect 3462 20271 3514 20323
rect 3942 20271 3994 20323
rect 4422 20271 4474 20323
rect 4902 20271 4954 20323
rect 5382 20271 5434 20323
rect 5910 20234 5962 20286
rect 6390 20234 6442 20286
rect 6870 20234 6922 20286
rect 7350 20271 7402 20323
rect 7830 20271 7882 20323
rect 8310 20271 8362 20323
rect 8790 20271 8842 20323
rect 1878 20160 1930 20212
rect 2358 20160 2410 20212
rect 2838 20160 2890 20212
rect 3318 20160 3370 20212
rect 3798 20160 3850 20212
rect 4278 20160 4330 20212
rect 4758 20160 4810 20212
rect 5284 20160 5336 20212
rect 5766 20160 5818 20212
rect 6246 20160 6298 20212
rect 6774 20160 6826 20212
rect 7254 20160 7306 20212
rect 7734 20160 7786 20212
rect 8214 20160 8266 20212
rect 8694 20160 8746 20212
rect 9174 20160 9226 20212
rect 6270 19494 6322 19546
rect 6334 19494 6386 19546
rect 6398 19494 6450 19546
rect 6462 19494 6514 19546
rect 5286 19013 5338 19065
rect 5910 19013 5962 19065
rect 6269 19013 6321 19065
rect 6870 19013 6922 19065
rect 4758 18939 4810 18991
rect 5382 18939 5434 18991
rect 5785 18939 5837 18991
rect 6390 18939 6442 18991
rect 6774 18939 6826 18991
rect 7350 18939 7402 18991
rect 8694 18939 8746 18991
rect 9270 18939 9322 18991
rect 1878 18828 1930 18880
rect 2406 18828 2458 18880
rect 2886 18828 2938 18880
rect 3366 18828 3418 18880
rect 3849 18828 3901 18880
rect 4333 18828 4385 18880
rect 4758 18828 4810 18880
rect 5286 18828 5338 18880
rect 5785 18828 5837 18880
rect 6269 18828 6321 18880
rect 6774 18828 6826 18880
rect 7254 18828 7306 18880
rect 7734 18828 7786 18880
rect 8214 18828 8266 18880
rect 8694 18828 8746 18880
rect 9174 18828 9226 18880
rect 2022 18717 2074 18769
rect 2982 18717 3034 18769
rect 3462 18717 3514 18769
rect 3942 18717 3994 18769
rect 4422 18717 4474 18769
rect 4902 18717 4954 18769
rect 5382 18717 5434 18769
rect 5910 18754 5962 18806
rect 6390 18754 6442 18806
rect 6870 18754 6922 18806
rect 7350 18717 7402 18769
rect 8310 18717 8362 18769
rect 8790 18717 8842 18769
rect 9270 18717 9322 18769
rect 2502 18643 2554 18695
rect 7830 18569 7882 18621
rect 3606 18162 3658 18214
rect 3670 18162 3722 18214
rect 3734 18162 3786 18214
rect 3798 18162 3850 18214
rect 8934 18162 8986 18214
rect 8998 18162 9050 18214
rect 9062 18162 9114 18214
rect 9126 18162 9178 18214
rect 9270 17829 9322 17881
rect 2022 17607 2074 17659
rect 2502 17607 2554 17659
rect 2982 17607 3034 17659
rect 3462 17607 3514 17659
rect 3942 17607 3994 17659
rect 4422 17607 4474 17659
rect 4902 17607 4954 17659
rect 5382 17607 5434 17659
rect 5910 17570 5962 17622
rect 6390 17570 6442 17622
rect 6870 17570 6922 17622
rect 7350 17607 7402 17659
rect 7830 17607 7882 17659
rect 8310 17607 8362 17659
rect 8790 17607 8842 17659
rect 1878 17496 1930 17548
rect 2358 17496 2410 17548
rect 2838 17496 2890 17548
rect 3318 17496 3370 17548
rect 3798 17496 3850 17548
rect 4278 17496 4330 17548
rect 4758 17496 4810 17548
rect 5284 17496 5336 17548
rect 5766 17496 5818 17548
rect 6246 17496 6298 17548
rect 6774 17496 6826 17548
rect 7254 17496 7306 17548
rect 7734 17496 7786 17548
rect 8214 17496 8266 17548
rect 8694 17496 8746 17548
rect 9174 17496 9226 17548
rect 6270 16830 6322 16882
rect 6334 16830 6386 16882
rect 6398 16830 6450 16882
rect 6462 16830 6514 16882
rect 5286 16349 5338 16401
rect 5910 16349 5962 16401
rect 6269 16349 6321 16401
rect 6870 16349 6922 16401
rect 4758 16275 4810 16327
rect 5382 16275 5434 16327
rect 5785 16275 5837 16327
rect 6390 16275 6442 16327
rect 6774 16275 6826 16327
rect 7350 16275 7402 16327
rect 8694 16275 8746 16327
rect 9270 16275 9322 16327
rect 1878 16164 1930 16216
rect 2406 16164 2458 16216
rect 2886 16164 2938 16216
rect 3366 16164 3418 16216
rect 3849 16164 3901 16216
rect 4333 16164 4385 16216
rect 4758 16164 4810 16216
rect 5286 16164 5338 16216
rect 5785 16164 5837 16216
rect 6269 16164 6321 16216
rect 6774 16164 6826 16216
rect 7254 16164 7306 16216
rect 7734 16164 7786 16216
rect 8214 16164 8266 16216
rect 8694 16164 8746 16216
rect 9174 16164 9226 16216
rect 2022 16053 2074 16105
rect 2982 16053 3034 16105
rect 3462 16053 3514 16105
rect 3942 16053 3994 16105
rect 4422 16053 4474 16105
rect 4902 16053 4954 16105
rect 5382 16053 5434 16105
rect 5910 16090 5962 16142
rect 6390 16090 6442 16142
rect 6870 16090 6922 16142
rect 7350 16053 7402 16105
rect 9270 16053 9322 16105
rect 2502 15979 2554 16031
rect 7830 15979 7882 16031
rect 8310 15979 8362 16031
rect 8790 15979 8842 16031
rect 3606 15498 3658 15550
rect 3670 15498 3722 15550
rect 3734 15498 3786 15550
rect 3798 15498 3850 15550
rect 8934 15498 8986 15550
rect 8998 15498 9050 15550
rect 9062 15498 9114 15550
rect 9126 15498 9178 15550
rect 9270 15165 9322 15217
rect 2022 14943 2074 14995
rect 2502 14943 2554 14995
rect 2982 14943 3034 14995
rect 3462 14943 3514 14995
rect 3942 14943 3994 14995
rect 4422 14943 4474 14995
rect 4902 14943 4954 14995
rect 5382 14943 5434 14995
rect 5910 14906 5962 14958
rect 6390 14906 6442 14958
rect 6870 14906 6922 14958
rect 7350 14943 7402 14995
rect 7830 14943 7882 14995
rect 8310 14943 8362 14995
rect 8790 14943 8842 14995
rect 1926 14832 1978 14884
rect 2358 14832 2410 14884
rect 2838 14832 2890 14884
rect 3318 14832 3370 14884
rect 3798 14832 3850 14884
rect 4278 14832 4330 14884
rect 4758 14832 4810 14884
rect 5284 14832 5336 14884
rect 5766 14832 5818 14884
rect 6246 14832 6298 14884
rect 6726 14832 6778 14884
rect 7206 14832 7258 14884
rect 7686 14832 7738 14884
rect 8166 14832 8218 14884
rect 8646 14832 8698 14884
rect 9126 14832 9178 14884
rect 6270 14166 6322 14218
rect 6334 14166 6386 14218
rect 6398 14166 6450 14218
rect 6462 14166 6514 14218
rect 5785 13611 5837 13663
rect 1878 13500 1930 13552
rect 2406 13500 2458 13552
rect 2886 13500 2938 13552
rect 3366 13500 3418 13552
rect 3849 13500 3901 13552
rect 4333 13500 4385 13552
rect 4817 13500 4869 13552
rect 5301 13500 5353 13552
rect 5785 13500 5837 13552
rect 6269 13500 6321 13552
rect 6390 13537 6442 13589
rect 6774 13500 6826 13552
rect 7254 13500 7306 13552
rect 7734 13500 7786 13552
rect 8214 13500 8266 13552
rect 8694 13500 8746 13552
rect 9174 13500 9226 13552
rect 2022 13389 2074 13441
rect 6390 13426 6442 13478
rect 9270 13389 9322 13441
rect 2502 13315 2554 13367
rect 2982 13315 3034 13367
rect 3462 13315 3514 13367
rect 3942 13315 3994 13367
rect 4422 13315 4474 13367
rect 4902 13315 4954 13367
rect 5382 13315 5434 13367
rect 7350 13315 7402 13367
rect 7830 13315 7882 13367
rect 8310 13315 8362 13367
rect 8790 13315 8842 13367
rect 5910 13130 5962 13182
rect 6870 13130 6922 13182
rect 6294 13019 6346 13071
rect 6870 13019 6922 13071
rect 3606 12834 3658 12886
rect 3670 12834 3722 12886
rect 3734 12834 3786 12886
rect 3798 12834 3850 12886
rect 8934 12834 8986 12886
rect 8998 12834 9050 12886
rect 9062 12834 9114 12886
rect 9126 12834 9178 12886
rect 3942 12501 3994 12553
rect 5382 12501 5434 12553
rect 6390 12538 6442 12590
rect 9270 12501 9322 12553
rect 2022 12279 2074 12331
rect 2502 12279 2554 12331
rect 2982 12279 3034 12331
rect 3462 12279 3514 12331
rect 4422 12279 4474 12331
rect 4902 12279 4954 12331
rect 5910 12242 5962 12294
rect 6870 12242 6922 12294
rect 7350 12279 7402 12331
rect 7830 12279 7882 12331
rect 8310 12279 8362 12331
rect 8790 12279 8842 12331
rect 1878 12168 1930 12220
rect 2358 12168 2410 12220
rect 2838 12168 2890 12220
rect 3318 12168 3370 12220
rect 3798 12168 3850 12220
rect 4278 12168 4330 12220
rect 4758 12168 4810 12220
rect 5284 12168 5336 12220
rect 5768 12168 5820 12220
rect 6246 12168 6298 12220
rect 6774 12168 6826 12220
rect 7206 12168 7258 12220
rect 7686 12168 7738 12220
rect 8166 12168 8218 12220
rect 8646 12168 8698 12220
rect 9126 12168 9178 12220
rect 6270 11502 6322 11554
rect 6334 11502 6386 11554
rect 6398 11502 6450 11554
rect 6462 11502 6514 11554
rect 5286 11021 5338 11073
rect 5910 11021 5962 11073
rect 6269 11021 6321 11073
rect 6870 11021 6922 11073
rect 4758 10947 4810 10999
rect 5382 10947 5434 10999
rect 5785 10947 5837 10999
rect 6390 10947 6442 10999
rect 6774 10947 6826 10999
rect 7350 10947 7402 10999
rect 8694 10947 8746 10999
rect 9270 10947 9322 10999
rect 1878 10836 1930 10888
rect 2406 10836 2458 10888
rect 2886 10836 2938 10888
rect 3366 10836 3418 10888
rect 3849 10836 3901 10888
rect 4333 10836 4385 10888
rect 4758 10836 4810 10888
rect 5286 10836 5338 10888
rect 5785 10836 5837 10888
rect 6269 10836 6321 10888
rect 6774 10836 6826 10888
rect 7254 10836 7306 10888
rect 7734 10836 7786 10888
rect 8214 10836 8266 10888
rect 8694 10836 8746 10888
rect 9174 10836 9226 10888
rect 2022 10725 2074 10777
rect 2982 10725 3034 10777
rect 3462 10725 3514 10777
rect 3942 10725 3994 10777
rect 4422 10725 4474 10777
rect 4902 10725 4954 10777
rect 5382 10725 5434 10777
rect 5910 10762 5962 10814
rect 6390 10762 6442 10814
rect 6870 10762 6922 10814
rect 7350 10725 7402 10777
rect 9270 10725 9322 10777
rect 2502 10651 2554 10703
rect 8310 10651 8362 10703
rect 8790 10651 8842 10703
rect 7830 10577 7882 10629
rect 3606 10170 3658 10222
rect 3670 10170 3722 10222
rect 3734 10170 3786 10222
rect 3798 10170 3850 10222
rect 8934 10170 8986 10222
rect 8998 10170 9050 10222
rect 9062 10170 9114 10222
rect 9126 10170 9178 10222
rect 9270 9837 9322 9889
rect 2022 9615 2074 9667
rect 2502 9615 2554 9667
rect 2982 9615 3034 9667
rect 3462 9615 3514 9667
rect 3942 9615 3994 9667
rect 4422 9615 4474 9667
rect 4902 9615 4954 9667
rect 5382 9615 5434 9667
rect 5910 9578 5962 9630
rect 6390 9578 6442 9630
rect 6870 9578 6922 9630
rect 7350 9615 7402 9667
rect 7830 9615 7882 9667
rect 8310 9615 8362 9667
rect 8790 9615 8842 9667
rect 1878 9504 1930 9556
rect 2358 9504 2410 9556
rect 2838 9504 2890 9556
rect 3318 9504 3370 9556
rect 3798 9504 3850 9556
rect 4278 9504 4330 9556
rect 4758 9504 4810 9556
rect 5284 9504 5336 9556
rect 5766 9504 5818 9556
rect 6246 9504 6298 9556
rect 6726 9504 6778 9556
rect 7206 9504 7258 9556
rect 7686 9504 7738 9556
rect 8166 9504 8218 9556
rect 8646 9504 8698 9556
rect 9126 9504 9178 9556
rect 6270 8838 6322 8890
rect 6334 8838 6386 8890
rect 6398 8838 6450 8890
rect 6462 8838 6514 8890
rect 5286 8357 5338 8409
rect 5910 8357 5962 8409
rect 6269 8357 6321 8409
rect 6870 8357 6922 8409
rect 4758 8283 4810 8335
rect 5382 8283 5434 8335
rect 5785 8283 5837 8335
rect 6390 8283 6442 8335
rect 6774 8283 6826 8335
rect 7350 8283 7402 8335
rect 8694 8283 8746 8335
rect 9270 8283 9322 8335
rect 1878 8172 1930 8224
rect 2406 8172 2458 8224
rect 2886 8172 2938 8224
rect 3366 8172 3418 8224
rect 3849 8172 3901 8224
rect 4333 8172 4385 8224
rect 4758 8172 4810 8224
rect 5286 8172 5338 8224
rect 5785 8172 5837 8224
rect 6269 8172 6321 8224
rect 6774 8172 6826 8224
rect 7254 8172 7306 8224
rect 7734 8172 7786 8224
rect 8214 8172 8266 8224
rect 8694 8172 8746 8224
rect 9174 8172 9226 8224
rect 2022 8061 2074 8113
rect 2982 8061 3034 8113
rect 3462 8061 3514 8113
rect 3942 8061 3994 8113
rect 4422 8061 4474 8113
rect 4902 8061 4954 8113
rect 5382 8061 5434 8113
rect 5910 8098 5962 8150
rect 6390 8098 6442 8150
rect 6870 8098 6922 8150
rect 7350 8061 7402 8113
rect 9270 8061 9322 8113
rect 2502 7987 2554 8039
rect 8310 7987 8362 8039
rect 8790 7987 8842 8039
rect 7830 7913 7882 7965
rect 3606 7506 3658 7558
rect 3670 7506 3722 7558
rect 3734 7506 3786 7558
rect 3798 7506 3850 7558
rect 8934 7506 8986 7558
rect 8998 7506 9050 7558
rect 9062 7506 9114 7558
rect 9126 7506 9178 7558
rect 9270 7173 9322 7225
rect 2022 6951 2074 7003
rect 2502 6951 2554 7003
rect 2982 6951 3034 7003
rect 3462 6951 3514 7003
rect 3942 6951 3994 7003
rect 4422 6951 4474 7003
rect 4902 6951 4954 7003
rect 5382 6951 5434 7003
rect 5910 6914 5962 6966
rect 6390 6914 6442 6966
rect 6870 6914 6922 6966
rect 7350 6951 7402 7003
rect 7830 6951 7882 7003
rect 8310 6951 8362 7003
rect 8790 6951 8842 7003
rect 1878 6840 1930 6892
rect 2358 6840 2410 6892
rect 2838 6840 2890 6892
rect 3318 6840 3370 6892
rect 3798 6840 3850 6892
rect 4278 6840 4330 6892
rect 4758 6840 4810 6892
rect 5284 6840 5336 6892
rect 5766 6840 5818 6892
rect 6246 6840 6298 6892
rect 6726 6840 6778 6892
rect 7206 6840 7258 6892
rect 7686 6840 7738 6892
rect 8166 6840 8218 6892
rect 8646 6840 8698 6892
rect 9126 6840 9178 6892
rect 6270 6174 6322 6226
rect 6334 6174 6386 6226
rect 6398 6174 6450 6226
rect 6462 6174 6514 6226
rect 5286 5693 5338 5745
rect 5910 5693 5962 5745
rect 6269 5693 6321 5745
rect 6870 5693 6922 5745
rect 4758 5619 4810 5671
rect 5382 5619 5434 5671
rect 5785 5619 5837 5671
rect 6390 5619 6442 5671
rect 6774 5619 6826 5671
rect 7350 5619 7402 5671
rect 8694 5619 8746 5671
rect 9270 5619 9322 5671
rect 1878 5508 1930 5560
rect 2406 5508 2458 5560
rect 2886 5508 2938 5560
rect 3366 5508 3418 5560
rect 3849 5508 3901 5560
rect 4333 5508 4385 5560
rect 4758 5508 4810 5560
rect 5286 5508 5338 5560
rect 5785 5508 5837 5560
rect 6269 5508 6321 5560
rect 6774 5508 6826 5560
rect 7254 5508 7306 5560
rect 7734 5508 7786 5560
rect 8214 5508 8266 5560
rect 8694 5508 8746 5560
rect 9174 5508 9226 5560
rect 2022 5397 2074 5449
rect 2982 5397 3034 5449
rect 3462 5397 3514 5449
rect 3942 5397 3994 5449
rect 4422 5397 4474 5449
rect 4902 5397 4954 5449
rect 5382 5397 5434 5449
rect 5910 5434 5962 5486
rect 6390 5434 6442 5486
rect 6870 5434 6922 5486
rect 7350 5397 7402 5449
rect 9270 5397 9322 5449
rect 2502 5323 2554 5375
rect 7830 5323 7882 5375
rect 8310 5323 8362 5375
rect 8790 5323 8842 5375
rect 3606 4842 3658 4894
rect 3670 4842 3722 4894
rect 3734 4842 3786 4894
rect 3798 4842 3850 4894
rect 8934 4842 8986 4894
rect 8998 4842 9050 4894
rect 9062 4842 9114 4894
rect 9126 4842 9178 4894
rect 9270 4509 9322 4561
rect 2022 4287 2074 4339
rect 2502 4287 2554 4339
rect 2982 4287 3034 4339
rect 3462 4287 3514 4339
rect 3942 4287 3994 4339
rect 4422 4287 4474 4339
rect 4902 4287 4954 4339
rect 5382 4287 5434 4339
rect 5910 4250 5962 4302
rect 6390 4250 6442 4302
rect 6870 4250 6922 4302
rect 7350 4287 7402 4339
rect 7830 4287 7882 4339
rect 8310 4287 8362 4339
rect 8790 4287 8842 4339
rect 1878 4176 1930 4228
rect 2358 4176 2410 4228
rect 2838 4176 2890 4228
rect 3318 4176 3370 4228
rect 3798 4176 3850 4228
rect 4278 4176 4330 4228
rect 4758 4176 4810 4228
rect 5284 4176 5336 4228
rect 5766 4176 5818 4228
rect 6246 4176 6298 4228
rect 6726 4176 6778 4228
rect 7206 4176 7258 4228
rect 7686 4176 7738 4228
rect 8166 4176 8218 4228
rect 8646 4176 8698 4228
rect 9126 4176 9178 4228
rect 6270 3510 6322 3562
rect 6334 3510 6386 3562
rect 6398 3510 6450 3562
rect 6462 3510 6514 3562
rect 5785 2955 5837 3007
rect 1878 2844 1930 2896
rect 2406 2844 2458 2896
rect 2886 2844 2938 2896
rect 3366 2844 3418 2896
rect 3849 2844 3901 2896
rect 4333 2844 4385 2896
rect 4817 2844 4869 2896
rect 5301 2844 5353 2896
rect 5785 2844 5837 2896
rect 6269 2844 6321 2896
rect 6390 2881 6442 2933
rect 6774 2844 6826 2896
rect 7254 2844 7306 2896
rect 7734 2844 7786 2896
rect 8214 2844 8266 2896
rect 8694 2844 8746 2896
rect 9174 2844 9226 2896
rect 2022 2733 2074 2785
rect 6390 2770 6442 2822
rect 7350 2733 7402 2785
rect 7830 2733 7882 2785
rect 8310 2733 8362 2785
rect 8790 2733 8842 2785
rect 9270 2733 9322 2785
rect 2502 2659 2554 2711
rect 2982 2659 3034 2711
rect 3462 2659 3514 2711
rect 3942 2659 3994 2711
rect 4422 2659 4474 2711
rect 4902 2659 4954 2711
rect 5382 2659 5434 2711
rect 5910 2474 5962 2526
rect 6870 2474 6922 2526
rect 6294 2363 6346 2415
rect 6870 2363 6922 2415
rect 3606 2178 3658 2230
rect 3670 2178 3722 2230
rect 3734 2178 3786 2230
rect 3798 2178 3850 2230
rect 8934 2178 8986 2230
rect 8998 2178 9050 2230
rect 9062 2178 9114 2230
rect 9126 2178 9178 2230
rect 6390 1882 6442 1934
rect 9270 1845 9322 1897
rect 3942 1771 3994 1823
rect 5382 1771 5434 1823
rect 2022 1623 2074 1675
rect 2502 1623 2554 1675
rect 2982 1623 3034 1675
rect 3462 1623 3514 1675
rect 4422 1623 4474 1675
rect 4902 1623 4954 1675
rect 5910 1586 5962 1638
rect 6870 1586 6922 1638
rect 7350 1623 7402 1675
rect 7830 1623 7882 1675
rect 8310 1623 8362 1675
rect 8790 1623 8842 1675
rect 1878 1512 1930 1564
rect 2358 1512 2410 1564
rect 2838 1512 2890 1564
rect 3318 1512 3370 1564
rect 3798 1512 3850 1564
rect 4333 1512 4385 1564
rect 4758 1512 4810 1564
rect 5284 1512 5336 1564
rect 5766 1512 5818 1564
rect 6246 1512 6298 1564
rect 6774 1512 6826 1564
rect 7206 1512 7258 1564
rect 7686 1512 7738 1564
rect 8166 1512 8218 1564
rect 8646 1512 8698 1564
rect 9126 1512 9178 1564
rect 6270 846 6322 898
rect 6334 846 6386 898
rect 6398 846 6450 898
rect 6462 846 6514 898
<< metal2 >>
rect 3580 52848 3876 52868
rect 3636 52846 3660 52848
rect 3716 52846 3740 52848
rect 3796 52846 3820 52848
rect 3658 52794 3660 52846
rect 3722 52794 3734 52846
rect 3796 52794 3798 52846
rect 3636 52792 3660 52794
rect 3716 52792 3740 52794
rect 3796 52792 3820 52794
rect 3580 52772 3876 52792
rect 8908 52848 9204 52868
rect 8964 52846 8988 52848
rect 9044 52846 9068 52848
rect 9124 52846 9148 52848
rect 8986 52794 8988 52846
rect 9050 52794 9062 52846
rect 9124 52794 9126 52846
rect 8964 52792 8988 52794
rect 9044 52792 9068 52794
rect 9124 52792 9148 52794
rect 8908 52772 9204 52792
rect 1350 52513 1402 52519
rect 1348 52478 1350 52487
rect 1402 52478 1404 52487
rect 1348 52413 1404 52422
rect 1452 52328 1504 52334
rect 1504 52297 2062 52316
rect 1504 52291 2074 52297
rect 1504 52288 2022 52291
rect 1452 52270 1504 52276
rect 1302 52254 1354 52260
rect 2022 52233 2074 52239
rect 1302 52196 1354 52202
rect 1110 52180 1162 52186
rect 1110 52122 1162 52128
rect 1122 52043 1150 52122
rect 1314 52075 1342 52196
rect 1878 52180 1930 52186
rect 1878 52122 1930 52128
rect 1890 52075 1918 52122
rect 1302 52069 1354 52075
rect 1108 52034 1164 52043
rect 1302 52011 1354 52017
rect 1878 52069 1930 52075
rect 1878 52011 1930 52017
rect 1108 51969 1164 51978
rect 1314 51576 1342 52011
rect 1218 51548 1342 51576
rect 1110 50848 1162 50854
rect 1110 50790 1162 50796
rect 1122 50711 1150 50790
rect 1108 50702 1164 50711
rect 1218 50688 1246 51548
rect 6244 51516 6540 51536
rect 6300 51514 6324 51516
rect 6380 51514 6404 51516
rect 6460 51514 6484 51516
rect 6322 51462 6324 51514
rect 6386 51462 6398 51514
rect 6460 51462 6462 51514
rect 6300 51460 6324 51462
rect 6380 51460 6404 51462
rect 6460 51460 6484 51462
rect 6244 51440 6540 51460
rect 1926 50848 1978 50854
rect 1314 50817 1438 50836
rect 1314 50811 1450 50817
rect 1314 50808 1398 50811
rect 1314 50780 1342 50808
rect 1302 50774 1354 50780
rect 1978 50808 2206 50836
rect 1926 50790 1978 50796
rect 1398 50753 1450 50759
rect 1302 50716 1354 50722
rect 1452 50700 1504 50706
rect 1218 50660 1390 50688
rect 1108 50637 1164 50646
rect 1362 50632 1390 50660
rect 1504 50669 2062 50688
rect 1504 50663 2074 50669
rect 1504 50660 2022 50663
rect 1452 50642 1504 50648
rect 1350 50626 1402 50632
rect 2022 50605 2074 50611
rect 1350 50568 1402 50574
rect 1782 50589 1834 50595
rect 1782 50531 1834 50537
rect 1794 49504 1822 50531
rect 2178 50174 2206 50808
rect 2034 50146 2206 50174
rect 3580 50184 3876 50204
rect 3636 50182 3660 50184
rect 3716 50182 3740 50184
rect 3796 50182 3820 50184
rect 2034 49855 2062 50146
rect 3658 50130 3660 50182
rect 3722 50130 3734 50182
rect 3796 50130 3798 50182
rect 3636 50128 3660 50130
rect 3716 50128 3740 50130
rect 3796 50128 3820 50130
rect 3580 50108 3876 50128
rect 8908 50184 9204 50204
rect 8964 50182 8988 50184
rect 9044 50182 9068 50184
rect 9124 50182 9148 50184
rect 8986 50130 8988 50182
rect 9050 50130 9062 50182
rect 9124 50130 9126 50182
rect 8964 50128 8988 50130
rect 9044 50128 9068 50130
rect 9124 50128 9148 50130
rect 8908 50108 9204 50128
rect 2022 49849 2074 49855
rect 2022 49791 2074 49797
rect 1878 49516 1930 49522
rect 1794 49476 1878 49504
rect 1110 48184 1162 48190
rect 1794 48153 1822 49476
rect 1878 49458 1930 49464
rect 6244 48852 6540 48872
rect 6300 48850 6324 48852
rect 6380 48850 6404 48852
rect 6460 48850 6484 48852
rect 6322 48798 6324 48850
rect 6386 48798 6398 48850
rect 6460 48798 6462 48850
rect 6300 48796 6324 48798
rect 6380 48796 6404 48798
rect 6460 48796 6484 48798
rect 6244 48776 6540 48796
rect 1878 48295 1930 48301
rect 1878 48237 1930 48243
rect 2502 48295 2554 48301
rect 2502 48237 2554 48243
rect 1890 48190 1918 48237
rect 1878 48184 1930 48190
rect 1110 48126 1162 48132
rect 1782 48147 1834 48153
rect 1122 48047 1150 48126
rect 1302 48110 1354 48116
rect 1878 48126 1930 48132
rect 2358 48184 2410 48190
rect 2358 48126 2410 48132
rect 1782 48089 1834 48095
rect 1302 48052 1354 48058
rect 1108 48038 1164 48047
rect 1314 48024 1342 48052
rect 1108 47973 1164 47982
rect 1218 47996 1342 48024
rect 1452 48036 1504 48042
rect 1218 46821 1246 47996
rect 1504 48005 2062 48024
rect 1504 47999 2074 48005
rect 1504 47996 2022 47999
rect 1452 47978 1504 47984
rect 2022 47941 2074 47947
rect 1494 47925 1546 47931
rect 1362 47873 1494 47876
rect 1362 47867 1546 47873
rect 1362 47857 1534 47867
rect 1350 47851 1534 47857
rect 1402 47848 1534 47851
rect 1350 47793 1402 47799
rect 2370 47454 2398 48126
rect 2514 48079 2542 48237
rect 2502 48073 2554 48079
rect 2502 48015 2554 48021
rect 3580 47520 3876 47540
rect 3636 47518 3660 47520
rect 3716 47518 3740 47520
rect 3796 47518 3820 47520
rect 3658 47466 3660 47518
rect 3722 47466 3734 47518
rect 3796 47466 3798 47518
rect 3636 47464 3660 47466
rect 3716 47464 3740 47466
rect 3796 47464 3820 47466
rect 2370 47426 2542 47454
rect 3580 47444 3876 47464
rect 8908 47520 9204 47540
rect 8964 47518 8988 47520
rect 9044 47518 9068 47520
rect 9124 47518 9148 47520
rect 8986 47466 8988 47518
rect 9050 47466 9062 47518
rect 9124 47466 9126 47518
rect 8964 47464 8988 47466
rect 9044 47464 9068 47466
rect 9124 47464 9148 47466
rect 8908 47444 9204 47464
rect 2514 47191 2542 47426
rect 2502 47185 2554 47191
rect 2502 47127 2554 47133
rect 2022 46963 2074 46969
rect 2022 46905 2074 46911
rect 1878 46852 1930 46858
rect 1794 46821 1878 46840
rect 1206 46815 1258 46821
rect 1206 46757 1258 46763
rect 1782 46815 1878 46821
rect 1834 46812 1878 46815
rect 2034 46840 2062 46905
rect 2358 46852 2410 46858
rect 2034 46812 2358 46840
rect 1878 46794 1930 46800
rect 2358 46794 2410 46800
rect 1782 46757 1834 46763
rect 1110 45520 1162 45526
rect 1110 45462 1162 45468
rect 1122 45383 1150 45462
rect 1108 45374 1164 45383
rect 1218 45360 1246 46757
rect 6244 46188 6540 46208
rect 6300 46186 6324 46188
rect 6380 46186 6404 46188
rect 6460 46186 6484 46188
rect 6322 46134 6324 46186
rect 6386 46134 6398 46186
rect 6460 46134 6462 46186
rect 6300 46132 6324 46134
rect 6380 46132 6404 46134
rect 6460 46132 6484 46134
rect 6244 46112 6540 46132
rect 1926 45520 1978 45526
rect 1314 45489 1438 45508
rect 1314 45483 1450 45489
rect 1314 45480 1398 45483
rect 1314 45452 1342 45480
rect 1302 45446 1354 45452
rect 2406 45520 2458 45526
rect 1978 45480 2302 45508
rect 1926 45462 1978 45468
rect 1398 45425 1450 45431
rect 1302 45388 1354 45394
rect 1452 45372 1504 45378
rect 1218 45332 1390 45360
rect 1108 45309 1164 45318
rect 1362 45304 1390 45332
rect 2274 45360 2302 45480
rect 2836 45522 2892 45531
rect 2458 45480 2782 45508
rect 2406 45462 2458 45468
rect 2754 45360 2782 45480
rect 2836 45457 2892 45466
rect 3318 45520 3370 45526
rect 3318 45462 3370 45468
rect 3460 45522 3516 45531
rect 1504 45341 2062 45360
rect 2274 45341 2542 45360
rect 2754 45341 3022 45360
rect 1504 45335 2074 45341
rect 1504 45332 2022 45335
rect 1452 45314 1504 45320
rect 1350 45298 1402 45304
rect 2274 45335 2554 45341
rect 2274 45332 2502 45335
rect 2022 45277 2074 45283
rect 2754 45335 3034 45341
rect 2754 45332 2982 45335
rect 2502 45277 2554 45283
rect 2982 45277 3034 45283
rect 1350 45240 1402 45246
rect 1782 45261 1834 45267
rect 1782 45203 1834 45209
rect 1794 44176 1822 45203
rect 3330 44768 3358 45462
rect 3460 45457 3516 45466
rect 3474 45415 3502 45457
rect 3462 45409 3514 45415
rect 3462 45351 3514 45357
rect 3580 44856 3876 44876
rect 3636 44854 3660 44856
rect 3716 44854 3740 44856
rect 3796 44854 3820 44856
rect 3658 44802 3660 44854
rect 3722 44802 3734 44854
rect 3796 44802 3798 44854
rect 3636 44800 3660 44802
rect 3716 44800 3740 44802
rect 3796 44800 3820 44802
rect 3580 44780 3876 44800
rect 8908 44856 9204 44876
rect 8964 44854 8988 44856
rect 9044 44854 9068 44856
rect 9124 44854 9148 44856
rect 8986 44802 8988 44854
rect 9050 44802 9062 44854
rect 9124 44802 9126 44854
rect 8964 44800 8988 44802
rect 9044 44800 9068 44802
rect 9124 44800 9148 44802
rect 8908 44780 9204 44800
rect 3330 44740 3502 44768
rect 3474 44527 3502 44740
rect 3462 44521 3514 44527
rect 2994 44453 3358 44472
rect 3462 44463 3514 44469
rect 2982 44447 3358 44453
rect 3034 44444 3358 44447
rect 2982 44389 3034 44395
rect 2022 44299 2074 44305
rect 2022 44241 2074 44247
rect 2502 44299 2554 44305
rect 2502 44241 2554 44247
rect 1878 44188 1930 44194
rect 1794 44148 1878 44176
rect 1110 42856 1162 42862
rect 1794 42825 1822 44148
rect 2034 44176 2062 44241
rect 2358 44188 2410 44194
rect 2034 44148 2358 44176
rect 1878 44130 1930 44136
rect 2514 44176 2542 44241
rect 3330 44194 3358 44444
rect 2838 44188 2890 44194
rect 2514 44148 2838 44176
rect 2358 44130 2410 44136
rect 2838 44130 2890 44136
rect 3318 44188 3370 44194
rect 3318 44130 3370 44136
rect 6244 43524 6540 43544
rect 6300 43522 6324 43524
rect 6380 43522 6404 43524
rect 6460 43522 6484 43524
rect 6322 43470 6324 43522
rect 6386 43470 6398 43522
rect 6460 43470 6462 43522
rect 6300 43468 6324 43470
rect 6380 43468 6404 43470
rect 6460 43468 6484 43470
rect 6244 43448 6540 43468
rect 4758 42967 4810 42973
rect 4758 42909 4810 42915
rect 5382 42967 5434 42973
rect 5382 42909 5434 42915
rect 4770 42862 4798 42909
rect 1926 42856 1978 42862
rect 1110 42798 1162 42804
rect 1782 42819 1834 42825
rect 1122 42719 1150 42798
rect 1302 42782 1354 42788
rect 2406 42856 2458 42862
rect 1978 42816 2302 42844
rect 1926 42798 1978 42804
rect 1782 42761 1834 42767
rect 1302 42724 1354 42730
rect 1108 42710 1164 42719
rect 1314 42696 1342 42724
rect 1108 42645 1164 42654
rect 1218 42668 1342 42696
rect 1452 42708 1504 42714
rect 1218 42381 1246 42668
rect 2274 42696 2302 42816
rect 2886 42856 2938 42862
rect 2458 42816 2782 42844
rect 2406 42798 2458 42804
rect 2754 42696 2782 42816
rect 3366 42856 3418 42862
rect 2938 42816 3262 42844
rect 2886 42798 2938 42804
rect 3234 42696 3262 42816
rect 3849 42856 3901 42862
rect 3418 42816 3742 42844
rect 3366 42798 3418 42804
rect 3714 42696 3742 42816
rect 4333 42856 4385 42862
rect 3901 42816 4222 42844
rect 3849 42798 3901 42804
rect 4194 42696 4222 42816
rect 4758 42856 4810 42862
rect 4385 42816 4702 42844
rect 4333 42798 4385 42804
rect 4674 42696 4702 42816
rect 4758 42798 4810 42804
rect 5301 42856 5353 42862
rect 5301 42798 5353 42804
rect 1504 42677 2062 42696
rect 2274 42677 2542 42696
rect 2754 42677 3022 42696
rect 3234 42677 3502 42696
rect 3714 42677 3982 42696
rect 4194 42677 4462 42696
rect 4674 42677 4942 42696
rect 1504 42671 2074 42677
rect 1504 42668 2022 42671
rect 1452 42650 1504 42656
rect 2274 42671 2554 42677
rect 2274 42668 2502 42671
rect 2022 42613 2074 42619
rect 2754 42671 3034 42677
rect 2754 42668 2982 42671
rect 2502 42613 2554 42619
rect 3234 42671 3514 42677
rect 3234 42668 3462 42671
rect 2982 42613 3034 42619
rect 3714 42671 3994 42677
rect 3714 42668 3942 42671
rect 3462 42613 3514 42619
rect 4194 42671 4474 42677
rect 4194 42668 4422 42671
rect 3942 42613 3994 42619
rect 4674 42671 4954 42677
rect 4674 42668 4902 42671
rect 4422 42613 4474 42619
rect 4902 42613 4954 42619
rect 1494 42597 1546 42603
rect 1362 42545 1494 42548
rect 1362 42539 1546 42545
rect 1362 42529 1534 42539
rect 1350 42523 1534 42529
rect 1402 42520 1534 42523
rect 1350 42465 1402 42471
rect 5313 42400 5341 42798
rect 5394 42751 5422 42909
rect 5382 42745 5434 42751
rect 5382 42687 5434 42693
rect 1206 42375 1258 42381
rect 1206 42317 1258 42323
rect 1782 42375 1834 42381
rect 5313 42372 5374 42400
rect 1782 42317 1834 42323
rect 1794 41512 1822 42317
rect 3580 42192 3876 42212
rect 3636 42190 3660 42192
rect 3716 42190 3740 42192
rect 3796 42190 3820 42192
rect 3658 42138 3660 42190
rect 3722 42138 3734 42190
rect 3796 42138 3798 42190
rect 3636 42136 3660 42138
rect 3716 42136 3740 42138
rect 3796 42136 3820 42138
rect 3580 42116 3876 42136
rect 5346 42150 5374 42372
rect 8908 42192 9204 42212
rect 8964 42190 8988 42192
rect 9044 42190 9068 42192
rect 9124 42190 9148 42192
rect 5346 42122 5422 42150
rect 5394 41863 5422 42122
rect 8986 42138 8988 42190
rect 9050 42138 9062 42190
rect 9124 42138 9126 42190
rect 8964 42136 8988 42138
rect 9044 42136 9068 42138
rect 9124 42136 9148 42138
rect 8908 42116 9204 42136
rect 5382 41857 5434 41863
rect 5382 41799 5434 41805
rect 2022 41635 2074 41641
rect 2022 41577 2074 41583
rect 2502 41635 2554 41641
rect 2502 41577 2554 41583
rect 2982 41635 3034 41641
rect 2982 41577 3034 41583
rect 3462 41635 3514 41641
rect 3462 41577 3514 41583
rect 3942 41635 3994 41641
rect 3942 41577 3994 41583
rect 4422 41635 4474 41641
rect 4422 41577 4474 41583
rect 4902 41635 4954 41641
rect 4902 41577 4954 41583
rect 1878 41524 1930 41530
rect 1794 41484 1878 41512
rect 1108 40194 1164 40203
rect 1794 40180 1822 41484
rect 2034 41512 2062 41577
rect 2358 41524 2410 41530
rect 2034 41484 2358 41512
rect 1878 41466 1930 41472
rect 2514 41512 2542 41577
rect 2838 41524 2890 41530
rect 2514 41484 2838 41512
rect 2358 41466 2410 41472
rect 2994 41512 3022 41577
rect 3318 41524 3370 41530
rect 2994 41484 3318 41512
rect 2838 41466 2890 41472
rect 3474 41512 3502 41577
rect 3798 41524 3850 41530
rect 3474 41484 3798 41512
rect 3318 41466 3370 41472
rect 3954 41512 3982 41577
rect 4278 41524 4330 41530
rect 3954 41484 4278 41512
rect 3798 41466 3850 41472
rect 4434 41512 4462 41577
rect 4758 41524 4810 41530
rect 4434 41484 4758 41512
rect 4278 41466 4330 41472
rect 4914 41512 4942 41577
rect 5284 41524 5336 41530
rect 4914 41484 5284 41512
rect 4758 41466 4810 41472
rect 5284 41466 5336 41472
rect 6244 40860 6540 40880
rect 6300 40858 6324 40860
rect 6380 40858 6404 40860
rect 6460 40858 6484 40860
rect 6322 40806 6324 40858
rect 6386 40806 6398 40858
rect 6460 40806 6462 40858
rect 6300 40804 6324 40806
rect 6380 40804 6404 40806
rect 6460 40804 6484 40806
rect 6244 40784 6540 40804
rect 5286 40377 5338 40383
rect 5286 40319 5338 40325
rect 5910 40377 5962 40383
rect 5910 40319 5962 40325
rect 6269 40377 6321 40383
rect 6269 40319 6321 40325
rect 6870 40377 6922 40383
rect 6870 40319 6922 40325
rect 4758 40303 4810 40309
rect 4758 40245 4810 40251
rect 4770 40198 4798 40245
rect 5298 40198 5326 40319
rect 5382 40303 5434 40309
rect 5382 40245 5434 40251
rect 5785 40303 5837 40309
rect 5785 40245 5837 40251
rect 1108 40129 1164 40138
rect 1362 40152 1822 40180
rect 1926 40192 1978 40198
rect 1274 40118 1326 40124
rect 1274 40060 1326 40066
rect 1286 40032 1314 40060
rect 1218 40004 1314 40032
rect 1218 38755 1246 40004
rect 1362 39976 1390 40152
rect 2406 40192 2458 40198
rect 1978 40152 2302 40180
rect 1926 40134 1978 40140
rect 2274 40106 2302 40152
rect 2886 40192 2938 40198
rect 2458 40152 2782 40180
rect 2406 40134 2458 40140
rect 2754 40106 2782 40152
rect 3366 40192 3418 40198
rect 2938 40152 3262 40180
rect 2886 40134 2938 40140
rect 3234 40106 3262 40152
rect 3849 40192 3901 40198
rect 3418 40152 3742 40180
rect 3366 40134 3418 40140
rect 3714 40106 3742 40152
rect 4333 40192 4385 40198
rect 3901 40152 4222 40180
rect 3849 40134 3901 40140
rect 4194 40106 4222 40152
rect 4758 40192 4810 40198
rect 4385 40152 4702 40180
rect 4333 40134 4385 40140
rect 4674 40106 4702 40152
rect 4758 40134 4810 40140
rect 5286 40192 5338 40198
rect 5286 40134 5338 40140
rect 2274 40087 2542 40106
rect 2754 40087 3022 40106
rect 3234 40087 3502 40106
rect 3714 40087 3982 40106
rect 4194 40087 4462 40106
rect 4674 40087 4942 40106
rect 5394 40087 5422 40245
rect 5797 40198 5825 40245
rect 5785 40192 5837 40198
rect 5785 40134 5837 40140
rect 5922 40124 5950 40319
rect 6281 40198 6309 40319
rect 6390 40303 6442 40309
rect 6390 40245 6442 40251
rect 6774 40303 6826 40309
rect 6774 40245 6826 40251
rect 6269 40192 6321 40198
rect 6269 40134 6321 40140
rect 6402 40124 6430 40245
rect 6786 40198 6814 40245
rect 6774 40192 6826 40198
rect 6774 40134 6826 40140
rect 6882 40124 6910 40319
rect 7350 40303 7402 40309
rect 7350 40245 7402 40251
rect 8694 40303 8746 40309
rect 8694 40245 8746 40251
rect 9270 40303 9322 40309
rect 9270 40245 9322 40251
rect 7254 40192 7306 40198
rect 7254 40134 7306 40140
rect 5910 40118 5962 40124
rect 2274 40081 2554 40087
rect 2274 40078 2502 40081
rect 1452 40044 1504 40050
rect 1504 40013 2062 40032
rect 2754 40081 3034 40087
rect 2754 40078 2982 40081
rect 2502 40023 2554 40029
rect 3234 40081 3514 40087
rect 3234 40078 3462 40081
rect 2982 40023 3034 40029
rect 3714 40081 3994 40087
rect 3714 40078 3942 40081
rect 3462 40023 3514 40029
rect 4194 40081 4474 40087
rect 4194 40078 4422 40081
rect 3942 40023 3994 40029
rect 4674 40081 4954 40087
rect 4674 40078 4902 40081
rect 4422 40023 4474 40029
rect 4902 40023 4954 40029
rect 5382 40081 5434 40087
rect 5910 40060 5962 40066
rect 6390 40118 6442 40124
rect 6390 40060 6442 40066
rect 6870 40118 6922 40124
rect 6870 40060 6922 40066
rect 5382 40023 5434 40029
rect 1504 40007 2074 40013
rect 1504 40004 2022 40007
rect 1452 39986 1504 39992
rect 1350 39970 1402 39976
rect 2022 39949 2074 39955
rect 1350 39912 1402 39918
rect 7266 39884 7294 40134
rect 7362 40087 7390 40245
rect 8706 40198 8734 40245
rect 7734 40192 7786 40198
rect 8214 40192 8266 40198
rect 7786 40152 8158 40180
rect 7734 40134 7786 40140
rect 8130 40106 8158 40152
rect 8694 40192 8746 40198
rect 8266 40152 8638 40180
rect 8214 40134 8266 40140
rect 8610 40106 8638 40152
rect 8694 40134 8746 40140
rect 9174 40192 9226 40198
rect 9174 40134 9226 40140
rect 8130 40087 8350 40106
rect 8610 40087 8830 40106
rect 7350 40081 7402 40087
rect 8130 40081 8362 40087
rect 8130 40078 8310 40081
rect 7350 40023 7402 40029
rect 8610 40081 8842 40087
rect 8610 40078 8790 40081
rect 8310 40023 8362 40029
rect 8790 40023 8842 40029
rect 7830 39933 7882 39939
rect 7266 39881 7830 39884
rect 7266 39875 7882 39881
rect 7266 39856 7870 39875
rect 9186 39736 9214 40134
rect 9282 40087 9310 40245
rect 9270 40081 9322 40087
rect 9270 40023 9322 40029
rect 9186 39708 9310 39736
rect 3580 39528 3876 39548
rect 3636 39526 3660 39528
rect 3716 39526 3740 39528
rect 3796 39526 3820 39528
rect 3658 39474 3660 39526
rect 3722 39474 3734 39526
rect 3796 39474 3798 39526
rect 3636 39472 3660 39474
rect 3716 39472 3740 39474
rect 3796 39472 3820 39474
rect 3580 39452 3876 39472
rect 8908 39528 9204 39548
rect 8964 39526 8988 39528
rect 9044 39526 9068 39528
rect 9124 39526 9148 39528
rect 8986 39474 8988 39526
rect 9050 39474 9062 39526
rect 9124 39474 9126 39526
rect 8964 39472 8988 39474
rect 9044 39472 9068 39474
rect 9124 39472 9148 39474
rect 8908 39452 9204 39472
rect 9282 39199 9310 39708
rect 9270 39193 9322 39199
rect 9270 39135 9322 39141
rect 2022 38971 2074 38977
rect 2502 38971 2554 38977
rect 2074 38919 2398 38922
rect 2022 38913 2398 38919
rect 2982 38971 3034 38977
rect 2554 38919 2878 38922
rect 2502 38913 2878 38919
rect 3462 38971 3514 38977
rect 3034 38919 3358 38922
rect 2982 38913 3358 38919
rect 3942 38971 3994 38977
rect 3514 38919 3838 38922
rect 3462 38913 3838 38919
rect 4422 38971 4474 38977
rect 3994 38919 4318 38922
rect 3942 38913 4318 38919
rect 4902 38971 4954 38977
rect 4474 38919 4798 38922
rect 4422 38913 4798 38919
rect 5382 38971 5434 38977
rect 4954 38919 5324 38922
rect 4902 38913 5324 38919
rect 7350 38971 7402 38977
rect 5910 38934 5962 38940
rect 5434 38919 5806 38922
rect 5382 38913 5806 38919
rect 2034 38894 2398 38913
rect 2514 38894 2878 38913
rect 2994 38894 3358 38913
rect 3474 38894 3838 38913
rect 3954 38894 4318 38913
rect 4434 38894 4798 38913
rect 4914 38894 5324 38913
rect 5394 38894 5806 38913
rect 2370 38866 2398 38894
rect 2850 38866 2878 38894
rect 3330 38866 3358 38894
rect 3810 38866 3838 38894
rect 4290 38866 4318 38894
rect 4770 38866 4798 38894
rect 5296 38866 5324 38894
rect 5778 38866 5806 38894
rect 6390 38934 6442 38940
rect 5962 38894 6286 38922
rect 5910 38876 5962 38882
rect 6258 38866 6286 38894
rect 6870 38934 6922 38940
rect 6442 38894 6622 38922
rect 6390 38876 6442 38882
rect 1878 38860 1930 38866
rect 1878 38802 1930 38808
rect 2358 38860 2410 38866
rect 2358 38802 2410 38808
rect 2838 38860 2890 38866
rect 2838 38802 2890 38808
rect 3318 38860 3370 38866
rect 3318 38802 3370 38808
rect 3798 38860 3850 38866
rect 3798 38802 3850 38808
rect 4278 38860 4330 38866
rect 4278 38802 4330 38808
rect 4758 38860 4810 38866
rect 4758 38802 4810 38808
rect 5284 38860 5336 38866
rect 5284 38802 5336 38808
rect 5766 38860 5818 38866
rect 5766 38802 5818 38808
rect 6246 38860 6298 38866
rect 6594 38848 6622 38894
rect 6922 38894 7294 38922
rect 7830 38971 7882 38977
rect 7402 38919 7774 38922
rect 7350 38913 7774 38919
rect 8310 38971 8362 38977
rect 7882 38919 8254 38922
rect 7830 38913 8254 38919
rect 8790 38971 8842 38977
rect 8362 38919 8734 38922
rect 8310 38913 8734 38919
rect 8842 38919 9214 38922
rect 8790 38913 9214 38919
rect 7362 38894 7774 38913
rect 7842 38894 8254 38913
rect 8322 38894 8734 38913
rect 8802 38894 9214 38913
rect 6870 38876 6922 38882
rect 7266 38866 7294 38894
rect 7746 38866 7774 38894
rect 8226 38866 8254 38894
rect 8706 38866 8734 38894
rect 9186 38866 9214 38894
rect 6726 38860 6778 38866
rect 6594 38820 6726 38848
rect 6246 38802 6298 38808
rect 6726 38802 6778 38808
rect 7254 38860 7306 38866
rect 7254 38802 7306 38808
rect 7734 38860 7786 38866
rect 7734 38802 7786 38808
rect 8214 38860 8266 38866
rect 8214 38802 8266 38808
rect 8694 38860 8746 38866
rect 8694 38802 8746 38808
rect 9174 38860 9226 38866
rect 9174 38802 9226 38808
rect 1890 38755 1918 38802
rect 1206 38749 1258 38755
rect 1206 38691 1258 38697
rect 1878 38749 1930 38755
rect 1878 38691 1930 38697
rect 1110 37528 1162 37534
rect 1110 37470 1162 37476
rect 1122 37391 1150 37470
rect 1108 37382 1164 37391
rect 1218 37368 1246 38691
rect 6244 38196 6540 38216
rect 6300 38194 6324 38196
rect 6380 38194 6404 38196
rect 6460 38194 6484 38196
rect 6322 38142 6324 38194
rect 6386 38142 6398 38194
rect 6460 38142 6462 38194
rect 6300 38140 6324 38142
rect 6380 38140 6404 38142
rect 6460 38140 6484 38142
rect 6244 38120 6540 38140
rect 5785 37713 5837 37719
rect 5785 37655 5837 37661
rect 6269 37713 6321 37719
rect 6269 37655 6321 37661
rect 6870 37713 6922 37719
rect 6870 37655 6922 37661
rect 5301 37639 5353 37645
rect 5301 37581 5353 37587
rect 5313 37534 5341 37581
rect 5797 37534 5825 37655
rect 5910 37639 5962 37645
rect 5910 37581 5962 37587
rect 1926 37528 1978 37534
rect 1398 37491 1450 37497
rect 1302 37454 1354 37460
rect 1354 37439 1398 37442
rect 2406 37528 2458 37534
rect 1978 37488 2302 37516
rect 1926 37470 1978 37476
rect 1354 37433 1450 37439
rect 2274 37442 2302 37488
rect 2886 37528 2938 37534
rect 2458 37488 2782 37516
rect 2406 37470 2458 37476
rect 2754 37442 2782 37488
rect 3366 37528 3418 37534
rect 2938 37488 3262 37516
rect 2886 37470 2938 37476
rect 3234 37442 3262 37488
rect 3849 37528 3901 37534
rect 3418 37488 3742 37516
rect 3366 37470 3418 37476
rect 3714 37442 3742 37488
rect 4333 37528 4385 37534
rect 3901 37488 4222 37516
rect 3849 37470 3901 37476
rect 4194 37442 4222 37488
rect 4817 37528 4869 37534
rect 4385 37488 4702 37516
rect 4333 37470 4385 37476
rect 4674 37442 4702 37488
rect 5301 37528 5353 37534
rect 4869 37488 5182 37516
rect 4817 37470 4869 37476
rect 5154 37442 5182 37488
rect 5301 37470 5353 37476
rect 5785 37528 5837 37534
rect 5785 37470 5837 37476
rect 5922 37460 5950 37581
rect 6281 37534 6309 37655
rect 6390 37639 6442 37645
rect 6390 37581 6442 37587
rect 6774 37639 6826 37645
rect 6774 37581 6826 37587
rect 6269 37528 6321 37534
rect 6269 37470 6321 37476
rect 6402 37460 6430 37581
rect 6786 37534 6814 37581
rect 6774 37528 6826 37534
rect 6774 37470 6826 37476
rect 6882 37460 6910 37655
rect 7350 37639 7402 37645
rect 7350 37581 7402 37587
rect 8694 37639 8746 37645
rect 8694 37581 8746 37587
rect 9270 37639 9322 37645
rect 9270 37581 9322 37587
rect 7254 37528 7306 37534
rect 7254 37470 7306 37476
rect 5910 37454 5962 37460
rect 1354 37414 1438 37433
rect 2274 37423 2542 37442
rect 2754 37423 3022 37442
rect 3234 37423 3502 37442
rect 3714 37423 3982 37442
rect 4194 37423 4462 37442
rect 4674 37423 4942 37442
rect 5154 37423 5422 37442
rect 2274 37417 2554 37423
rect 2274 37414 2502 37417
rect 1302 37396 1354 37402
rect 1452 37380 1504 37386
rect 1218 37340 1390 37368
rect 1108 37317 1164 37326
rect 1362 37312 1390 37340
rect 1504 37349 2062 37368
rect 2754 37417 3034 37423
rect 2754 37414 2982 37417
rect 2502 37359 2554 37365
rect 3234 37417 3514 37423
rect 3234 37414 3462 37417
rect 2982 37359 3034 37365
rect 3714 37417 3994 37423
rect 3714 37414 3942 37417
rect 3462 37359 3514 37365
rect 4194 37417 4474 37423
rect 4194 37414 4422 37417
rect 3942 37359 3994 37365
rect 4674 37417 4954 37423
rect 4674 37414 4902 37417
rect 4422 37359 4474 37365
rect 5154 37417 5434 37423
rect 5154 37414 5382 37417
rect 4902 37359 4954 37365
rect 5910 37396 5962 37402
rect 6390 37454 6442 37460
rect 6390 37396 6442 37402
rect 6870 37454 6922 37460
rect 6870 37396 6922 37402
rect 5382 37359 5434 37365
rect 1504 37343 2074 37349
rect 1504 37340 2022 37343
rect 1452 37322 1504 37328
rect 1350 37306 1402 37312
rect 2022 37285 2074 37291
rect 1350 37248 1402 37254
rect 1782 37269 1834 37275
rect 1782 37211 1834 37217
rect 7266 37220 7294 37470
rect 7362 37423 7390 37581
rect 8706 37534 8734 37581
rect 7734 37528 7786 37534
rect 8214 37528 8266 37534
rect 7786 37488 8158 37516
rect 7734 37470 7786 37476
rect 8130 37442 8158 37488
rect 8694 37528 8746 37534
rect 8266 37488 8638 37516
rect 8214 37470 8266 37476
rect 8610 37442 8638 37488
rect 8694 37470 8746 37476
rect 9174 37528 9226 37534
rect 9174 37470 9226 37476
rect 8130 37423 8350 37442
rect 8610 37423 8830 37442
rect 7350 37417 7402 37423
rect 8130 37417 8362 37423
rect 8130 37414 8310 37417
rect 7350 37359 7402 37365
rect 8610 37417 8842 37423
rect 8610 37414 8790 37417
rect 8310 37359 8362 37365
rect 8790 37359 8842 37365
rect 7830 37343 7882 37349
rect 7830 37285 7882 37291
rect 7842 37220 7870 37285
rect 1794 33520 1822 37211
rect 7266 37192 7870 37220
rect 9186 37072 9214 37470
rect 9282 37423 9310 37581
rect 9270 37417 9322 37423
rect 9270 37359 9322 37365
rect 9186 37044 9310 37072
rect 3580 36864 3876 36884
rect 3636 36862 3660 36864
rect 3716 36862 3740 36864
rect 3796 36862 3820 36864
rect 3658 36810 3660 36862
rect 3722 36810 3734 36862
rect 3796 36810 3798 36862
rect 3636 36808 3660 36810
rect 3716 36808 3740 36810
rect 3796 36808 3820 36810
rect 3580 36788 3876 36808
rect 8908 36864 9204 36884
rect 8964 36862 8988 36864
rect 9044 36862 9068 36864
rect 9124 36862 9148 36864
rect 8986 36810 8988 36862
rect 9050 36810 9062 36862
rect 9124 36810 9126 36862
rect 8964 36808 8988 36810
rect 9044 36808 9068 36810
rect 9124 36808 9148 36810
rect 8908 36788 9204 36808
rect 9282 36535 9310 37044
rect 9270 36529 9322 36535
rect 9270 36471 9322 36477
rect 2022 36307 2074 36313
rect 2502 36307 2554 36313
rect 2074 36255 2398 36258
rect 2022 36249 2398 36255
rect 2982 36307 3034 36313
rect 2554 36255 2878 36258
rect 2502 36249 2878 36255
rect 3462 36307 3514 36313
rect 3034 36255 3358 36258
rect 2982 36249 3358 36255
rect 3942 36307 3994 36313
rect 3514 36255 3838 36258
rect 3462 36249 3838 36255
rect 4422 36307 4474 36313
rect 3994 36255 4318 36258
rect 3942 36249 4318 36255
rect 4902 36307 4954 36313
rect 4474 36255 4798 36258
rect 4422 36249 4798 36255
rect 5382 36307 5434 36313
rect 4954 36255 5324 36258
rect 4902 36249 5324 36255
rect 7350 36307 7402 36313
rect 5910 36270 5962 36276
rect 5434 36255 5806 36258
rect 5382 36249 5806 36255
rect 2034 36230 2398 36249
rect 2514 36230 2878 36249
rect 2994 36230 3358 36249
rect 3474 36230 3838 36249
rect 3954 36230 4318 36249
rect 4434 36230 4798 36249
rect 4914 36230 5324 36249
rect 5394 36230 5806 36249
rect 2370 36202 2398 36230
rect 2850 36202 2878 36230
rect 3330 36202 3358 36230
rect 3810 36202 3838 36230
rect 4290 36202 4318 36230
rect 4770 36202 4798 36230
rect 5296 36202 5324 36230
rect 5778 36202 5806 36230
rect 6390 36270 6442 36276
rect 5962 36230 6286 36258
rect 5910 36212 5962 36218
rect 6258 36202 6286 36230
rect 6870 36270 6922 36276
rect 6442 36230 6622 36258
rect 6390 36212 6442 36218
rect 1926 36196 1978 36202
rect 2358 36196 2410 36202
rect 1978 36156 2110 36184
rect 1926 36138 1978 36144
rect 2082 35000 2110 36156
rect 2358 36138 2410 36144
rect 2838 36196 2890 36202
rect 2838 36138 2890 36144
rect 3318 36196 3370 36202
rect 3318 36138 3370 36144
rect 3798 36196 3850 36202
rect 3798 36138 3850 36144
rect 4278 36196 4330 36202
rect 4278 36138 4330 36144
rect 4758 36196 4810 36202
rect 4758 36138 4810 36144
rect 5284 36196 5336 36202
rect 5284 36138 5336 36144
rect 5766 36196 5818 36202
rect 5766 36138 5818 36144
rect 6246 36196 6298 36202
rect 6594 36184 6622 36230
rect 7350 36249 7402 36255
rect 7830 36307 7882 36313
rect 7830 36249 7882 36255
rect 8310 36307 8362 36313
rect 8310 36249 8362 36255
rect 8790 36307 8842 36313
rect 8790 36249 8842 36255
rect 6870 36212 6922 36218
rect 6726 36196 6778 36202
rect 6594 36156 6726 36184
rect 6246 36138 6298 36144
rect 6882 36184 6910 36212
rect 7206 36196 7258 36202
rect 6882 36156 7206 36184
rect 6726 36138 6778 36144
rect 7362 36184 7390 36249
rect 7686 36196 7738 36202
rect 7362 36156 7686 36184
rect 7206 36138 7258 36144
rect 7842 36184 7870 36249
rect 8166 36196 8218 36202
rect 7842 36156 8166 36184
rect 7686 36138 7738 36144
rect 8322 36184 8350 36249
rect 8646 36196 8698 36202
rect 8322 36156 8646 36184
rect 8166 36138 8218 36144
rect 8802 36184 8830 36249
rect 9126 36196 9178 36202
rect 8802 36156 9126 36184
rect 8646 36138 8698 36144
rect 9126 36138 9178 36144
rect 6244 35532 6540 35552
rect 6300 35530 6324 35532
rect 6380 35530 6404 35532
rect 6460 35530 6484 35532
rect 6322 35478 6324 35530
rect 6386 35478 6398 35530
rect 6460 35478 6462 35530
rect 6300 35476 6324 35478
rect 6380 35476 6404 35478
rect 6460 35476 6484 35478
rect 6244 35456 6540 35476
rect 2034 34972 2110 35000
rect 5785 34975 5837 34981
rect 1878 34864 1930 34870
rect 1878 34806 1930 34812
rect 1890 34727 1918 34806
rect 2034 34759 2062 34972
rect 5785 34917 5837 34923
rect 9090 34972 9310 35000
rect 2406 34864 2458 34870
rect 2886 34864 2938 34870
rect 2458 34824 2782 34852
rect 2406 34806 2458 34812
rect 2022 34753 2074 34759
rect 1876 34718 1932 34727
rect 2022 34695 2074 34701
rect 2500 34718 2556 34727
rect 1876 34653 1932 34662
rect 2754 34704 2782 34824
rect 3366 34864 3418 34870
rect 2938 34824 3262 34852
rect 2886 34806 2938 34812
rect 3234 34704 3262 34824
rect 3849 34864 3901 34870
rect 3418 34824 3742 34852
rect 3366 34806 3418 34812
rect 3714 34704 3742 34824
rect 4333 34864 4385 34870
rect 3901 34824 4222 34852
rect 3849 34806 3901 34812
rect 4194 34704 4222 34824
rect 4817 34864 4869 34870
rect 4385 34824 4702 34852
rect 4333 34806 4385 34812
rect 4674 34704 4702 34824
rect 5299 34866 5355 34875
rect 5797 34870 5825 34917
rect 6390 34901 6442 34907
rect 4869 34824 5182 34852
rect 4817 34806 4869 34812
rect 5154 34704 5182 34824
rect 5299 34801 5355 34810
rect 5785 34864 5837 34870
rect 5785 34806 5837 34812
rect 5908 34866 5964 34875
rect 5908 34801 5964 34810
rect 6269 34864 6321 34870
rect 6321 34812 6334 34852
rect 6390 34843 6442 34849
rect 6774 34864 6826 34870
rect 6269 34806 6334 34812
rect 2754 34685 3022 34704
rect 3234 34685 3502 34704
rect 3714 34685 3982 34704
rect 4194 34685 4462 34704
rect 4674 34685 4942 34704
rect 5154 34685 5422 34704
rect 2754 34679 3034 34685
rect 2754 34676 2982 34679
rect 2500 34653 2502 34662
rect 2554 34653 2556 34662
rect 2502 34621 2554 34627
rect 3234 34679 3514 34685
rect 3234 34676 3462 34679
rect 2982 34621 3034 34627
rect 3714 34679 3994 34685
rect 3714 34676 3942 34679
rect 3462 34621 3514 34627
rect 4194 34679 4474 34685
rect 4194 34676 4422 34679
rect 3942 34621 3994 34627
rect 4674 34679 4954 34685
rect 4674 34676 4902 34679
rect 4422 34621 4474 34627
rect 5154 34679 5434 34685
rect 5154 34676 5382 34679
rect 4902 34621 4954 34627
rect 5382 34621 5434 34627
rect 5922 34500 5950 34801
rect 5910 34494 5962 34500
rect 5910 34436 5962 34442
rect 6306 34389 6334 34806
rect 6402 34796 6430 34843
rect 7254 34864 7306 34870
rect 6826 34824 7198 34852
rect 6774 34806 6826 34812
rect 6390 34790 6442 34796
rect 6390 34732 6442 34738
rect 7170 34704 7198 34824
rect 7734 34864 7786 34870
rect 7306 34824 7678 34852
rect 7254 34806 7306 34812
rect 7650 34704 7678 34824
rect 8214 34864 8266 34870
rect 7786 34824 8158 34852
rect 7734 34806 7786 34812
rect 8130 34704 8158 34824
rect 8694 34864 8746 34870
rect 8266 34824 8638 34852
rect 8214 34806 8266 34812
rect 8610 34704 8638 34824
rect 9090 34852 9118 34972
rect 8746 34824 9118 34852
rect 9174 34864 9226 34870
rect 8694 34806 8746 34812
rect 9174 34806 9226 34812
rect 7170 34685 7390 34704
rect 7650 34685 7870 34704
rect 8130 34685 8350 34704
rect 8610 34685 8830 34704
rect 7170 34679 7402 34685
rect 7170 34676 7350 34679
rect 7650 34679 7882 34685
rect 7650 34676 7830 34679
rect 7350 34621 7402 34627
rect 8130 34679 8362 34685
rect 8130 34676 8310 34679
rect 7830 34621 7882 34627
rect 8610 34679 8842 34685
rect 8610 34676 8790 34679
rect 8310 34621 8362 34627
rect 8790 34621 8842 34627
rect 6870 34494 6922 34500
rect 6870 34436 6922 34442
rect 6882 34389 6910 34436
rect 9186 34408 9214 34806
rect 9282 34759 9310 34972
rect 9270 34753 9322 34759
rect 9270 34695 9322 34701
rect 6294 34383 6346 34389
rect 6294 34325 6346 34331
rect 6870 34383 6922 34389
rect 9186 34380 9310 34408
rect 6870 34325 6922 34331
rect 3580 34200 3876 34220
rect 3636 34198 3660 34200
rect 3716 34198 3740 34200
rect 3796 34198 3820 34200
rect 3658 34146 3660 34198
rect 3722 34146 3734 34198
rect 3796 34146 3798 34198
rect 3636 34144 3660 34146
rect 3716 34144 3740 34146
rect 3796 34144 3820 34146
rect 3580 34124 3876 34144
rect 8908 34200 9204 34220
rect 8964 34198 8988 34200
rect 9044 34198 9068 34200
rect 9124 34198 9148 34200
rect 8986 34146 8988 34198
rect 9050 34146 9062 34198
rect 9124 34146 9126 34198
rect 8964 34144 8988 34146
rect 9044 34144 9068 34146
rect 9124 34144 9148 34146
rect 8908 34124 9204 34144
rect 6390 33902 6442 33908
rect 9282 33871 9310 34380
rect 6390 33844 6442 33850
rect 9270 33865 9322 33871
rect 6402 33816 6430 33844
rect 2994 33797 3358 33816
rect 3954 33797 4318 33816
rect 5394 33797 5806 33816
rect 2982 33791 3358 33797
rect 3034 33788 3358 33791
rect 2982 33733 3034 33739
rect 2022 33643 2074 33649
rect 2502 33643 2554 33649
rect 2074 33591 2398 33594
rect 2022 33585 2398 33591
rect 2554 33591 2878 33594
rect 2502 33585 2878 33591
rect 2034 33566 2398 33585
rect 2514 33566 2878 33585
rect 2370 33538 2398 33566
rect 2850 33538 2878 33566
rect 3330 33538 3358 33788
rect 3942 33791 4318 33797
rect 3994 33788 4318 33791
rect 3942 33733 3994 33739
rect 3462 33643 3514 33649
rect 3514 33591 3838 33594
rect 3462 33585 3838 33591
rect 3474 33566 3838 33585
rect 3810 33538 3838 33566
rect 4290 33538 4318 33788
rect 5382 33791 5806 33797
rect 5434 33788 5806 33791
rect 6402 33788 6814 33816
rect 9270 33807 9322 33813
rect 5382 33733 5434 33739
rect 4422 33643 4474 33649
rect 4902 33643 4954 33649
rect 4474 33591 4798 33594
rect 4422 33585 4798 33591
rect 4954 33591 5324 33594
rect 4902 33585 5324 33591
rect 4434 33566 4798 33585
rect 4914 33566 5324 33585
rect 4770 33538 4798 33566
rect 5296 33538 5324 33566
rect 5778 33538 5806 33788
rect 5910 33606 5962 33612
rect 5962 33566 6286 33594
rect 5910 33548 5962 33554
rect 6258 33538 6286 33566
rect 6786 33538 6814 33788
rect 7350 33643 7402 33649
rect 6870 33606 6922 33612
rect 7830 33643 7882 33649
rect 7402 33603 7774 33631
rect 7350 33585 7402 33591
rect 6870 33548 6922 33554
rect 1878 33532 1930 33538
rect 1794 33492 1878 33520
rect 1110 32200 1162 32206
rect 1110 32142 1162 32148
rect 1122 32063 1150 32142
rect 1274 32126 1326 32132
rect 1794 32114 1822 33492
rect 1878 33474 1930 33480
rect 2358 33532 2410 33538
rect 2358 33474 2410 33480
rect 2838 33532 2890 33538
rect 2838 33474 2890 33480
rect 3318 33532 3370 33538
rect 3318 33474 3370 33480
rect 3798 33532 3850 33538
rect 3798 33474 3850 33480
rect 4278 33532 4330 33538
rect 4278 33474 4330 33480
rect 4758 33532 4810 33538
rect 4758 33474 4810 33480
rect 5284 33532 5336 33538
rect 5284 33474 5336 33480
rect 5766 33532 5818 33538
rect 5766 33474 5818 33480
rect 6246 33532 6298 33538
rect 6246 33474 6298 33480
rect 6774 33532 6826 33538
rect 6882 33520 6910 33548
rect 7746 33538 7774 33603
rect 8310 33643 8362 33649
rect 7882 33603 8254 33631
rect 7830 33585 7882 33591
rect 8226 33538 8254 33603
rect 8790 33643 8842 33649
rect 8362 33603 8734 33631
rect 8310 33585 8362 33591
rect 8706 33538 8734 33603
rect 8842 33603 9214 33631
rect 8790 33585 8842 33591
rect 9186 33538 9214 33603
rect 7206 33532 7258 33538
rect 6882 33492 7206 33520
rect 6774 33474 6826 33480
rect 7206 33474 7258 33480
rect 7734 33532 7786 33538
rect 7734 33474 7786 33480
rect 8214 33532 8266 33538
rect 8214 33474 8266 33480
rect 8694 33532 8746 33538
rect 8694 33474 8746 33480
rect 9174 33532 9226 33538
rect 9174 33474 9226 33480
rect 6244 32868 6540 32888
rect 6300 32866 6324 32868
rect 6380 32866 6404 32868
rect 6460 32866 6484 32868
rect 6322 32814 6324 32866
rect 6386 32814 6398 32866
rect 6460 32814 6462 32866
rect 6300 32812 6324 32814
rect 6380 32812 6404 32814
rect 6460 32812 6484 32814
rect 6244 32792 6540 32812
rect 5286 32385 5338 32391
rect 5286 32327 5338 32333
rect 5910 32385 5962 32391
rect 5910 32327 5962 32333
rect 6269 32385 6321 32391
rect 6269 32327 6321 32333
rect 6870 32385 6922 32391
rect 6870 32327 6922 32333
rect 4758 32311 4810 32317
rect 4758 32253 4810 32259
rect 4770 32206 4798 32253
rect 5298 32206 5326 32327
rect 5382 32311 5434 32317
rect 5382 32253 5434 32259
rect 5785 32311 5837 32317
rect 5785 32253 5837 32259
rect 1926 32200 1978 32206
rect 2406 32200 2458 32206
rect 1978 32160 2302 32188
rect 1926 32142 1978 32148
rect 1274 32068 1326 32074
rect 1362 32086 1822 32114
rect 2274 32114 2302 32160
rect 2886 32200 2938 32206
rect 2458 32160 2782 32188
rect 2406 32142 2458 32148
rect 2754 32114 2782 32160
rect 3366 32200 3418 32206
rect 2938 32160 3262 32188
rect 2886 32142 2938 32148
rect 3234 32114 3262 32160
rect 3849 32200 3901 32206
rect 3418 32160 3742 32188
rect 3366 32142 3418 32148
rect 3714 32114 3742 32160
rect 4333 32200 4385 32206
rect 3901 32160 4222 32188
rect 3849 32142 3901 32148
rect 4194 32114 4222 32160
rect 4758 32200 4810 32206
rect 4385 32160 4702 32188
rect 4333 32142 4385 32148
rect 4674 32114 4702 32160
rect 4758 32142 4810 32148
rect 5286 32200 5338 32206
rect 5286 32142 5338 32148
rect 2274 32095 2542 32114
rect 2754 32095 3022 32114
rect 3234 32095 3502 32114
rect 3714 32095 3982 32114
rect 4194 32095 4462 32114
rect 4674 32095 4942 32114
rect 5394 32095 5422 32253
rect 5797 32206 5825 32253
rect 5785 32200 5837 32206
rect 5785 32142 5837 32148
rect 5922 32132 5950 32327
rect 6281 32206 6309 32327
rect 6390 32311 6442 32317
rect 6390 32253 6442 32259
rect 6774 32311 6826 32317
rect 6774 32253 6826 32259
rect 6269 32200 6321 32206
rect 6269 32142 6321 32148
rect 6402 32132 6430 32253
rect 6786 32206 6814 32253
rect 6774 32200 6826 32206
rect 6774 32142 6826 32148
rect 6882 32132 6910 32327
rect 7350 32311 7402 32317
rect 7350 32253 7402 32259
rect 8694 32311 8746 32317
rect 8694 32253 8746 32259
rect 9270 32311 9322 32317
rect 9270 32253 9322 32259
rect 7254 32200 7306 32206
rect 7254 32142 7306 32148
rect 5910 32126 5962 32132
rect 2274 32089 2554 32095
rect 2274 32086 2502 32089
rect 1108 32054 1164 32063
rect 1108 31989 1164 31998
rect 1286 31892 1314 32068
rect 1362 31984 1390 32086
rect 1452 32052 1504 32058
rect 1504 32021 2062 32040
rect 2754 32089 3034 32095
rect 2754 32086 2982 32089
rect 2502 32031 2554 32037
rect 3234 32089 3514 32095
rect 3234 32086 3462 32089
rect 2982 32031 3034 32037
rect 3714 32089 3994 32095
rect 3714 32086 3942 32089
rect 3462 32031 3514 32037
rect 4194 32089 4474 32095
rect 4194 32086 4422 32089
rect 3942 32031 3994 32037
rect 4674 32089 4954 32095
rect 4674 32086 4902 32089
rect 4422 32031 4474 32037
rect 4902 32031 4954 32037
rect 5382 32089 5434 32095
rect 5910 32068 5962 32074
rect 6390 32126 6442 32132
rect 6390 32068 6442 32074
rect 6870 32126 6922 32132
rect 6870 32068 6922 32074
rect 5382 32031 5434 32037
rect 1504 32015 2074 32021
rect 1504 32012 2022 32015
rect 1452 31994 1504 32000
rect 1350 31978 1402 31984
rect 2022 31957 2074 31963
rect 1350 31920 1402 31926
rect 7266 31892 7294 32142
rect 7362 32095 7390 32253
rect 8706 32206 8734 32253
rect 7734 32200 7786 32206
rect 8214 32200 8266 32206
rect 7786 32160 8158 32188
rect 7734 32142 7786 32148
rect 8130 32114 8158 32160
rect 8694 32200 8746 32206
rect 8266 32160 8638 32188
rect 8214 32142 8266 32148
rect 8610 32114 8638 32160
rect 8694 32142 8746 32148
rect 9174 32200 9226 32206
rect 9174 32142 9226 32148
rect 8130 32095 8350 32114
rect 8610 32095 8830 32114
rect 7350 32089 7402 32095
rect 8130 32089 8362 32095
rect 8130 32086 8310 32089
rect 7350 32031 7402 32037
rect 8610 32089 8842 32095
rect 8610 32086 8790 32089
rect 8310 32031 8362 32037
rect 8790 32031 8842 32037
rect 7830 31941 7882 31947
rect 1286 31864 1342 31892
rect 7266 31889 7830 31892
rect 7266 31883 7882 31889
rect 7266 31864 7870 31883
rect 1314 31725 1342 31864
rect 9186 31744 9214 32142
rect 9282 32095 9310 32253
rect 9270 32089 9322 32095
rect 9270 32031 9322 32037
rect 1302 31719 1354 31725
rect 1302 31661 1354 31667
rect 1782 31719 1834 31725
rect 9186 31716 9310 31744
rect 1782 31661 1834 31667
rect 1794 22864 1822 31661
rect 3580 31536 3876 31556
rect 3636 31534 3660 31536
rect 3716 31534 3740 31536
rect 3796 31534 3820 31536
rect 3658 31482 3660 31534
rect 3722 31482 3734 31534
rect 3796 31482 3798 31534
rect 3636 31480 3660 31482
rect 3716 31480 3740 31482
rect 3796 31480 3820 31482
rect 3580 31460 3876 31480
rect 8908 31536 9204 31556
rect 8964 31534 8988 31536
rect 9044 31534 9068 31536
rect 9124 31534 9148 31536
rect 8986 31482 8988 31534
rect 9050 31482 9062 31534
rect 9124 31482 9126 31534
rect 8964 31480 8988 31482
rect 9044 31480 9068 31482
rect 9124 31480 9148 31482
rect 8908 31460 9204 31480
rect 9282 31207 9310 31716
rect 9270 31201 9322 31207
rect 9270 31143 9322 31149
rect 2022 30979 2074 30985
rect 2502 30979 2554 30985
rect 2074 30927 2398 30930
rect 2022 30921 2398 30927
rect 2982 30979 3034 30985
rect 2554 30927 2878 30930
rect 2502 30921 2878 30927
rect 3462 30979 3514 30985
rect 3034 30927 3262 30930
rect 2982 30921 3262 30927
rect 3942 30979 3994 30985
rect 3514 30939 3838 30967
rect 3462 30921 3514 30927
rect 2034 30902 2398 30921
rect 2514 30902 2878 30921
rect 2994 30902 3262 30921
rect 2370 30874 2398 30902
rect 2850 30874 2878 30902
rect 1878 30868 1930 30874
rect 1878 30810 1930 30816
rect 2358 30868 2410 30874
rect 2358 30810 2410 30816
rect 2838 30868 2890 30874
rect 3234 30856 3262 30902
rect 3810 30874 3838 30939
rect 4422 30979 4474 30985
rect 3994 30939 4318 30967
rect 3942 30921 3994 30927
rect 4290 30874 4318 30939
rect 4902 30979 4954 30985
rect 4474 30939 4798 30967
rect 4422 30921 4474 30927
rect 4770 30874 4798 30939
rect 5382 30979 5434 30985
rect 4954 30939 5324 30967
rect 4902 30921 4954 30927
rect 5296 30874 5324 30939
rect 7350 30979 7402 30985
rect 5434 30939 5806 30967
rect 5382 30921 5434 30927
rect 5778 30874 5806 30939
rect 5910 30942 5962 30948
rect 6390 30942 6442 30948
rect 5962 30902 6286 30930
rect 5910 30884 5962 30890
rect 6258 30874 6286 30902
rect 6870 30942 6922 30948
rect 6442 30902 6814 30930
rect 6390 30884 6442 30890
rect 6786 30874 6814 30902
rect 6922 30902 7294 30930
rect 7830 30979 7882 30985
rect 7402 30939 7774 30967
rect 7350 30921 7402 30927
rect 6870 30884 6922 30890
rect 7266 30874 7294 30902
rect 7746 30874 7774 30939
rect 8310 30979 8362 30985
rect 7882 30939 8254 30967
rect 7830 30921 7882 30927
rect 8226 30874 8254 30939
rect 8790 30979 8842 30985
rect 8362 30939 8734 30967
rect 8310 30921 8362 30927
rect 8706 30874 8734 30939
rect 8842 30939 9214 30967
rect 8790 30921 8842 30927
rect 9186 30874 9214 30939
rect 3318 30868 3370 30874
rect 3234 30828 3318 30856
rect 2838 30810 2890 30816
rect 3318 30810 3370 30816
rect 3798 30868 3850 30874
rect 3798 30810 3850 30816
rect 4278 30868 4330 30874
rect 4278 30810 4330 30816
rect 4758 30868 4810 30874
rect 4758 30810 4810 30816
rect 5284 30868 5336 30874
rect 5284 30810 5336 30816
rect 5766 30868 5818 30874
rect 5766 30810 5818 30816
rect 6246 30868 6298 30874
rect 6246 30810 6298 30816
rect 6774 30868 6826 30874
rect 6774 30810 6826 30816
rect 7254 30868 7306 30874
rect 7254 30810 7306 30816
rect 7734 30868 7786 30874
rect 7734 30810 7786 30816
rect 8214 30868 8266 30874
rect 8214 30810 8266 30816
rect 8694 30868 8746 30874
rect 8694 30810 8746 30816
rect 9174 30868 9226 30874
rect 9174 30810 9226 30816
rect 1890 30264 1918 30810
rect 1890 30236 2014 30264
rect 1986 29635 2014 30236
rect 6244 30204 6540 30224
rect 6300 30202 6324 30204
rect 6380 30202 6404 30204
rect 6460 30202 6484 30204
rect 6322 30150 6324 30202
rect 6386 30150 6398 30202
rect 6460 30150 6462 30202
rect 6300 30148 6324 30150
rect 6380 30148 6404 30150
rect 6460 30148 6484 30150
rect 6244 30128 6540 30148
rect 5286 29721 5338 29727
rect 5286 29663 5338 29669
rect 5910 29721 5962 29727
rect 5910 29663 5962 29669
rect 6269 29721 6321 29727
rect 6269 29663 6321 29669
rect 6870 29721 6922 29727
rect 6870 29663 6922 29669
rect 4758 29647 4810 29653
rect 1986 29607 2062 29635
rect 1878 29536 1930 29542
rect 1878 29478 1930 29484
rect 1890 29399 1918 29478
rect 2034 29431 2062 29607
rect 4758 29589 4810 29595
rect 4770 29542 4798 29589
rect 5298 29542 5326 29663
rect 5382 29647 5434 29653
rect 5382 29589 5434 29595
rect 5785 29647 5837 29653
rect 5785 29589 5837 29595
rect 2406 29536 2458 29542
rect 2886 29536 2938 29542
rect 2458 29496 2782 29524
rect 2406 29478 2458 29484
rect 2754 29450 2782 29496
rect 3366 29536 3418 29542
rect 2938 29496 3262 29524
rect 2886 29478 2938 29484
rect 3234 29450 3262 29496
rect 3849 29536 3901 29542
rect 3418 29496 3742 29524
rect 3366 29478 3418 29484
rect 2754 29431 3022 29450
rect 3234 29431 3502 29450
rect 2022 29425 2074 29431
rect 1876 29390 1932 29399
rect 2754 29425 3034 29431
rect 2754 29422 2982 29425
rect 2022 29367 2074 29373
rect 2500 29390 2556 29399
rect 1876 29325 1932 29334
rect 3234 29425 3514 29431
rect 3234 29422 3462 29425
rect 2982 29367 3034 29373
rect 3714 29413 3742 29496
rect 4333 29536 4385 29542
rect 3901 29496 4222 29524
rect 3849 29478 3901 29484
rect 4194 29450 4222 29496
rect 4758 29536 4810 29542
rect 4385 29496 4702 29524
rect 4333 29478 4385 29484
rect 4674 29450 4702 29496
rect 4758 29478 4810 29484
rect 5286 29536 5338 29542
rect 5286 29478 5338 29484
rect 4194 29431 4462 29450
rect 4674 29431 4942 29450
rect 5394 29431 5422 29589
rect 5797 29542 5825 29589
rect 5785 29536 5837 29542
rect 5785 29478 5837 29484
rect 5922 29468 5950 29663
rect 6281 29542 6309 29663
rect 6390 29647 6442 29653
rect 6390 29589 6442 29595
rect 6774 29647 6826 29653
rect 6774 29589 6826 29595
rect 6269 29536 6321 29542
rect 6269 29478 6321 29484
rect 6402 29468 6430 29589
rect 6786 29542 6814 29589
rect 6774 29536 6826 29542
rect 6774 29478 6826 29484
rect 6882 29468 6910 29663
rect 7350 29647 7402 29653
rect 7350 29589 7402 29595
rect 8694 29647 8746 29653
rect 8694 29589 8746 29595
rect 9270 29647 9322 29653
rect 9270 29589 9322 29595
rect 7254 29536 7306 29542
rect 7254 29478 7306 29484
rect 5910 29462 5962 29468
rect 3942 29425 3994 29431
rect 3714 29385 3942 29413
rect 3462 29367 3514 29373
rect 4194 29425 4474 29431
rect 4194 29422 4422 29425
rect 3942 29367 3994 29373
rect 4674 29425 4954 29431
rect 4674 29422 4902 29425
rect 4422 29367 4474 29373
rect 4902 29367 4954 29373
rect 5382 29425 5434 29431
rect 5910 29404 5962 29410
rect 6390 29462 6442 29468
rect 6390 29404 6442 29410
rect 6870 29462 6922 29468
rect 6870 29404 6922 29410
rect 5382 29367 5434 29373
rect 2500 29325 2502 29334
rect 2554 29325 2556 29334
rect 2502 29293 2554 29299
rect 7266 29228 7294 29478
rect 7362 29431 7390 29589
rect 8706 29542 8734 29589
rect 7734 29536 7786 29542
rect 8214 29536 8266 29542
rect 7786 29496 8158 29524
rect 7734 29478 7786 29484
rect 7350 29425 7402 29431
rect 8130 29413 8158 29496
rect 8694 29536 8746 29542
rect 8266 29496 8638 29524
rect 8214 29478 8266 29484
rect 8310 29425 8362 29431
rect 8130 29385 8310 29413
rect 7350 29367 7402 29373
rect 8610 29413 8638 29496
rect 8694 29478 8746 29484
rect 9174 29536 9226 29542
rect 9174 29478 9226 29484
rect 8790 29425 8842 29431
rect 8610 29385 8790 29413
rect 8310 29367 8362 29373
rect 8790 29367 8842 29373
rect 7830 29277 7882 29283
rect 7266 29225 7830 29228
rect 7266 29219 7882 29225
rect 7266 29200 7870 29219
rect 9186 29080 9214 29478
rect 9282 29431 9310 29589
rect 9270 29425 9322 29431
rect 9270 29367 9322 29373
rect 9186 29052 9310 29080
rect 3580 28872 3876 28892
rect 3636 28870 3660 28872
rect 3716 28870 3740 28872
rect 3796 28870 3820 28872
rect 3658 28818 3660 28870
rect 3722 28818 3734 28870
rect 3796 28818 3798 28870
rect 3636 28816 3660 28818
rect 3716 28816 3740 28818
rect 3796 28816 3820 28818
rect 3580 28796 3876 28816
rect 8908 28872 9204 28892
rect 8964 28870 8988 28872
rect 9044 28870 9068 28872
rect 9124 28870 9148 28872
rect 8986 28818 8988 28870
rect 9050 28818 9062 28870
rect 9124 28818 9126 28870
rect 8964 28816 8988 28818
rect 9044 28816 9068 28818
rect 9124 28816 9148 28818
rect 8908 28796 9204 28816
rect 9282 28543 9310 29052
rect 9270 28537 9322 28543
rect 9270 28479 9322 28485
rect 2022 28315 2074 28321
rect 2502 28315 2554 28321
rect 2074 28263 2398 28266
rect 2022 28257 2398 28263
rect 2982 28315 3034 28321
rect 2554 28263 2878 28266
rect 2502 28257 2878 28263
rect 3462 28315 3514 28321
rect 3034 28263 3262 28266
rect 2982 28257 3262 28263
rect 3942 28315 3994 28321
rect 3514 28275 3838 28303
rect 3462 28257 3514 28263
rect 2034 28238 2398 28257
rect 2514 28238 2878 28257
rect 2994 28238 3262 28257
rect 2370 28210 2398 28238
rect 2850 28210 2878 28238
rect 1878 28204 1930 28210
rect 1878 28146 1930 28152
rect 2358 28204 2410 28210
rect 2358 28146 2410 28152
rect 2838 28204 2890 28210
rect 3234 28192 3262 28238
rect 3810 28210 3838 28275
rect 4422 28315 4474 28321
rect 3994 28275 4318 28303
rect 3942 28257 3994 28263
rect 4290 28210 4318 28275
rect 4902 28315 4954 28321
rect 4474 28275 4798 28303
rect 4422 28257 4474 28263
rect 4770 28210 4798 28275
rect 5382 28315 5434 28321
rect 4954 28275 5324 28303
rect 4902 28257 4954 28263
rect 5296 28210 5324 28275
rect 7350 28315 7402 28321
rect 5434 28275 5806 28303
rect 5382 28257 5434 28263
rect 5778 28210 5806 28275
rect 5910 28278 5962 28284
rect 6390 28278 6442 28284
rect 5962 28238 6286 28266
rect 5910 28220 5962 28226
rect 6258 28210 6286 28238
rect 6870 28278 6922 28284
rect 6442 28238 6814 28266
rect 6390 28220 6442 28226
rect 6786 28210 6814 28238
rect 6922 28238 7294 28266
rect 7830 28315 7882 28321
rect 7402 28275 7774 28303
rect 7350 28257 7402 28263
rect 6870 28220 6922 28226
rect 7266 28210 7294 28238
rect 7746 28210 7774 28275
rect 8310 28315 8362 28321
rect 7882 28275 8254 28303
rect 7830 28257 7882 28263
rect 8226 28210 8254 28275
rect 8790 28315 8842 28321
rect 8362 28275 8734 28303
rect 8310 28257 8362 28263
rect 8706 28210 8734 28275
rect 8842 28275 9214 28303
rect 8790 28257 8842 28263
rect 9186 28210 9214 28275
rect 3318 28204 3370 28210
rect 3234 28164 3318 28192
rect 2838 28146 2890 28152
rect 3318 28146 3370 28152
rect 3798 28204 3850 28210
rect 3798 28146 3850 28152
rect 4278 28204 4330 28210
rect 4278 28146 4330 28152
rect 4758 28204 4810 28210
rect 4758 28146 4810 28152
rect 5284 28204 5336 28210
rect 5284 28146 5336 28152
rect 5766 28204 5818 28210
rect 5766 28146 5818 28152
rect 6246 28204 6298 28210
rect 6246 28146 6298 28152
rect 6774 28204 6826 28210
rect 6774 28146 6826 28152
rect 7254 28204 7306 28210
rect 7254 28146 7306 28152
rect 7734 28204 7786 28210
rect 7734 28146 7786 28152
rect 8214 28204 8266 28210
rect 8214 28146 8266 28152
rect 8694 28204 8746 28210
rect 8694 28146 8746 28152
rect 9174 28204 9226 28210
rect 9174 28146 9226 28152
rect 1890 27896 1918 28146
rect 1890 27868 2014 27896
rect 1986 26971 2014 27868
rect 6244 27540 6540 27560
rect 6300 27538 6324 27540
rect 6380 27538 6404 27540
rect 6460 27538 6484 27540
rect 6322 27486 6324 27538
rect 6386 27486 6398 27538
rect 6460 27486 6462 27538
rect 6300 27484 6324 27486
rect 6380 27484 6404 27486
rect 6460 27484 6484 27486
rect 6244 27464 6540 27484
rect 5286 27057 5338 27063
rect 5286 26999 5338 27005
rect 5910 27057 5962 27063
rect 5910 26999 5962 27005
rect 6269 27057 6321 27063
rect 6269 26999 6321 27005
rect 6870 27057 6922 27063
rect 6870 26999 6922 27005
rect 4758 26983 4810 26989
rect 1986 26943 2062 26971
rect 1878 26872 1930 26878
rect 1878 26814 1930 26820
rect 1890 26735 1918 26814
rect 2034 26767 2062 26943
rect 4758 26925 4810 26931
rect 4770 26878 4798 26925
rect 5298 26878 5326 26999
rect 5382 26983 5434 26989
rect 5382 26925 5434 26931
rect 5785 26983 5837 26989
rect 5785 26925 5837 26931
rect 2406 26872 2458 26878
rect 2886 26872 2938 26878
rect 2458 26832 2782 26860
rect 2406 26814 2458 26820
rect 2754 26786 2782 26832
rect 3366 26872 3418 26878
rect 2938 26832 3262 26860
rect 2886 26814 2938 26820
rect 3234 26786 3262 26832
rect 3849 26872 3901 26878
rect 3418 26832 3742 26860
rect 3366 26814 3418 26820
rect 2754 26767 3022 26786
rect 3234 26767 3502 26786
rect 2022 26761 2074 26767
rect 1876 26726 1932 26735
rect 2754 26761 3034 26767
rect 2754 26758 2982 26761
rect 2022 26703 2074 26709
rect 2500 26726 2556 26735
rect 1876 26661 1932 26670
rect 3234 26761 3514 26767
rect 3234 26758 3462 26761
rect 2982 26703 3034 26709
rect 3714 26749 3742 26832
rect 4333 26872 4385 26878
rect 3901 26832 4222 26860
rect 3849 26814 3901 26820
rect 3942 26761 3994 26767
rect 3714 26721 3942 26749
rect 3462 26703 3514 26709
rect 4194 26749 4222 26832
rect 4758 26872 4810 26878
rect 4385 26832 4702 26860
rect 4333 26814 4385 26820
rect 4674 26786 4702 26832
rect 4758 26814 4810 26820
rect 5286 26872 5338 26878
rect 5286 26814 5338 26820
rect 4674 26767 4942 26786
rect 5394 26767 5422 26925
rect 5797 26878 5825 26925
rect 5785 26872 5837 26878
rect 5785 26814 5837 26820
rect 5922 26804 5950 26999
rect 6281 26878 6309 26999
rect 6390 26983 6442 26989
rect 6390 26925 6442 26931
rect 6774 26983 6826 26989
rect 6774 26925 6826 26931
rect 6269 26872 6321 26878
rect 6269 26814 6321 26820
rect 6402 26804 6430 26925
rect 6786 26878 6814 26925
rect 6774 26872 6826 26878
rect 6774 26814 6826 26820
rect 6882 26804 6910 26999
rect 7350 26983 7402 26989
rect 7350 26925 7402 26931
rect 8694 26983 8746 26989
rect 8694 26925 8746 26931
rect 9270 26983 9322 26989
rect 9270 26925 9322 26931
rect 7254 26872 7306 26878
rect 7254 26814 7306 26820
rect 5910 26798 5962 26804
rect 4422 26761 4474 26767
rect 4194 26721 4422 26749
rect 3942 26703 3994 26709
rect 4674 26761 4954 26767
rect 4674 26758 4902 26761
rect 4422 26703 4474 26709
rect 4902 26703 4954 26709
rect 5382 26761 5434 26767
rect 5910 26740 5962 26746
rect 6390 26798 6442 26804
rect 6390 26740 6442 26746
rect 6870 26798 6922 26804
rect 6870 26740 6922 26746
rect 5382 26703 5434 26709
rect 2500 26661 2502 26670
rect 2554 26661 2556 26670
rect 2502 26629 2554 26635
rect 7266 26564 7294 26814
rect 7362 26767 7390 26925
rect 8706 26878 8734 26925
rect 7734 26872 7786 26878
rect 8214 26872 8266 26878
rect 7786 26832 8158 26860
rect 7734 26814 7786 26820
rect 7350 26761 7402 26767
rect 8130 26749 8158 26832
rect 8694 26872 8746 26878
rect 8266 26832 8638 26860
rect 8214 26814 8266 26820
rect 8610 26786 8638 26832
rect 8694 26814 8746 26820
rect 9174 26872 9226 26878
rect 9174 26814 9226 26820
rect 8610 26767 8830 26786
rect 8310 26761 8362 26767
rect 8130 26721 8310 26749
rect 7350 26703 7402 26709
rect 8610 26761 8842 26767
rect 8610 26758 8790 26761
rect 8310 26703 8362 26709
rect 8790 26703 8842 26709
rect 7830 26687 7882 26693
rect 7830 26629 7882 26635
rect 7842 26564 7870 26629
rect 7266 26536 7870 26564
rect 9186 26416 9214 26814
rect 9282 26767 9310 26925
rect 9270 26761 9322 26767
rect 9270 26703 9322 26709
rect 9186 26388 9310 26416
rect 3580 26208 3876 26228
rect 3636 26206 3660 26208
rect 3716 26206 3740 26208
rect 3796 26206 3820 26208
rect 3658 26154 3660 26206
rect 3722 26154 3734 26206
rect 3796 26154 3798 26206
rect 3636 26152 3660 26154
rect 3716 26152 3740 26154
rect 3796 26152 3820 26154
rect 3580 26132 3876 26152
rect 8908 26208 9204 26228
rect 8964 26206 8988 26208
rect 9044 26206 9068 26208
rect 9124 26206 9148 26208
rect 8986 26154 8988 26206
rect 9050 26154 9062 26206
rect 9124 26154 9126 26206
rect 8964 26152 8988 26154
rect 9044 26152 9068 26154
rect 9124 26152 9148 26154
rect 8908 26132 9204 26152
rect 9282 25879 9310 26388
rect 9270 25873 9322 25879
rect 9270 25815 9322 25821
rect 2022 25651 2074 25657
rect 2502 25651 2554 25657
rect 2074 25599 2398 25602
rect 2022 25593 2398 25599
rect 2982 25651 3034 25657
rect 2554 25599 2878 25602
rect 2502 25593 2878 25599
rect 3462 25651 3514 25657
rect 3034 25599 3262 25602
rect 2982 25593 3262 25599
rect 3942 25651 3994 25657
rect 3514 25611 3838 25639
rect 3462 25593 3514 25599
rect 2034 25574 2398 25593
rect 2514 25574 2878 25593
rect 2994 25574 3262 25593
rect 2370 25546 2398 25574
rect 2850 25546 2878 25574
rect 1926 25540 1978 25546
rect 2358 25540 2410 25546
rect 1978 25500 2110 25528
rect 1926 25482 1978 25488
rect 2082 24344 2110 25500
rect 2358 25482 2410 25488
rect 2838 25540 2890 25546
rect 3234 25528 3262 25574
rect 3810 25546 3838 25611
rect 4422 25651 4474 25657
rect 3994 25611 4318 25639
rect 3942 25593 3994 25599
rect 4290 25546 4318 25611
rect 4902 25651 4954 25657
rect 4474 25611 4798 25639
rect 4422 25593 4474 25599
rect 4770 25546 4798 25611
rect 5382 25651 5434 25657
rect 4954 25611 5324 25639
rect 4902 25593 4954 25599
rect 5296 25546 5324 25611
rect 7350 25651 7402 25657
rect 5434 25611 5806 25639
rect 5382 25593 5434 25599
rect 5778 25546 5806 25611
rect 5910 25614 5962 25620
rect 6390 25614 6442 25620
rect 5962 25574 6286 25602
rect 5910 25556 5962 25562
rect 6258 25546 6286 25574
rect 6870 25614 6922 25620
rect 6442 25574 6814 25602
rect 6390 25556 6442 25562
rect 6786 25546 6814 25574
rect 6922 25574 7294 25602
rect 7830 25651 7882 25657
rect 7402 25611 7774 25639
rect 7350 25593 7402 25599
rect 6870 25556 6922 25562
rect 7266 25546 7294 25574
rect 7746 25546 7774 25611
rect 8310 25651 8362 25657
rect 7882 25611 8254 25639
rect 7830 25593 7882 25599
rect 8226 25546 8254 25611
rect 8790 25651 8842 25657
rect 8362 25611 8734 25639
rect 8310 25593 8362 25599
rect 8706 25546 8734 25611
rect 8842 25611 9214 25639
rect 8790 25593 8842 25599
rect 9186 25546 9214 25611
rect 3318 25540 3370 25546
rect 3234 25500 3318 25528
rect 2838 25482 2890 25488
rect 3318 25482 3370 25488
rect 3798 25540 3850 25546
rect 3798 25482 3850 25488
rect 4278 25540 4330 25546
rect 4278 25482 4330 25488
rect 4758 25540 4810 25546
rect 4758 25482 4810 25488
rect 5284 25540 5336 25546
rect 5284 25482 5336 25488
rect 5766 25540 5818 25546
rect 5766 25482 5818 25488
rect 6246 25540 6298 25546
rect 6246 25482 6298 25488
rect 6774 25540 6826 25546
rect 6774 25482 6826 25488
rect 7254 25540 7306 25546
rect 7254 25482 7306 25488
rect 7734 25540 7786 25546
rect 7734 25482 7786 25488
rect 8214 25540 8266 25546
rect 8214 25482 8266 25488
rect 8694 25540 8746 25546
rect 8694 25482 8746 25488
rect 9174 25540 9226 25546
rect 9174 25482 9226 25488
rect 6244 24876 6540 24896
rect 6300 24874 6324 24876
rect 6380 24874 6404 24876
rect 6460 24874 6484 24876
rect 6322 24822 6324 24874
rect 6386 24822 6398 24874
rect 6460 24822 6462 24874
rect 6300 24820 6324 24822
rect 6380 24820 6404 24822
rect 6460 24820 6484 24822
rect 6244 24800 6540 24820
rect 2034 24316 2110 24344
rect 5785 24319 5837 24325
rect 1878 24208 1930 24214
rect 1878 24150 1930 24156
rect 1890 24071 1918 24150
rect 2034 24103 2062 24316
rect 5785 24261 5837 24267
rect 9090 24316 9310 24344
rect 2406 24208 2458 24214
rect 2886 24208 2938 24214
rect 2458 24168 2782 24196
rect 2406 24150 2458 24156
rect 2022 24097 2074 24103
rect 1876 24062 1932 24071
rect 2022 24039 2074 24045
rect 2500 24062 2556 24071
rect 1876 23997 1932 24006
rect 2754 24048 2782 24168
rect 3366 24208 3418 24214
rect 2938 24168 3262 24196
rect 2886 24150 2938 24156
rect 3234 24048 3262 24168
rect 3849 24208 3901 24214
rect 3418 24168 3742 24196
rect 3366 24150 3418 24156
rect 2754 24029 3022 24048
rect 3234 24029 3502 24048
rect 2754 24023 3034 24029
rect 2754 24020 2982 24023
rect 2500 23997 2502 24006
rect 2554 23997 2556 24006
rect 2502 23965 2554 23971
rect 3234 24023 3514 24029
rect 3234 24020 3462 24023
rect 2982 23965 3034 23971
rect 3714 24011 3742 24168
rect 4333 24208 4385 24214
rect 3901 24168 4222 24196
rect 3849 24150 3901 24156
rect 4194 24048 4222 24168
rect 4817 24208 4869 24214
rect 4385 24168 4606 24196
rect 4333 24150 4385 24156
rect 4194 24029 4462 24048
rect 3942 24023 3994 24029
rect 3714 23983 3942 24011
rect 3462 23965 3514 23971
rect 4194 24023 4474 24029
rect 4194 24020 4422 24023
rect 3942 23965 3994 23971
rect 4578 24011 4606 24168
rect 5299 24210 5355 24219
rect 5797 24214 5825 24261
rect 6390 24245 6442 24251
rect 4869 24168 5182 24196
rect 4817 24150 4869 24156
rect 4902 24023 4954 24029
rect 4578 23983 4902 24011
rect 4422 23965 4474 23971
rect 5154 24011 5182 24168
rect 5299 24145 5355 24154
rect 5785 24208 5837 24214
rect 5785 24150 5837 24156
rect 5908 24210 5964 24219
rect 5908 24145 5964 24154
rect 6269 24208 6321 24214
rect 6321 24156 6334 24196
rect 6390 24187 6442 24193
rect 6774 24208 6826 24214
rect 6269 24150 6334 24156
rect 5382 24023 5434 24029
rect 5154 23983 5382 24011
rect 4902 23965 4954 23971
rect 5382 23965 5434 23971
rect 5922 23844 5950 24145
rect 5910 23838 5962 23844
rect 5910 23780 5962 23786
rect 6306 23733 6334 24150
rect 6402 24140 6430 24187
rect 7254 24208 7306 24214
rect 6826 24168 7198 24196
rect 6774 24150 6826 24156
rect 6390 24134 6442 24140
rect 6390 24076 6442 24082
rect 7170 24048 7198 24168
rect 7732 24210 7788 24219
rect 7306 24168 7678 24196
rect 7254 24150 7306 24156
rect 7170 24029 7390 24048
rect 7170 24023 7402 24029
rect 7170 24020 7350 24023
rect 7650 24011 7678 24168
rect 7732 24145 7788 24154
rect 8214 24208 8266 24214
rect 8214 24150 8266 24156
rect 8308 24210 8364 24219
rect 7830 24023 7882 24029
rect 7650 23983 7830 24011
rect 7350 23965 7402 23971
rect 8226 24011 8254 24150
rect 8308 24145 8364 24154
rect 8694 24208 8746 24214
rect 9090 24196 9118 24316
rect 8746 24168 9118 24196
rect 9174 24208 9226 24214
rect 8694 24150 8746 24156
rect 9174 24150 9226 24156
rect 8322 24103 8350 24145
rect 8310 24097 8362 24103
rect 8310 24039 8362 24045
rect 8790 24023 8842 24029
rect 8226 23983 8790 24011
rect 7830 23965 7882 23971
rect 8790 23965 8842 23971
rect 6870 23838 6922 23844
rect 6870 23780 6922 23786
rect 6882 23733 6910 23780
rect 9186 23752 9214 24150
rect 9282 24103 9310 24316
rect 9270 24097 9322 24103
rect 9270 24039 9322 24045
rect 6294 23727 6346 23733
rect 6294 23669 6346 23675
rect 6870 23727 6922 23733
rect 9186 23724 9310 23752
rect 6870 23669 6922 23675
rect 3580 23544 3876 23564
rect 3636 23542 3660 23544
rect 3716 23542 3740 23544
rect 3796 23542 3820 23544
rect 3658 23490 3660 23542
rect 3722 23490 3734 23542
rect 3796 23490 3798 23542
rect 3636 23488 3660 23490
rect 3716 23488 3740 23490
rect 3796 23488 3820 23490
rect 3580 23468 3876 23488
rect 8908 23544 9204 23564
rect 8964 23542 8988 23544
rect 9044 23542 9068 23544
rect 9124 23542 9148 23544
rect 8986 23490 8988 23542
rect 9050 23490 9062 23542
rect 9124 23490 9126 23542
rect 8964 23488 8988 23490
rect 9044 23488 9068 23490
rect 9124 23488 9148 23490
rect 8908 23468 9204 23488
rect 6390 23246 6442 23252
rect 9282 23215 9310 23724
rect 6390 23188 6442 23194
rect 9270 23209 9322 23215
rect 6402 23160 6430 23188
rect 3954 23141 4318 23160
rect 5394 23141 5806 23160
rect 3942 23135 4318 23141
rect 3994 23132 4318 23135
rect 3942 23077 3994 23083
rect 2022 22987 2074 22993
rect 2502 22987 2554 22993
rect 2074 22935 2398 22938
rect 2022 22929 2398 22935
rect 2982 22987 3034 22993
rect 2554 22935 2878 22938
rect 2502 22929 2878 22935
rect 3462 22987 3514 22993
rect 3034 22935 3262 22938
rect 2982 22929 3262 22935
rect 3514 22947 3838 22975
rect 3462 22929 3514 22935
rect 2034 22910 2398 22929
rect 2514 22910 2878 22929
rect 2994 22910 3262 22929
rect 2370 22882 2398 22910
rect 2850 22882 2878 22910
rect 1878 22876 1930 22882
rect 1794 22836 1878 22864
rect 1108 21546 1164 21555
rect 1108 21481 1164 21490
rect 1274 21470 1326 21476
rect 1794 21458 1822 22836
rect 1878 22818 1930 22824
rect 2358 22876 2410 22882
rect 2358 22818 2410 22824
rect 2838 22876 2890 22882
rect 3234 22864 3262 22910
rect 3810 22882 3838 22947
rect 4290 22938 4318 23132
rect 5382 23135 5806 23141
rect 5434 23132 5806 23135
rect 6402 23132 6814 23160
rect 7842 23141 8158 23160
rect 9270 23151 9322 23157
rect 5382 23077 5434 23083
rect 4422 22987 4474 22993
rect 4290 22910 4356 22938
rect 4902 22987 4954 22993
rect 4474 22947 4798 22975
rect 4422 22929 4474 22935
rect 4328 22882 4356 22910
rect 4770 22882 4798 22947
rect 4954 22947 5324 22975
rect 4902 22929 4954 22935
rect 5296 22882 5324 22947
rect 5778 22882 5806 23132
rect 5910 22950 5962 22956
rect 5962 22910 6286 22938
rect 5910 22892 5962 22898
rect 6258 22882 6286 22910
rect 6786 22882 6814 23132
rect 7830 23135 8158 23141
rect 7882 23132 8158 23135
rect 7830 23077 7882 23083
rect 7350 22987 7402 22993
rect 6870 22950 6922 22956
rect 6922 22910 7294 22938
rect 7402 22947 7774 22975
rect 7350 22929 7402 22935
rect 6870 22892 6922 22898
rect 7266 22882 7294 22910
rect 7746 22882 7774 22947
rect 8130 22938 8158 23132
rect 8310 22987 8362 22993
rect 8130 22910 8206 22938
rect 8790 22987 8842 22993
rect 8362 22947 8734 22975
rect 8310 22929 8362 22935
rect 8178 22882 8206 22910
rect 8706 22882 8734 22947
rect 8842 22947 9214 22975
rect 8790 22929 8842 22935
rect 9186 22882 9214 22947
rect 3318 22876 3370 22882
rect 3234 22836 3318 22864
rect 2838 22818 2890 22824
rect 3318 22818 3370 22824
rect 3798 22876 3850 22882
rect 3798 22818 3850 22824
rect 4316 22876 4368 22882
rect 4316 22818 4368 22824
rect 4758 22876 4810 22882
rect 4758 22818 4810 22824
rect 5284 22876 5336 22882
rect 5284 22818 5336 22824
rect 5766 22876 5818 22882
rect 5766 22818 5818 22824
rect 6246 22876 6298 22882
rect 6246 22818 6298 22824
rect 6774 22876 6826 22882
rect 6774 22818 6826 22824
rect 7254 22876 7306 22882
rect 7254 22818 7306 22824
rect 7734 22876 7786 22882
rect 7734 22818 7786 22824
rect 8166 22876 8218 22882
rect 8166 22818 8218 22824
rect 8694 22876 8746 22882
rect 8694 22818 8746 22824
rect 9174 22876 9226 22882
rect 9174 22818 9226 22824
rect 6244 22212 6540 22232
rect 6300 22210 6324 22212
rect 6380 22210 6404 22212
rect 6460 22210 6484 22212
rect 6322 22158 6324 22210
rect 6386 22158 6398 22210
rect 6460 22158 6462 22210
rect 6300 22156 6324 22158
rect 6380 22156 6404 22158
rect 6460 22156 6484 22158
rect 6244 22136 6540 22156
rect 5286 21729 5338 21735
rect 5286 21671 5338 21677
rect 5910 21729 5962 21735
rect 5910 21671 5962 21677
rect 6269 21729 6321 21735
rect 6269 21671 6321 21677
rect 6870 21729 6922 21735
rect 6870 21671 6922 21677
rect 4758 21655 4810 21661
rect 4758 21597 4810 21603
rect 4770 21550 4798 21597
rect 5298 21550 5326 21671
rect 5382 21655 5434 21661
rect 5382 21597 5434 21603
rect 5785 21655 5837 21661
rect 5785 21597 5837 21603
rect 1926 21544 1978 21550
rect 2406 21544 2458 21550
rect 1978 21504 2302 21532
rect 1926 21486 1978 21492
rect 1274 21412 1326 21418
rect 1362 21430 1822 21458
rect 2274 21458 2302 21504
rect 2886 21544 2938 21550
rect 2458 21504 2782 21532
rect 2406 21486 2458 21492
rect 2754 21458 2782 21504
rect 3366 21544 3418 21550
rect 2938 21504 3262 21532
rect 2886 21486 2938 21492
rect 3234 21458 3262 21504
rect 3849 21544 3901 21550
rect 3418 21504 3742 21532
rect 3366 21486 3418 21492
rect 3714 21458 3742 21504
rect 4333 21544 4385 21550
rect 3901 21504 4222 21532
rect 3849 21486 3901 21492
rect 4194 21458 4222 21504
rect 4758 21544 4810 21550
rect 4385 21504 4702 21532
rect 4333 21486 4385 21492
rect 4674 21458 4702 21504
rect 4758 21486 4810 21492
rect 5286 21544 5338 21550
rect 5286 21486 5338 21492
rect 2274 21439 2542 21458
rect 2754 21439 3022 21458
rect 3234 21439 3502 21458
rect 3714 21439 3982 21458
rect 4194 21439 4462 21458
rect 4674 21439 4942 21458
rect 5394 21439 5422 21597
rect 5797 21550 5825 21597
rect 5785 21544 5837 21550
rect 5785 21486 5837 21492
rect 5922 21476 5950 21671
rect 6281 21550 6309 21671
rect 6390 21655 6442 21661
rect 6390 21597 6442 21603
rect 6774 21655 6826 21661
rect 6774 21597 6826 21603
rect 6269 21544 6321 21550
rect 6269 21486 6321 21492
rect 6402 21476 6430 21597
rect 6786 21550 6814 21597
rect 6774 21544 6826 21550
rect 6774 21486 6826 21492
rect 6882 21476 6910 21671
rect 7350 21655 7402 21661
rect 7350 21597 7402 21603
rect 8694 21655 8746 21661
rect 8694 21597 8746 21603
rect 9270 21655 9322 21661
rect 9270 21597 9322 21603
rect 7254 21544 7306 21550
rect 7254 21486 7306 21492
rect 5910 21470 5962 21476
rect 2274 21433 2554 21439
rect 2274 21430 2502 21433
rect 1286 21236 1314 21412
rect 1362 21328 1390 21430
rect 1452 21396 1504 21402
rect 1504 21365 2062 21384
rect 2754 21433 3034 21439
rect 2754 21430 2982 21433
rect 2502 21375 2554 21381
rect 3234 21433 3514 21439
rect 3234 21430 3462 21433
rect 2982 21375 3034 21381
rect 3714 21433 3994 21439
rect 3714 21430 3942 21433
rect 3462 21375 3514 21381
rect 4194 21433 4474 21439
rect 4194 21430 4422 21433
rect 3942 21375 3994 21381
rect 4674 21433 4954 21439
rect 4674 21430 4902 21433
rect 4422 21375 4474 21381
rect 4902 21375 4954 21381
rect 5382 21433 5434 21439
rect 5910 21412 5962 21418
rect 6390 21470 6442 21476
rect 6390 21412 6442 21418
rect 6870 21470 6922 21476
rect 6870 21412 6922 21418
rect 5382 21375 5434 21381
rect 1504 21359 2074 21365
rect 1504 21356 2022 21359
rect 1452 21338 1504 21344
rect 1350 21322 1402 21328
rect 2022 21301 2074 21307
rect 1350 21264 1402 21270
rect 7266 21236 7294 21486
rect 7362 21439 7390 21597
rect 8706 21550 8734 21597
rect 7734 21544 7786 21550
rect 8214 21544 8266 21550
rect 7786 21504 8158 21532
rect 7734 21486 7786 21492
rect 8130 21458 8158 21504
rect 8694 21544 8746 21550
rect 8266 21504 8638 21532
rect 8214 21486 8266 21492
rect 8610 21458 8638 21504
rect 8694 21486 8746 21492
rect 9174 21544 9226 21550
rect 9174 21486 9226 21492
rect 8130 21439 8350 21458
rect 8610 21439 8830 21458
rect 7350 21433 7402 21439
rect 8130 21433 8362 21439
rect 8130 21430 8310 21433
rect 7350 21375 7402 21381
rect 8610 21433 8842 21439
rect 8610 21430 8790 21433
rect 8310 21375 8362 21381
rect 8790 21375 8842 21381
rect 7830 21285 7882 21291
rect 1286 21208 1342 21236
rect 7266 21233 7830 21236
rect 7266 21227 7882 21233
rect 7266 21208 7870 21227
rect 1314 21069 1342 21208
rect 9186 21088 9214 21486
rect 9282 21439 9310 21597
rect 9270 21433 9322 21439
rect 9270 21375 9322 21381
rect 1302 21063 1354 21069
rect 1302 21005 1354 21011
rect 1782 21063 1834 21069
rect 9186 21060 9310 21088
rect 1782 21005 1834 21011
rect 1794 1552 1822 21005
rect 3580 20880 3876 20900
rect 3636 20878 3660 20880
rect 3716 20878 3740 20880
rect 3796 20878 3820 20880
rect 3658 20826 3660 20878
rect 3722 20826 3734 20878
rect 3796 20826 3798 20878
rect 3636 20824 3660 20826
rect 3716 20824 3740 20826
rect 3796 20824 3820 20826
rect 3580 20804 3876 20824
rect 8908 20880 9204 20900
rect 8964 20878 8988 20880
rect 9044 20878 9068 20880
rect 9124 20878 9148 20880
rect 8986 20826 8988 20878
rect 9050 20826 9062 20878
rect 9124 20826 9126 20878
rect 8964 20824 8988 20826
rect 9044 20824 9068 20826
rect 9124 20824 9148 20826
rect 8908 20804 9204 20824
rect 9282 20551 9310 21060
rect 9270 20545 9322 20551
rect 9270 20487 9322 20493
rect 2022 20323 2074 20329
rect 2502 20323 2554 20329
rect 2074 20271 2398 20274
rect 2022 20265 2398 20271
rect 2982 20323 3034 20329
rect 2554 20271 2878 20274
rect 2502 20265 2878 20271
rect 3462 20323 3514 20329
rect 3034 20271 3262 20274
rect 2982 20265 3262 20271
rect 3942 20323 3994 20329
rect 3514 20283 3838 20311
rect 3462 20265 3514 20271
rect 2034 20246 2398 20265
rect 2514 20246 2878 20265
rect 2994 20246 3262 20265
rect 2370 20218 2398 20246
rect 2850 20218 2878 20246
rect 1878 20212 1930 20218
rect 1878 20154 1930 20160
rect 2358 20212 2410 20218
rect 2358 20154 2410 20160
rect 2838 20212 2890 20218
rect 3234 20200 3262 20246
rect 3810 20218 3838 20283
rect 4422 20323 4474 20329
rect 3994 20283 4318 20311
rect 3942 20265 3994 20271
rect 4290 20218 4318 20283
rect 4902 20323 4954 20329
rect 4474 20283 4798 20311
rect 4422 20265 4474 20271
rect 4770 20218 4798 20283
rect 5382 20323 5434 20329
rect 4954 20283 5324 20311
rect 4902 20265 4954 20271
rect 5296 20218 5324 20283
rect 7350 20323 7402 20329
rect 5434 20283 5806 20311
rect 5382 20265 5434 20271
rect 5778 20218 5806 20283
rect 5910 20286 5962 20292
rect 6390 20286 6442 20292
rect 5962 20246 6286 20274
rect 5910 20228 5962 20234
rect 6258 20218 6286 20246
rect 6870 20286 6922 20292
rect 6442 20246 6814 20274
rect 6390 20228 6442 20234
rect 6786 20218 6814 20246
rect 6922 20246 7294 20274
rect 7830 20323 7882 20329
rect 7402 20283 7774 20311
rect 7350 20265 7402 20271
rect 6870 20228 6922 20234
rect 7266 20218 7294 20246
rect 7746 20218 7774 20283
rect 8310 20323 8362 20329
rect 7882 20283 8254 20311
rect 7830 20265 7882 20271
rect 8226 20218 8254 20283
rect 8790 20323 8842 20329
rect 8362 20283 8734 20311
rect 8310 20265 8362 20271
rect 8706 20218 8734 20283
rect 8842 20283 9214 20311
rect 8790 20265 8842 20271
rect 9186 20218 9214 20283
rect 3318 20212 3370 20218
rect 3234 20172 3318 20200
rect 2838 20154 2890 20160
rect 3318 20154 3370 20160
rect 3798 20212 3850 20218
rect 3798 20154 3850 20160
rect 4278 20212 4330 20218
rect 4278 20154 4330 20160
rect 4758 20212 4810 20218
rect 4758 20154 4810 20160
rect 5284 20212 5336 20218
rect 5284 20154 5336 20160
rect 5766 20212 5818 20218
rect 5766 20154 5818 20160
rect 6246 20212 6298 20218
rect 6246 20154 6298 20160
rect 6774 20212 6826 20218
rect 6774 20154 6826 20160
rect 7254 20212 7306 20218
rect 7254 20154 7306 20160
rect 7734 20212 7786 20218
rect 7734 20154 7786 20160
rect 8214 20212 8266 20218
rect 8214 20154 8266 20160
rect 8694 20212 8746 20218
rect 8694 20154 8746 20160
rect 9174 20212 9226 20218
rect 9174 20154 9226 20160
rect 1890 18979 1918 20154
rect 6244 19548 6540 19568
rect 6300 19546 6324 19548
rect 6380 19546 6404 19548
rect 6460 19546 6484 19548
rect 6322 19494 6324 19546
rect 6386 19494 6398 19546
rect 6460 19494 6462 19546
rect 6300 19492 6324 19494
rect 6380 19492 6404 19494
rect 6460 19492 6484 19494
rect 6244 19472 6540 19492
rect 5286 19065 5338 19071
rect 5286 19007 5338 19013
rect 5910 19065 5962 19071
rect 5910 19007 5962 19013
rect 6269 19065 6321 19071
rect 6269 19007 6321 19013
rect 6870 19065 6922 19071
rect 6870 19007 6922 19013
rect 4758 18991 4810 18997
rect 1890 18951 2062 18979
rect 1878 18880 1930 18886
rect 1878 18822 1930 18828
rect 1890 18743 1918 18822
rect 2034 18775 2062 18951
rect 4758 18933 4810 18939
rect 4770 18886 4798 18933
rect 5298 18886 5326 19007
rect 5382 18991 5434 18997
rect 5382 18933 5434 18939
rect 5785 18991 5837 18997
rect 5785 18933 5837 18939
rect 2406 18880 2458 18886
rect 2886 18880 2938 18886
rect 2458 18840 2782 18868
rect 2406 18822 2458 18828
rect 2754 18794 2782 18840
rect 3366 18880 3418 18886
rect 2938 18840 3262 18868
rect 2886 18822 2938 18828
rect 3234 18794 3262 18840
rect 3849 18880 3901 18886
rect 3418 18840 3742 18868
rect 3366 18822 3418 18828
rect 2754 18775 3022 18794
rect 3234 18775 3502 18794
rect 2022 18769 2074 18775
rect 1876 18734 1932 18743
rect 2754 18769 3034 18775
rect 2754 18766 2982 18769
rect 2022 18711 2074 18717
rect 2500 18734 2556 18743
rect 1876 18669 1932 18678
rect 3234 18769 3514 18775
rect 3234 18766 3462 18769
rect 2982 18711 3034 18717
rect 3714 18757 3742 18840
rect 4333 18880 4385 18886
rect 3901 18840 4222 18868
rect 3849 18822 3901 18828
rect 4194 18794 4222 18840
rect 4758 18880 4810 18886
rect 4385 18840 4702 18868
rect 4333 18822 4385 18828
rect 4674 18794 4702 18840
rect 4758 18822 4810 18828
rect 5286 18880 5338 18886
rect 5286 18822 5338 18828
rect 4194 18775 4462 18794
rect 4674 18775 4942 18794
rect 5394 18775 5422 18933
rect 5797 18886 5825 18933
rect 5785 18880 5837 18886
rect 5785 18822 5837 18828
rect 5922 18812 5950 19007
rect 6281 18886 6309 19007
rect 6390 18991 6442 18997
rect 6390 18933 6442 18939
rect 6774 18991 6826 18997
rect 6774 18933 6826 18939
rect 6269 18880 6321 18886
rect 6269 18822 6321 18828
rect 6402 18812 6430 18933
rect 6786 18886 6814 18933
rect 6774 18880 6826 18886
rect 6774 18822 6826 18828
rect 6882 18812 6910 19007
rect 7350 18991 7402 18997
rect 7350 18933 7402 18939
rect 8694 18991 8746 18997
rect 8694 18933 8746 18939
rect 9270 18991 9322 18997
rect 9270 18933 9322 18939
rect 7254 18880 7306 18886
rect 7254 18822 7306 18828
rect 5910 18806 5962 18812
rect 3942 18769 3994 18775
rect 3714 18729 3942 18757
rect 3462 18711 3514 18717
rect 4194 18769 4474 18775
rect 4194 18766 4422 18769
rect 3942 18711 3994 18717
rect 4674 18769 4954 18775
rect 4674 18766 4902 18769
rect 4422 18711 4474 18717
rect 4902 18711 4954 18717
rect 5382 18769 5434 18775
rect 5910 18748 5962 18754
rect 6390 18806 6442 18812
rect 6390 18748 6442 18754
rect 6870 18806 6922 18812
rect 6870 18748 6922 18754
rect 5382 18711 5434 18717
rect 2500 18669 2502 18678
rect 2554 18669 2556 18678
rect 2502 18637 2554 18643
rect 7266 18572 7294 18822
rect 7362 18775 7390 18933
rect 8706 18886 8734 18933
rect 7734 18880 7786 18886
rect 8214 18880 8266 18886
rect 7786 18840 8158 18868
rect 7734 18822 7786 18828
rect 7350 18769 7402 18775
rect 8130 18757 8158 18840
rect 8694 18880 8746 18886
rect 8266 18840 8638 18868
rect 8214 18822 8266 18828
rect 8310 18769 8362 18775
rect 8130 18729 8310 18757
rect 7350 18711 7402 18717
rect 8610 18757 8638 18840
rect 8694 18822 8746 18828
rect 9174 18880 9226 18886
rect 9174 18822 9226 18828
rect 8790 18769 8842 18775
rect 8610 18729 8790 18757
rect 8310 18711 8362 18717
rect 8790 18711 8842 18717
rect 7830 18621 7882 18627
rect 7266 18569 7830 18572
rect 7266 18563 7882 18569
rect 7266 18544 7870 18563
rect 9186 18424 9214 18822
rect 9282 18775 9310 18933
rect 9270 18769 9322 18775
rect 9270 18711 9322 18717
rect 9186 18396 9310 18424
rect 3580 18216 3876 18236
rect 3636 18214 3660 18216
rect 3716 18214 3740 18216
rect 3796 18214 3820 18216
rect 3658 18162 3660 18214
rect 3722 18162 3734 18214
rect 3796 18162 3798 18214
rect 3636 18160 3660 18162
rect 3716 18160 3740 18162
rect 3796 18160 3820 18162
rect 3580 18140 3876 18160
rect 8908 18216 9204 18236
rect 8964 18214 8988 18216
rect 9044 18214 9068 18216
rect 9124 18214 9148 18216
rect 8986 18162 8988 18214
rect 9050 18162 9062 18214
rect 9124 18162 9126 18214
rect 8964 18160 8988 18162
rect 9044 18160 9068 18162
rect 9124 18160 9148 18162
rect 8908 18140 9204 18160
rect 9282 17887 9310 18396
rect 9270 17881 9322 17887
rect 9270 17823 9322 17829
rect 2022 17659 2074 17665
rect 2502 17659 2554 17665
rect 2074 17607 2398 17610
rect 2022 17601 2398 17607
rect 2982 17659 3034 17665
rect 2554 17607 2878 17610
rect 2502 17601 2878 17607
rect 3462 17659 3514 17665
rect 3034 17607 3262 17610
rect 2982 17601 3262 17607
rect 3942 17659 3994 17665
rect 3514 17619 3838 17647
rect 3462 17601 3514 17607
rect 2034 17582 2398 17601
rect 2514 17582 2878 17601
rect 2994 17582 3262 17601
rect 2370 17554 2398 17582
rect 2850 17554 2878 17582
rect 1878 17548 1930 17554
rect 1878 17490 1930 17496
rect 2358 17548 2410 17554
rect 2358 17490 2410 17496
rect 2838 17548 2890 17554
rect 3234 17536 3262 17582
rect 3810 17554 3838 17619
rect 4422 17659 4474 17665
rect 3994 17619 4318 17647
rect 3942 17601 3994 17607
rect 4290 17554 4318 17619
rect 4902 17659 4954 17665
rect 4474 17619 4798 17647
rect 4422 17601 4474 17607
rect 4770 17554 4798 17619
rect 5382 17659 5434 17665
rect 4954 17619 5324 17647
rect 4902 17601 4954 17607
rect 5296 17554 5324 17619
rect 7350 17659 7402 17665
rect 5434 17619 5806 17647
rect 5382 17601 5434 17607
rect 5778 17554 5806 17619
rect 5910 17622 5962 17628
rect 6390 17622 6442 17628
rect 5962 17582 6286 17610
rect 5910 17564 5962 17570
rect 6258 17554 6286 17582
rect 6870 17622 6922 17628
rect 6442 17582 6814 17610
rect 6390 17564 6442 17570
rect 6786 17554 6814 17582
rect 6922 17582 7294 17610
rect 7830 17659 7882 17665
rect 7402 17619 7774 17647
rect 7350 17601 7402 17607
rect 6870 17564 6922 17570
rect 7266 17554 7294 17582
rect 7746 17554 7774 17619
rect 8310 17659 8362 17665
rect 7882 17619 8254 17647
rect 7830 17601 7882 17607
rect 8226 17554 8254 17619
rect 8790 17659 8842 17665
rect 8362 17619 8734 17647
rect 8310 17601 8362 17607
rect 8706 17554 8734 17619
rect 8842 17619 9214 17647
rect 8790 17601 8842 17607
rect 9186 17554 9214 17619
rect 3318 17548 3370 17554
rect 3234 17508 3318 17536
rect 2838 17490 2890 17496
rect 3318 17490 3370 17496
rect 3798 17548 3850 17554
rect 3798 17490 3850 17496
rect 4278 17548 4330 17554
rect 4278 17490 4330 17496
rect 4758 17548 4810 17554
rect 4758 17490 4810 17496
rect 5284 17548 5336 17554
rect 5284 17490 5336 17496
rect 5766 17548 5818 17554
rect 5766 17490 5818 17496
rect 6246 17548 6298 17554
rect 6246 17490 6298 17496
rect 6774 17548 6826 17554
rect 6774 17490 6826 17496
rect 7254 17548 7306 17554
rect 7254 17490 7306 17496
rect 7734 17548 7786 17554
rect 7734 17490 7786 17496
rect 8214 17548 8266 17554
rect 8214 17490 8266 17496
rect 8694 17548 8746 17554
rect 8694 17490 8746 17496
rect 9174 17548 9226 17554
rect 9174 17490 9226 17496
rect 1890 16315 1918 17490
rect 6244 16884 6540 16904
rect 6300 16882 6324 16884
rect 6380 16882 6404 16884
rect 6460 16882 6484 16884
rect 6322 16830 6324 16882
rect 6386 16830 6398 16882
rect 6460 16830 6462 16882
rect 6300 16828 6324 16830
rect 6380 16828 6404 16830
rect 6460 16828 6484 16830
rect 6244 16808 6540 16828
rect 5286 16401 5338 16407
rect 5286 16343 5338 16349
rect 5910 16401 5962 16407
rect 5910 16343 5962 16349
rect 6269 16401 6321 16407
rect 6269 16343 6321 16349
rect 6870 16401 6922 16407
rect 6870 16343 6922 16349
rect 4758 16327 4810 16333
rect 1890 16287 2062 16315
rect 1878 16216 1930 16222
rect 1878 16158 1930 16164
rect 1890 16079 1918 16158
rect 2034 16111 2062 16287
rect 4758 16269 4810 16275
rect 4770 16222 4798 16269
rect 5298 16222 5326 16343
rect 5382 16327 5434 16333
rect 5382 16269 5434 16275
rect 5785 16327 5837 16333
rect 5785 16269 5837 16275
rect 2406 16216 2458 16222
rect 2886 16216 2938 16222
rect 2458 16176 2782 16204
rect 2406 16158 2458 16164
rect 2754 16130 2782 16176
rect 3366 16216 3418 16222
rect 2938 16176 3262 16204
rect 2886 16158 2938 16164
rect 3234 16130 3262 16176
rect 3849 16216 3901 16222
rect 3418 16176 3742 16204
rect 3366 16158 3418 16164
rect 3714 16130 3742 16176
rect 4333 16216 4385 16222
rect 3901 16176 4222 16204
rect 3849 16158 3901 16164
rect 4194 16130 4222 16176
rect 4758 16216 4810 16222
rect 4385 16176 4702 16204
rect 4333 16158 4385 16164
rect 4674 16130 4702 16176
rect 4758 16158 4810 16164
rect 5286 16216 5338 16222
rect 5286 16158 5338 16164
rect 2754 16111 3022 16130
rect 3234 16111 3502 16130
rect 3714 16111 3982 16130
rect 4194 16111 4462 16130
rect 4674 16111 4942 16130
rect 5394 16111 5422 16269
rect 5797 16222 5825 16269
rect 5785 16216 5837 16222
rect 5785 16158 5837 16164
rect 5922 16148 5950 16343
rect 6281 16222 6309 16343
rect 6390 16327 6442 16333
rect 6390 16269 6442 16275
rect 6774 16327 6826 16333
rect 6774 16269 6826 16275
rect 6269 16216 6321 16222
rect 6269 16158 6321 16164
rect 6402 16148 6430 16269
rect 6786 16222 6814 16269
rect 6774 16216 6826 16222
rect 6774 16158 6826 16164
rect 6882 16148 6910 16343
rect 7350 16327 7402 16333
rect 7350 16269 7402 16275
rect 8694 16327 8746 16333
rect 8694 16269 8746 16275
rect 9270 16327 9322 16333
rect 9270 16269 9322 16275
rect 7254 16216 7306 16222
rect 7254 16158 7306 16164
rect 5910 16142 5962 16148
rect 2022 16105 2074 16111
rect 1876 16070 1932 16079
rect 2754 16105 3034 16111
rect 2754 16102 2982 16105
rect 2022 16047 2074 16053
rect 2500 16070 2556 16079
rect 1876 16005 1932 16014
rect 3234 16105 3514 16111
rect 3234 16102 3462 16105
rect 2982 16047 3034 16053
rect 3714 16105 3994 16111
rect 3714 16102 3942 16105
rect 3462 16047 3514 16053
rect 4194 16105 4474 16111
rect 4194 16102 4422 16105
rect 3942 16047 3994 16053
rect 4674 16105 4954 16111
rect 4674 16102 4902 16105
rect 4422 16047 4474 16053
rect 4902 16047 4954 16053
rect 5382 16105 5434 16111
rect 5910 16084 5962 16090
rect 6390 16142 6442 16148
rect 6390 16084 6442 16090
rect 6870 16142 6922 16148
rect 6870 16084 6922 16090
rect 5382 16047 5434 16053
rect 2500 16005 2502 16014
rect 2554 16005 2556 16014
rect 2502 15973 2554 15979
rect 7266 15908 7294 16158
rect 7362 16111 7390 16269
rect 8706 16222 8734 16269
rect 7734 16216 7786 16222
rect 8214 16216 8266 16222
rect 7786 16176 8158 16204
rect 7734 16158 7786 16164
rect 7350 16105 7402 16111
rect 7350 16047 7402 16053
rect 8130 16056 8158 16176
rect 8694 16216 8746 16222
rect 8266 16176 8638 16204
rect 8214 16158 8266 16164
rect 8610 16056 8638 16176
rect 8694 16158 8746 16164
rect 9174 16216 9226 16222
rect 9174 16158 9226 16164
rect 8130 16037 8350 16056
rect 8610 16037 8830 16056
rect 7830 16031 7882 16037
rect 8130 16031 8362 16037
rect 8130 16028 8310 16031
rect 7830 15973 7882 15979
rect 8610 16031 8842 16037
rect 8610 16028 8790 16031
rect 8310 15973 8362 15979
rect 8790 15973 8842 15979
rect 7842 15908 7870 15973
rect 7266 15880 7870 15908
rect 9186 15760 9214 16158
rect 9282 16111 9310 16269
rect 9270 16105 9322 16111
rect 9270 16047 9322 16053
rect 9186 15732 9310 15760
rect 3580 15552 3876 15572
rect 3636 15550 3660 15552
rect 3716 15550 3740 15552
rect 3796 15550 3820 15552
rect 3658 15498 3660 15550
rect 3722 15498 3734 15550
rect 3796 15498 3798 15550
rect 3636 15496 3660 15498
rect 3716 15496 3740 15498
rect 3796 15496 3820 15498
rect 3580 15476 3876 15496
rect 8908 15552 9204 15572
rect 8964 15550 8988 15552
rect 9044 15550 9068 15552
rect 9124 15550 9148 15552
rect 8986 15498 8988 15550
rect 9050 15498 9062 15550
rect 9124 15498 9126 15550
rect 8964 15496 8988 15498
rect 9044 15496 9068 15498
rect 9124 15496 9148 15498
rect 8908 15476 9204 15496
rect 9282 15223 9310 15732
rect 9270 15217 9322 15223
rect 9270 15159 9322 15165
rect 2022 14995 2074 15001
rect 2502 14995 2554 15001
rect 2074 14943 2398 14946
rect 2022 14937 2398 14943
rect 2982 14995 3034 15001
rect 2554 14943 2878 14946
rect 2502 14937 2878 14943
rect 3462 14995 3514 15001
rect 3034 14943 3358 14946
rect 2982 14937 3358 14943
rect 3942 14995 3994 15001
rect 3514 14943 3838 14946
rect 3462 14937 3838 14943
rect 4422 14995 4474 15001
rect 3994 14943 4318 14946
rect 3942 14937 4318 14943
rect 4902 14995 4954 15001
rect 4474 14943 4798 14946
rect 4422 14937 4798 14943
rect 5382 14995 5434 15001
rect 4954 14943 5324 14946
rect 4902 14937 5324 14943
rect 7350 14995 7402 15001
rect 5910 14958 5962 14964
rect 5434 14943 5806 14946
rect 5382 14937 5806 14943
rect 2034 14918 2398 14937
rect 2514 14918 2878 14937
rect 2994 14918 3358 14937
rect 3474 14918 3838 14937
rect 3954 14918 4318 14937
rect 4434 14918 4798 14937
rect 4914 14918 5324 14937
rect 5394 14918 5806 14937
rect 2370 14890 2398 14918
rect 2850 14890 2878 14918
rect 3330 14890 3358 14918
rect 3810 14890 3838 14918
rect 4290 14890 4318 14918
rect 4770 14890 4798 14918
rect 5296 14890 5324 14918
rect 5778 14890 5806 14918
rect 6390 14958 6442 14964
rect 5962 14918 6286 14946
rect 5910 14900 5962 14906
rect 6258 14890 6286 14918
rect 6870 14958 6922 14964
rect 6442 14918 6622 14946
rect 6390 14900 6442 14906
rect 1926 14884 1978 14890
rect 2358 14884 2410 14890
rect 1978 14844 2110 14872
rect 1926 14826 1978 14832
rect 2082 13688 2110 14844
rect 2358 14826 2410 14832
rect 2838 14884 2890 14890
rect 2838 14826 2890 14832
rect 3318 14884 3370 14890
rect 3318 14826 3370 14832
rect 3798 14884 3850 14890
rect 3798 14826 3850 14832
rect 4278 14884 4330 14890
rect 4278 14826 4330 14832
rect 4758 14884 4810 14890
rect 4758 14826 4810 14832
rect 5284 14884 5336 14890
rect 5284 14826 5336 14832
rect 5766 14884 5818 14890
rect 5766 14826 5818 14832
rect 6246 14884 6298 14890
rect 6594 14872 6622 14918
rect 7350 14937 7402 14943
rect 7830 14995 7882 15001
rect 7830 14937 7882 14943
rect 8310 14995 8362 15001
rect 8310 14937 8362 14943
rect 8790 14995 8842 15001
rect 8790 14937 8842 14943
rect 6870 14900 6922 14906
rect 6726 14884 6778 14890
rect 6594 14844 6726 14872
rect 6246 14826 6298 14832
rect 6882 14872 6910 14900
rect 7206 14884 7258 14890
rect 6882 14844 7206 14872
rect 6726 14826 6778 14832
rect 7362 14872 7390 14937
rect 7686 14884 7738 14890
rect 7362 14844 7686 14872
rect 7206 14826 7258 14832
rect 7842 14872 7870 14937
rect 8166 14884 8218 14890
rect 7842 14844 8166 14872
rect 7686 14826 7738 14832
rect 8322 14872 8350 14937
rect 8646 14884 8698 14890
rect 8322 14844 8646 14872
rect 8166 14826 8218 14832
rect 8802 14872 8830 14937
rect 9126 14884 9178 14890
rect 8802 14844 9126 14872
rect 8646 14826 8698 14832
rect 9126 14826 9178 14832
rect 6244 14220 6540 14240
rect 6300 14218 6324 14220
rect 6380 14218 6404 14220
rect 6460 14218 6484 14220
rect 6322 14166 6324 14218
rect 6386 14166 6398 14218
rect 6460 14166 6462 14218
rect 6300 14164 6324 14166
rect 6380 14164 6404 14166
rect 6460 14164 6484 14166
rect 6244 14144 6540 14164
rect 2034 13660 2110 13688
rect 5785 13663 5837 13669
rect 1878 13552 1930 13558
rect 1878 13494 1930 13500
rect 1890 13415 1918 13494
rect 2034 13447 2062 13660
rect 5785 13605 5837 13611
rect 9090 13660 9310 13688
rect 2406 13552 2458 13558
rect 2886 13552 2938 13558
rect 2458 13512 2782 13540
rect 2406 13494 2458 13500
rect 2022 13441 2074 13447
rect 1876 13406 1932 13415
rect 2022 13383 2074 13389
rect 2500 13406 2556 13415
rect 1876 13341 1932 13350
rect 2754 13392 2782 13512
rect 3366 13552 3418 13558
rect 2938 13512 3262 13540
rect 2886 13494 2938 13500
rect 3234 13392 3262 13512
rect 3849 13552 3901 13558
rect 3418 13512 3742 13540
rect 3366 13494 3418 13500
rect 3714 13392 3742 13512
rect 4333 13552 4385 13558
rect 3901 13512 4222 13540
rect 3849 13494 3901 13500
rect 4194 13392 4222 13512
rect 4817 13552 4869 13558
rect 4385 13512 4702 13540
rect 4333 13494 4385 13500
rect 4674 13392 4702 13512
rect 5299 13554 5355 13563
rect 5797 13558 5825 13605
rect 6390 13589 6442 13595
rect 4869 13512 5182 13540
rect 4817 13494 4869 13500
rect 5154 13392 5182 13512
rect 5299 13489 5355 13498
rect 5785 13552 5837 13558
rect 5785 13494 5837 13500
rect 5908 13554 5964 13563
rect 5908 13489 5964 13498
rect 6269 13552 6321 13558
rect 6321 13500 6334 13540
rect 6390 13531 6442 13537
rect 6774 13552 6826 13558
rect 6269 13494 6334 13500
rect 2754 13373 3022 13392
rect 3234 13373 3502 13392
rect 3714 13373 3982 13392
rect 4194 13373 4462 13392
rect 4674 13373 4942 13392
rect 5154 13373 5422 13392
rect 2754 13367 3034 13373
rect 2754 13364 2982 13367
rect 2500 13341 2502 13350
rect 2554 13341 2556 13350
rect 2502 13309 2554 13315
rect 3234 13367 3514 13373
rect 3234 13364 3462 13367
rect 2982 13309 3034 13315
rect 3714 13367 3994 13373
rect 3714 13364 3942 13367
rect 3462 13309 3514 13315
rect 4194 13367 4474 13373
rect 4194 13364 4422 13367
rect 3942 13309 3994 13315
rect 4674 13367 4954 13373
rect 4674 13364 4902 13367
rect 4422 13309 4474 13315
rect 5154 13367 5434 13373
rect 5154 13364 5382 13367
rect 4902 13309 4954 13315
rect 5382 13309 5434 13315
rect 5922 13188 5950 13489
rect 5910 13182 5962 13188
rect 5910 13124 5962 13130
rect 6306 13077 6334 13494
rect 6402 13484 6430 13531
rect 7254 13552 7306 13558
rect 6826 13512 7198 13540
rect 6774 13494 6826 13500
rect 6390 13478 6442 13484
rect 6390 13420 6442 13426
rect 7170 13392 7198 13512
rect 7734 13552 7786 13558
rect 7306 13512 7678 13540
rect 7254 13494 7306 13500
rect 7650 13392 7678 13512
rect 8214 13552 8266 13558
rect 7786 13512 8158 13540
rect 7734 13494 7786 13500
rect 8130 13392 8158 13512
rect 8694 13552 8746 13558
rect 8266 13512 8638 13540
rect 8214 13494 8266 13500
rect 8610 13392 8638 13512
rect 9090 13540 9118 13660
rect 8746 13512 9118 13540
rect 9174 13552 9226 13558
rect 8694 13494 8746 13500
rect 9174 13494 9226 13500
rect 7170 13373 7390 13392
rect 7650 13373 7870 13392
rect 8130 13373 8350 13392
rect 8610 13373 8830 13392
rect 7170 13367 7402 13373
rect 7170 13364 7350 13367
rect 7650 13367 7882 13373
rect 7650 13364 7830 13367
rect 7350 13309 7402 13315
rect 8130 13367 8362 13373
rect 8130 13364 8310 13367
rect 7830 13309 7882 13315
rect 8610 13367 8842 13373
rect 8610 13364 8790 13367
rect 8310 13309 8362 13315
rect 8790 13309 8842 13315
rect 6870 13182 6922 13188
rect 6870 13124 6922 13130
rect 6882 13077 6910 13124
rect 9186 13096 9214 13494
rect 9282 13447 9310 13660
rect 9270 13441 9322 13447
rect 9270 13383 9322 13389
rect 6294 13071 6346 13077
rect 6294 13013 6346 13019
rect 6870 13071 6922 13077
rect 9186 13068 9310 13096
rect 6870 13013 6922 13019
rect 3580 12888 3876 12908
rect 3636 12886 3660 12888
rect 3716 12886 3740 12888
rect 3796 12886 3820 12888
rect 3658 12834 3660 12886
rect 3722 12834 3734 12886
rect 3796 12834 3798 12886
rect 3636 12832 3660 12834
rect 3716 12832 3740 12834
rect 3796 12832 3820 12834
rect 3580 12812 3876 12832
rect 8908 12888 9204 12908
rect 8964 12886 8988 12888
rect 9044 12886 9068 12888
rect 9124 12886 9148 12888
rect 8986 12834 8988 12886
rect 9050 12834 9062 12886
rect 9124 12834 9126 12886
rect 8964 12832 8988 12834
rect 9044 12832 9068 12834
rect 9124 12832 9148 12834
rect 8908 12812 9204 12832
rect 6390 12590 6442 12596
rect 3942 12553 3994 12559
rect 5382 12553 5434 12559
rect 3994 12501 4318 12504
rect 3942 12495 4318 12501
rect 9282 12559 9310 13068
rect 6390 12532 6442 12538
rect 9270 12553 9322 12559
rect 6402 12504 6430 12532
rect 5434 12501 5808 12504
rect 5382 12495 5808 12501
rect 3954 12476 4318 12495
rect 5394 12476 5808 12495
rect 6402 12476 6814 12504
rect 9270 12495 9322 12501
rect 2022 12331 2074 12337
rect 2502 12331 2554 12337
rect 2074 12279 2398 12282
rect 2022 12273 2398 12279
rect 2982 12331 3034 12337
rect 2554 12279 2878 12282
rect 2502 12273 2878 12279
rect 3462 12331 3514 12337
rect 3034 12279 3358 12282
rect 2982 12273 3358 12279
rect 3514 12279 3838 12282
rect 3462 12273 3838 12279
rect 2034 12254 2398 12273
rect 2514 12254 2878 12273
rect 2994 12254 3358 12273
rect 3474 12254 3838 12273
rect 2370 12226 2398 12254
rect 2850 12226 2878 12254
rect 3330 12226 3358 12254
rect 3810 12226 3838 12254
rect 4290 12226 4318 12476
rect 4422 12331 4474 12337
rect 4902 12331 4954 12337
rect 4474 12279 4798 12282
rect 4422 12273 4798 12279
rect 4954 12279 5324 12282
rect 4902 12273 5324 12279
rect 4434 12254 4798 12273
rect 4914 12254 5324 12273
rect 4770 12226 4798 12254
rect 5296 12226 5324 12254
rect 5780 12226 5808 12476
rect 5910 12294 5962 12300
rect 5962 12254 6286 12282
rect 5910 12236 5962 12242
rect 6258 12226 6286 12254
rect 6786 12226 6814 12476
rect 7350 12331 7402 12337
rect 6870 12294 6922 12300
rect 7350 12273 7402 12279
rect 7830 12331 7882 12337
rect 7830 12273 7882 12279
rect 8310 12331 8362 12337
rect 8310 12273 8362 12279
rect 8790 12331 8842 12337
rect 8790 12273 8842 12279
rect 6870 12236 6922 12242
rect 1878 12220 1930 12226
rect 1878 12162 1930 12168
rect 2358 12220 2410 12226
rect 2358 12162 2410 12168
rect 2838 12220 2890 12226
rect 2838 12162 2890 12168
rect 3318 12220 3370 12226
rect 3318 12162 3370 12168
rect 3798 12220 3850 12226
rect 3798 12162 3850 12168
rect 4278 12220 4330 12226
rect 4278 12162 4330 12168
rect 4758 12220 4810 12226
rect 4758 12162 4810 12168
rect 5284 12220 5336 12226
rect 5284 12162 5336 12168
rect 5768 12220 5820 12226
rect 5768 12162 5820 12168
rect 6246 12220 6298 12226
rect 6246 12162 6298 12168
rect 6774 12220 6826 12226
rect 6882 12208 6910 12236
rect 7206 12220 7258 12226
rect 6882 12180 7206 12208
rect 6774 12162 6826 12168
rect 7362 12208 7390 12273
rect 7686 12220 7738 12226
rect 7362 12180 7686 12208
rect 7206 12162 7258 12168
rect 7842 12208 7870 12273
rect 8166 12220 8218 12226
rect 7842 12180 8166 12208
rect 7686 12162 7738 12168
rect 8322 12208 8350 12273
rect 8646 12220 8698 12226
rect 8322 12180 8646 12208
rect 8166 12162 8218 12168
rect 8802 12208 8830 12273
rect 9126 12220 9178 12226
rect 8802 12180 9126 12208
rect 8646 12162 8698 12168
rect 9126 12162 9178 12168
rect 1890 10987 1918 12162
rect 6244 11556 6540 11576
rect 6300 11554 6324 11556
rect 6380 11554 6404 11556
rect 6460 11554 6484 11556
rect 6322 11502 6324 11554
rect 6386 11502 6398 11554
rect 6460 11502 6462 11554
rect 6300 11500 6324 11502
rect 6380 11500 6404 11502
rect 6460 11500 6484 11502
rect 6244 11480 6540 11500
rect 5286 11073 5338 11079
rect 5286 11015 5338 11021
rect 5910 11073 5962 11079
rect 5910 11015 5962 11021
rect 6269 11073 6321 11079
rect 6269 11015 6321 11021
rect 6870 11073 6922 11079
rect 6870 11015 6922 11021
rect 4758 10999 4810 11005
rect 1890 10959 2062 10987
rect 1878 10888 1930 10894
rect 1878 10830 1930 10836
rect 1890 10751 1918 10830
rect 2034 10783 2062 10959
rect 4758 10941 4810 10947
rect 4770 10894 4798 10941
rect 5298 10894 5326 11015
rect 5382 10999 5434 11005
rect 5382 10941 5434 10947
rect 5785 10999 5837 11005
rect 5785 10941 5837 10947
rect 2406 10888 2458 10894
rect 2886 10888 2938 10894
rect 2458 10848 2782 10876
rect 2406 10830 2458 10836
rect 2754 10802 2782 10848
rect 3366 10888 3418 10894
rect 2938 10848 3262 10876
rect 2886 10830 2938 10836
rect 3234 10802 3262 10848
rect 3849 10888 3901 10894
rect 3418 10848 3742 10876
rect 3366 10830 3418 10836
rect 3714 10802 3742 10848
rect 4333 10888 4385 10894
rect 3901 10848 4222 10876
rect 3849 10830 3901 10836
rect 4194 10802 4222 10848
rect 4758 10888 4810 10894
rect 4385 10848 4702 10876
rect 4333 10830 4385 10836
rect 4674 10802 4702 10848
rect 4758 10830 4810 10836
rect 5286 10888 5338 10894
rect 5286 10830 5338 10836
rect 2754 10783 3022 10802
rect 3234 10783 3502 10802
rect 3714 10783 3982 10802
rect 4194 10783 4462 10802
rect 4674 10783 4942 10802
rect 5394 10783 5422 10941
rect 5797 10894 5825 10941
rect 5785 10888 5837 10894
rect 5785 10830 5837 10836
rect 5922 10820 5950 11015
rect 6281 10894 6309 11015
rect 6390 10999 6442 11005
rect 6390 10941 6442 10947
rect 6774 10999 6826 11005
rect 6774 10941 6826 10947
rect 6269 10888 6321 10894
rect 6269 10830 6321 10836
rect 6402 10820 6430 10941
rect 6786 10894 6814 10941
rect 6774 10888 6826 10894
rect 6774 10830 6826 10836
rect 6882 10820 6910 11015
rect 7350 10999 7402 11005
rect 7350 10941 7402 10947
rect 8694 10999 8746 11005
rect 8694 10941 8746 10947
rect 9270 10999 9322 11005
rect 9270 10941 9322 10947
rect 7254 10888 7306 10894
rect 7254 10830 7306 10836
rect 5910 10814 5962 10820
rect 2022 10777 2074 10783
rect 1876 10742 1932 10751
rect 2754 10777 3034 10783
rect 2754 10774 2982 10777
rect 2022 10719 2074 10725
rect 2500 10742 2556 10751
rect 1876 10677 1932 10686
rect 3234 10777 3514 10783
rect 3234 10774 3462 10777
rect 2982 10719 3034 10725
rect 3714 10777 3994 10783
rect 3714 10774 3942 10777
rect 3462 10719 3514 10725
rect 4194 10777 4474 10783
rect 4194 10774 4422 10777
rect 3942 10719 3994 10725
rect 4674 10777 4954 10783
rect 4674 10774 4902 10777
rect 4422 10719 4474 10725
rect 4902 10719 4954 10725
rect 5382 10777 5434 10783
rect 5910 10756 5962 10762
rect 6390 10814 6442 10820
rect 6390 10756 6442 10762
rect 6870 10814 6922 10820
rect 6870 10756 6922 10762
rect 5382 10719 5434 10725
rect 2500 10677 2502 10686
rect 2554 10677 2556 10686
rect 2502 10645 2554 10651
rect 7266 10580 7294 10830
rect 7362 10783 7390 10941
rect 8706 10894 8734 10941
rect 7734 10888 7786 10894
rect 8214 10888 8266 10894
rect 7786 10848 8158 10876
rect 7734 10830 7786 10836
rect 7350 10777 7402 10783
rect 7350 10719 7402 10725
rect 8130 10728 8158 10848
rect 8694 10888 8746 10894
rect 8266 10848 8638 10876
rect 8214 10830 8266 10836
rect 8610 10728 8638 10848
rect 8694 10830 8746 10836
rect 9174 10888 9226 10894
rect 9174 10830 9226 10836
rect 8130 10709 8350 10728
rect 8610 10709 8830 10728
rect 8130 10703 8362 10709
rect 8130 10700 8310 10703
rect 8610 10703 8842 10709
rect 8610 10700 8790 10703
rect 8310 10645 8362 10651
rect 8790 10645 8842 10651
rect 7830 10629 7882 10635
rect 7266 10577 7830 10580
rect 7266 10571 7882 10577
rect 7266 10552 7870 10571
rect 9186 10432 9214 10830
rect 9282 10783 9310 10941
rect 9270 10777 9322 10783
rect 9270 10719 9322 10725
rect 9186 10404 9310 10432
rect 3580 10224 3876 10244
rect 3636 10222 3660 10224
rect 3716 10222 3740 10224
rect 3796 10222 3820 10224
rect 3658 10170 3660 10222
rect 3722 10170 3734 10222
rect 3796 10170 3798 10222
rect 3636 10168 3660 10170
rect 3716 10168 3740 10170
rect 3796 10168 3820 10170
rect 3580 10148 3876 10168
rect 8908 10224 9204 10244
rect 8964 10222 8988 10224
rect 9044 10222 9068 10224
rect 9124 10222 9148 10224
rect 8986 10170 8988 10222
rect 9050 10170 9062 10222
rect 9124 10170 9126 10222
rect 8964 10168 8988 10170
rect 9044 10168 9068 10170
rect 9124 10168 9148 10170
rect 8908 10148 9204 10168
rect 9282 9895 9310 10404
rect 9270 9889 9322 9895
rect 9270 9831 9322 9837
rect 2022 9667 2074 9673
rect 2502 9667 2554 9673
rect 2074 9615 2398 9618
rect 2022 9609 2398 9615
rect 2982 9667 3034 9673
rect 2554 9615 2878 9618
rect 2502 9609 2878 9615
rect 3462 9667 3514 9673
rect 3034 9615 3358 9618
rect 2982 9609 3358 9615
rect 3942 9667 3994 9673
rect 3514 9615 3838 9618
rect 3462 9609 3838 9615
rect 4422 9667 4474 9673
rect 3994 9615 4318 9618
rect 3942 9609 4318 9615
rect 4902 9667 4954 9673
rect 4474 9615 4798 9618
rect 4422 9609 4798 9615
rect 5382 9667 5434 9673
rect 4954 9615 5324 9618
rect 4902 9609 5324 9615
rect 7350 9667 7402 9673
rect 5910 9630 5962 9636
rect 5434 9615 5806 9618
rect 5382 9609 5806 9615
rect 2034 9590 2398 9609
rect 2514 9590 2878 9609
rect 2994 9590 3358 9609
rect 3474 9590 3838 9609
rect 3954 9590 4318 9609
rect 4434 9590 4798 9609
rect 4914 9590 5324 9609
rect 5394 9590 5806 9609
rect 2370 9562 2398 9590
rect 2850 9562 2878 9590
rect 3330 9562 3358 9590
rect 3810 9562 3838 9590
rect 4290 9562 4318 9590
rect 4770 9562 4798 9590
rect 5296 9562 5324 9590
rect 5778 9562 5806 9590
rect 6390 9630 6442 9636
rect 5962 9590 6286 9618
rect 5910 9572 5962 9578
rect 6258 9562 6286 9590
rect 6870 9630 6922 9636
rect 6442 9590 6622 9618
rect 6390 9572 6442 9578
rect 1878 9556 1930 9562
rect 1878 9498 1930 9504
rect 2358 9556 2410 9562
rect 2358 9498 2410 9504
rect 2838 9556 2890 9562
rect 2838 9498 2890 9504
rect 3318 9556 3370 9562
rect 3318 9498 3370 9504
rect 3798 9556 3850 9562
rect 3798 9498 3850 9504
rect 4278 9556 4330 9562
rect 4278 9498 4330 9504
rect 4758 9556 4810 9562
rect 4758 9498 4810 9504
rect 5284 9556 5336 9562
rect 5284 9498 5336 9504
rect 5766 9556 5818 9562
rect 5766 9498 5818 9504
rect 6246 9556 6298 9562
rect 6594 9544 6622 9590
rect 7350 9609 7402 9615
rect 7830 9667 7882 9673
rect 7830 9609 7882 9615
rect 8310 9667 8362 9673
rect 8310 9609 8362 9615
rect 8790 9667 8842 9673
rect 8790 9609 8842 9615
rect 6870 9572 6922 9578
rect 6726 9556 6778 9562
rect 6594 9516 6726 9544
rect 6246 9498 6298 9504
rect 6882 9544 6910 9572
rect 7206 9556 7258 9562
rect 6882 9516 7206 9544
rect 6726 9498 6778 9504
rect 7362 9544 7390 9609
rect 7686 9556 7738 9562
rect 7362 9516 7686 9544
rect 7206 9498 7258 9504
rect 7842 9544 7870 9609
rect 8166 9556 8218 9562
rect 7842 9516 8166 9544
rect 7686 9498 7738 9504
rect 8322 9544 8350 9609
rect 8646 9556 8698 9562
rect 8322 9516 8646 9544
rect 8166 9498 8218 9504
rect 8802 9544 8830 9609
rect 9126 9556 9178 9562
rect 8802 9516 9126 9544
rect 8646 9498 8698 9504
rect 9126 9498 9178 9504
rect 1890 8323 1918 9498
rect 6244 8892 6540 8912
rect 6300 8890 6324 8892
rect 6380 8890 6404 8892
rect 6460 8890 6484 8892
rect 6322 8838 6324 8890
rect 6386 8838 6398 8890
rect 6460 8838 6462 8890
rect 6300 8836 6324 8838
rect 6380 8836 6404 8838
rect 6460 8836 6484 8838
rect 6244 8816 6540 8836
rect 5286 8409 5338 8415
rect 5286 8351 5338 8357
rect 5910 8409 5962 8415
rect 5910 8351 5962 8357
rect 6269 8409 6321 8415
rect 6269 8351 6321 8357
rect 6870 8409 6922 8415
rect 6870 8351 6922 8357
rect 4758 8335 4810 8341
rect 1890 8295 2062 8323
rect 1878 8224 1930 8230
rect 1878 8166 1930 8172
rect 1890 8087 1918 8166
rect 2034 8119 2062 8295
rect 4758 8277 4810 8283
rect 4770 8230 4798 8277
rect 5298 8230 5326 8351
rect 5382 8335 5434 8341
rect 5382 8277 5434 8283
rect 5785 8335 5837 8341
rect 5785 8277 5837 8283
rect 2406 8224 2458 8230
rect 2886 8224 2938 8230
rect 2458 8184 2782 8212
rect 2406 8166 2458 8172
rect 2754 8138 2782 8184
rect 3366 8224 3418 8230
rect 2938 8184 3262 8212
rect 2886 8166 2938 8172
rect 3234 8138 3262 8184
rect 3849 8224 3901 8230
rect 3418 8184 3742 8212
rect 3366 8166 3418 8172
rect 3714 8138 3742 8184
rect 4333 8224 4385 8230
rect 3901 8184 4222 8212
rect 3849 8166 3901 8172
rect 4194 8138 4222 8184
rect 4758 8224 4810 8230
rect 4385 8184 4702 8212
rect 4333 8166 4385 8172
rect 4674 8138 4702 8184
rect 4758 8166 4810 8172
rect 5286 8224 5338 8230
rect 5286 8166 5338 8172
rect 2754 8119 3022 8138
rect 3234 8119 3502 8138
rect 3714 8119 3982 8138
rect 4194 8119 4462 8138
rect 4674 8119 4942 8138
rect 5394 8119 5422 8277
rect 5797 8230 5825 8277
rect 5785 8224 5837 8230
rect 5785 8166 5837 8172
rect 5922 8156 5950 8351
rect 6281 8230 6309 8351
rect 6390 8335 6442 8341
rect 6390 8277 6442 8283
rect 6774 8335 6826 8341
rect 6774 8277 6826 8283
rect 6269 8224 6321 8230
rect 6269 8166 6321 8172
rect 6402 8156 6430 8277
rect 6786 8230 6814 8277
rect 6774 8224 6826 8230
rect 6774 8166 6826 8172
rect 6882 8156 6910 8351
rect 7350 8335 7402 8341
rect 7350 8277 7402 8283
rect 8694 8335 8746 8341
rect 8694 8277 8746 8283
rect 9270 8335 9322 8341
rect 9270 8277 9322 8283
rect 7254 8224 7306 8230
rect 7254 8166 7306 8172
rect 5910 8150 5962 8156
rect 2022 8113 2074 8119
rect 1876 8078 1932 8087
rect 2754 8113 3034 8119
rect 2754 8110 2982 8113
rect 2022 8055 2074 8061
rect 2500 8078 2556 8087
rect 1876 8013 1932 8022
rect 3234 8113 3514 8119
rect 3234 8110 3462 8113
rect 2982 8055 3034 8061
rect 3714 8113 3994 8119
rect 3714 8110 3942 8113
rect 3462 8055 3514 8061
rect 4194 8113 4474 8119
rect 4194 8110 4422 8113
rect 3942 8055 3994 8061
rect 4674 8113 4954 8119
rect 4674 8110 4902 8113
rect 4422 8055 4474 8061
rect 4902 8055 4954 8061
rect 5382 8113 5434 8119
rect 5910 8092 5962 8098
rect 6390 8150 6442 8156
rect 6390 8092 6442 8098
rect 6870 8150 6922 8156
rect 6870 8092 6922 8098
rect 5382 8055 5434 8061
rect 2500 8013 2502 8022
rect 2554 8013 2556 8022
rect 2502 7981 2554 7987
rect 7266 7916 7294 8166
rect 7362 8119 7390 8277
rect 8706 8230 8734 8277
rect 7734 8224 7786 8230
rect 8214 8224 8266 8230
rect 7786 8184 8158 8212
rect 7734 8166 7786 8172
rect 7350 8113 7402 8119
rect 7350 8055 7402 8061
rect 8130 8064 8158 8184
rect 8694 8224 8746 8230
rect 8266 8184 8638 8212
rect 8214 8166 8266 8172
rect 8610 8064 8638 8184
rect 8694 8166 8746 8172
rect 9174 8224 9226 8230
rect 9174 8166 9226 8172
rect 8130 8045 8350 8064
rect 8610 8045 8830 8064
rect 8130 8039 8362 8045
rect 8130 8036 8310 8039
rect 8610 8039 8842 8045
rect 8610 8036 8790 8039
rect 8310 7981 8362 7987
rect 8790 7981 8842 7987
rect 7830 7965 7882 7971
rect 7266 7913 7830 7916
rect 7266 7907 7882 7913
rect 7266 7888 7870 7907
rect 9186 7768 9214 8166
rect 9282 8119 9310 8277
rect 9270 8113 9322 8119
rect 9270 8055 9322 8061
rect 9186 7740 9310 7768
rect 3580 7560 3876 7580
rect 3636 7558 3660 7560
rect 3716 7558 3740 7560
rect 3796 7558 3820 7560
rect 3658 7506 3660 7558
rect 3722 7506 3734 7558
rect 3796 7506 3798 7558
rect 3636 7504 3660 7506
rect 3716 7504 3740 7506
rect 3796 7504 3820 7506
rect 3580 7484 3876 7504
rect 8908 7560 9204 7580
rect 8964 7558 8988 7560
rect 9044 7558 9068 7560
rect 9124 7558 9148 7560
rect 8986 7506 8988 7558
rect 9050 7506 9062 7558
rect 9124 7506 9126 7558
rect 8964 7504 8988 7506
rect 9044 7504 9068 7506
rect 9124 7504 9148 7506
rect 8908 7484 9204 7504
rect 9282 7231 9310 7740
rect 9270 7225 9322 7231
rect 9270 7167 9322 7173
rect 2022 7003 2074 7009
rect 2502 7003 2554 7009
rect 2074 6951 2398 6954
rect 2022 6945 2398 6951
rect 2982 7003 3034 7009
rect 2554 6951 2878 6954
rect 2502 6945 2878 6951
rect 3462 7003 3514 7009
rect 3034 6951 3358 6954
rect 2982 6945 3358 6951
rect 3942 7003 3994 7009
rect 3514 6951 3838 6954
rect 3462 6945 3838 6951
rect 4422 7003 4474 7009
rect 3994 6951 4318 6954
rect 3942 6945 4318 6951
rect 4902 7003 4954 7009
rect 4474 6951 4798 6954
rect 4422 6945 4798 6951
rect 5382 7003 5434 7009
rect 4954 6951 5324 6954
rect 4902 6945 5324 6951
rect 7350 7003 7402 7009
rect 5910 6966 5962 6972
rect 5434 6951 5806 6954
rect 5382 6945 5806 6951
rect 2034 6926 2398 6945
rect 2514 6926 2878 6945
rect 2994 6926 3358 6945
rect 3474 6926 3838 6945
rect 3954 6926 4318 6945
rect 4434 6926 4798 6945
rect 4914 6926 5324 6945
rect 5394 6926 5806 6945
rect 2370 6898 2398 6926
rect 2850 6898 2878 6926
rect 3330 6898 3358 6926
rect 3810 6898 3838 6926
rect 4290 6898 4318 6926
rect 4770 6898 4798 6926
rect 5296 6898 5324 6926
rect 5778 6898 5806 6926
rect 6390 6966 6442 6972
rect 5962 6926 6286 6954
rect 5910 6908 5962 6914
rect 6258 6898 6286 6926
rect 6870 6966 6922 6972
rect 6442 6926 6622 6954
rect 6390 6908 6442 6914
rect 1878 6892 1930 6898
rect 1878 6834 1930 6840
rect 2358 6892 2410 6898
rect 2358 6834 2410 6840
rect 2838 6892 2890 6898
rect 2838 6834 2890 6840
rect 3318 6892 3370 6898
rect 3318 6834 3370 6840
rect 3798 6892 3850 6898
rect 3798 6834 3850 6840
rect 4278 6892 4330 6898
rect 4278 6834 4330 6840
rect 4758 6892 4810 6898
rect 4758 6834 4810 6840
rect 5284 6892 5336 6898
rect 5284 6834 5336 6840
rect 5766 6892 5818 6898
rect 5766 6834 5818 6840
rect 6246 6892 6298 6898
rect 6594 6880 6622 6926
rect 7350 6945 7402 6951
rect 7830 7003 7882 7009
rect 7830 6945 7882 6951
rect 8310 7003 8362 7009
rect 8310 6945 8362 6951
rect 8790 7003 8842 7009
rect 8790 6945 8842 6951
rect 6870 6908 6922 6914
rect 6726 6892 6778 6898
rect 6594 6852 6726 6880
rect 6246 6834 6298 6840
rect 6882 6880 6910 6908
rect 7206 6892 7258 6898
rect 6882 6852 7206 6880
rect 6726 6834 6778 6840
rect 7362 6880 7390 6945
rect 7686 6892 7738 6898
rect 7362 6852 7686 6880
rect 7206 6834 7258 6840
rect 7842 6880 7870 6945
rect 8166 6892 8218 6898
rect 7842 6852 8166 6880
rect 7686 6834 7738 6840
rect 8322 6880 8350 6945
rect 8646 6892 8698 6898
rect 8322 6852 8646 6880
rect 8166 6834 8218 6840
rect 8802 6880 8830 6945
rect 9126 6892 9178 6898
rect 8802 6852 9126 6880
rect 8646 6834 8698 6840
rect 9126 6834 9178 6840
rect 1890 5659 1918 6834
rect 6244 6228 6540 6248
rect 6300 6226 6324 6228
rect 6380 6226 6404 6228
rect 6460 6226 6484 6228
rect 6322 6174 6324 6226
rect 6386 6174 6398 6226
rect 6460 6174 6462 6226
rect 6300 6172 6324 6174
rect 6380 6172 6404 6174
rect 6460 6172 6484 6174
rect 6244 6152 6540 6172
rect 5286 5745 5338 5751
rect 5286 5687 5338 5693
rect 5910 5745 5962 5751
rect 5910 5687 5962 5693
rect 6269 5745 6321 5751
rect 6269 5687 6321 5693
rect 6870 5745 6922 5751
rect 6870 5687 6922 5693
rect 4758 5671 4810 5677
rect 1890 5631 2062 5659
rect 1878 5560 1930 5566
rect 1878 5502 1930 5508
rect 1890 5423 1918 5502
rect 2034 5455 2062 5631
rect 4758 5613 4810 5619
rect 4770 5566 4798 5613
rect 5298 5566 5326 5687
rect 5382 5671 5434 5677
rect 5382 5613 5434 5619
rect 5785 5671 5837 5677
rect 5785 5613 5837 5619
rect 2406 5560 2458 5566
rect 2886 5560 2938 5566
rect 2458 5520 2782 5548
rect 2406 5502 2458 5508
rect 2754 5474 2782 5520
rect 3366 5560 3418 5566
rect 2938 5520 3262 5548
rect 2886 5502 2938 5508
rect 3234 5474 3262 5520
rect 3849 5560 3901 5566
rect 3418 5520 3742 5548
rect 3366 5502 3418 5508
rect 3714 5474 3742 5520
rect 4333 5560 4385 5566
rect 3901 5520 4222 5548
rect 3849 5502 3901 5508
rect 4194 5474 4222 5520
rect 4758 5560 4810 5566
rect 4385 5520 4702 5548
rect 4333 5502 4385 5508
rect 4674 5474 4702 5520
rect 4758 5502 4810 5508
rect 5286 5560 5338 5566
rect 5286 5502 5338 5508
rect 2754 5455 3022 5474
rect 3234 5455 3502 5474
rect 3714 5455 3982 5474
rect 4194 5455 4462 5474
rect 4674 5455 4942 5474
rect 5394 5455 5422 5613
rect 5797 5566 5825 5613
rect 5785 5560 5837 5566
rect 5785 5502 5837 5508
rect 5922 5492 5950 5687
rect 6281 5566 6309 5687
rect 6390 5671 6442 5677
rect 6390 5613 6442 5619
rect 6774 5671 6826 5677
rect 6774 5613 6826 5619
rect 6269 5560 6321 5566
rect 6269 5502 6321 5508
rect 6402 5492 6430 5613
rect 6786 5566 6814 5613
rect 6774 5560 6826 5566
rect 6774 5502 6826 5508
rect 6882 5492 6910 5687
rect 7350 5671 7402 5677
rect 7350 5613 7402 5619
rect 8694 5671 8746 5677
rect 8694 5613 8746 5619
rect 9270 5671 9322 5677
rect 9270 5613 9322 5619
rect 7254 5560 7306 5566
rect 7254 5502 7306 5508
rect 5910 5486 5962 5492
rect 2022 5449 2074 5455
rect 1876 5414 1932 5423
rect 2754 5449 3034 5455
rect 2754 5446 2982 5449
rect 2022 5391 2074 5397
rect 2500 5414 2556 5423
rect 1876 5349 1932 5358
rect 3234 5449 3514 5455
rect 3234 5446 3462 5449
rect 2982 5391 3034 5397
rect 3714 5449 3994 5455
rect 3714 5446 3942 5449
rect 3462 5391 3514 5397
rect 4194 5449 4474 5455
rect 4194 5446 4422 5449
rect 3942 5391 3994 5397
rect 4674 5449 4954 5455
rect 4674 5446 4902 5449
rect 4422 5391 4474 5397
rect 4902 5391 4954 5397
rect 5382 5449 5434 5455
rect 5910 5428 5962 5434
rect 6390 5486 6442 5492
rect 6390 5428 6442 5434
rect 6870 5486 6922 5492
rect 6870 5428 6922 5434
rect 5382 5391 5434 5397
rect 2500 5349 2502 5358
rect 2554 5349 2556 5358
rect 2502 5317 2554 5323
rect 7266 5252 7294 5502
rect 7362 5455 7390 5613
rect 8706 5566 8734 5613
rect 7734 5560 7786 5566
rect 8214 5560 8266 5566
rect 7786 5520 8158 5548
rect 7734 5502 7786 5508
rect 7350 5449 7402 5455
rect 7350 5391 7402 5397
rect 8130 5400 8158 5520
rect 8694 5560 8746 5566
rect 8266 5520 8638 5548
rect 8214 5502 8266 5508
rect 8610 5400 8638 5520
rect 8694 5502 8746 5508
rect 9174 5560 9226 5566
rect 9174 5502 9226 5508
rect 8130 5381 8350 5400
rect 8610 5381 8830 5400
rect 7830 5375 7882 5381
rect 8130 5375 8362 5381
rect 8130 5372 8310 5375
rect 7830 5317 7882 5323
rect 8610 5375 8842 5381
rect 8610 5372 8790 5375
rect 8310 5317 8362 5323
rect 8790 5317 8842 5323
rect 7842 5252 7870 5317
rect 7266 5224 7870 5252
rect 9186 5104 9214 5502
rect 9282 5455 9310 5613
rect 9270 5449 9322 5455
rect 9270 5391 9322 5397
rect 9186 5076 9310 5104
rect 3580 4896 3876 4916
rect 3636 4894 3660 4896
rect 3716 4894 3740 4896
rect 3796 4894 3820 4896
rect 3658 4842 3660 4894
rect 3722 4842 3734 4894
rect 3796 4842 3798 4894
rect 3636 4840 3660 4842
rect 3716 4840 3740 4842
rect 3796 4840 3820 4842
rect 3580 4820 3876 4840
rect 8908 4896 9204 4916
rect 8964 4894 8988 4896
rect 9044 4894 9068 4896
rect 9124 4894 9148 4896
rect 8986 4842 8988 4894
rect 9050 4842 9062 4894
rect 9124 4842 9126 4894
rect 8964 4840 8988 4842
rect 9044 4840 9068 4842
rect 9124 4840 9148 4842
rect 8908 4820 9204 4840
rect 9282 4567 9310 5076
rect 9270 4561 9322 4567
rect 9270 4503 9322 4509
rect 2022 4339 2074 4345
rect 2502 4339 2554 4345
rect 2074 4287 2398 4290
rect 2022 4281 2398 4287
rect 2982 4339 3034 4345
rect 2554 4287 2878 4290
rect 2502 4281 2878 4287
rect 3462 4339 3514 4345
rect 3034 4287 3358 4290
rect 2982 4281 3358 4287
rect 3942 4339 3994 4345
rect 3514 4287 3838 4290
rect 3462 4281 3838 4287
rect 4422 4339 4474 4345
rect 3994 4287 4318 4290
rect 3942 4281 4318 4287
rect 4902 4339 4954 4345
rect 4474 4287 4798 4290
rect 4422 4281 4798 4287
rect 5382 4339 5434 4345
rect 4954 4287 5324 4290
rect 4902 4281 5324 4287
rect 7350 4339 7402 4345
rect 5910 4302 5962 4308
rect 5434 4287 5806 4290
rect 5382 4281 5806 4287
rect 2034 4262 2398 4281
rect 2514 4262 2878 4281
rect 2994 4262 3358 4281
rect 3474 4262 3838 4281
rect 3954 4262 4318 4281
rect 4434 4262 4798 4281
rect 4914 4262 5324 4281
rect 5394 4262 5806 4281
rect 2370 4234 2398 4262
rect 2850 4234 2878 4262
rect 3330 4234 3358 4262
rect 3810 4234 3838 4262
rect 4290 4234 4318 4262
rect 4770 4234 4798 4262
rect 5296 4234 5324 4262
rect 5778 4234 5806 4262
rect 6390 4302 6442 4308
rect 5962 4262 6286 4290
rect 5910 4244 5962 4250
rect 6258 4234 6286 4262
rect 6870 4302 6922 4308
rect 6442 4262 6622 4290
rect 6390 4244 6442 4250
rect 1878 4228 1930 4234
rect 1878 4170 1930 4176
rect 2358 4228 2410 4234
rect 2358 4170 2410 4176
rect 2838 4228 2890 4234
rect 2838 4170 2890 4176
rect 3318 4228 3370 4234
rect 3318 4170 3370 4176
rect 3798 4228 3850 4234
rect 3798 4170 3850 4176
rect 4278 4228 4330 4234
rect 4278 4170 4330 4176
rect 4758 4228 4810 4234
rect 4758 4170 4810 4176
rect 5284 4228 5336 4234
rect 5284 4170 5336 4176
rect 5766 4228 5818 4234
rect 5766 4170 5818 4176
rect 6246 4228 6298 4234
rect 6594 4216 6622 4262
rect 7350 4281 7402 4287
rect 7830 4339 7882 4345
rect 7830 4281 7882 4287
rect 8310 4339 8362 4345
rect 8310 4281 8362 4287
rect 8790 4339 8842 4345
rect 8790 4281 8842 4287
rect 6870 4244 6922 4250
rect 6726 4228 6778 4234
rect 6594 4188 6726 4216
rect 6246 4170 6298 4176
rect 6882 4216 6910 4244
rect 7206 4228 7258 4234
rect 6882 4188 7206 4216
rect 6726 4170 6778 4176
rect 7362 4216 7390 4281
rect 7686 4228 7738 4234
rect 7362 4188 7686 4216
rect 7206 4170 7258 4176
rect 7842 4216 7870 4281
rect 8166 4228 8218 4234
rect 7842 4188 8166 4216
rect 7686 4170 7738 4176
rect 8322 4216 8350 4281
rect 8646 4228 8698 4234
rect 8322 4188 8646 4216
rect 8166 4170 8218 4176
rect 8802 4216 8830 4281
rect 9126 4228 9178 4234
rect 8802 4188 9126 4216
rect 8646 4170 8698 4176
rect 9126 4170 9178 4176
rect 1890 4068 1918 4170
rect 1890 4040 2110 4068
rect 1878 2896 1930 2902
rect 2082 2884 2110 4040
rect 6244 3564 6540 3584
rect 6300 3562 6324 3564
rect 6380 3562 6404 3564
rect 6460 3562 6484 3564
rect 6322 3510 6324 3562
rect 6386 3510 6398 3562
rect 6460 3510 6462 3562
rect 6300 3508 6324 3510
rect 6380 3508 6404 3510
rect 6460 3508 6484 3510
rect 6244 3488 6540 3508
rect 5785 3007 5837 3013
rect 5785 2949 5837 2955
rect 9090 3004 9310 3032
rect 1878 2838 1930 2844
rect 2034 2856 2110 2884
rect 2406 2896 2458 2902
rect 1890 2759 1918 2838
rect 2034 2791 2062 2856
rect 2886 2896 2938 2902
rect 2458 2856 2782 2884
rect 2406 2838 2458 2844
rect 2022 2785 2074 2791
rect 1876 2750 1932 2759
rect 2022 2727 2074 2733
rect 2500 2750 2556 2759
rect 1876 2685 1932 2694
rect 2754 2736 2782 2856
rect 3366 2896 3418 2902
rect 2938 2856 3262 2884
rect 2886 2838 2938 2844
rect 3234 2736 3262 2856
rect 3849 2896 3901 2902
rect 3418 2856 3742 2884
rect 3366 2838 3418 2844
rect 3714 2736 3742 2856
rect 4333 2896 4385 2902
rect 3901 2856 4222 2884
rect 3849 2838 3901 2844
rect 4194 2736 4222 2856
rect 4817 2896 4869 2902
rect 4385 2856 4702 2884
rect 4333 2838 4385 2844
rect 4674 2736 4702 2856
rect 5299 2898 5355 2907
rect 5797 2902 5825 2949
rect 6390 2933 6442 2939
rect 4869 2856 5182 2884
rect 4817 2838 4869 2844
rect 5154 2736 5182 2856
rect 5299 2833 5355 2842
rect 5785 2896 5837 2902
rect 5785 2838 5837 2844
rect 5908 2898 5964 2907
rect 5908 2833 5964 2842
rect 6269 2896 6321 2902
rect 6321 2844 6334 2884
rect 6390 2875 6442 2881
rect 6774 2896 6826 2902
rect 6269 2838 6334 2844
rect 2754 2717 3022 2736
rect 3234 2717 3502 2736
rect 3714 2717 3982 2736
rect 4194 2717 4462 2736
rect 4674 2717 4942 2736
rect 5154 2717 5422 2736
rect 2754 2711 3034 2717
rect 2754 2708 2982 2711
rect 2500 2685 2502 2694
rect 2554 2685 2556 2694
rect 2502 2653 2554 2659
rect 3234 2711 3514 2717
rect 3234 2708 3462 2711
rect 2982 2653 3034 2659
rect 3714 2711 3994 2717
rect 3714 2708 3942 2711
rect 3462 2653 3514 2659
rect 4194 2711 4474 2717
rect 4194 2708 4422 2711
rect 3942 2653 3994 2659
rect 4674 2711 4954 2717
rect 4674 2708 4902 2711
rect 4422 2653 4474 2659
rect 5154 2711 5434 2717
rect 5154 2708 5382 2711
rect 4902 2653 4954 2659
rect 5382 2653 5434 2659
rect 5922 2532 5950 2833
rect 5910 2526 5962 2532
rect 5910 2468 5962 2474
rect 6306 2421 6334 2838
rect 6402 2828 6430 2875
rect 7254 2896 7306 2902
rect 6826 2856 7198 2884
rect 6774 2838 6826 2844
rect 6390 2822 6442 2828
rect 7170 2810 7198 2856
rect 7734 2896 7786 2902
rect 7306 2856 7678 2884
rect 7254 2838 7306 2844
rect 7650 2810 7678 2856
rect 8214 2896 8266 2902
rect 7786 2856 8158 2884
rect 7734 2838 7786 2844
rect 8130 2810 8158 2856
rect 8694 2896 8746 2902
rect 8266 2856 8638 2884
rect 8214 2838 8266 2844
rect 8610 2810 8638 2856
rect 9090 2884 9118 3004
rect 8746 2856 9118 2884
rect 9174 2896 9226 2902
rect 8694 2838 8746 2844
rect 9174 2838 9226 2844
rect 7170 2791 7390 2810
rect 7650 2791 7870 2810
rect 8130 2791 8350 2810
rect 8610 2791 8830 2810
rect 7170 2785 7402 2791
rect 7170 2782 7350 2785
rect 6390 2764 6442 2770
rect 7650 2785 7882 2791
rect 7650 2782 7830 2785
rect 7350 2727 7402 2733
rect 8130 2785 8362 2791
rect 8130 2782 8310 2785
rect 7830 2727 7882 2733
rect 8610 2785 8842 2791
rect 8610 2782 8790 2785
rect 8310 2727 8362 2733
rect 8790 2727 8842 2733
rect 6870 2526 6922 2532
rect 6870 2468 6922 2474
rect 6882 2421 6910 2468
rect 6294 2415 6346 2421
rect 6294 2357 6346 2363
rect 6870 2415 6922 2421
rect 9186 2403 9214 2838
rect 9282 2791 9310 3004
rect 9270 2785 9322 2791
rect 9270 2727 9322 2733
rect 9186 2375 9310 2403
rect 6870 2357 6922 2363
rect 3580 2232 3876 2252
rect 3636 2230 3660 2232
rect 3716 2230 3740 2232
rect 3796 2230 3820 2232
rect 3658 2178 3660 2230
rect 3722 2178 3734 2230
rect 3796 2178 3798 2230
rect 3636 2176 3660 2178
rect 3716 2176 3740 2178
rect 3796 2176 3820 2178
rect 3580 2156 3876 2176
rect 8908 2232 9204 2252
rect 8964 2230 8988 2232
rect 9044 2230 9068 2232
rect 9124 2230 9148 2232
rect 8986 2178 8988 2230
rect 9050 2178 9062 2230
rect 9124 2178 9126 2230
rect 8964 2176 8988 2178
rect 9044 2176 9068 2178
rect 9124 2176 9148 2178
rect 8908 2156 9204 2176
rect 6390 1934 6442 1940
rect 9282 1903 9310 2375
rect 6390 1876 6442 1882
rect 9270 1897 9322 1903
rect 6402 1848 6430 1876
rect 3954 1829 4318 1848
rect 5394 1829 5806 1848
rect 3942 1823 4318 1829
rect 3994 1820 4318 1823
rect 3942 1765 3994 1771
rect 2022 1675 2074 1681
rect 2502 1675 2554 1681
rect 2074 1623 2398 1626
rect 2022 1617 2398 1623
rect 2982 1675 3034 1681
rect 2554 1623 2878 1626
rect 2502 1617 2878 1623
rect 3462 1675 3514 1681
rect 3034 1623 3358 1626
rect 2982 1617 3358 1623
rect 4290 1626 4318 1820
rect 5382 1823 5806 1829
rect 5434 1820 5806 1823
rect 6402 1820 6814 1848
rect 9270 1839 9322 1845
rect 5382 1765 5434 1771
rect 4422 1675 4474 1681
rect 3514 1623 3838 1626
rect 3462 1617 3838 1623
rect 2034 1598 2398 1617
rect 2514 1598 2878 1617
rect 2994 1598 3358 1617
rect 3474 1598 3838 1617
rect 4290 1598 4373 1626
rect 4902 1675 4954 1681
rect 4474 1623 4798 1626
rect 4422 1617 4798 1623
rect 4954 1623 5324 1626
rect 4902 1617 5324 1623
rect 4434 1598 4798 1617
rect 4914 1598 5324 1617
rect 1876 1566 1932 1575
rect 2370 1570 2398 1598
rect 2850 1570 2878 1598
rect 3330 1570 3358 1598
rect 3810 1570 3838 1598
rect 4345 1570 4373 1598
rect 4770 1570 4798 1598
rect 5296 1570 5324 1598
rect 5778 1570 5806 1820
rect 5910 1638 5962 1644
rect 5962 1598 6286 1626
rect 5910 1580 5962 1586
rect 6258 1570 6286 1598
rect 6786 1570 6814 1820
rect 7350 1675 7402 1681
rect 6870 1638 6922 1644
rect 7350 1617 7402 1623
rect 7830 1675 7882 1681
rect 7830 1617 7882 1623
rect 8310 1675 8362 1681
rect 8310 1617 8362 1623
rect 8790 1675 8842 1681
rect 8790 1617 8842 1623
rect 6870 1580 6922 1586
rect 1794 1524 1876 1552
rect 1876 1501 1932 1510
rect 2358 1564 2410 1570
rect 2358 1506 2410 1512
rect 2838 1564 2890 1570
rect 2838 1506 2890 1512
rect 3318 1564 3370 1570
rect 3318 1506 3370 1512
rect 3798 1564 3850 1570
rect 3798 1506 3850 1512
rect 4333 1564 4385 1570
rect 4333 1506 4385 1512
rect 4758 1564 4810 1570
rect 4758 1506 4810 1512
rect 5284 1564 5336 1570
rect 5284 1506 5336 1512
rect 5766 1564 5818 1570
rect 5766 1506 5818 1512
rect 6246 1564 6298 1570
rect 6246 1506 6298 1512
rect 6774 1564 6826 1570
rect 6882 1552 6910 1580
rect 7206 1564 7258 1570
rect 6882 1524 7206 1552
rect 6774 1506 6826 1512
rect 7362 1552 7390 1617
rect 7686 1564 7738 1570
rect 7362 1524 7686 1552
rect 7206 1506 7258 1512
rect 7842 1552 7870 1617
rect 8166 1564 8218 1570
rect 7842 1524 8166 1552
rect 7686 1506 7738 1512
rect 8322 1552 8350 1617
rect 8646 1564 8698 1570
rect 8322 1524 8646 1552
rect 8166 1506 8218 1512
rect 8802 1552 8830 1617
rect 9126 1564 9178 1570
rect 8802 1524 9126 1552
rect 8646 1506 8698 1512
rect 9126 1506 9178 1512
rect 6244 900 6540 920
rect 6300 898 6324 900
rect 6380 898 6404 900
rect 6460 898 6484 900
rect 6322 846 6324 898
rect 6386 846 6398 898
rect 6460 846 6462 898
rect 6300 844 6324 846
rect 6380 844 6404 846
rect 6460 844 6484 846
rect 6244 824 6540 844
<< via2 >>
rect 3580 52846 3636 52848
rect 3660 52846 3716 52848
rect 3740 52846 3796 52848
rect 3820 52846 3876 52848
rect 3580 52794 3606 52846
rect 3606 52794 3636 52846
rect 3660 52794 3670 52846
rect 3670 52794 3716 52846
rect 3740 52794 3786 52846
rect 3786 52794 3796 52846
rect 3820 52794 3850 52846
rect 3850 52794 3876 52846
rect 3580 52792 3636 52794
rect 3660 52792 3716 52794
rect 3740 52792 3796 52794
rect 3820 52792 3876 52794
rect 8908 52846 8964 52848
rect 8988 52846 9044 52848
rect 9068 52846 9124 52848
rect 9148 52846 9204 52848
rect 8908 52794 8934 52846
rect 8934 52794 8964 52846
rect 8988 52794 8998 52846
rect 8998 52794 9044 52846
rect 9068 52794 9114 52846
rect 9114 52794 9124 52846
rect 9148 52794 9178 52846
rect 9178 52794 9204 52846
rect 8908 52792 8964 52794
rect 8988 52792 9044 52794
rect 9068 52792 9124 52794
rect 9148 52792 9204 52794
rect 1348 52461 1350 52478
rect 1350 52461 1402 52478
rect 1402 52461 1404 52478
rect 1348 52422 1404 52461
rect 1108 51978 1164 52034
rect 1108 50646 1164 50702
rect 6244 51514 6300 51516
rect 6324 51514 6380 51516
rect 6404 51514 6460 51516
rect 6484 51514 6540 51516
rect 6244 51462 6270 51514
rect 6270 51462 6300 51514
rect 6324 51462 6334 51514
rect 6334 51462 6380 51514
rect 6404 51462 6450 51514
rect 6450 51462 6460 51514
rect 6484 51462 6514 51514
rect 6514 51462 6540 51514
rect 6244 51460 6300 51462
rect 6324 51460 6380 51462
rect 6404 51460 6460 51462
rect 6484 51460 6540 51462
rect 3580 50182 3636 50184
rect 3660 50182 3716 50184
rect 3740 50182 3796 50184
rect 3820 50182 3876 50184
rect 3580 50130 3606 50182
rect 3606 50130 3636 50182
rect 3660 50130 3670 50182
rect 3670 50130 3716 50182
rect 3740 50130 3786 50182
rect 3786 50130 3796 50182
rect 3820 50130 3850 50182
rect 3850 50130 3876 50182
rect 3580 50128 3636 50130
rect 3660 50128 3716 50130
rect 3740 50128 3796 50130
rect 3820 50128 3876 50130
rect 8908 50182 8964 50184
rect 8988 50182 9044 50184
rect 9068 50182 9124 50184
rect 9148 50182 9204 50184
rect 8908 50130 8934 50182
rect 8934 50130 8964 50182
rect 8988 50130 8998 50182
rect 8998 50130 9044 50182
rect 9068 50130 9114 50182
rect 9114 50130 9124 50182
rect 9148 50130 9178 50182
rect 9178 50130 9204 50182
rect 8908 50128 8964 50130
rect 8988 50128 9044 50130
rect 9068 50128 9124 50130
rect 9148 50128 9204 50130
rect 6244 48850 6300 48852
rect 6324 48850 6380 48852
rect 6404 48850 6460 48852
rect 6484 48850 6540 48852
rect 6244 48798 6270 48850
rect 6270 48798 6300 48850
rect 6324 48798 6334 48850
rect 6334 48798 6380 48850
rect 6404 48798 6450 48850
rect 6450 48798 6460 48850
rect 6484 48798 6514 48850
rect 6514 48798 6540 48850
rect 6244 48796 6300 48798
rect 6324 48796 6380 48798
rect 6404 48796 6460 48798
rect 6484 48796 6540 48798
rect 1108 47982 1164 48038
rect 3580 47518 3636 47520
rect 3660 47518 3716 47520
rect 3740 47518 3796 47520
rect 3820 47518 3876 47520
rect 3580 47466 3606 47518
rect 3606 47466 3636 47518
rect 3660 47466 3670 47518
rect 3670 47466 3716 47518
rect 3740 47466 3786 47518
rect 3786 47466 3796 47518
rect 3820 47466 3850 47518
rect 3850 47466 3876 47518
rect 3580 47464 3636 47466
rect 3660 47464 3716 47466
rect 3740 47464 3796 47466
rect 3820 47464 3876 47466
rect 8908 47518 8964 47520
rect 8988 47518 9044 47520
rect 9068 47518 9124 47520
rect 9148 47518 9204 47520
rect 8908 47466 8934 47518
rect 8934 47466 8964 47518
rect 8988 47466 8998 47518
rect 8998 47466 9044 47518
rect 9068 47466 9114 47518
rect 9114 47466 9124 47518
rect 9148 47466 9178 47518
rect 9178 47466 9204 47518
rect 8908 47464 8964 47466
rect 8988 47464 9044 47466
rect 9068 47464 9124 47466
rect 9148 47464 9204 47466
rect 1108 45318 1164 45374
rect 6244 46186 6300 46188
rect 6324 46186 6380 46188
rect 6404 46186 6460 46188
rect 6484 46186 6540 46188
rect 6244 46134 6270 46186
rect 6270 46134 6300 46186
rect 6324 46134 6334 46186
rect 6334 46134 6380 46186
rect 6404 46134 6450 46186
rect 6450 46134 6460 46186
rect 6484 46134 6514 46186
rect 6514 46134 6540 46186
rect 6244 46132 6300 46134
rect 6324 46132 6380 46134
rect 6404 46132 6460 46134
rect 6484 46132 6540 46134
rect 2836 45520 2892 45522
rect 2836 45468 2838 45520
rect 2838 45468 2890 45520
rect 2890 45468 2892 45520
rect 2836 45466 2892 45468
rect 3460 45466 3516 45522
rect 3580 44854 3636 44856
rect 3660 44854 3716 44856
rect 3740 44854 3796 44856
rect 3820 44854 3876 44856
rect 3580 44802 3606 44854
rect 3606 44802 3636 44854
rect 3660 44802 3670 44854
rect 3670 44802 3716 44854
rect 3740 44802 3786 44854
rect 3786 44802 3796 44854
rect 3820 44802 3850 44854
rect 3850 44802 3876 44854
rect 3580 44800 3636 44802
rect 3660 44800 3716 44802
rect 3740 44800 3796 44802
rect 3820 44800 3876 44802
rect 8908 44854 8964 44856
rect 8988 44854 9044 44856
rect 9068 44854 9124 44856
rect 9148 44854 9204 44856
rect 8908 44802 8934 44854
rect 8934 44802 8964 44854
rect 8988 44802 8998 44854
rect 8998 44802 9044 44854
rect 9068 44802 9114 44854
rect 9114 44802 9124 44854
rect 9148 44802 9178 44854
rect 9178 44802 9204 44854
rect 8908 44800 8964 44802
rect 8988 44800 9044 44802
rect 9068 44800 9124 44802
rect 9148 44800 9204 44802
rect 6244 43522 6300 43524
rect 6324 43522 6380 43524
rect 6404 43522 6460 43524
rect 6484 43522 6540 43524
rect 6244 43470 6270 43522
rect 6270 43470 6300 43522
rect 6324 43470 6334 43522
rect 6334 43470 6380 43522
rect 6404 43470 6450 43522
rect 6450 43470 6460 43522
rect 6484 43470 6514 43522
rect 6514 43470 6540 43522
rect 6244 43468 6300 43470
rect 6324 43468 6380 43470
rect 6404 43468 6460 43470
rect 6484 43468 6540 43470
rect 1108 42654 1164 42710
rect 3580 42190 3636 42192
rect 3660 42190 3716 42192
rect 3740 42190 3796 42192
rect 3820 42190 3876 42192
rect 3580 42138 3606 42190
rect 3606 42138 3636 42190
rect 3660 42138 3670 42190
rect 3670 42138 3716 42190
rect 3740 42138 3786 42190
rect 3786 42138 3796 42190
rect 3820 42138 3850 42190
rect 3850 42138 3876 42190
rect 3580 42136 3636 42138
rect 3660 42136 3716 42138
rect 3740 42136 3796 42138
rect 3820 42136 3876 42138
rect 8908 42190 8964 42192
rect 8988 42190 9044 42192
rect 9068 42190 9124 42192
rect 9148 42190 9204 42192
rect 8908 42138 8934 42190
rect 8934 42138 8964 42190
rect 8988 42138 8998 42190
rect 8998 42138 9044 42190
rect 9068 42138 9114 42190
rect 9114 42138 9124 42190
rect 9148 42138 9178 42190
rect 9178 42138 9204 42190
rect 8908 42136 8964 42138
rect 8988 42136 9044 42138
rect 9068 42136 9124 42138
rect 9148 42136 9204 42138
rect 1108 40192 1164 40194
rect 1108 40140 1110 40192
rect 1110 40140 1162 40192
rect 1162 40140 1164 40192
rect 6244 40858 6300 40860
rect 6324 40858 6380 40860
rect 6404 40858 6460 40860
rect 6484 40858 6540 40860
rect 6244 40806 6270 40858
rect 6270 40806 6300 40858
rect 6324 40806 6334 40858
rect 6334 40806 6380 40858
rect 6404 40806 6450 40858
rect 6450 40806 6460 40858
rect 6484 40806 6514 40858
rect 6514 40806 6540 40858
rect 6244 40804 6300 40806
rect 6324 40804 6380 40806
rect 6404 40804 6460 40806
rect 6484 40804 6540 40806
rect 1108 40138 1164 40140
rect 3580 39526 3636 39528
rect 3660 39526 3716 39528
rect 3740 39526 3796 39528
rect 3820 39526 3876 39528
rect 3580 39474 3606 39526
rect 3606 39474 3636 39526
rect 3660 39474 3670 39526
rect 3670 39474 3716 39526
rect 3740 39474 3786 39526
rect 3786 39474 3796 39526
rect 3820 39474 3850 39526
rect 3850 39474 3876 39526
rect 3580 39472 3636 39474
rect 3660 39472 3716 39474
rect 3740 39472 3796 39474
rect 3820 39472 3876 39474
rect 8908 39526 8964 39528
rect 8988 39526 9044 39528
rect 9068 39526 9124 39528
rect 9148 39526 9204 39528
rect 8908 39474 8934 39526
rect 8934 39474 8964 39526
rect 8988 39474 8998 39526
rect 8998 39474 9044 39526
rect 9068 39474 9114 39526
rect 9114 39474 9124 39526
rect 9148 39474 9178 39526
rect 9178 39474 9204 39526
rect 8908 39472 8964 39474
rect 8988 39472 9044 39474
rect 9068 39472 9124 39474
rect 9148 39472 9204 39474
rect 1108 37326 1164 37382
rect 6244 38194 6300 38196
rect 6324 38194 6380 38196
rect 6404 38194 6460 38196
rect 6484 38194 6540 38196
rect 6244 38142 6270 38194
rect 6270 38142 6300 38194
rect 6324 38142 6334 38194
rect 6334 38142 6380 38194
rect 6404 38142 6450 38194
rect 6450 38142 6460 38194
rect 6484 38142 6514 38194
rect 6514 38142 6540 38194
rect 6244 38140 6300 38142
rect 6324 38140 6380 38142
rect 6404 38140 6460 38142
rect 6484 38140 6540 38142
rect 3580 36862 3636 36864
rect 3660 36862 3716 36864
rect 3740 36862 3796 36864
rect 3820 36862 3876 36864
rect 3580 36810 3606 36862
rect 3606 36810 3636 36862
rect 3660 36810 3670 36862
rect 3670 36810 3716 36862
rect 3740 36810 3786 36862
rect 3786 36810 3796 36862
rect 3820 36810 3850 36862
rect 3850 36810 3876 36862
rect 3580 36808 3636 36810
rect 3660 36808 3716 36810
rect 3740 36808 3796 36810
rect 3820 36808 3876 36810
rect 8908 36862 8964 36864
rect 8988 36862 9044 36864
rect 9068 36862 9124 36864
rect 9148 36862 9204 36864
rect 8908 36810 8934 36862
rect 8934 36810 8964 36862
rect 8988 36810 8998 36862
rect 8998 36810 9044 36862
rect 9068 36810 9114 36862
rect 9114 36810 9124 36862
rect 9148 36810 9178 36862
rect 9178 36810 9204 36862
rect 8908 36808 8964 36810
rect 8988 36808 9044 36810
rect 9068 36808 9124 36810
rect 9148 36808 9204 36810
rect 6244 35530 6300 35532
rect 6324 35530 6380 35532
rect 6404 35530 6460 35532
rect 6484 35530 6540 35532
rect 6244 35478 6270 35530
rect 6270 35478 6300 35530
rect 6324 35478 6334 35530
rect 6334 35478 6380 35530
rect 6404 35478 6450 35530
rect 6450 35478 6460 35530
rect 6484 35478 6514 35530
rect 6514 35478 6540 35530
rect 6244 35476 6300 35478
rect 6324 35476 6380 35478
rect 6404 35476 6460 35478
rect 6484 35476 6540 35478
rect 1876 34662 1932 34718
rect 2500 34679 2556 34718
rect 2500 34662 2502 34679
rect 2502 34662 2554 34679
rect 2554 34662 2556 34679
rect 5299 34864 5355 34866
rect 5299 34812 5301 34864
rect 5301 34812 5353 34864
rect 5353 34812 5355 34864
rect 5299 34810 5355 34812
rect 5908 34810 5964 34866
rect 3580 34198 3636 34200
rect 3660 34198 3716 34200
rect 3740 34198 3796 34200
rect 3820 34198 3876 34200
rect 3580 34146 3606 34198
rect 3606 34146 3636 34198
rect 3660 34146 3670 34198
rect 3670 34146 3716 34198
rect 3740 34146 3786 34198
rect 3786 34146 3796 34198
rect 3820 34146 3850 34198
rect 3850 34146 3876 34198
rect 3580 34144 3636 34146
rect 3660 34144 3716 34146
rect 3740 34144 3796 34146
rect 3820 34144 3876 34146
rect 8908 34198 8964 34200
rect 8988 34198 9044 34200
rect 9068 34198 9124 34200
rect 9148 34198 9204 34200
rect 8908 34146 8934 34198
rect 8934 34146 8964 34198
rect 8988 34146 8998 34198
rect 8998 34146 9044 34198
rect 9068 34146 9114 34198
rect 9114 34146 9124 34198
rect 9148 34146 9178 34198
rect 9178 34146 9204 34198
rect 8908 34144 8964 34146
rect 8988 34144 9044 34146
rect 9068 34144 9124 34146
rect 9148 34144 9204 34146
rect 6244 32866 6300 32868
rect 6324 32866 6380 32868
rect 6404 32866 6460 32868
rect 6484 32866 6540 32868
rect 6244 32814 6270 32866
rect 6270 32814 6300 32866
rect 6324 32814 6334 32866
rect 6334 32814 6380 32866
rect 6404 32814 6450 32866
rect 6450 32814 6460 32866
rect 6484 32814 6514 32866
rect 6514 32814 6540 32866
rect 6244 32812 6300 32814
rect 6324 32812 6380 32814
rect 6404 32812 6460 32814
rect 6484 32812 6540 32814
rect 1108 31998 1164 32054
rect 3580 31534 3636 31536
rect 3660 31534 3716 31536
rect 3740 31534 3796 31536
rect 3820 31534 3876 31536
rect 3580 31482 3606 31534
rect 3606 31482 3636 31534
rect 3660 31482 3670 31534
rect 3670 31482 3716 31534
rect 3740 31482 3786 31534
rect 3786 31482 3796 31534
rect 3820 31482 3850 31534
rect 3850 31482 3876 31534
rect 3580 31480 3636 31482
rect 3660 31480 3716 31482
rect 3740 31480 3796 31482
rect 3820 31480 3876 31482
rect 8908 31534 8964 31536
rect 8988 31534 9044 31536
rect 9068 31534 9124 31536
rect 9148 31534 9204 31536
rect 8908 31482 8934 31534
rect 8934 31482 8964 31534
rect 8988 31482 8998 31534
rect 8998 31482 9044 31534
rect 9068 31482 9114 31534
rect 9114 31482 9124 31534
rect 9148 31482 9178 31534
rect 9178 31482 9204 31534
rect 8908 31480 8964 31482
rect 8988 31480 9044 31482
rect 9068 31480 9124 31482
rect 9148 31480 9204 31482
rect 6244 30202 6300 30204
rect 6324 30202 6380 30204
rect 6404 30202 6460 30204
rect 6484 30202 6540 30204
rect 6244 30150 6270 30202
rect 6270 30150 6300 30202
rect 6324 30150 6334 30202
rect 6334 30150 6380 30202
rect 6404 30150 6450 30202
rect 6450 30150 6460 30202
rect 6484 30150 6514 30202
rect 6514 30150 6540 30202
rect 6244 30148 6300 30150
rect 6324 30148 6380 30150
rect 6404 30148 6460 30150
rect 6484 30148 6540 30150
rect 1876 29334 1932 29390
rect 2500 29351 2556 29390
rect 2500 29334 2502 29351
rect 2502 29334 2554 29351
rect 2554 29334 2556 29351
rect 3580 28870 3636 28872
rect 3660 28870 3716 28872
rect 3740 28870 3796 28872
rect 3820 28870 3876 28872
rect 3580 28818 3606 28870
rect 3606 28818 3636 28870
rect 3660 28818 3670 28870
rect 3670 28818 3716 28870
rect 3740 28818 3786 28870
rect 3786 28818 3796 28870
rect 3820 28818 3850 28870
rect 3850 28818 3876 28870
rect 3580 28816 3636 28818
rect 3660 28816 3716 28818
rect 3740 28816 3796 28818
rect 3820 28816 3876 28818
rect 8908 28870 8964 28872
rect 8988 28870 9044 28872
rect 9068 28870 9124 28872
rect 9148 28870 9204 28872
rect 8908 28818 8934 28870
rect 8934 28818 8964 28870
rect 8988 28818 8998 28870
rect 8998 28818 9044 28870
rect 9068 28818 9114 28870
rect 9114 28818 9124 28870
rect 9148 28818 9178 28870
rect 9178 28818 9204 28870
rect 8908 28816 8964 28818
rect 8988 28816 9044 28818
rect 9068 28816 9124 28818
rect 9148 28816 9204 28818
rect 6244 27538 6300 27540
rect 6324 27538 6380 27540
rect 6404 27538 6460 27540
rect 6484 27538 6540 27540
rect 6244 27486 6270 27538
rect 6270 27486 6300 27538
rect 6324 27486 6334 27538
rect 6334 27486 6380 27538
rect 6404 27486 6450 27538
rect 6450 27486 6460 27538
rect 6484 27486 6514 27538
rect 6514 27486 6540 27538
rect 6244 27484 6300 27486
rect 6324 27484 6380 27486
rect 6404 27484 6460 27486
rect 6484 27484 6540 27486
rect 1876 26670 1932 26726
rect 2500 26687 2556 26726
rect 2500 26670 2502 26687
rect 2502 26670 2554 26687
rect 2554 26670 2556 26687
rect 3580 26206 3636 26208
rect 3660 26206 3716 26208
rect 3740 26206 3796 26208
rect 3820 26206 3876 26208
rect 3580 26154 3606 26206
rect 3606 26154 3636 26206
rect 3660 26154 3670 26206
rect 3670 26154 3716 26206
rect 3740 26154 3786 26206
rect 3786 26154 3796 26206
rect 3820 26154 3850 26206
rect 3850 26154 3876 26206
rect 3580 26152 3636 26154
rect 3660 26152 3716 26154
rect 3740 26152 3796 26154
rect 3820 26152 3876 26154
rect 8908 26206 8964 26208
rect 8988 26206 9044 26208
rect 9068 26206 9124 26208
rect 9148 26206 9204 26208
rect 8908 26154 8934 26206
rect 8934 26154 8964 26206
rect 8988 26154 8998 26206
rect 8998 26154 9044 26206
rect 9068 26154 9114 26206
rect 9114 26154 9124 26206
rect 9148 26154 9178 26206
rect 9178 26154 9204 26206
rect 8908 26152 8964 26154
rect 8988 26152 9044 26154
rect 9068 26152 9124 26154
rect 9148 26152 9204 26154
rect 6244 24874 6300 24876
rect 6324 24874 6380 24876
rect 6404 24874 6460 24876
rect 6484 24874 6540 24876
rect 6244 24822 6270 24874
rect 6270 24822 6300 24874
rect 6324 24822 6334 24874
rect 6334 24822 6380 24874
rect 6404 24822 6450 24874
rect 6450 24822 6460 24874
rect 6484 24822 6514 24874
rect 6514 24822 6540 24874
rect 6244 24820 6300 24822
rect 6324 24820 6380 24822
rect 6404 24820 6460 24822
rect 6484 24820 6540 24822
rect 1876 24006 1932 24062
rect 2500 24023 2556 24062
rect 2500 24006 2502 24023
rect 2502 24006 2554 24023
rect 2554 24006 2556 24023
rect 5299 24208 5355 24210
rect 5299 24156 5301 24208
rect 5301 24156 5353 24208
rect 5353 24156 5355 24208
rect 5299 24154 5355 24156
rect 5908 24154 5964 24210
rect 7732 24208 7788 24210
rect 7732 24156 7734 24208
rect 7734 24156 7786 24208
rect 7786 24156 7788 24208
rect 7732 24154 7788 24156
rect 8308 24154 8364 24210
rect 3580 23542 3636 23544
rect 3660 23542 3716 23544
rect 3740 23542 3796 23544
rect 3820 23542 3876 23544
rect 3580 23490 3606 23542
rect 3606 23490 3636 23542
rect 3660 23490 3670 23542
rect 3670 23490 3716 23542
rect 3740 23490 3786 23542
rect 3786 23490 3796 23542
rect 3820 23490 3850 23542
rect 3850 23490 3876 23542
rect 3580 23488 3636 23490
rect 3660 23488 3716 23490
rect 3740 23488 3796 23490
rect 3820 23488 3876 23490
rect 8908 23542 8964 23544
rect 8988 23542 9044 23544
rect 9068 23542 9124 23544
rect 9148 23542 9204 23544
rect 8908 23490 8934 23542
rect 8934 23490 8964 23542
rect 8988 23490 8998 23542
rect 8998 23490 9044 23542
rect 9068 23490 9114 23542
rect 9114 23490 9124 23542
rect 9148 23490 9178 23542
rect 9178 23490 9204 23542
rect 8908 23488 8964 23490
rect 8988 23488 9044 23490
rect 9068 23488 9124 23490
rect 9148 23488 9204 23490
rect 1108 21544 1164 21546
rect 1108 21492 1110 21544
rect 1110 21492 1162 21544
rect 1162 21492 1164 21544
rect 1108 21490 1164 21492
rect 6244 22210 6300 22212
rect 6324 22210 6380 22212
rect 6404 22210 6460 22212
rect 6484 22210 6540 22212
rect 6244 22158 6270 22210
rect 6270 22158 6300 22210
rect 6324 22158 6334 22210
rect 6334 22158 6380 22210
rect 6404 22158 6450 22210
rect 6450 22158 6460 22210
rect 6484 22158 6514 22210
rect 6514 22158 6540 22210
rect 6244 22156 6300 22158
rect 6324 22156 6380 22158
rect 6404 22156 6460 22158
rect 6484 22156 6540 22158
rect 3580 20878 3636 20880
rect 3660 20878 3716 20880
rect 3740 20878 3796 20880
rect 3820 20878 3876 20880
rect 3580 20826 3606 20878
rect 3606 20826 3636 20878
rect 3660 20826 3670 20878
rect 3670 20826 3716 20878
rect 3740 20826 3786 20878
rect 3786 20826 3796 20878
rect 3820 20826 3850 20878
rect 3850 20826 3876 20878
rect 3580 20824 3636 20826
rect 3660 20824 3716 20826
rect 3740 20824 3796 20826
rect 3820 20824 3876 20826
rect 8908 20878 8964 20880
rect 8988 20878 9044 20880
rect 9068 20878 9124 20880
rect 9148 20878 9204 20880
rect 8908 20826 8934 20878
rect 8934 20826 8964 20878
rect 8988 20826 8998 20878
rect 8998 20826 9044 20878
rect 9068 20826 9114 20878
rect 9114 20826 9124 20878
rect 9148 20826 9178 20878
rect 9178 20826 9204 20878
rect 8908 20824 8964 20826
rect 8988 20824 9044 20826
rect 9068 20824 9124 20826
rect 9148 20824 9204 20826
rect 6244 19546 6300 19548
rect 6324 19546 6380 19548
rect 6404 19546 6460 19548
rect 6484 19546 6540 19548
rect 6244 19494 6270 19546
rect 6270 19494 6300 19546
rect 6324 19494 6334 19546
rect 6334 19494 6380 19546
rect 6404 19494 6450 19546
rect 6450 19494 6460 19546
rect 6484 19494 6514 19546
rect 6514 19494 6540 19546
rect 6244 19492 6300 19494
rect 6324 19492 6380 19494
rect 6404 19492 6460 19494
rect 6484 19492 6540 19494
rect 1876 18678 1932 18734
rect 2500 18695 2556 18734
rect 2500 18678 2502 18695
rect 2502 18678 2554 18695
rect 2554 18678 2556 18695
rect 3580 18214 3636 18216
rect 3660 18214 3716 18216
rect 3740 18214 3796 18216
rect 3820 18214 3876 18216
rect 3580 18162 3606 18214
rect 3606 18162 3636 18214
rect 3660 18162 3670 18214
rect 3670 18162 3716 18214
rect 3740 18162 3786 18214
rect 3786 18162 3796 18214
rect 3820 18162 3850 18214
rect 3850 18162 3876 18214
rect 3580 18160 3636 18162
rect 3660 18160 3716 18162
rect 3740 18160 3796 18162
rect 3820 18160 3876 18162
rect 8908 18214 8964 18216
rect 8988 18214 9044 18216
rect 9068 18214 9124 18216
rect 9148 18214 9204 18216
rect 8908 18162 8934 18214
rect 8934 18162 8964 18214
rect 8988 18162 8998 18214
rect 8998 18162 9044 18214
rect 9068 18162 9114 18214
rect 9114 18162 9124 18214
rect 9148 18162 9178 18214
rect 9178 18162 9204 18214
rect 8908 18160 8964 18162
rect 8988 18160 9044 18162
rect 9068 18160 9124 18162
rect 9148 18160 9204 18162
rect 6244 16882 6300 16884
rect 6324 16882 6380 16884
rect 6404 16882 6460 16884
rect 6484 16882 6540 16884
rect 6244 16830 6270 16882
rect 6270 16830 6300 16882
rect 6324 16830 6334 16882
rect 6334 16830 6380 16882
rect 6404 16830 6450 16882
rect 6450 16830 6460 16882
rect 6484 16830 6514 16882
rect 6514 16830 6540 16882
rect 6244 16828 6300 16830
rect 6324 16828 6380 16830
rect 6404 16828 6460 16830
rect 6484 16828 6540 16830
rect 1876 16014 1932 16070
rect 2500 16031 2556 16070
rect 2500 16014 2502 16031
rect 2502 16014 2554 16031
rect 2554 16014 2556 16031
rect 3580 15550 3636 15552
rect 3660 15550 3716 15552
rect 3740 15550 3796 15552
rect 3820 15550 3876 15552
rect 3580 15498 3606 15550
rect 3606 15498 3636 15550
rect 3660 15498 3670 15550
rect 3670 15498 3716 15550
rect 3740 15498 3786 15550
rect 3786 15498 3796 15550
rect 3820 15498 3850 15550
rect 3850 15498 3876 15550
rect 3580 15496 3636 15498
rect 3660 15496 3716 15498
rect 3740 15496 3796 15498
rect 3820 15496 3876 15498
rect 8908 15550 8964 15552
rect 8988 15550 9044 15552
rect 9068 15550 9124 15552
rect 9148 15550 9204 15552
rect 8908 15498 8934 15550
rect 8934 15498 8964 15550
rect 8988 15498 8998 15550
rect 8998 15498 9044 15550
rect 9068 15498 9114 15550
rect 9114 15498 9124 15550
rect 9148 15498 9178 15550
rect 9178 15498 9204 15550
rect 8908 15496 8964 15498
rect 8988 15496 9044 15498
rect 9068 15496 9124 15498
rect 9148 15496 9204 15498
rect 6244 14218 6300 14220
rect 6324 14218 6380 14220
rect 6404 14218 6460 14220
rect 6484 14218 6540 14220
rect 6244 14166 6270 14218
rect 6270 14166 6300 14218
rect 6324 14166 6334 14218
rect 6334 14166 6380 14218
rect 6404 14166 6450 14218
rect 6450 14166 6460 14218
rect 6484 14166 6514 14218
rect 6514 14166 6540 14218
rect 6244 14164 6300 14166
rect 6324 14164 6380 14166
rect 6404 14164 6460 14166
rect 6484 14164 6540 14166
rect 1876 13350 1932 13406
rect 2500 13367 2556 13406
rect 2500 13350 2502 13367
rect 2502 13350 2554 13367
rect 2554 13350 2556 13367
rect 5299 13552 5355 13554
rect 5299 13500 5301 13552
rect 5301 13500 5353 13552
rect 5353 13500 5355 13552
rect 5299 13498 5355 13500
rect 5908 13498 5964 13554
rect 3580 12886 3636 12888
rect 3660 12886 3716 12888
rect 3740 12886 3796 12888
rect 3820 12886 3876 12888
rect 3580 12834 3606 12886
rect 3606 12834 3636 12886
rect 3660 12834 3670 12886
rect 3670 12834 3716 12886
rect 3740 12834 3786 12886
rect 3786 12834 3796 12886
rect 3820 12834 3850 12886
rect 3850 12834 3876 12886
rect 3580 12832 3636 12834
rect 3660 12832 3716 12834
rect 3740 12832 3796 12834
rect 3820 12832 3876 12834
rect 8908 12886 8964 12888
rect 8988 12886 9044 12888
rect 9068 12886 9124 12888
rect 9148 12886 9204 12888
rect 8908 12834 8934 12886
rect 8934 12834 8964 12886
rect 8988 12834 8998 12886
rect 8998 12834 9044 12886
rect 9068 12834 9114 12886
rect 9114 12834 9124 12886
rect 9148 12834 9178 12886
rect 9178 12834 9204 12886
rect 8908 12832 8964 12834
rect 8988 12832 9044 12834
rect 9068 12832 9124 12834
rect 9148 12832 9204 12834
rect 6244 11554 6300 11556
rect 6324 11554 6380 11556
rect 6404 11554 6460 11556
rect 6484 11554 6540 11556
rect 6244 11502 6270 11554
rect 6270 11502 6300 11554
rect 6324 11502 6334 11554
rect 6334 11502 6380 11554
rect 6404 11502 6450 11554
rect 6450 11502 6460 11554
rect 6484 11502 6514 11554
rect 6514 11502 6540 11554
rect 6244 11500 6300 11502
rect 6324 11500 6380 11502
rect 6404 11500 6460 11502
rect 6484 11500 6540 11502
rect 1876 10686 1932 10742
rect 2500 10703 2556 10742
rect 2500 10686 2502 10703
rect 2502 10686 2554 10703
rect 2554 10686 2556 10703
rect 3580 10222 3636 10224
rect 3660 10222 3716 10224
rect 3740 10222 3796 10224
rect 3820 10222 3876 10224
rect 3580 10170 3606 10222
rect 3606 10170 3636 10222
rect 3660 10170 3670 10222
rect 3670 10170 3716 10222
rect 3740 10170 3786 10222
rect 3786 10170 3796 10222
rect 3820 10170 3850 10222
rect 3850 10170 3876 10222
rect 3580 10168 3636 10170
rect 3660 10168 3716 10170
rect 3740 10168 3796 10170
rect 3820 10168 3876 10170
rect 8908 10222 8964 10224
rect 8988 10222 9044 10224
rect 9068 10222 9124 10224
rect 9148 10222 9204 10224
rect 8908 10170 8934 10222
rect 8934 10170 8964 10222
rect 8988 10170 8998 10222
rect 8998 10170 9044 10222
rect 9068 10170 9114 10222
rect 9114 10170 9124 10222
rect 9148 10170 9178 10222
rect 9178 10170 9204 10222
rect 8908 10168 8964 10170
rect 8988 10168 9044 10170
rect 9068 10168 9124 10170
rect 9148 10168 9204 10170
rect 6244 8890 6300 8892
rect 6324 8890 6380 8892
rect 6404 8890 6460 8892
rect 6484 8890 6540 8892
rect 6244 8838 6270 8890
rect 6270 8838 6300 8890
rect 6324 8838 6334 8890
rect 6334 8838 6380 8890
rect 6404 8838 6450 8890
rect 6450 8838 6460 8890
rect 6484 8838 6514 8890
rect 6514 8838 6540 8890
rect 6244 8836 6300 8838
rect 6324 8836 6380 8838
rect 6404 8836 6460 8838
rect 6484 8836 6540 8838
rect 1876 8022 1932 8078
rect 2500 8039 2556 8078
rect 2500 8022 2502 8039
rect 2502 8022 2554 8039
rect 2554 8022 2556 8039
rect 3580 7558 3636 7560
rect 3660 7558 3716 7560
rect 3740 7558 3796 7560
rect 3820 7558 3876 7560
rect 3580 7506 3606 7558
rect 3606 7506 3636 7558
rect 3660 7506 3670 7558
rect 3670 7506 3716 7558
rect 3740 7506 3786 7558
rect 3786 7506 3796 7558
rect 3820 7506 3850 7558
rect 3850 7506 3876 7558
rect 3580 7504 3636 7506
rect 3660 7504 3716 7506
rect 3740 7504 3796 7506
rect 3820 7504 3876 7506
rect 8908 7558 8964 7560
rect 8988 7558 9044 7560
rect 9068 7558 9124 7560
rect 9148 7558 9204 7560
rect 8908 7506 8934 7558
rect 8934 7506 8964 7558
rect 8988 7506 8998 7558
rect 8998 7506 9044 7558
rect 9068 7506 9114 7558
rect 9114 7506 9124 7558
rect 9148 7506 9178 7558
rect 9178 7506 9204 7558
rect 8908 7504 8964 7506
rect 8988 7504 9044 7506
rect 9068 7504 9124 7506
rect 9148 7504 9204 7506
rect 6244 6226 6300 6228
rect 6324 6226 6380 6228
rect 6404 6226 6460 6228
rect 6484 6226 6540 6228
rect 6244 6174 6270 6226
rect 6270 6174 6300 6226
rect 6324 6174 6334 6226
rect 6334 6174 6380 6226
rect 6404 6174 6450 6226
rect 6450 6174 6460 6226
rect 6484 6174 6514 6226
rect 6514 6174 6540 6226
rect 6244 6172 6300 6174
rect 6324 6172 6380 6174
rect 6404 6172 6460 6174
rect 6484 6172 6540 6174
rect 1876 5358 1932 5414
rect 2500 5375 2556 5414
rect 2500 5358 2502 5375
rect 2502 5358 2554 5375
rect 2554 5358 2556 5375
rect 3580 4894 3636 4896
rect 3660 4894 3716 4896
rect 3740 4894 3796 4896
rect 3820 4894 3876 4896
rect 3580 4842 3606 4894
rect 3606 4842 3636 4894
rect 3660 4842 3670 4894
rect 3670 4842 3716 4894
rect 3740 4842 3786 4894
rect 3786 4842 3796 4894
rect 3820 4842 3850 4894
rect 3850 4842 3876 4894
rect 3580 4840 3636 4842
rect 3660 4840 3716 4842
rect 3740 4840 3796 4842
rect 3820 4840 3876 4842
rect 8908 4894 8964 4896
rect 8988 4894 9044 4896
rect 9068 4894 9124 4896
rect 9148 4894 9204 4896
rect 8908 4842 8934 4894
rect 8934 4842 8964 4894
rect 8988 4842 8998 4894
rect 8998 4842 9044 4894
rect 9068 4842 9114 4894
rect 9114 4842 9124 4894
rect 9148 4842 9178 4894
rect 9178 4842 9204 4894
rect 8908 4840 8964 4842
rect 8988 4840 9044 4842
rect 9068 4840 9124 4842
rect 9148 4840 9204 4842
rect 6244 3562 6300 3564
rect 6324 3562 6380 3564
rect 6404 3562 6460 3564
rect 6484 3562 6540 3564
rect 6244 3510 6270 3562
rect 6270 3510 6300 3562
rect 6324 3510 6334 3562
rect 6334 3510 6380 3562
rect 6404 3510 6450 3562
rect 6450 3510 6460 3562
rect 6484 3510 6514 3562
rect 6514 3510 6540 3562
rect 6244 3508 6300 3510
rect 6324 3508 6380 3510
rect 6404 3508 6460 3510
rect 6484 3508 6540 3510
rect 1876 2694 1932 2750
rect 2500 2711 2556 2750
rect 2500 2694 2502 2711
rect 2502 2694 2554 2711
rect 2554 2694 2556 2711
rect 5299 2896 5355 2898
rect 5299 2844 5301 2896
rect 5301 2844 5353 2896
rect 5353 2844 5355 2896
rect 5299 2842 5355 2844
rect 5908 2842 5964 2898
rect 3580 2230 3636 2232
rect 3660 2230 3716 2232
rect 3740 2230 3796 2232
rect 3820 2230 3876 2232
rect 3580 2178 3606 2230
rect 3606 2178 3636 2230
rect 3660 2178 3670 2230
rect 3670 2178 3716 2230
rect 3740 2178 3786 2230
rect 3786 2178 3796 2230
rect 3820 2178 3850 2230
rect 3850 2178 3876 2230
rect 3580 2176 3636 2178
rect 3660 2176 3716 2178
rect 3740 2176 3796 2178
rect 3820 2176 3876 2178
rect 8908 2230 8964 2232
rect 8988 2230 9044 2232
rect 9068 2230 9124 2232
rect 9148 2230 9204 2232
rect 8908 2178 8934 2230
rect 8934 2178 8964 2230
rect 8988 2178 8998 2230
rect 8998 2178 9044 2230
rect 9068 2178 9114 2230
rect 9114 2178 9124 2230
rect 9148 2178 9178 2230
rect 9178 2178 9204 2230
rect 8908 2176 8964 2178
rect 8988 2176 9044 2178
rect 9068 2176 9124 2178
rect 9148 2176 9204 2178
rect 1876 1564 1932 1566
rect 1876 1512 1878 1564
rect 1878 1512 1930 1564
rect 1930 1512 1932 1564
rect 1876 1510 1932 1512
rect 6244 898 6300 900
rect 6324 898 6380 900
rect 6404 898 6460 900
rect 6484 898 6540 900
rect 6244 846 6270 898
rect 6270 846 6300 898
rect 6324 846 6334 898
rect 6334 846 6380 898
rect 6404 846 6450 898
rect 6450 846 6460 898
rect 6484 846 6514 898
rect 6514 846 6540 898
rect 6244 844 6300 846
rect 6324 844 6380 846
rect 6404 844 6460 846
rect 6484 844 6540 846
<< metal3 >>
rect 800 52752 920 53008
rect 3568 52852 3888 52853
rect 3568 52788 3576 52852
rect 3640 52788 3656 52852
rect 3720 52788 3736 52852
rect 3800 52788 3816 52852
rect 3880 52788 3888 52852
rect 3568 52787 3888 52788
rect 8896 52852 9216 52853
rect 8896 52788 8904 52852
rect 8968 52788 8984 52852
rect 9048 52788 9064 52852
rect 9128 52788 9144 52852
rect 9208 52788 9216 52852
rect 8896 52787 9216 52788
rect 830 52480 890 52752
rect 1343 52480 1409 52483
rect 830 52478 1409 52480
rect 830 52422 1348 52478
rect 1404 52422 1409 52478
rect 830 52420 1409 52422
rect 1343 52417 1409 52420
rect 1103 52036 1169 52039
rect 830 52034 1169 52036
rect 830 51978 1108 52034
rect 1164 51978 1169 52034
rect 830 51976 1169 51978
rect 830 51648 890 51976
rect 1103 51973 1169 51976
rect 800 51392 920 51648
rect 6232 51520 6552 51521
rect 6232 51456 6240 51520
rect 6304 51456 6320 51520
rect 6384 51456 6400 51520
rect 6464 51456 6480 51520
rect 6544 51456 6552 51520
rect 6232 51455 6552 51456
rect 1103 50704 1169 50707
rect 830 50702 1169 50704
rect 830 50646 1108 50702
rect 1164 50646 1169 50702
rect 830 50644 1169 50646
rect 830 50288 890 50644
rect 1103 50641 1169 50644
rect 800 50032 920 50288
rect 3568 50188 3888 50189
rect 3568 50124 3576 50188
rect 3640 50124 3656 50188
rect 3720 50124 3736 50188
rect 3800 50124 3816 50188
rect 3880 50124 3888 50188
rect 3568 50123 3888 50124
rect 8896 50188 9216 50189
rect 8896 50124 8904 50188
rect 8968 50124 8984 50188
rect 9048 50124 9064 50188
rect 9128 50124 9144 50188
rect 9208 50124 9216 50188
rect 8896 50123 9216 50124
rect 6232 48856 6552 48857
rect 6232 48792 6240 48856
rect 6304 48792 6320 48856
rect 6384 48792 6400 48856
rect 6464 48792 6480 48856
rect 6544 48792 6552 48856
rect 6232 48791 6552 48792
rect 1103 48040 1169 48043
rect 830 48038 1169 48040
rect 830 47982 1108 48038
rect 1164 47982 1169 48038
rect 830 47980 1169 47982
rect 830 47568 890 47980
rect 1103 47977 1169 47980
rect 800 47312 920 47568
rect 3568 47524 3888 47525
rect 3568 47460 3576 47524
rect 3640 47460 3656 47524
rect 3720 47460 3736 47524
rect 3800 47460 3816 47524
rect 3880 47460 3888 47524
rect 3568 47459 3888 47460
rect 8896 47524 9216 47525
rect 8896 47460 8904 47524
rect 8968 47460 8984 47524
rect 9048 47460 9064 47524
rect 9128 47460 9144 47524
rect 9208 47460 9216 47524
rect 8896 47459 9216 47460
rect 6232 46192 6552 46193
rect 6232 46128 6240 46192
rect 6304 46128 6320 46192
rect 6384 46128 6400 46192
rect 6464 46128 6480 46192
rect 6544 46128 6552 46192
rect 6232 46127 6552 46128
rect 2831 45524 2897 45527
rect 3455 45524 3521 45527
rect 2831 45522 3521 45524
rect 2831 45466 2836 45522
rect 2892 45466 3460 45522
rect 3516 45466 3521 45522
rect 2831 45464 3521 45466
rect 2831 45461 2897 45464
rect 3455 45461 3521 45464
rect 1103 45376 1169 45379
rect 830 45374 1169 45376
rect 830 45318 1108 45374
rect 1164 45318 1169 45374
rect 830 45316 1169 45318
rect 830 44984 890 45316
rect 1103 45313 1169 45316
rect 800 44728 920 44984
rect 3568 44860 3888 44861
rect 3568 44796 3576 44860
rect 3640 44796 3656 44860
rect 3720 44796 3736 44860
rect 3800 44796 3816 44860
rect 3880 44796 3888 44860
rect 3568 44795 3888 44796
rect 8896 44860 9216 44861
rect 8896 44796 8904 44860
rect 8968 44796 8984 44860
rect 9048 44796 9064 44860
rect 9128 44796 9144 44860
rect 9208 44796 9216 44860
rect 8896 44795 9216 44796
rect 6232 43528 6552 43529
rect 6232 43464 6240 43528
rect 6304 43464 6320 43528
rect 6384 43464 6400 43528
rect 6464 43464 6480 43528
rect 6544 43464 6552 43528
rect 6232 43463 6552 43464
rect 1103 42712 1169 42715
rect 830 42710 1169 42712
rect 830 42654 1108 42710
rect 1164 42654 1169 42710
rect 830 42652 1169 42654
rect 830 42264 890 42652
rect 1103 42649 1169 42652
rect 800 42008 920 42264
rect 3568 42196 3888 42197
rect 3568 42132 3576 42196
rect 3640 42132 3656 42196
rect 3720 42132 3736 42196
rect 3800 42132 3816 42196
rect 3880 42132 3888 42196
rect 3568 42131 3888 42132
rect 8896 42196 9216 42197
rect 8896 42132 8904 42196
rect 8968 42132 8984 42196
rect 9048 42132 9064 42196
rect 9128 42132 9144 42196
rect 9208 42132 9216 42196
rect 8896 42131 9216 42132
rect 6232 40864 6552 40865
rect 6232 40800 6240 40864
rect 6304 40800 6320 40864
rect 6384 40800 6400 40864
rect 6464 40800 6480 40864
rect 6544 40800 6552 40864
rect 6232 40799 6552 40800
rect 1103 40196 1169 40199
rect 830 40194 1169 40196
rect 830 40138 1108 40194
rect 1164 40138 1169 40194
rect 830 40136 1169 40138
rect 830 39680 890 40136
rect 1103 40133 1169 40136
rect 800 39424 920 39680
rect 3568 39532 3888 39533
rect 3568 39468 3576 39532
rect 3640 39468 3656 39532
rect 3720 39468 3736 39532
rect 3800 39468 3816 39532
rect 3880 39468 3888 39532
rect 3568 39467 3888 39468
rect 8896 39532 9216 39533
rect 8896 39468 8904 39532
rect 8968 39468 8984 39532
rect 9048 39468 9064 39532
rect 9128 39468 9144 39532
rect 9208 39468 9216 39532
rect 8896 39467 9216 39468
rect 6232 38200 6552 38201
rect 6232 38136 6240 38200
rect 6304 38136 6320 38200
rect 6384 38136 6400 38200
rect 6464 38136 6480 38200
rect 6544 38136 6552 38200
rect 6232 38135 6552 38136
rect 1103 37384 1169 37387
rect 830 37382 1169 37384
rect 830 37326 1108 37382
rect 1164 37326 1169 37382
rect 830 37324 1169 37326
rect 830 36960 890 37324
rect 1103 37321 1169 37324
rect 800 36704 920 36960
rect 3568 36868 3888 36869
rect 3568 36804 3576 36868
rect 3640 36804 3656 36868
rect 3720 36804 3736 36868
rect 3800 36804 3816 36868
rect 3880 36804 3888 36868
rect 3568 36803 3888 36804
rect 8896 36868 9216 36869
rect 8896 36804 8904 36868
rect 8968 36804 8984 36868
rect 9048 36804 9064 36868
rect 9128 36804 9144 36868
rect 9208 36804 9216 36868
rect 8896 36803 9216 36804
rect 6232 35536 6552 35537
rect 6232 35472 6240 35536
rect 6304 35472 6320 35536
rect 6384 35472 6400 35536
rect 6464 35472 6480 35536
rect 6544 35472 6552 35536
rect 6232 35471 6552 35472
rect 5294 34868 5360 34871
rect 5903 34868 5969 34871
rect 5294 34866 5969 34868
rect 5294 34810 5299 34866
rect 5355 34810 5908 34866
rect 5964 34810 5969 34866
rect 5294 34808 5969 34810
rect 5294 34805 5360 34808
rect 5903 34805 5969 34808
rect 1871 34720 1937 34723
rect 2495 34720 2561 34723
rect 1871 34718 2561 34720
rect 1871 34662 1876 34718
rect 1932 34662 2500 34718
rect 2556 34662 2561 34718
rect 1871 34660 2561 34662
rect 1871 34657 1937 34660
rect 2495 34657 2561 34660
rect 3568 34204 3888 34205
rect 3568 34140 3576 34204
rect 3640 34140 3656 34204
rect 3720 34140 3736 34204
rect 3800 34140 3816 34204
rect 3880 34140 3888 34204
rect 3568 34139 3888 34140
rect 8896 34204 9216 34205
rect 8896 34140 8904 34204
rect 8968 34140 8984 34204
rect 9048 34140 9064 34204
rect 9128 34140 9144 34204
rect 9208 34140 9216 34204
rect 8896 34139 9216 34140
rect 6232 32872 6552 32873
rect 6232 32808 6240 32872
rect 6304 32808 6320 32872
rect 6384 32808 6400 32872
rect 6464 32808 6480 32872
rect 6544 32808 6552 32872
rect 6232 32807 6552 32808
rect 1103 32056 1169 32059
rect 830 32054 1169 32056
rect 830 31998 1108 32054
rect 1164 31998 1169 32054
rect 830 31996 1169 31998
rect 830 31656 890 31996
rect 1103 31993 1169 31996
rect 800 31400 920 31656
rect 3568 31540 3888 31541
rect 3568 31476 3576 31540
rect 3640 31476 3656 31540
rect 3720 31476 3736 31540
rect 3800 31476 3816 31540
rect 3880 31476 3888 31540
rect 3568 31475 3888 31476
rect 8896 31540 9216 31541
rect 8896 31476 8904 31540
rect 8968 31476 8984 31540
rect 9048 31476 9064 31540
rect 9128 31476 9144 31540
rect 9208 31476 9216 31540
rect 8896 31475 9216 31476
rect 6232 30208 6552 30209
rect 6232 30144 6240 30208
rect 6304 30144 6320 30208
rect 6384 30144 6400 30208
rect 6464 30144 6480 30208
rect 6544 30144 6552 30208
rect 6232 30143 6552 30144
rect 1871 29392 1937 29395
rect 2495 29392 2561 29395
rect 1871 29390 2561 29392
rect 1871 29334 1876 29390
rect 1932 29334 2500 29390
rect 2556 29334 2561 29390
rect 1871 29332 2561 29334
rect 1871 29329 1937 29332
rect 2495 29329 2561 29332
rect 3568 28876 3888 28877
rect 3568 28812 3576 28876
rect 3640 28812 3656 28876
rect 3720 28812 3736 28876
rect 3800 28812 3816 28876
rect 3880 28812 3888 28876
rect 3568 28811 3888 28812
rect 8896 28876 9216 28877
rect 8896 28812 8904 28876
rect 8968 28812 8984 28876
rect 9048 28812 9064 28876
rect 9128 28812 9144 28876
rect 9208 28812 9216 28876
rect 8896 28811 9216 28812
rect 6232 27544 6552 27545
rect 6232 27480 6240 27544
rect 6304 27480 6320 27544
rect 6384 27480 6400 27544
rect 6464 27480 6480 27544
rect 6544 27480 6552 27544
rect 6232 27479 6552 27480
rect 1871 26728 1937 26731
rect 2495 26728 2561 26731
rect 1871 26726 2561 26728
rect 1871 26670 1876 26726
rect 1932 26670 2500 26726
rect 2556 26670 2561 26726
rect 1871 26668 2561 26670
rect 1871 26665 1937 26668
rect 2495 26665 2561 26668
rect 3568 26212 3888 26213
rect 3568 26148 3576 26212
rect 3640 26148 3656 26212
rect 3720 26148 3736 26212
rect 3800 26148 3816 26212
rect 3880 26148 3888 26212
rect 3568 26147 3888 26148
rect 8896 26212 9216 26213
rect 8896 26148 8904 26212
rect 8968 26148 8984 26212
rect 9048 26148 9064 26212
rect 9128 26148 9144 26212
rect 9208 26148 9216 26212
rect 8896 26147 9216 26148
rect 6232 24880 6552 24881
rect 6232 24816 6240 24880
rect 6304 24816 6320 24880
rect 6384 24816 6400 24880
rect 6464 24816 6480 24880
rect 6544 24816 6552 24880
rect 6232 24815 6552 24816
rect 5294 24212 5360 24215
rect 5903 24212 5969 24215
rect 5294 24210 5969 24212
rect 5294 24154 5299 24210
rect 5355 24154 5908 24210
rect 5964 24154 5969 24210
rect 5294 24152 5969 24154
rect 5294 24149 5360 24152
rect 5903 24149 5969 24152
rect 7727 24212 7793 24215
rect 8303 24212 8369 24215
rect 7727 24210 8369 24212
rect 7727 24154 7732 24210
rect 7788 24154 8308 24210
rect 8364 24154 8369 24210
rect 7727 24152 8369 24154
rect 7727 24149 7793 24152
rect 8303 24149 8369 24152
rect 1871 24064 1937 24067
rect 2495 24064 2561 24067
rect 1871 24062 2561 24064
rect 1871 24006 1876 24062
rect 1932 24006 2500 24062
rect 2556 24006 2561 24062
rect 1871 24004 2561 24006
rect 1871 24001 1937 24004
rect 2495 24001 2561 24004
rect 3568 23548 3888 23549
rect 3568 23484 3576 23548
rect 3640 23484 3656 23548
rect 3720 23484 3736 23548
rect 3800 23484 3816 23548
rect 3880 23484 3888 23548
rect 3568 23483 3888 23484
rect 8896 23548 9216 23549
rect 8896 23484 8904 23548
rect 8968 23484 8984 23548
rect 9048 23484 9064 23548
rect 9128 23484 9144 23548
rect 9208 23484 9216 23548
rect 8896 23483 9216 23484
rect 6232 22216 6552 22217
rect 6232 22152 6240 22216
rect 6304 22152 6320 22216
rect 6384 22152 6400 22216
rect 6464 22152 6480 22216
rect 6544 22152 6552 22216
rect 6232 22151 6552 22152
rect 1103 21548 1169 21551
rect 830 21546 1169 21548
rect 830 21490 1108 21546
rect 1164 21490 1169 21546
rect 830 21488 1169 21490
rect 830 21048 890 21488
rect 1103 21485 1169 21488
rect 800 20792 920 21048
rect 3568 20884 3888 20885
rect 3568 20820 3576 20884
rect 3640 20820 3656 20884
rect 3720 20820 3736 20884
rect 3800 20820 3816 20884
rect 3880 20820 3888 20884
rect 3568 20819 3888 20820
rect 8896 20884 9216 20885
rect 8896 20820 8904 20884
rect 8968 20820 8984 20884
rect 9048 20820 9064 20884
rect 9128 20820 9144 20884
rect 9208 20820 9216 20884
rect 8896 20819 9216 20820
rect 6232 19552 6552 19553
rect 6232 19488 6240 19552
rect 6304 19488 6320 19552
rect 6384 19488 6400 19552
rect 6464 19488 6480 19552
rect 6544 19488 6552 19552
rect 6232 19487 6552 19488
rect 1871 18736 1937 18739
rect 2495 18736 2561 18739
rect 1871 18734 2561 18736
rect 1871 18678 1876 18734
rect 1932 18678 2500 18734
rect 2556 18678 2561 18734
rect 1871 18676 2561 18678
rect 1871 18673 1937 18676
rect 2495 18673 2561 18676
rect 3568 18220 3888 18221
rect 3568 18156 3576 18220
rect 3640 18156 3656 18220
rect 3720 18156 3736 18220
rect 3800 18156 3816 18220
rect 3880 18156 3888 18220
rect 3568 18155 3888 18156
rect 8896 18220 9216 18221
rect 8896 18156 8904 18220
rect 8968 18156 8984 18220
rect 9048 18156 9064 18220
rect 9128 18156 9144 18220
rect 9208 18156 9216 18220
rect 8896 18155 9216 18156
rect 6232 16888 6552 16889
rect 6232 16824 6240 16888
rect 6304 16824 6320 16888
rect 6384 16824 6400 16888
rect 6464 16824 6480 16888
rect 6544 16824 6552 16888
rect 6232 16823 6552 16824
rect 1871 16072 1937 16075
rect 2495 16072 2561 16075
rect 1871 16070 2561 16072
rect 1871 16014 1876 16070
rect 1932 16014 2500 16070
rect 2556 16014 2561 16070
rect 1871 16012 2561 16014
rect 1871 16009 1937 16012
rect 2495 16009 2561 16012
rect 3568 15556 3888 15557
rect 3568 15492 3576 15556
rect 3640 15492 3656 15556
rect 3720 15492 3736 15556
rect 3800 15492 3816 15556
rect 3880 15492 3888 15556
rect 3568 15491 3888 15492
rect 8896 15556 9216 15557
rect 8896 15492 8904 15556
rect 8968 15492 8984 15556
rect 9048 15492 9064 15556
rect 9128 15492 9144 15556
rect 9208 15492 9216 15556
rect 8896 15491 9216 15492
rect 6232 14224 6552 14225
rect 6232 14160 6240 14224
rect 6304 14160 6320 14224
rect 6384 14160 6400 14224
rect 6464 14160 6480 14224
rect 6544 14160 6552 14224
rect 6232 14159 6552 14160
rect 5294 13556 5360 13559
rect 5903 13556 5969 13559
rect 5294 13554 5969 13556
rect 5294 13498 5299 13554
rect 5355 13498 5908 13554
rect 5964 13498 5969 13554
rect 5294 13496 5969 13498
rect 5294 13493 5360 13496
rect 5903 13493 5969 13496
rect 1871 13408 1937 13411
rect 2495 13408 2561 13411
rect 1871 13406 2561 13408
rect 1871 13350 1876 13406
rect 1932 13350 2500 13406
rect 2556 13350 2561 13406
rect 1871 13348 2561 13350
rect 1871 13345 1937 13348
rect 2495 13345 2561 13348
rect 3568 12892 3888 12893
rect 3568 12828 3576 12892
rect 3640 12828 3656 12892
rect 3720 12828 3736 12892
rect 3800 12828 3816 12892
rect 3880 12828 3888 12892
rect 3568 12827 3888 12828
rect 8896 12892 9216 12893
rect 8896 12828 8904 12892
rect 8968 12828 8984 12892
rect 9048 12828 9064 12892
rect 9128 12828 9144 12892
rect 9208 12828 9216 12892
rect 8896 12827 9216 12828
rect 6232 11560 6552 11561
rect 6232 11496 6240 11560
rect 6304 11496 6320 11560
rect 6384 11496 6400 11560
rect 6464 11496 6480 11560
rect 6544 11496 6552 11560
rect 6232 11495 6552 11496
rect 1871 10744 1937 10747
rect 2495 10744 2561 10747
rect 1871 10742 2561 10744
rect 1871 10686 1876 10742
rect 1932 10686 2500 10742
rect 2556 10686 2561 10742
rect 1871 10684 2561 10686
rect 1871 10681 1937 10684
rect 2495 10681 2561 10684
rect 3568 10228 3888 10229
rect 3568 10164 3576 10228
rect 3640 10164 3656 10228
rect 3720 10164 3736 10228
rect 3800 10164 3816 10228
rect 3880 10164 3888 10228
rect 3568 10163 3888 10164
rect 8896 10228 9216 10229
rect 8896 10164 8904 10228
rect 8968 10164 8984 10228
rect 9048 10164 9064 10228
rect 9128 10164 9144 10228
rect 9208 10164 9216 10228
rect 8896 10163 9216 10164
rect 6232 8896 6552 8897
rect 6232 8832 6240 8896
rect 6304 8832 6320 8896
rect 6384 8832 6400 8896
rect 6464 8832 6480 8896
rect 6544 8832 6552 8896
rect 6232 8831 6552 8832
rect 1871 8080 1937 8083
rect 2495 8080 2561 8083
rect 1871 8078 2561 8080
rect 1871 8022 1876 8078
rect 1932 8022 2500 8078
rect 2556 8022 2561 8078
rect 1871 8020 2561 8022
rect 1871 8017 1937 8020
rect 2495 8017 2561 8020
rect 3568 7564 3888 7565
rect 3568 7500 3576 7564
rect 3640 7500 3656 7564
rect 3720 7500 3736 7564
rect 3800 7500 3816 7564
rect 3880 7500 3888 7564
rect 3568 7499 3888 7500
rect 8896 7564 9216 7565
rect 8896 7500 8904 7564
rect 8968 7500 8984 7564
rect 9048 7500 9064 7564
rect 9128 7500 9144 7564
rect 9208 7500 9216 7564
rect 8896 7499 9216 7500
rect 6232 6232 6552 6233
rect 6232 6168 6240 6232
rect 6304 6168 6320 6232
rect 6384 6168 6400 6232
rect 6464 6168 6480 6232
rect 6544 6168 6552 6232
rect 6232 6167 6552 6168
rect 1871 5416 1937 5419
rect 2495 5416 2561 5419
rect 1871 5414 2561 5416
rect 1871 5358 1876 5414
rect 1932 5358 2500 5414
rect 2556 5358 2561 5414
rect 1871 5356 2561 5358
rect 1871 5353 1937 5356
rect 2495 5353 2561 5356
rect 3568 4900 3888 4901
rect 3568 4836 3576 4900
rect 3640 4836 3656 4900
rect 3720 4836 3736 4900
rect 3800 4836 3816 4900
rect 3880 4836 3888 4900
rect 3568 4835 3888 4836
rect 8896 4900 9216 4901
rect 8896 4836 8904 4900
rect 8968 4836 8984 4900
rect 9048 4836 9064 4900
rect 9128 4836 9144 4900
rect 9208 4836 9216 4900
rect 8896 4835 9216 4836
rect 6232 3568 6552 3569
rect 6232 3504 6240 3568
rect 6304 3504 6320 3568
rect 6384 3504 6400 3568
rect 6464 3504 6480 3568
rect 6544 3504 6552 3568
rect 6232 3503 6552 3504
rect 5294 2900 5360 2903
rect 5903 2900 5969 2903
rect 5294 2898 5969 2900
rect 5294 2842 5299 2898
rect 5355 2842 5908 2898
rect 5964 2842 5969 2898
rect 5294 2840 5969 2842
rect 5294 2837 5360 2840
rect 5903 2837 5969 2840
rect 1871 2752 1937 2755
rect 2495 2752 2561 2755
rect 1871 2750 2561 2752
rect 1871 2694 1876 2750
rect 1932 2694 2500 2750
rect 2556 2694 2561 2750
rect 1871 2692 2561 2694
rect 1871 2689 1937 2692
rect 2495 2689 2561 2692
rect 3568 2236 3888 2237
rect 3568 2172 3576 2236
rect 3640 2172 3656 2236
rect 3720 2172 3736 2236
rect 3800 2172 3816 2236
rect 3880 2172 3888 2236
rect 3568 2171 3888 2172
rect 8896 2236 9216 2237
rect 8896 2172 8904 2236
rect 8968 2172 8984 2236
rect 9048 2172 9064 2236
rect 9128 2172 9144 2236
rect 9208 2172 9216 2236
rect 8896 2171 9216 2172
rect 1871 1568 1937 1571
rect 830 1566 1937 1568
rect 830 1510 1876 1566
rect 1932 1510 1937 1566
rect 830 1508 1937 1510
rect 830 1056 890 1508
rect 1871 1505 1937 1508
rect 800 800 920 1056
rect 6232 904 6552 905
rect 6232 840 6240 904
rect 6304 840 6320 904
rect 6384 840 6400 904
rect 6464 840 6480 904
rect 6544 840 6552 904
rect 6232 839 6552 840
<< via3 >>
rect 3576 52848 3640 52852
rect 3576 52792 3580 52848
rect 3580 52792 3636 52848
rect 3636 52792 3640 52848
rect 3576 52788 3640 52792
rect 3656 52848 3720 52852
rect 3656 52792 3660 52848
rect 3660 52792 3716 52848
rect 3716 52792 3720 52848
rect 3656 52788 3720 52792
rect 3736 52848 3800 52852
rect 3736 52792 3740 52848
rect 3740 52792 3796 52848
rect 3796 52792 3800 52848
rect 3736 52788 3800 52792
rect 3816 52848 3880 52852
rect 3816 52792 3820 52848
rect 3820 52792 3876 52848
rect 3876 52792 3880 52848
rect 3816 52788 3880 52792
rect 8904 52848 8968 52852
rect 8904 52792 8908 52848
rect 8908 52792 8964 52848
rect 8964 52792 8968 52848
rect 8904 52788 8968 52792
rect 8984 52848 9048 52852
rect 8984 52792 8988 52848
rect 8988 52792 9044 52848
rect 9044 52792 9048 52848
rect 8984 52788 9048 52792
rect 9064 52848 9128 52852
rect 9064 52792 9068 52848
rect 9068 52792 9124 52848
rect 9124 52792 9128 52848
rect 9064 52788 9128 52792
rect 9144 52848 9208 52852
rect 9144 52792 9148 52848
rect 9148 52792 9204 52848
rect 9204 52792 9208 52848
rect 9144 52788 9208 52792
rect 6240 51516 6304 51520
rect 6240 51460 6244 51516
rect 6244 51460 6300 51516
rect 6300 51460 6304 51516
rect 6240 51456 6304 51460
rect 6320 51516 6384 51520
rect 6320 51460 6324 51516
rect 6324 51460 6380 51516
rect 6380 51460 6384 51516
rect 6320 51456 6384 51460
rect 6400 51516 6464 51520
rect 6400 51460 6404 51516
rect 6404 51460 6460 51516
rect 6460 51460 6464 51516
rect 6400 51456 6464 51460
rect 6480 51516 6544 51520
rect 6480 51460 6484 51516
rect 6484 51460 6540 51516
rect 6540 51460 6544 51516
rect 6480 51456 6544 51460
rect 3576 50184 3640 50188
rect 3576 50128 3580 50184
rect 3580 50128 3636 50184
rect 3636 50128 3640 50184
rect 3576 50124 3640 50128
rect 3656 50184 3720 50188
rect 3656 50128 3660 50184
rect 3660 50128 3716 50184
rect 3716 50128 3720 50184
rect 3656 50124 3720 50128
rect 3736 50184 3800 50188
rect 3736 50128 3740 50184
rect 3740 50128 3796 50184
rect 3796 50128 3800 50184
rect 3736 50124 3800 50128
rect 3816 50184 3880 50188
rect 3816 50128 3820 50184
rect 3820 50128 3876 50184
rect 3876 50128 3880 50184
rect 3816 50124 3880 50128
rect 8904 50184 8968 50188
rect 8904 50128 8908 50184
rect 8908 50128 8964 50184
rect 8964 50128 8968 50184
rect 8904 50124 8968 50128
rect 8984 50184 9048 50188
rect 8984 50128 8988 50184
rect 8988 50128 9044 50184
rect 9044 50128 9048 50184
rect 8984 50124 9048 50128
rect 9064 50184 9128 50188
rect 9064 50128 9068 50184
rect 9068 50128 9124 50184
rect 9124 50128 9128 50184
rect 9064 50124 9128 50128
rect 9144 50184 9208 50188
rect 9144 50128 9148 50184
rect 9148 50128 9204 50184
rect 9204 50128 9208 50184
rect 9144 50124 9208 50128
rect 6240 48852 6304 48856
rect 6240 48796 6244 48852
rect 6244 48796 6300 48852
rect 6300 48796 6304 48852
rect 6240 48792 6304 48796
rect 6320 48852 6384 48856
rect 6320 48796 6324 48852
rect 6324 48796 6380 48852
rect 6380 48796 6384 48852
rect 6320 48792 6384 48796
rect 6400 48852 6464 48856
rect 6400 48796 6404 48852
rect 6404 48796 6460 48852
rect 6460 48796 6464 48852
rect 6400 48792 6464 48796
rect 6480 48852 6544 48856
rect 6480 48796 6484 48852
rect 6484 48796 6540 48852
rect 6540 48796 6544 48852
rect 6480 48792 6544 48796
rect 3576 47520 3640 47524
rect 3576 47464 3580 47520
rect 3580 47464 3636 47520
rect 3636 47464 3640 47520
rect 3576 47460 3640 47464
rect 3656 47520 3720 47524
rect 3656 47464 3660 47520
rect 3660 47464 3716 47520
rect 3716 47464 3720 47520
rect 3656 47460 3720 47464
rect 3736 47520 3800 47524
rect 3736 47464 3740 47520
rect 3740 47464 3796 47520
rect 3796 47464 3800 47520
rect 3736 47460 3800 47464
rect 3816 47520 3880 47524
rect 3816 47464 3820 47520
rect 3820 47464 3876 47520
rect 3876 47464 3880 47520
rect 3816 47460 3880 47464
rect 8904 47520 8968 47524
rect 8904 47464 8908 47520
rect 8908 47464 8964 47520
rect 8964 47464 8968 47520
rect 8904 47460 8968 47464
rect 8984 47520 9048 47524
rect 8984 47464 8988 47520
rect 8988 47464 9044 47520
rect 9044 47464 9048 47520
rect 8984 47460 9048 47464
rect 9064 47520 9128 47524
rect 9064 47464 9068 47520
rect 9068 47464 9124 47520
rect 9124 47464 9128 47520
rect 9064 47460 9128 47464
rect 9144 47520 9208 47524
rect 9144 47464 9148 47520
rect 9148 47464 9204 47520
rect 9204 47464 9208 47520
rect 9144 47460 9208 47464
rect 6240 46188 6304 46192
rect 6240 46132 6244 46188
rect 6244 46132 6300 46188
rect 6300 46132 6304 46188
rect 6240 46128 6304 46132
rect 6320 46188 6384 46192
rect 6320 46132 6324 46188
rect 6324 46132 6380 46188
rect 6380 46132 6384 46188
rect 6320 46128 6384 46132
rect 6400 46188 6464 46192
rect 6400 46132 6404 46188
rect 6404 46132 6460 46188
rect 6460 46132 6464 46188
rect 6400 46128 6464 46132
rect 6480 46188 6544 46192
rect 6480 46132 6484 46188
rect 6484 46132 6540 46188
rect 6540 46132 6544 46188
rect 6480 46128 6544 46132
rect 3576 44856 3640 44860
rect 3576 44800 3580 44856
rect 3580 44800 3636 44856
rect 3636 44800 3640 44856
rect 3576 44796 3640 44800
rect 3656 44856 3720 44860
rect 3656 44800 3660 44856
rect 3660 44800 3716 44856
rect 3716 44800 3720 44856
rect 3656 44796 3720 44800
rect 3736 44856 3800 44860
rect 3736 44800 3740 44856
rect 3740 44800 3796 44856
rect 3796 44800 3800 44856
rect 3736 44796 3800 44800
rect 3816 44856 3880 44860
rect 3816 44800 3820 44856
rect 3820 44800 3876 44856
rect 3876 44800 3880 44856
rect 3816 44796 3880 44800
rect 8904 44856 8968 44860
rect 8904 44800 8908 44856
rect 8908 44800 8964 44856
rect 8964 44800 8968 44856
rect 8904 44796 8968 44800
rect 8984 44856 9048 44860
rect 8984 44800 8988 44856
rect 8988 44800 9044 44856
rect 9044 44800 9048 44856
rect 8984 44796 9048 44800
rect 9064 44856 9128 44860
rect 9064 44800 9068 44856
rect 9068 44800 9124 44856
rect 9124 44800 9128 44856
rect 9064 44796 9128 44800
rect 9144 44856 9208 44860
rect 9144 44800 9148 44856
rect 9148 44800 9204 44856
rect 9204 44800 9208 44856
rect 9144 44796 9208 44800
rect 6240 43524 6304 43528
rect 6240 43468 6244 43524
rect 6244 43468 6300 43524
rect 6300 43468 6304 43524
rect 6240 43464 6304 43468
rect 6320 43524 6384 43528
rect 6320 43468 6324 43524
rect 6324 43468 6380 43524
rect 6380 43468 6384 43524
rect 6320 43464 6384 43468
rect 6400 43524 6464 43528
rect 6400 43468 6404 43524
rect 6404 43468 6460 43524
rect 6460 43468 6464 43524
rect 6400 43464 6464 43468
rect 6480 43524 6544 43528
rect 6480 43468 6484 43524
rect 6484 43468 6540 43524
rect 6540 43468 6544 43524
rect 6480 43464 6544 43468
rect 3576 42192 3640 42196
rect 3576 42136 3580 42192
rect 3580 42136 3636 42192
rect 3636 42136 3640 42192
rect 3576 42132 3640 42136
rect 3656 42192 3720 42196
rect 3656 42136 3660 42192
rect 3660 42136 3716 42192
rect 3716 42136 3720 42192
rect 3656 42132 3720 42136
rect 3736 42192 3800 42196
rect 3736 42136 3740 42192
rect 3740 42136 3796 42192
rect 3796 42136 3800 42192
rect 3736 42132 3800 42136
rect 3816 42192 3880 42196
rect 3816 42136 3820 42192
rect 3820 42136 3876 42192
rect 3876 42136 3880 42192
rect 3816 42132 3880 42136
rect 8904 42192 8968 42196
rect 8904 42136 8908 42192
rect 8908 42136 8964 42192
rect 8964 42136 8968 42192
rect 8904 42132 8968 42136
rect 8984 42192 9048 42196
rect 8984 42136 8988 42192
rect 8988 42136 9044 42192
rect 9044 42136 9048 42192
rect 8984 42132 9048 42136
rect 9064 42192 9128 42196
rect 9064 42136 9068 42192
rect 9068 42136 9124 42192
rect 9124 42136 9128 42192
rect 9064 42132 9128 42136
rect 9144 42192 9208 42196
rect 9144 42136 9148 42192
rect 9148 42136 9204 42192
rect 9204 42136 9208 42192
rect 9144 42132 9208 42136
rect 6240 40860 6304 40864
rect 6240 40804 6244 40860
rect 6244 40804 6300 40860
rect 6300 40804 6304 40860
rect 6240 40800 6304 40804
rect 6320 40860 6384 40864
rect 6320 40804 6324 40860
rect 6324 40804 6380 40860
rect 6380 40804 6384 40860
rect 6320 40800 6384 40804
rect 6400 40860 6464 40864
rect 6400 40804 6404 40860
rect 6404 40804 6460 40860
rect 6460 40804 6464 40860
rect 6400 40800 6464 40804
rect 6480 40860 6544 40864
rect 6480 40804 6484 40860
rect 6484 40804 6540 40860
rect 6540 40804 6544 40860
rect 6480 40800 6544 40804
rect 3576 39528 3640 39532
rect 3576 39472 3580 39528
rect 3580 39472 3636 39528
rect 3636 39472 3640 39528
rect 3576 39468 3640 39472
rect 3656 39528 3720 39532
rect 3656 39472 3660 39528
rect 3660 39472 3716 39528
rect 3716 39472 3720 39528
rect 3656 39468 3720 39472
rect 3736 39528 3800 39532
rect 3736 39472 3740 39528
rect 3740 39472 3796 39528
rect 3796 39472 3800 39528
rect 3736 39468 3800 39472
rect 3816 39528 3880 39532
rect 3816 39472 3820 39528
rect 3820 39472 3876 39528
rect 3876 39472 3880 39528
rect 3816 39468 3880 39472
rect 8904 39528 8968 39532
rect 8904 39472 8908 39528
rect 8908 39472 8964 39528
rect 8964 39472 8968 39528
rect 8904 39468 8968 39472
rect 8984 39528 9048 39532
rect 8984 39472 8988 39528
rect 8988 39472 9044 39528
rect 9044 39472 9048 39528
rect 8984 39468 9048 39472
rect 9064 39528 9128 39532
rect 9064 39472 9068 39528
rect 9068 39472 9124 39528
rect 9124 39472 9128 39528
rect 9064 39468 9128 39472
rect 9144 39528 9208 39532
rect 9144 39472 9148 39528
rect 9148 39472 9204 39528
rect 9204 39472 9208 39528
rect 9144 39468 9208 39472
rect 6240 38196 6304 38200
rect 6240 38140 6244 38196
rect 6244 38140 6300 38196
rect 6300 38140 6304 38196
rect 6240 38136 6304 38140
rect 6320 38196 6384 38200
rect 6320 38140 6324 38196
rect 6324 38140 6380 38196
rect 6380 38140 6384 38196
rect 6320 38136 6384 38140
rect 6400 38196 6464 38200
rect 6400 38140 6404 38196
rect 6404 38140 6460 38196
rect 6460 38140 6464 38196
rect 6400 38136 6464 38140
rect 6480 38196 6544 38200
rect 6480 38140 6484 38196
rect 6484 38140 6540 38196
rect 6540 38140 6544 38196
rect 6480 38136 6544 38140
rect 3576 36864 3640 36868
rect 3576 36808 3580 36864
rect 3580 36808 3636 36864
rect 3636 36808 3640 36864
rect 3576 36804 3640 36808
rect 3656 36864 3720 36868
rect 3656 36808 3660 36864
rect 3660 36808 3716 36864
rect 3716 36808 3720 36864
rect 3656 36804 3720 36808
rect 3736 36864 3800 36868
rect 3736 36808 3740 36864
rect 3740 36808 3796 36864
rect 3796 36808 3800 36864
rect 3736 36804 3800 36808
rect 3816 36864 3880 36868
rect 3816 36808 3820 36864
rect 3820 36808 3876 36864
rect 3876 36808 3880 36864
rect 3816 36804 3880 36808
rect 8904 36864 8968 36868
rect 8904 36808 8908 36864
rect 8908 36808 8964 36864
rect 8964 36808 8968 36864
rect 8904 36804 8968 36808
rect 8984 36864 9048 36868
rect 8984 36808 8988 36864
rect 8988 36808 9044 36864
rect 9044 36808 9048 36864
rect 8984 36804 9048 36808
rect 9064 36864 9128 36868
rect 9064 36808 9068 36864
rect 9068 36808 9124 36864
rect 9124 36808 9128 36864
rect 9064 36804 9128 36808
rect 9144 36864 9208 36868
rect 9144 36808 9148 36864
rect 9148 36808 9204 36864
rect 9204 36808 9208 36864
rect 9144 36804 9208 36808
rect 6240 35532 6304 35536
rect 6240 35476 6244 35532
rect 6244 35476 6300 35532
rect 6300 35476 6304 35532
rect 6240 35472 6304 35476
rect 6320 35532 6384 35536
rect 6320 35476 6324 35532
rect 6324 35476 6380 35532
rect 6380 35476 6384 35532
rect 6320 35472 6384 35476
rect 6400 35532 6464 35536
rect 6400 35476 6404 35532
rect 6404 35476 6460 35532
rect 6460 35476 6464 35532
rect 6400 35472 6464 35476
rect 6480 35532 6544 35536
rect 6480 35476 6484 35532
rect 6484 35476 6540 35532
rect 6540 35476 6544 35532
rect 6480 35472 6544 35476
rect 3576 34200 3640 34204
rect 3576 34144 3580 34200
rect 3580 34144 3636 34200
rect 3636 34144 3640 34200
rect 3576 34140 3640 34144
rect 3656 34200 3720 34204
rect 3656 34144 3660 34200
rect 3660 34144 3716 34200
rect 3716 34144 3720 34200
rect 3656 34140 3720 34144
rect 3736 34200 3800 34204
rect 3736 34144 3740 34200
rect 3740 34144 3796 34200
rect 3796 34144 3800 34200
rect 3736 34140 3800 34144
rect 3816 34200 3880 34204
rect 3816 34144 3820 34200
rect 3820 34144 3876 34200
rect 3876 34144 3880 34200
rect 3816 34140 3880 34144
rect 8904 34200 8968 34204
rect 8904 34144 8908 34200
rect 8908 34144 8964 34200
rect 8964 34144 8968 34200
rect 8904 34140 8968 34144
rect 8984 34200 9048 34204
rect 8984 34144 8988 34200
rect 8988 34144 9044 34200
rect 9044 34144 9048 34200
rect 8984 34140 9048 34144
rect 9064 34200 9128 34204
rect 9064 34144 9068 34200
rect 9068 34144 9124 34200
rect 9124 34144 9128 34200
rect 9064 34140 9128 34144
rect 9144 34200 9208 34204
rect 9144 34144 9148 34200
rect 9148 34144 9204 34200
rect 9204 34144 9208 34200
rect 9144 34140 9208 34144
rect 6240 32868 6304 32872
rect 6240 32812 6244 32868
rect 6244 32812 6300 32868
rect 6300 32812 6304 32868
rect 6240 32808 6304 32812
rect 6320 32868 6384 32872
rect 6320 32812 6324 32868
rect 6324 32812 6380 32868
rect 6380 32812 6384 32868
rect 6320 32808 6384 32812
rect 6400 32868 6464 32872
rect 6400 32812 6404 32868
rect 6404 32812 6460 32868
rect 6460 32812 6464 32868
rect 6400 32808 6464 32812
rect 6480 32868 6544 32872
rect 6480 32812 6484 32868
rect 6484 32812 6540 32868
rect 6540 32812 6544 32868
rect 6480 32808 6544 32812
rect 3576 31536 3640 31540
rect 3576 31480 3580 31536
rect 3580 31480 3636 31536
rect 3636 31480 3640 31536
rect 3576 31476 3640 31480
rect 3656 31536 3720 31540
rect 3656 31480 3660 31536
rect 3660 31480 3716 31536
rect 3716 31480 3720 31536
rect 3656 31476 3720 31480
rect 3736 31536 3800 31540
rect 3736 31480 3740 31536
rect 3740 31480 3796 31536
rect 3796 31480 3800 31536
rect 3736 31476 3800 31480
rect 3816 31536 3880 31540
rect 3816 31480 3820 31536
rect 3820 31480 3876 31536
rect 3876 31480 3880 31536
rect 3816 31476 3880 31480
rect 8904 31536 8968 31540
rect 8904 31480 8908 31536
rect 8908 31480 8964 31536
rect 8964 31480 8968 31536
rect 8904 31476 8968 31480
rect 8984 31536 9048 31540
rect 8984 31480 8988 31536
rect 8988 31480 9044 31536
rect 9044 31480 9048 31536
rect 8984 31476 9048 31480
rect 9064 31536 9128 31540
rect 9064 31480 9068 31536
rect 9068 31480 9124 31536
rect 9124 31480 9128 31536
rect 9064 31476 9128 31480
rect 9144 31536 9208 31540
rect 9144 31480 9148 31536
rect 9148 31480 9204 31536
rect 9204 31480 9208 31536
rect 9144 31476 9208 31480
rect 6240 30204 6304 30208
rect 6240 30148 6244 30204
rect 6244 30148 6300 30204
rect 6300 30148 6304 30204
rect 6240 30144 6304 30148
rect 6320 30204 6384 30208
rect 6320 30148 6324 30204
rect 6324 30148 6380 30204
rect 6380 30148 6384 30204
rect 6320 30144 6384 30148
rect 6400 30204 6464 30208
rect 6400 30148 6404 30204
rect 6404 30148 6460 30204
rect 6460 30148 6464 30204
rect 6400 30144 6464 30148
rect 6480 30204 6544 30208
rect 6480 30148 6484 30204
rect 6484 30148 6540 30204
rect 6540 30148 6544 30204
rect 6480 30144 6544 30148
rect 3576 28872 3640 28876
rect 3576 28816 3580 28872
rect 3580 28816 3636 28872
rect 3636 28816 3640 28872
rect 3576 28812 3640 28816
rect 3656 28872 3720 28876
rect 3656 28816 3660 28872
rect 3660 28816 3716 28872
rect 3716 28816 3720 28872
rect 3656 28812 3720 28816
rect 3736 28872 3800 28876
rect 3736 28816 3740 28872
rect 3740 28816 3796 28872
rect 3796 28816 3800 28872
rect 3736 28812 3800 28816
rect 3816 28872 3880 28876
rect 3816 28816 3820 28872
rect 3820 28816 3876 28872
rect 3876 28816 3880 28872
rect 3816 28812 3880 28816
rect 8904 28872 8968 28876
rect 8904 28816 8908 28872
rect 8908 28816 8964 28872
rect 8964 28816 8968 28872
rect 8904 28812 8968 28816
rect 8984 28872 9048 28876
rect 8984 28816 8988 28872
rect 8988 28816 9044 28872
rect 9044 28816 9048 28872
rect 8984 28812 9048 28816
rect 9064 28872 9128 28876
rect 9064 28816 9068 28872
rect 9068 28816 9124 28872
rect 9124 28816 9128 28872
rect 9064 28812 9128 28816
rect 9144 28872 9208 28876
rect 9144 28816 9148 28872
rect 9148 28816 9204 28872
rect 9204 28816 9208 28872
rect 9144 28812 9208 28816
rect 6240 27540 6304 27544
rect 6240 27484 6244 27540
rect 6244 27484 6300 27540
rect 6300 27484 6304 27540
rect 6240 27480 6304 27484
rect 6320 27540 6384 27544
rect 6320 27484 6324 27540
rect 6324 27484 6380 27540
rect 6380 27484 6384 27540
rect 6320 27480 6384 27484
rect 6400 27540 6464 27544
rect 6400 27484 6404 27540
rect 6404 27484 6460 27540
rect 6460 27484 6464 27540
rect 6400 27480 6464 27484
rect 6480 27540 6544 27544
rect 6480 27484 6484 27540
rect 6484 27484 6540 27540
rect 6540 27484 6544 27540
rect 6480 27480 6544 27484
rect 3576 26208 3640 26212
rect 3576 26152 3580 26208
rect 3580 26152 3636 26208
rect 3636 26152 3640 26208
rect 3576 26148 3640 26152
rect 3656 26208 3720 26212
rect 3656 26152 3660 26208
rect 3660 26152 3716 26208
rect 3716 26152 3720 26208
rect 3656 26148 3720 26152
rect 3736 26208 3800 26212
rect 3736 26152 3740 26208
rect 3740 26152 3796 26208
rect 3796 26152 3800 26208
rect 3736 26148 3800 26152
rect 3816 26208 3880 26212
rect 3816 26152 3820 26208
rect 3820 26152 3876 26208
rect 3876 26152 3880 26208
rect 3816 26148 3880 26152
rect 8904 26208 8968 26212
rect 8904 26152 8908 26208
rect 8908 26152 8964 26208
rect 8964 26152 8968 26208
rect 8904 26148 8968 26152
rect 8984 26208 9048 26212
rect 8984 26152 8988 26208
rect 8988 26152 9044 26208
rect 9044 26152 9048 26208
rect 8984 26148 9048 26152
rect 9064 26208 9128 26212
rect 9064 26152 9068 26208
rect 9068 26152 9124 26208
rect 9124 26152 9128 26208
rect 9064 26148 9128 26152
rect 9144 26208 9208 26212
rect 9144 26152 9148 26208
rect 9148 26152 9204 26208
rect 9204 26152 9208 26208
rect 9144 26148 9208 26152
rect 6240 24876 6304 24880
rect 6240 24820 6244 24876
rect 6244 24820 6300 24876
rect 6300 24820 6304 24876
rect 6240 24816 6304 24820
rect 6320 24876 6384 24880
rect 6320 24820 6324 24876
rect 6324 24820 6380 24876
rect 6380 24820 6384 24876
rect 6320 24816 6384 24820
rect 6400 24876 6464 24880
rect 6400 24820 6404 24876
rect 6404 24820 6460 24876
rect 6460 24820 6464 24876
rect 6400 24816 6464 24820
rect 6480 24876 6544 24880
rect 6480 24820 6484 24876
rect 6484 24820 6540 24876
rect 6540 24820 6544 24876
rect 6480 24816 6544 24820
rect 3576 23544 3640 23548
rect 3576 23488 3580 23544
rect 3580 23488 3636 23544
rect 3636 23488 3640 23544
rect 3576 23484 3640 23488
rect 3656 23544 3720 23548
rect 3656 23488 3660 23544
rect 3660 23488 3716 23544
rect 3716 23488 3720 23544
rect 3656 23484 3720 23488
rect 3736 23544 3800 23548
rect 3736 23488 3740 23544
rect 3740 23488 3796 23544
rect 3796 23488 3800 23544
rect 3736 23484 3800 23488
rect 3816 23544 3880 23548
rect 3816 23488 3820 23544
rect 3820 23488 3876 23544
rect 3876 23488 3880 23544
rect 3816 23484 3880 23488
rect 8904 23544 8968 23548
rect 8904 23488 8908 23544
rect 8908 23488 8964 23544
rect 8964 23488 8968 23544
rect 8904 23484 8968 23488
rect 8984 23544 9048 23548
rect 8984 23488 8988 23544
rect 8988 23488 9044 23544
rect 9044 23488 9048 23544
rect 8984 23484 9048 23488
rect 9064 23544 9128 23548
rect 9064 23488 9068 23544
rect 9068 23488 9124 23544
rect 9124 23488 9128 23544
rect 9064 23484 9128 23488
rect 9144 23544 9208 23548
rect 9144 23488 9148 23544
rect 9148 23488 9204 23544
rect 9204 23488 9208 23544
rect 9144 23484 9208 23488
rect 6240 22212 6304 22216
rect 6240 22156 6244 22212
rect 6244 22156 6300 22212
rect 6300 22156 6304 22212
rect 6240 22152 6304 22156
rect 6320 22212 6384 22216
rect 6320 22156 6324 22212
rect 6324 22156 6380 22212
rect 6380 22156 6384 22212
rect 6320 22152 6384 22156
rect 6400 22212 6464 22216
rect 6400 22156 6404 22212
rect 6404 22156 6460 22212
rect 6460 22156 6464 22212
rect 6400 22152 6464 22156
rect 6480 22212 6544 22216
rect 6480 22156 6484 22212
rect 6484 22156 6540 22212
rect 6540 22156 6544 22212
rect 6480 22152 6544 22156
rect 3576 20880 3640 20884
rect 3576 20824 3580 20880
rect 3580 20824 3636 20880
rect 3636 20824 3640 20880
rect 3576 20820 3640 20824
rect 3656 20880 3720 20884
rect 3656 20824 3660 20880
rect 3660 20824 3716 20880
rect 3716 20824 3720 20880
rect 3656 20820 3720 20824
rect 3736 20880 3800 20884
rect 3736 20824 3740 20880
rect 3740 20824 3796 20880
rect 3796 20824 3800 20880
rect 3736 20820 3800 20824
rect 3816 20880 3880 20884
rect 3816 20824 3820 20880
rect 3820 20824 3876 20880
rect 3876 20824 3880 20880
rect 3816 20820 3880 20824
rect 8904 20880 8968 20884
rect 8904 20824 8908 20880
rect 8908 20824 8964 20880
rect 8964 20824 8968 20880
rect 8904 20820 8968 20824
rect 8984 20880 9048 20884
rect 8984 20824 8988 20880
rect 8988 20824 9044 20880
rect 9044 20824 9048 20880
rect 8984 20820 9048 20824
rect 9064 20880 9128 20884
rect 9064 20824 9068 20880
rect 9068 20824 9124 20880
rect 9124 20824 9128 20880
rect 9064 20820 9128 20824
rect 9144 20880 9208 20884
rect 9144 20824 9148 20880
rect 9148 20824 9204 20880
rect 9204 20824 9208 20880
rect 9144 20820 9208 20824
rect 6240 19548 6304 19552
rect 6240 19492 6244 19548
rect 6244 19492 6300 19548
rect 6300 19492 6304 19548
rect 6240 19488 6304 19492
rect 6320 19548 6384 19552
rect 6320 19492 6324 19548
rect 6324 19492 6380 19548
rect 6380 19492 6384 19548
rect 6320 19488 6384 19492
rect 6400 19548 6464 19552
rect 6400 19492 6404 19548
rect 6404 19492 6460 19548
rect 6460 19492 6464 19548
rect 6400 19488 6464 19492
rect 6480 19548 6544 19552
rect 6480 19492 6484 19548
rect 6484 19492 6540 19548
rect 6540 19492 6544 19548
rect 6480 19488 6544 19492
rect 3576 18216 3640 18220
rect 3576 18160 3580 18216
rect 3580 18160 3636 18216
rect 3636 18160 3640 18216
rect 3576 18156 3640 18160
rect 3656 18216 3720 18220
rect 3656 18160 3660 18216
rect 3660 18160 3716 18216
rect 3716 18160 3720 18216
rect 3656 18156 3720 18160
rect 3736 18216 3800 18220
rect 3736 18160 3740 18216
rect 3740 18160 3796 18216
rect 3796 18160 3800 18216
rect 3736 18156 3800 18160
rect 3816 18216 3880 18220
rect 3816 18160 3820 18216
rect 3820 18160 3876 18216
rect 3876 18160 3880 18216
rect 3816 18156 3880 18160
rect 8904 18216 8968 18220
rect 8904 18160 8908 18216
rect 8908 18160 8964 18216
rect 8964 18160 8968 18216
rect 8904 18156 8968 18160
rect 8984 18216 9048 18220
rect 8984 18160 8988 18216
rect 8988 18160 9044 18216
rect 9044 18160 9048 18216
rect 8984 18156 9048 18160
rect 9064 18216 9128 18220
rect 9064 18160 9068 18216
rect 9068 18160 9124 18216
rect 9124 18160 9128 18216
rect 9064 18156 9128 18160
rect 9144 18216 9208 18220
rect 9144 18160 9148 18216
rect 9148 18160 9204 18216
rect 9204 18160 9208 18216
rect 9144 18156 9208 18160
rect 6240 16884 6304 16888
rect 6240 16828 6244 16884
rect 6244 16828 6300 16884
rect 6300 16828 6304 16884
rect 6240 16824 6304 16828
rect 6320 16884 6384 16888
rect 6320 16828 6324 16884
rect 6324 16828 6380 16884
rect 6380 16828 6384 16884
rect 6320 16824 6384 16828
rect 6400 16884 6464 16888
rect 6400 16828 6404 16884
rect 6404 16828 6460 16884
rect 6460 16828 6464 16884
rect 6400 16824 6464 16828
rect 6480 16884 6544 16888
rect 6480 16828 6484 16884
rect 6484 16828 6540 16884
rect 6540 16828 6544 16884
rect 6480 16824 6544 16828
rect 3576 15552 3640 15556
rect 3576 15496 3580 15552
rect 3580 15496 3636 15552
rect 3636 15496 3640 15552
rect 3576 15492 3640 15496
rect 3656 15552 3720 15556
rect 3656 15496 3660 15552
rect 3660 15496 3716 15552
rect 3716 15496 3720 15552
rect 3656 15492 3720 15496
rect 3736 15552 3800 15556
rect 3736 15496 3740 15552
rect 3740 15496 3796 15552
rect 3796 15496 3800 15552
rect 3736 15492 3800 15496
rect 3816 15552 3880 15556
rect 3816 15496 3820 15552
rect 3820 15496 3876 15552
rect 3876 15496 3880 15552
rect 3816 15492 3880 15496
rect 8904 15552 8968 15556
rect 8904 15496 8908 15552
rect 8908 15496 8964 15552
rect 8964 15496 8968 15552
rect 8904 15492 8968 15496
rect 8984 15552 9048 15556
rect 8984 15496 8988 15552
rect 8988 15496 9044 15552
rect 9044 15496 9048 15552
rect 8984 15492 9048 15496
rect 9064 15552 9128 15556
rect 9064 15496 9068 15552
rect 9068 15496 9124 15552
rect 9124 15496 9128 15552
rect 9064 15492 9128 15496
rect 9144 15552 9208 15556
rect 9144 15496 9148 15552
rect 9148 15496 9204 15552
rect 9204 15496 9208 15552
rect 9144 15492 9208 15496
rect 6240 14220 6304 14224
rect 6240 14164 6244 14220
rect 6244 14164 6300 14220
rect 6300 14164 6304 14220
rect 6240 14160 6304 14164
rect 6320 14220 6384 14224
rect 6320 14164 6324 14220
rect 6324 14164 6380 14220
rect 6380 14164 6384 14220
rect 6320 14160 6384 14164
rect 6400 14220 6464 14224
rect 6400 14164 6404 14220
rect 6404 14164 6460 14220
rect 6460 14164 6464 14220
rect 6400 14160 6464 14164
rect 6480 14220 6544 14224
rect 6480 14164 6484 14220
rect 6484 14164 6540 14220
rect 6540 14164 6544 14220
rect 6480 14160 6544 14164
rect 3576 12888 3640 12892
rect 3576 12832 3580 12888
rect 3580 12832 3636 12888
rect 3636 12832 3640 12888
rect 3576 12828 3640 12832
rect 3656 12888 3720 12892
rect 3656 12832 3660 12888
rect 3660 12832 3716 12888
rect 3716 12832 3720 12888
rect 3656 12828 3720 12832
rect 3736 12888 3800 12892
rect 3736 12832 3740 12888
rect 3740 12832 3796 12888
rect 3796 12832 3800 12888
rect 3736 12828 3800 12832
rect 3816 12888 3880 12892
rect 3816 12832 3820 12888
rect 3820 12832 3876 12888
rect 3876 12832 3880 12888
rect 3816 12828 3880 12832
rect 8904 12888 8968 12892
rect 8904 12832 8908 12888
rect 8908 12832 8964 12888
rect 8964 12832 8968 12888
rect 8904 12828 8968 12832
rect 8984 12888 9048 12892
rect 8984 12832 8988 12888
rect 8988 12832 9044 12888
rect 9044 12832 9048 12888
rect 8984 12828 9048 12832
rect 9064 12888 9128 12892
rect 9064 12832 9068 12888
rect 9068 12832 9124 12888
rect 9124 12832 9128 12888
rect 9064 12828 9128 12832
rect 9144 12888 9208 12892
rect 9144 12832 9148 12888
rect 9148 12832 9204 12888
rect 9204 12832 9208 12888
rect 9144 12828 9208 12832
rect 6240 11556 6304 11560
rect 6240 11500 6244 11556
rect 6244 11500 6300 11556
rect 6300 11500 6304 11556
rect 6240 11496 6304 11500
rect 6320 11556 6384 11560
rect 6320 11500 6324 11556
rect 6324 11500 6380 11556
rect 6380 11500 6384 11556
rect 6320 11496 6384 11500
rect 6400 11556 6464 11560
rect 6400 11500 6404 11556
rect 6404 11500 6460 11556
rect 6460 11500 6464 11556
rect 6400 11496 6464 11500
rect 6480 11556 6544 11560
rect 6480 11500 6484 11556
rect 6484 11500 6540 11556
rect 6540 11500 6544 11556
rect 6480 11496 6544 11500
rect 3576 10224 3640 10228
rect 3576 10168 3580 10224
rect 3580 10168 3636 10224
rect 3636 10168 3640 10224
rect 3576 10164 3640 10168
rect 3656 10224 3720 10228
rect 3656 10168 3660 10224
rect 3660 10168 3716 10224
rect 3716 10168 3720 10224
rect 3656 10164 3720 10168
rect 3736 10224 3800 10228
rect 3736 10168 3740 10224
rect 3740 10168 3796 10224
rect 3796 10168 3800 10224
rect 3736 10164 3800 10168
rect 3816 10224 3880 10228
rect 3816 10168 3820 10224
rect 3820 10168 3876 10224
rect 3876 10168 3880 10224
rect 3816 10164 3880 10168
rect 8904 10224 8968 10228
rect 8904 10168 8908 10224
rect 8908 10168 8964 10224
rect 8964 10168 8968 10224
rect 8904 10164 8968 10168
rect 8984 10224 9048 10228
rect 8984 10168 8988 10224
rect 8988 10168 9044 10224
rect 9044 10168 9048 10224
rect 8984 10164 9048 10168
rect 9064 10224 9128 10228
rect 9064 10168 9068 10224
rect 9068 10168 9124 10224
rect 9124 10168 9128 10224
rect 9064 10164 9128 10168
rect 9144 10224 9208 10228
rect 9144 10168 9148 10224
rect 9148 10168 9204 10224
rect 9204 10168 9208 10224
rect 9144 10164 9208 10168
rect 6240 8892 6304 8896
rect 6240 8836 6244 8892
rect 6244 8836 6300 8892
rect 6300 8836 6304 8892
rect 6240 8832 6304 8836
rect 6320 8892 6384 8896
rect 6320 8836 6324 8892
rect 6324 8836 6380 8892
rect 6380 8836 6384 8892
rect 6320 8832 6384 8836
rect 6400 8892 6464 8896
rect 6400 8836 6404 8892
rect 6404 8836 6460 8892
rect 6460 8836 6464 8892
rect 6400 8832 6464 8836
rect 6480 8892 6544 8896
rect 6480 8836 6484 8892
rect 6484 8836 6540 8892
rect 6540 8836 6544 8892
rect 6480 8832 6544 8836
rect 3576 7560 3640 7564
rect 3576 7504 3580 7560
rect 3580 7504 3636 7560
rect 3636 7504 3640 7560
rect 3576 7500 3640 7504
rect 3656 7560 3720 7564
rect 3656 7504 3660 7560
rect 3660 7504 3716 7560
rect 3716 7504 3720 7560
rect 3656 7500 3720 7504
rect 3736 7560 3800 7564
rect 3736 7504 3740 7560
rect 3740 7504 3796 7560
rect 3796 7504 3800 7560
rect 3736 7500 3800 7504
rect 3816 7560 3880 7564
rect 3816 7504 3820 7560
rect 3820 7504 3876 7560
rect 3876 7504 3880 7560
rect 3816 7500 3880 7504
rect 8904 7560 8968 7564
rect 8904 7504 8908 7560
rect 8908 7504 8964 7560
rect 8964 7504 8968 7560
rect 8904 7500 8968 7504
rect 8984 7560 9048 7564
rect 8984 7504 8988 7560
rect 8988 7504 9044 7560
rect 9044 7504 9048 7560
rect 8984 7500 9048 7504
rect 9064 7560 9128 7564
rect 9064 7504 9068 7560
rect 9068 7504 9124 7560
rect 9124 7504 9128 7560
rect 9064 7500 9128 7504
rect 9144 7560 9208 7564
rect 9144 7504 9148 7560
rect 9148 7504 9204 7560
rect 9204 7504 9208 7560
rect 9144 7500 9208 7504
rect 6240 6228 6304 6232
rect 6240 6172 6244 6228
rect 6244 6172 6300 6228
rect 6300 6172 6304 6228
rect 6240 6168 6304 6172
rect 6320 6228 6384 6232
rect 6320 6172 6324 6228
rect 6324 6172 6380 6228
rect 6380 6172 6384 6228
rect 6320 6168 6384 6172
rect 6400 6228 6464 6232
rect 6400 6172 6404 6228
rect 6404 6172 6460 6228
rect 6460 6172 6464 6228
rect 6400 6168 6464 6172
rect 6480 6228 6544 6232
rect 6480 6172 6484 6228
rect 6484 6172 6540 6228
rect 6540 6172 6544 6228
rect 6480 6168 6544 6172
rect 3576 4896 3640 4900
rect 3576 4840 3580 4896
rect 3580 4840 3636 4896
rect 3636 4840 3640 4896
rect 3576 4836 3640 4840
rect 3656 4896 3720 4900
rect 3656 4840 3660 4896
rect 3660 4840 3716 4896
rect 3716 4840 3720 4896
rect 3656 4836 3720 4840
rect 3736 4896 3800 4900
rect 3736 4840 3740 4896
rect 3740 4840 3796 4896
rect 3796 4840 3800 4896
rect 3736 4836 3800 4840
rect 3816 4896 3880 4900
rect 3816 4840 3820 4896
rect 3820 4840 3876 4896
rect 3876 4840 3880 4896
rect 3816 4836 3880 4840
rect 8904 4896 8968 4900
rect 8904 4840 8908 4896
rect 8908 4840 8964 4896
rect 8964 4840 8968 4896
rect 8904 4836 8968 4840
rect 8984 4896 9048 4900
rect 8984 4840 8988 4896
rect 8988 4840 9044 4896
rect 9044 4840 9048 4896
rect 8984 4836 9048 4840
rect 9064 4896 9128 4900
rect 9064 4840 9068 4896
rect 9068 4840 9124 4896
rect 9124 4840 9128 4896
rect 9064 4836 9128 4840
rect 9144 4896 9208 4900
rect 9144 4840 9148 4896
rect 9148 4840 9204 4896
rect 9204 4840 9208 4896
rect 9144 4836 9208 4840
rect 6240 3564 6304 3568
rect 6240 3508 6244 3564
rect 6244 3508 6300 3564
rect 6300 3508 6304 3564
rect 6240 3504 6304 3508
rect 6320 3564 6384 3568
rect 6320 3508 6324 3564
rect 6324 3508 6380 3564
rect 6380 3508 6384 3564
rect 6320 3504 6384 3508
rect 6400 3564 6464 3568
rect 6400 3508 6404 3564
rect 6404 3508 6460 3564
rect 6460 3508 6464 3564
rect 6400 3504 6464 3508
rect 6480 3564 6544 3568
rect 6480 3508 6484 3564
rect 6484 3508 6540 3564
rect 6540 3508 6544 3564
rect 6480 3504 6544 3508
rect 3576 2232 3640 2236
rect 3576 2176 3580 2232
rect 3580 2176 3636 2232
rect 3636 2176 3640 2232
rect 3576 2172 3640 2176
rect 3656 2232 3720 2236
rect 3656 2176 3660 2232
rect 3660 2176 3716 2232
rect 3716 2176 3720 2232
rect 3656 2172 3720 2176
rect 3736 2232 3800 2236
rect 3736 2176 3740 2232
rect 3740 2176 3796 2232
rect 3796 2176 3800 2232
rect 3736 2172 3800 2176
rect 3816 2232 3880 2236
rect 3816 2176 3820 2232
rect 3820 2176 3876 2232
rect 3876 2176 3880 2232
rect 3816 2172 3880 2176
rect 8904 2232 8968 2236
rect 8904 2176 8908 2232
rect 8908 2176 8964 2232
rect 8964 2176 8968 2232
rect 8904 2172 8968 2176
rect 8984 2232 9048 2236
rect 8984 2176 8988 2232
rect 8988 2176 9044 2232
rect 9044 2176 9048 2232
rect 8984 2172 9048 2176
rect 9064 2232 9128 2236
rect 9064 2176 9068 2232
rect 9068 2176 9124 2232
rect 9124 2176 9128 2232
rect 9064 2172 9128 2176
rect 9144 2232 9208 2236
rect 9144 2176 9148 2232
rect 9148 2176 9204 2232
rect 9204 2176 9208 2232
rect 9144 2172 9208 2176
rect 6240 900 6304 904
rect 6240 844 6244 900
rect 6244 844 6300 900
rect 6300 844 6304 900
rect 6240 840 6304 844
rect 6320 900 6384 904
rect 6320 844 6324 900
rect 6324 844 6380 900
rect 6380 844 6384 900
rect 6320 840 6384 844
rect 6400 900 6464 904
rect 6400 844 6404 900
rect 6404 844 6460 900
rect 6460 844 6464 900
rect 6400 840 6464 844
rect 6480 900 6544 904
rect 6480 844 6484 900
rect 6484 844 6540 900
rect 6540 844 6544 900
rect 6480 840 6544 844
<< metal4 >>
rect 3568 52852 3888 52868
rect 3568 52788 3576 52852
rect 3640 52788 3656 52852
rect 3720 52788 3736 52852
rect 3800 52788 3816 52852
rect 3880 52788 3888 52852
rect 3568 50188 3888 52788
rect 3568 50124 3576 50188
rect 3640 50124 3656 50188
rect 3720 50124 3736 50188
rect 3800 50124 3816 50188
rect 3880 50124 3888 50188
rect 3568 47524 3888 50124
rect 3568 47460 3576 47524
rect 3640 47460 3656 47524
rect 3720 47460 3736 47524
rect 3800 47460 3816 47524
rect 3880 47460 3888 47524
rect 3568 44860 3888 47460
rect 3568 44796 3576 44860
rect 3640 44796 3656 44860
rect 3720 44796 3736 44860
rect 3800 44796 3816 44860
rect 3880 44796 3888 44860
rect 3568 42196 3888 44796
rect 3568 42132 3576 42196
rect 3640 42132 3656 42196
rect 3720 42132 3736 42196
rect 3800 42132 3816 42196
rect 3880 42132 3888 42196
rect 3568 39532 3888 42132
rect 3568 39468 3576 39532
rect 3640 39468 3656 39532
rect 3720 39468 3736 39532
rect 3800 39468 3816 39532
rect 3880 39468 3888 39532
rect 3568 36868 3888 39468
rect 3568 36804 3576 36868
rect 3640 36804 3656 36868
rect 3720 36804 3736 36868
rect 3800 36804 3816 36868
rect 3880 36804 3888 36868
rect 3568 34204 3888 36804
rect 3568 34140 3576 34204
rect 3640 34140 3656 34204
rect 3720 34140 3736 34204
rect 3800 34140 3816 34204
rect 3880 34140 3888 34204
rect 3568 31540 3888 34140
rect 3568 31476 3576 31540
rect 3640 31476 3656 31540
rect 3720 31476 3736 31540
rect 3800 31476 3816 31540
rect 3880 31476 3888 31540
rect 3568 28876 3888 31476
rect 3568 28812 3576 28876
rect 3640 28812 3656 28876
rect 3720 28812 3736 28876
rect 3800 28812 3816 28876
rect 3880 28812 3888 28876
rect 3568 26212 3888 28812
rect 3568 26148 3576 26212
rect 3640 26148 3656 26212
rect 3720 26148 3736 26212
rect 3800 26148 3816 26212
rect 3880 26148 3888 26212
rect 3568 23548 3888 26148
rect 3568 23484 3576 23548
rect 3640 23484 3656 23548
rect 3720 23484 3736 23548
rect 3800 23484 3816 23548
rect 3880 23484 3888 23548
rect 3568 20884 3888 23484
rect 3568 20820 3576 20884
rect 3640 20820 3656 20884
rect 3720 20820 3736 20884
rect 3800 20820 3816 20884
rect 3880 20820 3888 20884
rect 3568 20782 3888 20820
rect 3568 20546 3610 20782
rect 3846 20546 3888 20782
rect 3568 18220 3888 20546
rect 3568 18156 3576 18220
rect 3640 18156 3656 18220
rect 3720 18156 3736 18220
rect 3800 18156 3816 18220
rect 3880 18156 3888 18220
rect 3568 15556 3888 18156
rect 3568 15492 3576 15556
rect 3640 15492 3656 15556
rect 3720 15492 3736 15556
rect 3800 15492 3816 15556
rect 3880 15492 3888 15556
rect 3568 12892 3888 15492
rect 3568 12828 3576 12892
rect 3640 12828 3656 12892
rect 3720 12828 3736 12892
rect 3800 12828 3816 12892
rect 3880 12828 3888 12892
rect 3568 10228 3888 12828
rect 3568 10164 3576 10228
rect 3640 10164 3656 10228
rect 3720 10164 3736 10228
rect 3800 10164 3816 10228
rect 3880 10164 3888 10228
rect 3568 7564 3888 10164
rect 3568 7500 3576 7564
rect 3640 7500 3656 7564
rect 3720 7500 3736 7564
rect 3800 7500 3816 7564
rect 3880 7500 3888 7564
rect 3568 4900 3888 7500
rect 3568 4836 3576 4900
rect 3640 4836 3656 4900
rect 3720 4836 3736 4900
rect 3800 4836 3816 4900
rect 3880 4836 3888 4900
rect 3568 2236 3888 4836
rect 3568 2172 3576 2236
rect 3640 2172 3656 2236
rect 3720 2172 3736 2236
rect 3800 2172 3816 2236
rect 3880 2172 3888 2236
rect 3568 824 3888 2172
rect 6232 51520 6552 52868
rect 6232 51456 6240 51520
rect 6304 51456 6320 51520
rect 6384 51456 6400 51520
rect 6464 51456 6480 51520
rect 6544 51456 6552 51520
rect 6232 48856 6552 51456
rect 6232 48792 6240 48856
rect 6304 48792 6320 48856
rect 6384 48792 6400 48856
rect 6464 48792 6480 48856
rect 6544 48792 6552 48856
rect 6232 46192 6552 48792
rect 6232 46128 6240 46192
rect 6304 46128 6320 46192
rect 6384 46128 6400 46192
rect 6464 46128 6480 46192
rect 6544 46128 6552 46192
rect 6232 43528 6552 46128
rect 6232 43464 6240 43528
rect 6304 43464 6320 43528
rect 6384 43464 6400 43528
rect 6464 43464 6480 43528
rect 6544 43464 6552 43528
rect 6232 40864 6552 43464
rect 6232 40800 6240 40864
rect 6304 40800 6320 40864
rect 6384 40800 6400 40864
rect 6464 40800 6480 40864
rect 6544 40800 6552 40864
rect 6232 38782 6552 40800
rect 6232 38546 6274 38782
rect 6510 38546 6552 38782
rect 6232 38200 6552 38546
rect 6232 38136 6240 38200
rect 6304 38136 6320 38200
rect 6384 38136 6400 38200
rect 6464 38136 6480 38200
rect 6544 38136 6552 38200
rect 6232 35536 6552 38136
rect 6232 35472 6240 35536
rect 6304 35472 6320 35536
rect 6384 35472 6400 35536
rect 6464 35472 6480 35536
rect 6544 35472 6552 35536
rect 6232 32872 6552 35472
rect 6232 32808 6240 32872
rect 6304 32808 6320 32872
rect 6384 32808 6400 32872
rect 6464 32808 6480 32872
rect 6544 32808 6552 32872
rect 6232 30208 6552 32808
rect 6232 30144 6240 30208
rect 6304 30144 6320 30208
rect 6384 30144 6400 30208
rect 6464 30144 6480 30208
rect 6544 30144 6552 30208
rect 6232 27544 6552 30144
rect 6232 27480 6240 27544
rect 6304 27480 6320 27544
rect 6384 27480 6400 27544
rect 6464 27480 6480 27544
rect 6544 27480 6552 27544
rect 6232 24880 6552 27480
rect 6232 24816 6240 24880
rect 6304 24816 6320 24880
rect 6384 24816 6400 24880
rect 6464 24816 6480 24880
rect 6544 24816 6552 24880
rect 6232 22216 6552 24816
rect 6232 22152 6240 22216
rect 6304 22152 6320 22216
rect 6384 22152 6400 22216
rect 6464 22152 6480 22216
rect 6544 22152 6552 22216
rect 6232 19552 6552 22152
rect 6232 19488 6240 19552
rect 6304 19488 6320 19552
rect 6384 19488 6400 19552
rect 6464 19488 6480 19552
rect 6544 19488 6552 19552
rect 6232 16888 6552 19488
rect 6232 16824 6240 16888
rect 6304 16824 6320 16888
rect 6384 16824 6400 16888
rect 6464 16824 6480 16888
rect 6544 16824 6552 16888
rect 6232 14224 6552 16824
rect 6232 14160 6240 14224
rect 6304 14160 6320 14224
rect 6384 14160 6400 14224
rect 6464 14160 6480 14224
rect 6544 14160 6552 14224
rect 6232 11560 6552 14160
rect 6232 11496 6240 11560
rect 6304 11496 6320 11560
rect 6384 11496 6400 11560
rect 6464 11496 6480 11560
rect 6544 11496 6552 11560
rect 6232 8896 6552 11496
rect 6232 8832 6240 8896
rect 6304 8832 6320 8896
rect 6384 8832 6400 8896
rect 6464 8832 6480 8896
rect 6544 8832 6552 8896
rect 6232 6232 6552 8832
rect 6232 6168 6240 6232
rect 6304 6168 6320 6232
rect 6384 6168 6400 6232
rect 6464 6168 6480 6232
rect 6544 6168 6552 6232
rect 6232 3568 6552 6168
rect 6232 3504 6240 3568
rect 6304 3504 6320 3568
rect 6384 3504 6400 3568
rect 6464 3504 6480 3568
rect 6544 3504 6552 3568
rect 6232 2782 6552 3504
rect 6232 2546 6274 2782
rect 6510 2546 6552 2782
rect 6232 904 6552 2546
rect 6232 840 6240 904
rect 6304 840 6320 904
rect 6384 840 6400 904
rect 6464 840 6480 904
rect 6544 840 6552 904
rect 6232 824 6552 840
rect 8896 52852 9216 52868
rect 8896 52788 8904 52852
rect 8968 52788 8984 52852
rect 9048 52788 9064 52852
rect 9128 52788 9144 52852
rect 9208 52788 9216 52852
rect 8896 50188 9216 52788
rect 8896 50124 8904 50188
rect 8968 50124 8984 50188
rect 9048 50124 9064 50188
rect 9128 50124 9144 50188
rect 9208 50124 9216 50188
rect 8896 47524 9216 50124
rect 8896 47460 8904 47524
rect 8968 47460 8984 47524
rect 9048 47460 9064 47524
rect 9128 47460 9144 47524
rect 9208 47460 9216 47524
rect 8896 44860 9216 47460
rect 8896 44796 8904 44860
rect 8968 44796 8984 44860
rect 9048 44796 9064 44860
rect 9128 44796 9144 44860
rect 9208 44796 9216 44860
rect 8896 42196 9216 44796
rect 8896 42132 8904 42196
rect 8968 42132 8984 42196
rect 9048 42132 9064 42196
rect 9128 42132 9144 42196
rect 9208 42132 9216 42196
rect 8896 39532 9216 42132
rect 8896 39468 8904 39532
rect 8968 39468 8984 39532
rect 9048 39468 9064 39532
rect 9128 39468 9144 39532
rect 9208 39468 9216 39532
rect 8896 36868 9216 39468
rect 8896 36804 8904 36868
rect 8968 36804 8984 36868
rect 9048 36804 9064 36868
rect 9128 36804 9144 36868
rect 9208 36804 9216 36868
rect 8896 34204 9216 36804
rect 8896 34140 8904 34204
rect 8968 34140 8984 34204
rect 9048 34140 9064 34204
rect 9128 34140 9144 34204
rect 9208 34140 9216 34204
rect 8896 31540 9216 34140
rect 8896 31476 8904 31540
rect 8968 31476 8984 31540
rect 9048 31476 9064 31540
rect 9128 31476 9144 31540
rect 9208 31476 9216 31540
rect 8896 28876 9216 31476
rect 8896 28812 8904 28876
rect 8968 28812 8984 28876
rect 9048 28812 9064 28876
rect 9128 28812 9144 28876
rect 9208 28812 9216 28876
rect 8896 26212 9216 28812
rect 8896 26148 8904 26212
rect 8968 26148 8984 26212
rect 9048 26148 9064 26212
rect 9128 26148 9144 26212
rect 9208 26148 9216 26212
rect 8896 23548 9216 26148
rect 8896 23484 8904 23548
rect 8968 23484 8984 23548
rect 9048 23484 9064 23548
rect 9128 23484 9144 23548
rect 9208 23484 9216 23548
rect 8896 20884 9216 23484
rect 8896 20820 8904 20884
rect 8968 20820 8984 20884
rect 9048 20820 9064 20884
rect 9128 20820 9144 20884
rect 9208 20820 9216 20884
rect 8896 20782 9216 20820
rect 8896 20546 8938 20782
rect 9174 20546 9216 20782
rect 8896 18220 9216 20546
rect 8896 18156 8904 18220
rect 8968 18156 8984 18220
rect 9048 18156 9064 18220
rect 9128 18156 9144 18220
rect 9208 18156 9216 18220
rect 8896 15556 9216 18156
rect 8896 15492 8904 15556
rect 8968 15492 8984 15556
rect 9048 15492 9064 15556
rect 9128 15492 9144 15556
rect 9208 15492 9216 15556
rect 8896 12892 9216 15492
rect 8896 12828 8904 12892
rect 8968 12828 8984 12892
rect 9048 12828 9064 12892
rect 9128 12828 9144 12892
rect 9208 12828 9216 12892
rect 8896 10228 9216 12828
rect 8896 10164 8904 10228
rect 8968 10164 8984 10228
rect 9048 10164 9064 10228
rect 9128 10164 9144 10228
rect 9208 10164 9216 10228
rect 8896 7564 9216 10164
rect 8896 7500 8904 7564
rect 8968 7500 8984 7564
rect 9048 7500 9064 7564
rect 9128 7500 9144 7564
rect 9208 7500 9216 7564
rect 8896 4900 9216 7500
rect 8896 4836 8904 4900
rect 8968 4836 8984 4900
rect 9048 4836 9064 4900
rect 9128 4836 9144 4900
rect 9208 4836 9216 4900
rect 8896 2236 9216 4836
rect 8896 2172 8904 2236
rect 8968 2172 8984 2236
rect 9048 2172 9064 2236
rect 9128 2172 9144 2236
rect 9208 2172 9216 2236
rect 8896 824 9216 2172
<< via4 >>
rect 3610 20546 3846 20782
rect 6274 38546 6510 38782
rect 6274 2546 6510 2782
rect 8938 20546 9174 20782
<< metal5 >>
rect 1064 38782 9556 38824
rect 1064 38546 6274 38782
rect 6510 38546 9556 38782
rect 1064 38504 9556 38546
rect 1064 20782 9556 20824
rect 1064 20546 3610 20782
rect 3846 20546 8938 20782
rect 9174 20546 9556 20782
rect 1064 20504 9556 20546
rect 1064 2782 9556 2824
rect 1064 2546 6274 2782
rect 6510 2546 9556 2782
rect 1064 2504 9556 2546
use sky130_osu_sc_18T_hs__decap_1  decap1_0 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 1614 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_5 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 1592 0 1 2204
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_4 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 1416 0 1 2204
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_3 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 1064 0 1 2204
box 0 0 352 1332
use sky130_osu_sc_18T_hs__decap_1  decap0_0
timestamp 1607194151
transform 1 0 1614 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_2
timestamp 1607194151
transform 1 0 1592 0 -1 2204
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_1
timestamp 1607194151
transform 1 0 1416 0 -1 2204
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_0
timestamp 1607194151
transform 1 0 1064 0 -1 2204
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_30 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 2296 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_1
timestamp 1607194151
transform 1 0 2098 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_31
timestamp 1607194151
transform 1 0 1812 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_1
timestamp 1607194151
transform 1 0 2296 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_1
timestamp 1607194151
transform 1 0 2098 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_0
timestamp 1607194151
transform 1 0 1812 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_3
timestamp 1607194151
transform 1 0 3066 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_29
timestamp 1607194151
transform 1 0 2780 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_2
timestamp 1607194151
transform 1 0 2582 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_3
timestamp 1607194151
transform 1 0 3066 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_2
timestamp 1607194151
transform 1 0 2780 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_2
timestamp 1607194151
transform 1 0 2582 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_27
timestamp 1607194151
transform 1 0 3748 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_4
timestamp 1607194151
transform 1 0 3550 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_28
timestamp 1607194151
transform 1 0 3264 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_4
timestamp 1607194151
transform 1 0 3748 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_4
timestamp 1607194151
transform 1 0 3550 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_3
timestamp 1607194151
transform 1 0 3264 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_6
timestamp 1607194151
transform 1 0 4518 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_26
timestamp 1607194151
transform 1 0 4232 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_5
timestamp 1607194151
transform 1 0 4034 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_6
timestamp 1607194151
transform 1 0 4518 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_5
timestamp 1607194151
transform 1 0 4232 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_5
timestamp 1607194151
transform 1 0 4034 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_24
timestamp 1607194151
transform 1 0 5200 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_7
timestamp 1607194151
transform 1 0 5002 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_25
timestamp 1607194151
transform 1 0 4716 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_7
timestamp 1607194151
transform 1 0 5200 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_7
timestamp 1607194151
transform 1 0 5002 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_6
timestamp 1607194151
transform 1 0 4716 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_9
timestamp 1607194151
transform 1 0 5970 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_23
timestamp 1607194151
transform 1 0 5684 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_8
timestamp 1607194151
transform 1 0 5486 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_9
timestamp 1607194151
transform 1 0 5970 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_8
timestamp 1607194151
transform 1 0 5684 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_8
timestamp 1607194151
transform 1 0 5486 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_21
timestamp 1607194151
transform 1 0 6652 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_10
timestamp 1607194151
transform 1 0 6454 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_22
timestamp 1607194151
transform 1 0 6168 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_10
timestamp 1607194151
transform 1 0 6652 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_10
timestamp 1607194151
transform 1 0 6454 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_9
timestamp 1607194151
transform 1 0 6168 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_20
timestamp 1607194151
transform 1 0 7136 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_11
timestamp 1607194151
transform 1 0 6938 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_11
timestamp 1607194151
transform 1 0 7136 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_11
timestamp 1607194151
transform 1 0 6938 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_18
timestamp 1607194151
transform 1 0 8104 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_13
timestamp 1607194151
transform 1 0 7906 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_19
timestamp 1607194151
transform 1 0 7620 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_12
timestamp 1607194151
transform 1 0 7422 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_13
timestamp 1607194151
transform 1 0 8104 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_13
timestamp 1607194151
transform 1 0 7906 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_12
timestamp 1607194151
transform 1 0 7620 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_12
timestamp 1607194151
transform 1 0 7422 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_17
timestamp 1607194151
transform 1 0 8588 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_14
timestamp 1607194151
transform 1 0 8390 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_14
timestamp 1607194151
transform 1 0 8588 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_14
timestamp 1607194151
transform 1 0 8390 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_16
timestamp 1607194151
transform 1 0 9358 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_16
timestamp 1607194151
transform 1 0 9072 0 1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap1_15
timestamp 1607194151
transform 1 0 8874 0 1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_16
timestamp 1607194151
transform 1 0 9358 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_15
timestamp 1607194151
transform 1 0 9072 0 -1 2204
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap0_15
timestamp 1607194151
transform 1 0 8874 0 -1 2204
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_0
timestamp 1607194151
transform 1 0 1614 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_8
timestamp 1607194151
transform 1 0 1592 0 -1 4868
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_7
timestamp 1607194151
transform 1 0 1416 0 -1 4868
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_6
timestamp 1607194151
transform 1 0 1064 0 -1 4868
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_33
timestamp 1607194151
transform 1 0 2296 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_1
timestamp 1607194151
transform 1 0 2098 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_32
timestamp 1607194151
transform 1 0 1812 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_3
timestamp 1607194151
transform 1 0 3066 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_34
timestamp 1607194151
transform 1 0 2780 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_2
timestamp 1607194151
transform 1 0 2582 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_36
timestamp 1607194151
transform 1 0 3748 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_4
timestamp 1607194151
transform 1 0 3550 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_35
timestamp 1607194151
transform 1 0 3264 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_6
timestamp 1607194151
transform 1 0 4518 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_37
timestamp 1607194151
transform 1 0 4232 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_5
timestamp 1607194151
transform 1 0 4034 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_39
timestamp 1607194151
transform 1 0 5200 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_7
timestamp 1607194151
transform 1 0 5002 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_38
timestamp 1607194151
transform 1 0 4716 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_9
timestamp 1607194151
transform 1 0 5970 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_40
timestamp 1607194151
transform 1 0 5684 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_8
timestamp 1607194151
transform 1 0 5486 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_42
timestamp 1607194151
transform 1 0 6652 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_10
timestamp 1607194151
transform 1 0 6454 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_41
timestamp 1607194151
transform 1 0 6168 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_43
timestamp 1607194151
transform 1 0 7136 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_11
timestamp 1607194151
transform 1 0 6938 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_45
timestamp 1607194151
transform 1 0 8104 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_13
timestamp 1607194151
transform 1 0 7906 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_44
timestamp 1607194151
transform 1 0 7620 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_12
timestamp 1607194151
transform 1 0 7422 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_46
timestamp 1607194151
transform 1 0 8588 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_14
timestamp 1607194151
transform 1 0 8390 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_16
timestamp 1607194151
transform 1 0 9358 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_47
timestamp 1607194151
transform 1 0 9072 0 -1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap2_15
timestamp 1607194151
transform 1 0 8874 0 -1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_0
timestamp 1607194151
transform 1 0 1614 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_11
timestamp 1607194151
transform 1 0 1592 0 1 4868
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_10
timestamp 1607194151
transform 1 0 1416 0 1 4868
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_9
timestamp 1607194151
transform 1 0 1064 0 1 4868
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_62
timestamp 1607194151
transform 1 0 2296 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_1
timestamp 1607194151
transform 1 0 2098 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_63
timestamp 1607194151
transform 1 0 1812 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_3
timestamp 1607194151
transform 1 0 3066 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_61
timestamp 1607194151
transform 1 0 2780 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_2
timestamp 1607194151
transform 1 0 2582 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_59
timestamp 1607194151
transform 1 0 3748 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_4
timestamp 1607194151
transform 1 0 3550 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_60
timestamp 1607194151
transform 1 0 3264 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_6
timestamp 1607194151
transform 1 0 4518 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_58
timestamp 1607194151
transform 1 0 4232 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_5
timestamp 1607194151
transform 1 0 4034 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_56
timestamp 1607194151
transform 1 0 5200 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_7
timestamp 1607194151
transform 1 0 5002 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_57
timestamp 1607194151
transform 1 0 4716 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_9
timestamp 1607194151
transform 1 0 5970 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_55
timestamp 1607194151
transform 1 0 5684 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_8
timestamp 1607194151
transform 1 0 5486 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_53
timestamp 1607194151
transform 1 0 6652 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_10
timestamp 1607194151
transform 1 0 6454 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_54
timestamp 1607194151
transform 1 0 6168 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_52
timestamp 1607194151
transform 1 0 7136 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_11
timestamp 1607194151
transform 1 0 6938 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_50
timestamp 1607194151
transform 1 0 8104 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_13
timestamp 1607194151
transform 1 0 7906 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_51
timestamp 1607194151
transform 1 0 7620 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_12
timestamp 1607194151
transform 1 0 7422 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_49
timestamp 1607194151
transform 1 0 8588 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_14
timestamp 1607194151
transform 1 0 8390 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_16
timestamp 1607194151
transform 1 0 9358 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_48
timestamp 1607194151
transform 1 0 9072 0 1 4868
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap3_15
timestamp 1607194151
transform 1 0 8874 0 1 4868
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_0
timestamp 1607194151
transform 1 0 1614 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_14
timestamp 1607194151
transform 1 0 1592 0 -1 7532
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_13
timestamp 1607194151
transform 1 0 1416 0 -1 7532
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_12
timestamp 1607194151
transform 1 0 1064 0 -1 7532
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_65
timestamp 1607194151
transform 1 0 2296 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_1
timestamp 1607194151
transform 1 0 2098 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_64
timestamp 1607194151
transform 1 0 1812 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_3
timestamp 1607194151
transform 1 0 3066 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_66
timestamp 1607194151
transform 1 0 2780 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_2
timestamp 1607194151
transform 1 0 2582 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_68
timestamp 1607194151
transform 1 0 3748 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_4
timestamp 1607194151
transform 1 0 3550 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_67
timestamp 1607194151
transform 1 0 3264 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_6
timestamp 1607194151
transform 1 0 4518 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_69
timestamp 1607194151
transform 1 0 4232 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_5
timestamp 1607194151
transform 1 0 4034 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_71
timestamp 1607194151
transform 1 0 5200 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_7
timestamp 1607194151
transform 1 0 5002 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_70
timestamp 1607194151
transform 1 0 4716 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_9
timestamp 1607194151
transform 1 0 5970 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_72
timestamp 1607194151
transform 1 0 5684 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_8
timestamp 1607194151
transform 1 0 5486 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_74
timestamp 1607194151
transform 1 0 6652 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_10
timestamp 1607194151
transform 1 0 6454 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_73
timestamp 1607194151
transform 1 0 6168 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_75
timestamp 1607194151
transform 1 0 7136 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_11
timestamp 1607194151
transform 1 0 6938 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_77
timestamp 1607194151
transform 1 0 8104 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_13
timestamp 1607194151
transform 1 0 7906 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_76
timestamp 1607194151
transform 1 0 7620 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_12
timestamp 1607194151
transform 1 0 7422 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_78
timestamp 1607194151
transform 1 0 8588 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_14
timestamp 1607194151
transform 1 0 8390 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_16
timestamp 1607194151
transform 1 0 9358 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_79
timestamp 1607194151
transform 1 0 9072 0 -1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap4_15
timestamp 1607194151
transform 1 0 8874 0 -1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_0
timestamp 1607194151
transform 1 0 1614 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_17
timestamp 1607194151
transform 1 0 1592 0 1 7532
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_16
timestamp 1607194151
transform 1 0 1416 0 1 7532
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_15
timestamp 1607194151
transform 1 0 1064 0 1 7532
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_94
timestamp 1607194151
transform 1 0 2296 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_1
timestamp 1607194151
transform 1 0 2098 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_95
timestamp 1607194151
transform 1 0 1812 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_3
timestamp 1607194151
transform 1 0 3066 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_93
timestamp 1607194151
transform 1 0 2780 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_2
timestamp 1607194151
transform 1 0 2582 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_91
timestamp 1607194151
transform 1 0 3748 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_4
timestamp 1607194151
transform 1 0 3550 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_92
timestamp 1607194151
transform 1 0 3264 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_6
timestamp 1607194151
transform 1 0 4518 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_90
timestamp 1607194151
transform 1 0 4232 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_5
timestamp 1607194151
transform 1 0 4034 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_88
timestamp 1607194151
transform 1 0 5200 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_7
timestamp 1607194151
transform 1 0 5002 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_89
timestamp 1607194151
transform 1 0 4716 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_9
timestamp 1607194151
transform 1 0 5970 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_87
timestamp 1607194151
transform 1 0 5684 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_8
timestamp 1607194151
transform 1 0 5486 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_85
timestamp 1607194151
transform 1 0 6652 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_10
timestamp 1607194151
transform 1 0 6454 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_86
timestamp 1607194151
transform 1 0 6168 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_84
timestamp 1607194151
transform 1 0 7136 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_11
timestamp 1607194151
transform 1 0 6938 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_82
timestamp 1607194151
transform 1 0 8104 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_13
timestamp 1607194151
transform 1 0 7906 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_83
timestamp 1607194151
transform 1 0 7620 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_12
timestamp 1607194151
transform 1 0 7422 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_81
timestamp 1607194151
transform 1 0 8588 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_14
timestamp 1607194151
transform 1 0 8390 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_16
timestamp 1607194151
transform 1 0 9358 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_80
timestamp 1607194151
transform 1 0 9072 0 1 7532
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap5_15
timestamp 1607194151
transform 1 0 8874 0 1 7532
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_0
timestamp 1607194151
transform 1 0 1614 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_20
timestamp 1607194151
transform 1 0 1592 0 -1 10196
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_19
timestamp 1607194151
transform 1 0 1416 0 -1 10196
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_18
timestamp 1607194151
transform 1 0 1064 0 -1 10196
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_97
timestamp 1607194151
transform 1 0 2296 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_1
timestamp 1607194151
transform 1 0 2098 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_96
timestamp 1607194151
transform 1 0 1812 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_3
timestamp 1607194151
transform 1 0 3066 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_98
timestamp 1607194151
transform 1 0 2780 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_2
timestamp 1607194151
transform 1 0 2582 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_100
timestamp 1607194151
transform 1 0 3748 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_4
timestamp 1607194151
transform 1 0 3550 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_99
timestamp 1607194151
transform 1 0 3264 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_6
timestamp 1607194151
transform 1 0 4518 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_101
timestamp 1607194151
transform 1 0 4232 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_5
timestamp 1607194151
transform 1 0 4034 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_103
timestamp 1607194151
transform 1 0 5200 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_7
timestamp 1607194151
transform 1 0 5002 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_102
timestamp 1607194151
transform 1 0 4716 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_9
timestamp 1607194151
transform 1 0 5970 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_104
timestamp 1607194151
transform 1 0 5684 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_8
timestamp 1607194151
transform 1 0 5486 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_106
timestamp 1607194151
transform 1 0 6652 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_10
timestamp 1607194151
transform 1 0 6454 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_105
timestamp 1607194151
transform 1 0 6168 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_107
timestamp 1607194151
transform 1 0 7136 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_11
timestamp 1607194151
transform 1 0 6938 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_109
timestamp 1607194151
transform 1 0 8104 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_13
timestamp 1607194151
transform 1 0 7906 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_108
timestamp 1607194151
transform 1 0 7620 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_12
timestamp 1607194151
transform 1 0 7422 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_110
timestamp 1607194151
transform 1 0 8588 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_14
timestamp 1607194151
transform 1 0 8390 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_16
timestamp 1607194151
transform 1 0 9358 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_111
timestamp 1607194151
transform 1 0 9072 0 -1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap6_15
timestamp 1607194151
transform 1 0 8874 0 -1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_0
timestamp 1607194151
transform 1 0 1614 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_23
timestamp 1607194151
transform 1 0 1592 0 1 10196
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_22
timestamp 1607194151
transform 1 0 1416 0 1 10196
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_21
timestamp 1607194151
transform 1 0 1064 0 1 10196
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_126
timestamp 1607194151
transform 1 0 2296 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_1
timestamp 1607194151
transform 1 0 2098 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_127
timestamp 1607194151
transform 1 0 1812 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_3
timestamp 1607194151
transform 1 0 3066 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_125
timestamp 1607194151
transform 1 0 2780 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_2
timestamp 1607194151
transform 1 0 2582 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_123
timestamp 1607194151
transform 1 0 3748 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_4
timestamp 1607194151
transform 1 0 3550 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_124
timestamp 1607194151
transform 1 0 3264 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_6
timestamp 1607194151
transform 1 0 4518 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_122
timestamp 1607194151
transform 1 0 4232 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_5
timestamp 1607194151
transform 1 0 4034 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_120
timestamp 1607194151
transform 1 0 5200 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_7
timestamp 1607194151
transform 1 0 5002 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_121
timestamp 1607194151
transform 1 0 4716 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_9
timestamp 1607194151
transform 1 0 5970 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_119
timestamp 1607194151
transform 1 0 5684 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_8
timestamp 1607194151
transform 1 0 5486 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_117
timestamp 1607194151
transform 1 0 6652 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_10
timestamp 1607194151
transform 1 0 6454 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_118
timestamp 1607194151
transform 1 0 6168 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_116
timestamp 1607194151
transform 1 0 7136 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_11
timestamp 1607194151
transform 1 0 6938 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_114
timestamp 1607194151
transform 1 0 8104 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_13
timestamp 1607194151
transform 1 0 7906 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_115
timestamp 1607194151
transform 1 0 7620 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_12
timestamp 1607194151
transform 1 0 7422 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_113
timestamp 1607194151
transform 1 0 8588 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_14
timestamp 1607194151
transform 1 0 8390 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_16
timestamp 1607194151
transform 1 0 9358 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_112
timestamp 1607194151
transform 1 0 9072 0 1 10196
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap7_15
timestamp 1607194151
transform 1 0 8874 0 1 10196
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_0
timestamp 1607194151
transform 1 0 1614 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_26
timestamp 1607194151
transform 1 0 1592 0 -1 12860
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_25
timestamp 1607194151
transform 1 0 1416 0 -1 12860
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_24
timestamp 1607194151
transform 1 0 1064 0 -1 12860
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_129
timestamp 1607194151
transform 1 0 2296 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_1
timestamp 1607194151
transform 1 0 2098 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_128
timestamp 1607194151
transform 1 0 1812 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_3
timestamp 1607194151
transform 1 0 3066 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_130
timestamp 1607194151
transform 1 0 2780 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_2
timestamp 1607194151
transform 1 0 2582 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_132
timestamp 1607194151
transform 1 0 3748 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_4
timestamp 1607194151
transform 1 0 3550 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_131
timestamp 1607194151
transform 1 0 3264 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_6
timestamp 1607194151
transform 1 0 4518 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_133
timestamp 1607194151
transform 1 0 4232 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_5
timestamp 1607194151
transform 1 0 4034 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_135
timestamp 1607194151
transform 1 0 5200 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_7
timestamp 1607194151
transform 1 0 5002 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_134
timestamp 1607194151
transform 1 0 4716 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_9
timestamp 1607194151
transform 1 0 5970 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_136
timestamp 1607194151
transform 1 0 5684 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_8
timestamp 1607194151
transform 1 0 5486 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_138
timestamp 1607194151
transform 1 0 6652 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_10
timestamp 1607194151
transform 1 0 6454 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_137
timestamp 1607194151
transform 1 0 6168 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_139
timestamp 1607194151
transform 1 0 7136 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_11
timestamp 1607194151
transform 1 0 6938 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_141
timestamp 1607194151
transform 1 0 8104 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_13
timestamp 1607194151
transform 1 0 7906 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_140
timestamp 1607194151
transform 1 0 7620 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_12
timestamp 1607194151
transform 1 0 7422 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_142
timestamp 1607194151
transform 1 0 8588 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_14
timestamp 1607194151
transform 1 0 8390 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_16
timestamp 1607194151
transform 1 0 9358 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_143
timestamp 1607194151
transform 1 0 9072 0 -1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap8_15
timestamp 1607194151
transform 1 0 8874 0 -1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_0
timestamp 1607194151
transform 1 0 1614 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_29
timestamp 1607194151
transform 1 0 1592 0 1 12860
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_28
timestamp 1607194151
transform 1 0 1416 0 1 12860
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_27
timestamp 1607194151
transform 1 0 1064 0 1 12860
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_158
timestamp 1607194151
transform 1 0 2296 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_1
timestamp 1607194151
transform 1 0 2098 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_159
timestamp 1607194151
transform 1 0 1812 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_3
timestamp 1607194151
transform 1 0 3066 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_157
timestamp 1607194151
transform 1 0 2780 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_2
timestamp 1607194151
transform 1 0 2582 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_155
timestamp 1607194151
transform 1 0 3748 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_4
timestamp 1607194151
transform 1 0 3550 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_156
timestamp 1607194151
transform 1 0 3264 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_6
timestamp 1607194151
transform 1 0 4518 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_154
timestamp 1607194151
transform 1 0 4232 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_5
timestamp 1607194151
transform 1 0 4034 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_152
timestamp 1607194151
transform 1 0 5200 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_7
timestamp 1607194151
transform 1 0 5002 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_153
timestamp 1607194151
transform 1 0 4716 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_9
timestamp 1607194151
transform 1 0 5970 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_151
timestamp 1607194151
transform 1 0 5684 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_8
timestamp 1607194151
transform 1 0 5486 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_149
timestamp 1607194151
transform 1 0 6652 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_10
timestamp 1607194151
transform 1 0 6454 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_150
timestamp 1607194151
transform 1 0 6168 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_148
timestamp 1607194151
transform 1 0 7136 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_11
timestamp 1607194151
transform 1 0 6938 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_146
timestamp 1607194151
transform 1 0 8104 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_13
timestamp 1607194151
transform 1 0 7906 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_147
timestamp 1607194151
transform 1 0 7620 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_12
timestamp 1607194151
transform 1 0 7422 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_145
timestamp 1607194151
transform 1 0 8588 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_14
timestamp 1607194151
transform 1 0 8390 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_16
timestamp 1607194151
transform 1 0 9358 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_144
timestamp 1607194151
transform 1 0 9072 0 1 12860
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap9_15
timestamp 1607194151
transform 1 0 8874 0 1 12860
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_0
timestamp 1607194151
transform 1 0 1614 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_32
timestamp 1607194151
transform 1 0 1592 0 -1 15524
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_31
timestamp 1607194151
transform 1 0 1416 0 -1 15524
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_30
timestamp 1607194151
transform 1 0 1064 0 -1 15524
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_161
timestamp 1607194151
transform 1 0 2296 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_1
timestamp 1607194151
transform 1 0 2098 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_160
timestamp 1607194151
transform 1 0 1812 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_3
timestamp 1607194151
transform 1 0 3066 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_162
timestamp 1607194151
transform 1 0 2780 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_2
timestamp 1607194151
transform 1 0 2582 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_164
timestamp 1607194151
transform 1 0 3748 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_4
timestamp 1607194151
transform 1 0 3550 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_163
timestamp 1607194151
transform 1 0 3264 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_6
timestamp 1607194151
transform 1 0 4518 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_165
timestamp 1607194151
transform 1 0 4232 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_5
timestamp 1607194151
transform 1 0 4034 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_167
timestamp 1607194151
transform 1 0 5200 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_7
timestamp 1607194151
transform 1 0 5002 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_166
timestamp 1607194151
transform 1 0 4716 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_9
timestamp 1607194151
transform 1 0 5970 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_168
timestamp 1607194151
transform 1 0 5684 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_8
timestamp 1607194151
transform 1 0 5486 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_170
timestamp 1607194151
transform 1 0 6652 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_10
timestamp 1607194151
transform 1 0 6454 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_169
timestamp 1607194151
transform 1 0 6168 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_171
timestamp 1607194151
transform 1 0 7136 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_11
timestamp 1607194151
transform 1 0 6938 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_173
timestamp 1607194151
transform 1 0 8104 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_13
timestamp 1607194151
transform 1 0 7906 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_172
timestamp 1607194151
transform 1 0 7620 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_12
timestamp 1607194151
transform 1 0 7422 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_174
timestamp 1607194151
transform 1 0 8588 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_14
timestamp 1607194151
transform 1 0 8390 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_16
timestamp 1607194151
transform 1 0 9358 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_175
timestamp 1607194151
transform 1 0 9072 0 -1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap10_15
timestamp 1607194151
transform 1 0 8874 0 -1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_0
timestamp 1607194151
transform 1 0 1614 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_35
timestamp 1607194151
transform 1 0 1592 0 1 15524
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_34
timestamp 1607194151
transform 1 0 1416 0 1 15524
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_33
timestamp 1607194151
transform 1 0 1064 0 1 15524
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_190
timestamp 1607194151
transform 1 0 2296 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_1
timestamp 1607194151
transform 1 0 2098 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_191
timestamp 1607194151
transform 1 0 1812 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_3
timestamp 1607194151
transform 1 0 3066 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_189
timestamp 1607194151
transform 1 0 2780 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_2
timestamp 1607194151
transform 1 0 2582 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_187
timestamp 1607194151
transform 1 0 3748 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_4
timestamp 1607194151
transform 1 0 3550 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_188
timestamp 1607194151
transform 1 0 3264 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_6
timestamp 1607194151
transform 1 0 4518 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_186
timestamp 1607194151
transform 1 0 4232 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_5
timestamp 1607194151
transform 1 0 4034 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_184
timestamp 1607194151
transform 1 0 5200 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_7
timestamp 1607194151
transform 1 0 5002 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_185
timestamp 1607194151
transform 1 0 4716 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_9
timestamp 1607194151
transform 1 0 5970 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_183
timestamp 1607194151
transform 1 0 5684 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_8
timestamp 1607194151
transform 1 0 5486 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_181
timestamp 1607194151
transform 1 0 6652 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_10
timestamp 1607194151
transform 1 0 6454 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_182
timestamp 1607194151
transform 1 0 6168 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_180
timestamp 1607194151
transform 1 0 7136 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_11
timestamp 1607194151
transform 1 0 6938 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_178
timestamp 1607194151
transform 1 0 8104 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_13
timestamp 1607194151
transform 1 0 7906 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_179
timestamp 1607194151
transform 1 0 7620 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_12
timestamp 1607194151
transform 1 0 7422 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_177
timestamp 1607194151
transform 1 0 8588 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_14
timestamp 1607194151
transform 1 0 8390 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_16
timestamp 1607194151
transform 1 0 9358 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_176
timestamp 1607194151
transform 1 0 9072 0 1 15524
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap11_15
timestamp 1607194151
transform 1 0 8874 0 1 15524
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_0
timestamp 1607194151
transform 1 0 1614 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_38
timestamp 1607194151
transform 1 0 1592 0 -1 18188
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_37
timestamp 1607194151
transform 1 0 1416 0 -1 18188
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_36
timestamp 1607194151
transform 1 0 1064 0 -1 18188
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_193
timestamp 1607194151
transform 1 0 2296 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_1
timestamp 1607194151
transform 1 0 2098 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_192
timestamp 1607194151
transform 1 0 1812 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_3
timestamp 1607194151
transform 1 0 3066 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_194
timestamp 1607194151
transform 1 0 2780 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_2
timestamp 1607194151
transform 1 0 2582 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_196
timestamp 1607194151
transform 1 0 3748 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_4
timestamp 1607194151
transform 1 0 3550 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_195
timestamp 1607194151
transform 1 0 3264 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_6
timestamp 1607194151
transform 1 0 4518 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_197
timestamp 1607194151
transform 1 0 4232 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_5
timestamp 1607194151
transform 1 0 4034 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_199
timestamp 1607194151
transform 1 0 5200 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_7
timestamp 1607194151
transform 1 0 5002 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_198
timestamp 1607194151
transform 1 0 4716 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_9
timestamp 1607194151
transform 1 0 5970 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_200
timestamp 1607194151
transform 1 0 5684 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_8
timestamp 1607194151
transform 1 0 5486 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_202
timestamp 1607194151
transform 1 0 6652 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_10
timestamp 1607194151
transform 1 0 6454 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_201
timestamp 1607194151
transform 1 0 6168 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_203
timestamp 1607194151
transform 1 0 7136 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_11
timestamp 1607194151
transform 1 0 6938 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_205
timestamp 1607194151
transform 1 0 8104 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_13
timestamp 1607194151
transform 1 0 7906 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_204
timestamp 1607194151
transform 1 0 7620 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_12
timestamp 1607194151
transform 1 0 7422 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_206
timestamp 1607194151
transform 1 0 8588 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_14
timestamp 1607194151
transform 1 0 8390 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_16
timestamp 1607194151
transform 1 0 9358 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_207
timestamp 1607194151
transform 1 0 9072 0 -1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap12_15
timestamp 1607194151
transform 1 0 8874 0 -1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_0
timestamp 1607194151
transform 1 0 1614 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_41
timestamp 1607194151
transform 1 0 1592 0 1 18188
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_40
timestamp 1607194151
transform 1 0 1416 0 1 18188
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_39
timestamp 1607194151
transform 1 0 1064 0 1 18188
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_222
timestamp 1607194151
transform 1 0 2296 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_1
timestamp 1607194151
transform 1 0 2098 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_223
timestamp 1607194151
transform 1 0 1812 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_3
timestamp 1607194151
transform 1 0 3066 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_221
timestamp 1607194151
transform 1 0 2780 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_2
timestamp 1607194151
transform 1 0 2582 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_219
timestamp 1607194151
transform 1 0 3748 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_4
timestamp 1607194151
transform 1 0 3550 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_220
timestamp 1607194151
transform 1 0 3264 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_6
timestamp 1607194151
transform 1 0 4518 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_218
timestamp 1607194151
transform 1 0 4232 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_5
timestamp 1607194151
transform 1 0 4034 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_216
timestamp 1607194151
transform 1 0 5200 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_7
timestamp 1607194151
transform 1 0 5002 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_217
timestamp 1607194151
transform 1 0 4716 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_9
timestamp 1607194151
transform 1 0 5970 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_215
timestamp 1607194151
transform 1 0 5684 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_8
timestamp 1607194151
transform 1 0 5486 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_213
timestamp 1607194151
transform 1 0 6652 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_10
timestamp 1607194151
transform 1 0 6454 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_214
timestamp 1607194151
transform 1 0 6168 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_212
timestamp 1607194151
transform 1 0 7136 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_11
timestamp 1607194151
transform 1 0 6938 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_210
timestamp 1607194151
transform 1 0 8104 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_13
timestamp 1607194151
transform 1 0 7906 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_211
timestamp 1607194151
transform 1 0 7620 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_12
timestamp 1607194151
transform 1 0 7422 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_209
timestamp 1607194151
transform 1 0 8588 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_14
timestamp 1607194151
transform 1 0 8390 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_16
timestamp 1607194151
transform 1 0 9358 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_208
timestamp 1607194151
transform 1 0 9072 0 1 18188
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap13_15
timestamp 1607194151
transform 1 0 8874 0 1 18188
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_0
timestamp 1607194151
transform 1 0 1614 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_44
timestamp 1607194151
transform 1 0 1592 0 -1 20852
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_43
timestamp 1607194151
transform 1 0 1416 0 -1 20852
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_42
timestamp 1607194151
transform 1 0 1064 0 -1 20852
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_8_225
timestamp 1607194151
transform 1 0 2296 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_1
timestamp 1607194151
transform 1 0 2098 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_224
timestamp 1607194151
transform 1 0 1812 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_3
timestamp 1607194151
transform 1 0 3066 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_226
timestamp 1607194151
transform 1 0 2780 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_2
timestamp 1607194151
transform 1 0 2582 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_228
timestamp 1607194151
transform 1 0 3748 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_4
timestamp 1607194151
transform 1 0 3550 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_227
timestamp 1607194151
transform 1 0 3264 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_6
timestamp 1607194151
transform 1 0 4518 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_229
timestamp 1607194151
transform 1 0 4232 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_5
timestamp 1607194151
transform 1 0 4034 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_231
timestamp 1607194151
transform 1 0 5200 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_7
timestamp 1607194151
transform 1 0 5002 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_230
timestamp 1607194151
transform 1 0 4716 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_9
timestamp 1607194151
transform 1 0 5970 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_232
timestamp 1607194151
transform 1 0 5684 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_8
timestamp 1607194151
transform 1 0 5486 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_234
timestamp 1607194151
transform 1 0 6652 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_10
timestamp 1607194151
transform 1 0 6454 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_233
timestamp 1607194151
transform 1 0 6168 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_235
timestamp 1607194151
transform 1 0 7136 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_11
timestamp 1607194151
transform 1 0 6938 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_237
timestamp 1607194151
transform 1 0 8104 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_13
timestamp 1607194151
transform 1 0 7906 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_236
timestamp 1607194151
transform 1 0 7620 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_12
timestamp 1607194151
transform 1 0 7422 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_238
timestamp 1607194151
transform 1 0 8588 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_14
timestamp 1607194151
transform 1 0 8390 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_16
timestamp 1607194151
transform 1 0 9358 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_239
timestamp 1607194151
transform 1 0 9072 0 -1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap14_15
timestamp 1607194151
transform 1 0 8874 0 -1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_0
timestamp 1607194151
transform 1 0 1614 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_8 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 1064 0 1 20852
box -9 0 553 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_254
timestamp 1607194151
transform 1 0 2296 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_1
timestamp 1607194151
transform 1 0 2098 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_255
timestamp 1607194151
transform 1 0 1812 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_3
timestamp 1607194151
transform 1 0 3066 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_253
timestamp 1607194151
transform 1 0 2780 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_2
timestamp 1607194151
transform 1 0 2582 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_251
timestamp 1607194151
transform 1 0 3748 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_4
timestamp 1607194151
transform 1 0 3550 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_252
timestamp 1607194151
transform 1 0 3264 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_6
timestamp 1607194151
transform 1 0 4518 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_250
timestamp 1607194151
transform 1 0 4232 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_5
timestamp 1607194151
transform 1 0 4034 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_248
timestamp 1607194151
transform 1 0 5200 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_7
timestamp 1607194151
transform 1 0 5002 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_249
timestamp 1607194151
transform 1 0 4716 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_9
timestamp 1607194151
transform 1 0 5970 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_247
timestamp 1607194151
transform 1 0 5684 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_8
timestamp 1607194151
transform 1 0 5486 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_245
timestamp 1607194151
transform 1 0 6652 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_10
timestamp 1607194151
transform 1 0 6454 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_246
timestamp 1607194151
transform 1 0 6168 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_244
timestamp 1607194151
transform 1 0 7136 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_11
timestamp 1607194151
transform 1 0 6938 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_242
timestamp 1607194151
transform 1 0 8104 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_13
timestamp 1607194151
transform 1 0 7906 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_243
timestamp 1607194151
transform 1 0 7620 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_12
timestamp 1607194151
transform 1 0 7422 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_241
timestamp 1607194151
transform 1 0 8588 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_14
timestamp 1607194151
transform 1 0 8390 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_16
timestamp 1607194151
transform 1 0 9358 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_8_240
timestamp 1607194151
transform 1 0 9072 0 1 20852
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap15_15
timestamp 1607194151
transform 1 0 8874 0 1 20852
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_0
timestamp 1607194151
transform 1 0 1614 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_47
timestamp 1607194151
transform 1 0 1592 0 -1 23516
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_46
timestamp 1607194151
transform 1 0 1416 0 -1 23516
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_45
timestamp 1607194151
transform 1 0 1064 0 -1 23516
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_7_1
timestamp 1607194151
transform 1 0 2296 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_1
timestamp 1607194151
transform 1 0 2098 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_0
timestamp 1607194151
transform 1 0 1812 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_3
timestamp 1607194151
transform 1 0 3066 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_2
timestamp 1607194151
transform 1 0 2780 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_2
timestamp 1607194151
transform 1 0 2582 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_4
timestamp 1607194151
transform 1 0 3748 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_4
timestamp 1607194151
transform 1 0 3550 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_3
timestamp 1607194151
transform 1 0 3264 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_6
timestamp 1607194151
transform 1 0 4518 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_5
timestamp 1607194151
transform 1 0 4232 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_5
timestamp 1607194151
transform 1 0 4034 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_7
timestamp 1607194151
transform 1 0 5200 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_7
timestamp 1607194151
transform 1 0 5002 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_6
timestamp 1607194151
transform 1 0 4716 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_9
timestamp 1607194151
transform 1 0 5970 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_8
timestamp 1607194151
transform 1 0 5684 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_8
timestamp 1607194151
transform 1 0 5486 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_10
timestamp 1607194151
transform 1 0 6652 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_10
timestamp 1607194151
transform 1 0 6454 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_9
timestamp 1607194151
transform 1 0 6168 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_11
timestamp 1607194151
transform 1 0 7136 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_11
timestamp 1607194151
transform 1 0 6938 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_13
timestamp 1607194151
transform 1 0 8104 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_13
timestamp 1607194151
transform 1 0 7906 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_12
timestamp 1607194151
transform 1 0 7620 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_12
timestamp 1607194151
transform 1 0 7422 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_14
timestamp 1607194151
transform 1 0 8588 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_14
timestamp 1607194151
transform 1 0 8390 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_16
timestamp 1607194151
transform 1 0 9358 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_15
timestamp 1607194151
transform 1 0 9072 0 -1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap16_15
timestamp 1607194151
transform 1 0 8874 0 -1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_0
timestamp 1607194151
transform 1 0 1614 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_50
timestamp 1607194151
transform 1 0 1592 0 1 23516
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_49
timestamp 1607194151
transform 1 0 1416 0 1 23516
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_48
timestamp 1607194151
transform 1 0 1064 0 1 23516
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_7_30
timestamp 1607194151
transform 1 0 2296 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_1
timestamp 1607194151
transform 1 0 2098 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_31
timestamp 1607194151
transform 1 0 1812 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_3
timestamp 1607194151
transform 1 0 3066 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_29
timestamp 1607194151
transform 1 0 2780 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_2
timestamp 1607194151
transform 1 0 2582 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_27
timestamp 1607194151
transform 1 0 3748 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_4
timestamp 1607194151
transform 1 0 3550 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_28
timestamp 1607194151
transform 1 0 3264 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_6
timestamp 1607194151
transform 1 0 4518 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_26
timestamp 1607194151
transform 1 0 4232 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_5
timestamp 1607194151
transform 1 0 4034 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_24
timestamp 1607194151
transform 1 0 5200 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_7
timestamp 1607194151
transform 1 0 5002 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_25
timestamp 1607194151
transform 1 0 4716 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_9
timestamp 1607194151
transform 1 0 5970 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_23
timestamp 1607194151
transform 1 0 5684 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_8
timestamp 1607194151
transform 1 0 5486 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_21
timestamp 1607194151
transform 1 0 6652 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_10
timestamp 1607194151
transform 1 0 6454 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_22
timestamp 1607194151
transform 1 0 6168 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_20
timestamp 1607194151
transform 1 0 7136 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_11
timestamp 1607194151
transform 1 0 6938 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_18
timestamp 1607194151
transform 1 0 8104 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_13
timestamp 1607194151
transform 1 0 7906 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_19
timestamp 1607194151
transform 1 0 7620 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_12
timestamp 1607194151
transform 1 0 7422 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_17
timestamp 1607194151
transform 1 0 8588 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_14
timestamp 1607194151
transform 1 0 8390 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_16
timestamp 1607194151
transform 1 0 9358 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_16
timestamp 1607194151
transform 1 0 9072 0 1 23516
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap17_15
timestamp 1607194151
transform 1 0 8874 0 1 23516
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_0
timestamp 1607194151
transform 1 0 1614 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_53
timestamp 1607194151
transform 1 0 1592 0 -1 26180
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_52
timestamp 1607194151
transform 1 0 1416 0 -1 26180
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_51
timestamp 1607194151
transform 1 0 1064 0 -1 26180
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_7_33
timestamp 1607194151
transform 1 0 2296 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_1
timestamp 1607194151
transform 1 0 2098 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_32
timestamp 1607194151
transform 1 0 1812 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_3
timestamp 1607194151
transform 1 0 3066 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_34
timestamp 1607194151
transform 1 0 2780 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_2
timestamp 1607194151
transform 1 0 2582 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_36
timestamp 1607194151
transform 1 0 3748 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_4
timestamp 1607194151
transform 1 0 3550 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_35
timestamp 1607194151
transform 1 0 3264 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_6
timestamp 1607194151
transform 1 0 4518 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_37
timestamp 1607194151
transform 1 0 4232 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_5
timestamp 1607194151
transform 1 0 4034 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_39
timestamp 1607194151
transform 1 0 5200 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_7
timestamp 1607194151
transform 1 0 5002 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_38
timestamp 1607194151
transform 1 0 4716 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_9
timestamp 1607194151
transform 1 0 5970 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_40
timestamp 1607194151
transform 1 0 5684 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_8
timestamp 1607194151
transform 1 0 5486 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_42
timestamp 1607194151
transform 1 0 6652 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_10
timestamp 1607194151
transform 1 0 6454 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_41
timestamp 1607194151
transform 1 0 6168 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_43
timestamp 1607194151
transform 1 0 7136 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_11
timestamp 1607194151
transform 1 0 6938 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_45
timestamp 1607194151
transform 1 0 8104 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_13
timestamp 1607194151
transform 1 0 7906 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_44
timestamp 1607194151
transform 1 0 7620 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_12
timestamp 1607194151
transform 1 0 7422 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_46
timestamp 1607194151
transform 1 0 8588 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_14
timestamp 1607194151
transform 1 0 8390 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_16
timestamp 1607194151
transform 1 0 9358 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_47
timestamp 1607194151
transform 1 0 9072 0 -1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap18_15
timestamp 1607194151
transform 1 0 8874 0 -1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_0
timestamp 1607194151
transform 1 0 1614 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_56
timestamp 1607194151
transform 1 0 1592 0 1 26180
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_55
timestamp 1607194151
transform 1 0 1416 0 1 26180
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_54
timestamp 1607194151
transform 1 0 1064 0 1 26180
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_7_62
timestamp 1607194151
transform 1 0 2296 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_1
timestamp 1607194151
transform 1 0 2098 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_63
timestamp 1607194151
transform 1 0 1812 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_3
timestamp 1607194151
transform 1 0 3066 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_61
timestamp 1607194151
transform 1 0 2780 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_2
timestamp 1607194151
transform 1 0 2582 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_59
timestamp 1607194151
transform 1 0 3748 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_4
timestamp 1607194151
transform 1 0 3550 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_60
timestamp 1607194151
transform 1 0 3264 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_6
timestamp 1607194151
transform 1 0 4518 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_58
timestamp 1607194151
transform 1 0 4232 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_5
timestamp 1607194151
transform 1 0 4034 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_56
timestamp 1607194151
transform 1 0 5200 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_7
timestamp 1607194151
transform 1 0 5002 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_57
timestamp 1607194151
transform 1 0 4716 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_9
timestamp 1607194151
transform 1 0 5970 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_55
timestamp 1607194151
transform 1 0 5684 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_8
timestamp 1607194151
transform 1 0 5486 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_53
timestamp 1607194151
transform 1 0 6652 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_10
timestamp 1607194151
transform 1 0 6454 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_54
timestamp 1607194151
transform 1 0 6168 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_52
timestamp 1607194151
transform 1 0 7136 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_11
timestamp 1607194151
transform 1 0 6938 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_50
timestamp 1607194151
transform 1 0 8104 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_13
timestamp 1607194151
transform 1 0 7906 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_51
timestamp 1607194151
transform 1 0 7620 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_12
timestamp 1607194151
transform 1 0 7422 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_49
timestamp 1607194151
transform 1 0 8588 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_14
timestamp 1607194151
transform 1 0 8390 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_16
timestamp 1607194151
transform 1 0 9358 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_48
timestamp 1607194151
transform 1 0 9072 0 1 26180
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap19_15
timestamp 1607194151
transform 1 0 8874 0 1 26180
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_0
timestamp 1607194151
transform 1 0 1614 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_59
timestamp 1607194151
transform 1 0 1592 0 -1 28844
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_58
timestamp 1607194151
transform 1 0 1416 0 -1 28844
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_57
timestamp 1607194151
transform 1 0 1064 0 -1 28844
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_7_65
timestamp 1607194151
transform 1 0 2296 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_1
timestamp 1607194151
transform 1 0 2098 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_64
timestamp 1607194151
transform 1 0 1812 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_3
timestamp 1607194151
transform 1 0 3066 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_66
timestamp 1607194151
transform 1 0 2780 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_2
timestamp 1607194151
transform 1 0 2582 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_68
timestamp 1607194151
transform 1 0 3748 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_4
timestamp 1607194151
transform 1 0 3550 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_67
timestamp 1607194151
transform 1 0 3264 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_6
timestamp 1607194151
transform 1 0 4518 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_69
timestamp 1607194151
transform 1 0 4232 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_5
timestamp 1607194151
transform 1 0 4034 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_71
timestamp 1607194151
transform 1 0 5200 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_7
timestamp 1607194151
transform 1 0 5002 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_70
timestamp 1607194151
transform 1 0 4716 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_9
timestamp 1607194151
transform 1 0 5970 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_72
timestamp 1607194151
transform 1 0 5684 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_8
timestamp 1607194151
transform 1 0 5486 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_74
timestamp 1607194151
transform 1 0 6652 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_10
timestamp 1607194151
transform 1 0 6454 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_73
timestamp 1607194151
transform 1 0 6168 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_75
timestamp 1607194151
transform 1 0 7136 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_11
timestamp 1607194151
transform 1 0 6938 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_77
timestamp 1607194151
transform 1 0 8104 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_13
timestamp 1607194151
transform 1 0 7906 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_76
timestamp 1607194151
transform 1 0 7620 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_12
timestamp 1607194151
transform 1 0 7422 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_78
timestamp 1607194151
transform 1 0 8588 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_14
timestamp 1607194151
transform 1 0 8390 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_16
timestamp 1607194151
transform 1 0 9358 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_79
timestamp 1607194151
transform 1 0 9072 0 -1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap20_15
timestamp 1607194151
transform 1 0 8874 0 -1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_0
timestamp 1607194151
transform 1 0 1614 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_62
timestamp 1607194151
transform 1 0 1592 0 1 28844
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_61
timestamp 1607194151
transform 1 0 1416 0 1 28844
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_60
timestamp 1607194151
transform 1 0 1064 0 1 28844
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_7_94
timestamp 1607194151
transform 1 0 2296 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_1
timestamp 1607194151
transform 1 0 2098 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_95
timestamp 1607194151
transform 1 0 1812 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_3
timestamp 1607194151
transform 1 0 3066 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_93
timestamp 1607194151
transform 1 0 2780 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_2
timestamp 1607194151
transform 1 0 2582 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_91
timestamp 1607194151
transform 1 0 3748 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_4
timestamp 1607194151
transform 1 0 3550 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_92
timestamp 1607194151
transform 1 0 3264 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_6
timestamp 1607194151
transform 1 0 4518 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_90
timestamp 1607194151
transform 1 0 4232 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_5
timestamp 1607194151
transform 1 0 4034 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_88
timestamp 1607194151
transform 1 0 5200 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_7
timestamp 1607194151
transform 1 0 5002 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_89
timestamp 1607194151
transform 1 0 4716 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_9
timestamp 1607194151
transform 1 0 5970 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_87
timestamp 1607194151
transform 1 0 5684 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_8
timestamp 1607194151
transform 1 0 5486 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_85
timestamp 1607194151
transform 1 0 6652 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_10
timestamp 1607194151
transform 1 0 6454 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_86
timestamp 1607194151
transform 1 0 6168 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_84
timestamp 1607194151
transform 1 0 7136 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_11
timestamp 1607194151
transform 1 0 6938 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_82
timestamp 1607194151
transform 1 0 8104 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_13
timestamp 1607194151
transform 1 0 7906 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_83
timestamp 1607194151
transform 1 0 7620 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_12
timestamp 1607194151
transform 1 0 7422 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_81
timestamp 1607194151
transform 1 0 8588 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_14
timestamp 1607194151
transform 1 0 8390 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_16
timestamp 1607194151
transform 1 0 9358 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_80
timestamp 1607194151
transform 1 0 9072 0 1 28844
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap21_15
timestamp 1607194151
transform 1 0 8874 0 1 28844
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_0
timestamp 1607194151
transform 1 0 1614 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_65
timestamp 1607194151
transform 1 0 1592 0 -1 31508
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_64
timestamp 1607194151
transform 1 0 1416 0 -1 31508
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_63
timestamp 1607194151
transform 1 0 1064 0 -1 31508
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_7_97
timestamp 1607194151
transform 1 0 2296 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_1
timestamp 1607194151
transform 1 0 2098 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_96
timestamp 1607194151
transform 1 0 1812 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_3
timestamp 1607194151
transform 1 0 3066 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_98
timestamp 1607194151
transform 1 0 2780 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_2
timestamp 1607194151
transform 1 0 2582 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_100
timestamp 1607194151
transform 1 0 3748 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_4
timestamp 1607194151
transform 1 0 3550 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_99
timestamp 1607194151
transform 1 0 3264 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_6
timestamp 1607194151
transform 1 0 4518 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_101
timestamp 1607194151
transform 1 0 4232 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_5
timestamp 1607194151
transform 1 0 4034 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_103
timestamp 1607194151
transform 1 0 5200 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_7
timestamp 1607194151
transform 1 0 5002 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_102
timestamp 1607194151
transform 1 0 4716 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_9
timestamp 1607194151
transform 1 0 5970 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_104
timestamp 1607194151
transform 1 0 5684 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_8
timestamp 1607194151
transform 1 0 5486 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_106
timestamp 1607194151
transform 1 0 6652 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_10
timestamp 1607194151
transform 1 0 6454 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_105
timestamp 1607194151
transform 1 0 6168 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_107
timestamp 1607194151
transform 1 0 7136 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_11
timestamp 1607194151
transform 1 0 6938 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_109
timestamp 1607194151
transform 1 0 8104 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_13
timestamp 1607194151
transform 1 0 7906 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_108
timestamp 1607194151
transform 1 0 7620 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_12
timestamp 1607194151
transform 1 0 7422 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_110
timestamp 1607194151
transform 1 0 8588 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_14
timestamp 1607194151
transform 1 0 8390 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_16
timestamp 1607194151
transform 1 0 9358 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_111
timestamp 1607194151
transform 1 0 9072 0 -1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap22_15
timestamp 1607194151
transform 1 0 8874 0 -1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_0
timestamp 1607194151
transform 1 0 1614 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_7
timestamp 1607194151
transform 1 0 1064 0 1 31508
box -9 0 553 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_126
timestamp 1607194151
transform 1 0 2296 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_1
timestamp 1607194151
transform 1 0 2098 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_127
timestamp 1607194151
transform 1 0 1812 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_3
timestamp 1607194151
transform 1 0 3066 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_125
timestamp 1607194151
transform 1 0 2780 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_2
timestamp 1607194151
transform 1 0 2582 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_123
timestamp 1607194151
transform 1 0 3748 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_4
timestamp 1607194151
transform 1 0 3550 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_124
timestamp 1607194151
transform 1 0 3264 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_6
timestamp 1607194151
transform 1 0 4518 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_122
timestamp 1607194151
transform 1 0 4232 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_5
timestamp 1607194151
transform 1 0 4034 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_120
timestamp 1607194151
transform 1 0 5200 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_7
timestamp 1607194151
transform 1 0 5002 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_121
timestamp 1607194151
transform 1 0 4716 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_9
timestamp 1607194151
transform 1 0 5970 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_119
timestamp 1607194151
transform 1 0 5684 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_8
timestamp 1607194151
transform 1 0 5486 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_117
timestamp 1607194151
transform 1 0 6652 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_10
timestamp 1607194151
transform 1 0 6454 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_118
timestamp 1607194151
transform 1 0 6168 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_116
timestamp 1607194151
transform 1 0 7136 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_11
timestamp 1607194151
transform 1 0 6938 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_114
timestamp 1607194151
transform 1 0 8104 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_13
timestamp 1607194151
transform 1 0 7906 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_115
timestamp 1607194151
transform 1 0 7620 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_12
timestamp 1607194151
transform 1 0 7422 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_113
timestamp 1607194151
transform 1 0 8588 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_14
timestamp 1607194151
transform 1 0 8390 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_16
timestamp 1607194151
transform 1 0 9358 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_7_112
timestamp 1607194151
transform 1 0 9072 0 1 31508
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap23_15
timestamp 1607194151
transform 1 0 8874 0 1 31508
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_0
timestamp 1607194151
transform 1 0 1614 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_68
timestamp 1607194151
transform 1 0 1592 0 -1 34172
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_67
timestamp 1607194151
transform 1 0 1416 0 -1 34172
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_66
timestamp 1607194151
transform 1 0 1064 0 -1 34172
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_6_1
timestamp 1607194151
transform 1 0 2296 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_1
timestamp 1607194151
transform 1 0 2098 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_0
timestamp 1607194151
transform 1 0 1812 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_3
timestamp 1607194151
transform 1 0 3066 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_2
timestamp 1607194151
transform 1 0 2780 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_2
timestamp 1607194151
transform 1 0 2582 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_4
timestamp 1607194151
transform 1 0 3748 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_4
timestamp 1607194151
transform 1 0 3550 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_3
timestamp 1607194151
transform 1 0 3264 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_6
timestamp 1607194151
transform 1 0 4518 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_5
timestamp 1607194151
transform 1 0 4232 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_5
timestamp 1607194151
transform 1 0 4034 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_7
timestamp 1607194151
transform 1 0 5200 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_7
timestamp 1607194151
transform 1 0 5002 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_6
timestamp 1607194151
transform 1 0 4716 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_9
timestamp 1607194151
transform 1 0 5970 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_8
timestamp 1607194151
transform 1 0 5684 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_8
timestamp 1607194151
transform 1 0 5486 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_10
timestamp 1607194151
transform 1 0 6652 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_10
timestamp 1607194151
transform 1 0 6454 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_9
timestamp 1607194151
transform 1 0 6168 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_11
timestamp 1607194151
transform 1 0 7136 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_11
timestamp 1607194151
transform 1 0 6938 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_13
timestamp 1607194151
transform 1 0 8104 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_13
timestamp 1607194151
transform 1 0 7906 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_12
timestamp 1607194151
transform 1 0 7620 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_12
timestamp 1607194151
transform 1 0 7422 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_14
timestamp 1607194151
transform 1 0 8588 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_14
timestamp 1607194151
transform 1 0 8390 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_16
timestamp 1607194151
transform 1 0 9358 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_15
timestamp 1607194151
transform 1 0 9072 0 -1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap24_15
timestamp 1607194151
transform 1 0 8874 0 -1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_0
timestamp 1607194151
transform 1 0 1614 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_71
timestamp 1607194151
transform 1 0 1592 0 1 34172
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_70
timestamp 1607194151
transform 1 0 1416 0 1 34172
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_69
timestamp 1607194151
transform 1 0 1064 0 1 34172
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_6_30
timestamp 1607194151
transform 1 0 2296 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_1
timestamp 1607194151
transform 1 0 2098 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_31
timestamp 1607194151
transform 1 0 1812 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_3
timestamp 1607194151
transform 1 0 3066 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_29
timestamp 1607194151
transform 1 0 2780 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_2
timestamp 1607194151
transform 1 0 2582 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_27
timestamp 1607194151
transform 1 0 3748 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_4
timestamp 1607194151
transform 1 0 3550 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_28
timestamp 1607194151
transform 1 0 3264 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_6
timestamp 1607194151
transform 1 0 4518 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_26
timestamp 1607194151
transform 1 0 4232 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_5
timestamp 1607194151
transform 1 0 4034 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_24
timestamp 1607194151
transform 1 0 5200 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_7
timestamp 1607194151
transform 1 0 5002 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_25
timestamp 1607194151
transform 1 0 4716 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_9
timestamp 1607194151
transform 1 0 5970 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_23
timestamp 1607194151
transform 1 0 5684 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_8
timestamp 1607194151
transform 1 0 5486 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_21
timestamp 1607194151
transform 1 0 6652 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_10
timestamp 1607194151
transform 1 0 6454 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_22
timestamp 1607194151
transform 1 0 6168 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_20
timestamp 1607194151
transform 1 0 7136 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_11
timestamp 1607194151
transform 1 0 6938 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_18
timestamp 1607194151
transform 1 0 8104 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_13
timestamp 1607194151
transform 1 0 7906 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_19
timestamp 1607194151
transform 1 0 7620 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_12
timestamp 1607194151
transform 1 0 7422 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_17
timestamp 1607194151
transform 1 0 8588 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_14
timestamp 1607194151
transform 1 0 8390 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_16
timestamp 1607194151
transform 1 0 9358 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_16
timestamp 1607194151
transform 1 0 9072 0 1 34172
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap25_15
timestamp 1607194151
transform 1 0 8874 0 1 34172
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_0
timestamp 1607194151
transform 1 0 1614 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_74
timestamp 1607194151
transform 1 0 1592 0 -1 36836
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_73
timestamp 1607194151
transform 1 0 1416 0 -1 36836
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_72
timestamp 1607194151
transform 1 0 1064 0 -1 36836
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_6_33
timestamp 1607194151
transform 1 0 2296 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_1
timestamp 1607194151
transform 1 0 2098 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_32
timestamp 1607194151
transform 1 0 1812 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_3
timestamp 1607194151
transform 1 0 3066 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_34
timestamp 1607194151
transform 1 0 2780 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_2
timestamp 1607194151
transform 1 0 2582 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_36
timestamp 1607194151
transform 1 0 3748 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_4
timestamp 1607194151
transform 1 0 3550 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_35
timestamp 1607194151
transform 1 0 3264 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_6
timestamp 1607194151
transform 1 0 4518 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_37
timestamp 1607194151
transform 1 0 4232 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_5
timestamp 1607194151
transform 1 0 4034 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_39
timestamp 1607194151
transform 1 0 5200 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_7
timestamp 1607194151
transform 1 0 5002 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_38
timestamp 1607194151
transform 1 0 4716 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_9
timestamp 1607194151
transform 1 0 5970 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_40
timestamp 1607194151
transform 1 0 5684 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_8
timestamp 1607194151
transform 1 0 5486 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_42
timestamp 1607194151
transform 1 0 6652 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_10
timestamp 1607194151
transform 1 0 6454 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_41
timestamp 1607194151
transform 1 0 6168 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_43
timestamp 1607194151
transform 1 0 7136 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_11
timestamp 1607194151
transform 1 0 6938 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_45
timestamp 1607194151
transform 1 0 8104 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_13
timestamp 1607194151
transform 1 0 7906 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_44
timestamp 1607194151
transform 1 0 7620 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_12
timestamp 1607194151
transform 1 0 7422 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_46
timestamp 1607194151
transform 1 0 8588 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_14
timestamp 1607194151
transform 1 0 8390 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_16
timestamp 1607194151
transform 1 0 9358 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_47
timestamp 1607194151
transform 1 0 9072 0 -1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap26_15
timestamp 1607194151
transform 1 0 8874 0 -1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_0
timestamp 1607194151
transform 1 0 1614 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_6
timestamp 1607194151
transform 1 0 1064 0 1 36836
box -9 0 553 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_62
timestamp 1607194151
transform 1 0 2296 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_1
timestamp 1607194151
transform 1 0 2098 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_63
timestamp 1607194151
transform 1 0 1812 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_3
timestamp 1607194151
transform 1 0 3066 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_61
timestamp 1607194151
transform 1 0 2780 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_2
timestamp 1607194151
transform 1 0 2582 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_59
timestamp 1607194151
transform 1 0 3748 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_4
timestamp 1607194151
transform 1 0 3550 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_60
timestamp 1607194151
transform 1 0 3264 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_6
timestamp 1607194151
transform 1 0 4518 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_58
timestamp 1607194151
transform 1 0 4232 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_5
timestamp 1607194151
transform 1 0 4034 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_56
timestamp 1607194151
transform 1 0 5200 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_7
timestamp 1607194151
transform 1 0 5002 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_57
timestamp 1607194151
transform 1 0 4716 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_9
timestamp 1607194151
transform 1 0 5970 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_55
timestamp 1607194151
transform 1 0 5684 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_8
timestamp 1607194151
transform 1 0 5486 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_53
timestamp 1607194151
transform 1 0 6652 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_10
timestamp 1607194151
transform 1 0 6454 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_54
timestamp 1607194151
transform 1 0 6168 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_52
timestamp 1607194151
transform 1 0 7136 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_11
timestamp 1607194151
transform 1 0 6938 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_50
timestamp 1607194151
transform 1 0 8104 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_13
timestamp 1607194151
transform 1 0 7906 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_51
timestamp 1607194151
transform 1 0 7620 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_12
timestamp 1607194151
transform 1 0 7422 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_49
timestamp 1607194151
transform 1 0 8588 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_14
timestamp 1607194151
transform 1 0 8390 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_16
timestamp 1607194151
transform 1 0 9358 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_6_48
timestamp 1607194151
transform 1 0 9072 0 1 36836
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap27_15
timestamp 1607194151
transform 1 0 8874 0 1 36836
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_0
timestamp 1607194151
transform 1 0 1614 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_77
timestamp 1607194151
transform 1 0 1592 0 -1 39500
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_76
timestamp 1607194151
transform 1 0 1416 0 -1 39500
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_75
timestamp 1607194151
transform 1 0 1064 0 -1 39500
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_5_1
timestamp 1607194151
transform 1 0 2296 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_1
timestamp 1607194151
transform 1 0 2098 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_0
timestamp 1607194151
transform 1 0 1812 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_3
timestamp 1607194151
transform 1 0 3066 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_2
timestamp 1607194151
transform 1 0 2780 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_2
timestamp 1607194151
transform 1 0 2582 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_4
timestamp 1607194151
transform 1 0 3748 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_4
timestamp 1607194151
transform 1 0 3550 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_3
timestamp 1607194151
transform 1 0 3264 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_6
timestamp 1607194151
transform 1 0 4518 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_5
timestamp 1607194151
transform 1 0 4232 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_5
timestamp 1607194151
transform 1 0 4034 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_7
timestamp 1607194151
transform 1 0 5200 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_7
timestamp 1607194151
transform 1 0 5002 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_6
timestamp 1607194151
transform 1 0 4716 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_9
timestamp 1607194151
transform 1 0 5970 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_8
timestamp 1607194151
transform 1 0 5684 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_8
timestamp 1607194151
transform 1 0 5486 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_10
timestamp 1607194151
transform 1 0 6652 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_10
timestamp 1607194151
transform 1 0 6454 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_9
timestamp 1607194151
transform 1 0 6168 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_11
timestamp 1607194151
transform 1 0 7136 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_11
timestamp 1607194151
transform 1 0 6938 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_13
timestamp 1607194151
transform 1 0 8104 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_13
timestamp 1607194151
transform 1 0 7906 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_12
timestamp 1607194151
transform 1 0 7620 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_12
timestamp 1607194151
transform 1 0 7422 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_14
timestamp 1607194151
transform 1 0 8588 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_14
timestamp 1607194151
transform 1 0 8390 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_16
timestamp 1607194151
transform 1 0 9358 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_15
timestamp 1607194151
transform 1 0 9072 0 -1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap28_15
timestamp 1607194151
transform 1 0 8874 0 -1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_0
timestamp 1607194151
transform 1 0 1614 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_5
timestamp 1607194151
transform 1 0 1064 0 1 39500
box -9 0 553 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_30
timestamp 1607194151
transform 1 0 2296 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_1
timestamp 1607194151
transform 1 0 2098 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_31
timestamp 1607194151
transform 1 0 1812 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_3
timestamp 1607194151
transform 1 0 3066 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_29
timestamp 1607194151
transform 1 0 2780 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_2
timestamp 1607194151
transform 1 0 2582 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_27
timestamp 1607194151
transform 1 0 3748 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_4
timestamp 1607194151
transform 1 0 3550 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_28
timestamp 1607194151
transform 1 0 3264 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_6
timestamp 1607194151
transform 1 0 4518 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_26
timestamp 1607194151
transform 1 0 4232 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_5
timestamp 1607194151
transform 1 0 4034 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_24
timestamp 1607194151
transform 1 0 5200 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_7
timestamp 1607194151
transform 1 0 5002 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_25
timestamp 1607194151
transform 1 0 4716 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_9
timestamp 1607194151
transform 1 0 5970 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_23
timestamp 1607194151
transform 1 0 5684 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_8
timestamp 1607194151
transform 1 0 5486 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_21
timestamp 1607194151
transform 1 0 6652 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_10
timestamp 1607194151
transform 1 0 6454 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_22
timestamp 1607194151
transform 1 0 6168 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_20
timestamp 1607194151
transform 1 0 7136 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_11
timestamp 1607194151
transform 1 0 6938 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_18
timestamp 1607194151
transform 1 0 8104 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_13
timestamp 1607194151
transform 1 0 7906 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_19
timestamp 1607194151
transform 1 0 7620 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_12
timestamp 1607194151
transform 1 0 7422 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_17
timestamp 1607194151
transform 1 0 8588 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_14
timestamp 1607194151
transform 1 0 8390 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_16
timestamp 1607194151
transform 1 0 9358 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_5_16
timestamp 1607194151
transform 1 0 9072 0 1 39500
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap29_15
timestamp 1607194151
transform 1 0 8874 0 1 39500
box -9 0 199 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_0
timestamp 1607194151
transform 1 0 1614 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_80
timestamp 1607194151
transform 1 0 1592 0 -1 42164
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_79
timestamp 1607194151
transform 1 0 1416 0 -1 42164
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_78
timestamp 1607194151
transform 1 0 1064 0 -1 42164
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_4_1
timestamp 1607194151
transform 1 0 2296 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_1
timestamp 1607194151
transform 1 0 2098 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_0
timestamp 1607194151
transform 1 0 1812 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_3
timestamp 1607194151
transform 1 0 3066 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_2
timestamp 1607194151
transform 1 0 2780 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_2
timestamp 1607194151
transform 1 0 2582 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_4
timestamp 1607194151
transform 1 0 3748 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_4
timestamp 1607194151
transform 1 0 3550 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_3
timestamp 1607194151
transform 1 0 3264 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_6
timestamp 1607194151
transform 1 0 4518 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_5
timestamp 1607194151
transform 1 0 4232 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_5
timestamp 1607194151
transform 1 0 4034 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_7
timestamp 1607194151
transform 1 0 5200 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap30_7
timestamp 1607194151
transform 1 0 5002 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_6
timestamp 1607194151
transform 1 0 4716 0 -1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_90 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 5684 0 -1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap30_8
timestamp 1607194151
transform 1 0 5486 0 -1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_91
timestamp 1607194151
transform 1 0 6388 0 -1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_92
timestamp 1607194151
transform 1 0 7092 0 -1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_93
timestamp 1607194151
transform 1 0 7796 0 -1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_94
timestamp 1607194151
transform 1 0 8500 0 -1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_95
timestamp 1607194151
transform 1 0 9204 0 -1 42164
box 0 0 352 1332
use sky130_osu_sc_18T_hs__decap_1  decap31_0
timestamp 1607194151
transform 1 0 1614 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_4
timestamp 1607194151
transform 1 0 1064 0 1 42164
box -9 0 553 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_14
timestamp 1607194151
transform 1 0 2296 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap31_1
timestamp 1607194151
transform 1 0 2098 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_15
timestamp 1607194151
transform 1 0 1812 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap31_3
timestamp 1607194151
transform 1 0 3066 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_13
timestamp 1607194151
transform 1 0 2780 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap31_2
timestamp 1607194151
transform 1 0 2582 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_11
timestamp 1607194151
transform 1 0 3748 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap31_4
timestamp 1607194151
transform 1 0 3550 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_12
timestamp 1607194151
transform 1 0 3264 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap31_6
timestamp 1607194151
transform 1 0 4518 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_10
timestamp 1607194151
transform 1 0 4232 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap31_5
timestamp 1607194151
transform 1 0 4034 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_8
timestamp 1607194151
transform 1 0 5200 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap31_7
timestamp 1607194151
transform 1 0 5002 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_4_9
timestamp 1607194151
transform 1 0 4716 0 1 42164
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_96
timestamp 1607194151
transform 1 0 5684 0 1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap31_8
timestamp 1607194151
transform 1 0 5486 0 1 42164
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_97
timestamp 1607194151
transform 1 0 6388 0 1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_98
timestamp 1607194151
transform 1 0 7092 0 1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_99
timestamp 1607194151
transform 1 0 7796 0 1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_100
timestamp 1607194151
transform 1 0 8500 0 1 42164
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_101
timestamp 1607194151
transform 1 0 9204 0 1 42164
box 0 0 352 1332
use sky130_osu_sc_18T_hs__decap_1  decap32_0
timestamp 1607194151
transform 1 0 1614 0 -1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_83
timestamp 1607194151
transform 1 0 1592 0 -1 44828
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_82
timestamp 1607194151
transform 1 0 1416 0 -1 44828
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_81
timestamp 1607194151
transform 1 0 1064 0 -1 44828
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_3_1
timestamp 1607194151
transform 1 0 2296 0 -1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap32_1
timestamp 1607194151
transform 1 0 2098 0 -1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_3_0
timestamp 1607194151
transform 1 0 1812 0 -1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap32_3
timestamp 1607194151
transform 1 0 3066 0 -1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_3_2
timestamp 1607194151
transform 1 0 2780 0 -1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap32_2
timestamp 1607194151
transform 1 0 2582 0 -1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_102
timestamp 1607194151
transform 1 0 3748 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap32_4
timestamp 1607194151
transform 1 0 3550 0 -1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_3_3
timestamp 1607194151
transform 1 0 3264 0 -1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_103
timestamp 1607194151
transform 1 0 4452 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_104
timestamp 1607194151
transform 1 0 5156 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_105
timestamp 1607194151
transform 1 0 5860 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_106
timestamp 1607194151
transform 1 0 6564 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_107
timestamp 1607194151
transform 1 0 7268 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_108
timestamp 1607194151
transform 1 0 7972 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_109
timestamp 1607194151
transform 1 0 8676 0 -1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_110
timestamp 1607194151
transform 1 0 9380 0 -1 44828
box 0 0 176 1332
use sky130_osu_sc_18T_hs__decap_1  decap33_0
timestamp 1607194151
transform 1 0 1614 0 1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_3
timestamp 1607194151
transform 1 0 1064 0 1 44828
box -9 0 553 1341
use sky130_osu_sc_18T_hs__buf_1  delay_3_6
timestamp 1607194151
transform 1 0 2296 0 1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap33_1
timestamp 1607194151
transform 1 0 2098 0 1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_3_7
timestamp 1607194151
transform 1 0 1812 0 1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap33_3
timestamp 1607194151
transform 1 0 3066 0 1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_3_5
timestamp 1607194151
transform 1 0 2780 0 1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap33_2
timestamp 1607194151
transform 1 0 2582 0 1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_111
timestamp 1607194151
transform 1 0 3748 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap33_4
timestamp 1607194151
transform 1 0 3550 0 1 44828
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_3_4
timestamp 1607194151
transform 1 0 3264 0 1 44828
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_112
timestamp 1607194151
transform 1 0 4452 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_113
timestamp 1607194151
transform 1 0 5156 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_114
timestamp 1607194151
transform 1 0 5860 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_115
timestamp 1607194151
transform 1 0 6564 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_116
timestamp 1607194151
transform 1 0 7268 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_117
timestamp 1607194151
transform 1 0 7972 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_118
timestamp 1607194151
transform 1 0 8676 0 1 44828
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_119
timestamp 1607194151
transform 1 0 9380 0 1 44828
box 0 0 176 1332
use sky130_osu_sc_18T_hs__decap_1  decap34_0
timestamp 1607194151
transform 1 0 1614 0 -1 47492
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_86
timestamp 1607194151
transform 1 0 1592 0 -1 47492
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_85
timestamp 1607194151
transform 1 0 1416 0 -1 47492
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_84
timestamp 1607194151
transform 1 0 1064 0 -1 47492
box 0 0 352 1332
use sky130_osu_sc_18T_hs__buf_1  delay_2_1
timestamp 1607194151
transform 1 0 2296 0 -1 47492
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap34_1
timestamp 1607194151
transform 1 0 2098 0 -1 47492
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_2_0
timestamp 1607194151
transform 1 0 1812 0 -1 47492
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_120
timestamp 1607194151
transform 1 0 2780 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap34_2
timestamp 1607194151
transform 1 0 2582 0 -1 47492
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_121
timestamp 1607194151
transform 1 0 3484 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_122
timestamp 1607194151
transform 1 0 4188 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_123
timestamp 1607194151
transform 1 0 4892 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_124
timestamp 1607194151
transform 1 0 5596 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_125
timestamp 1607194151
transform 1 0 6300 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_126
timestamp 1607194151
transform 1 0 7004 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_127
timestamp 1607194151
transform 1 0 7708 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_128
timestamp 1607194151
transform 1 0 8412 0 -1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_4  FILL_130 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 9468 0 -1 47492
box 0 0 88 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_129
timestamp 1607194151
transform 1 0 9116 0 -1 47492
box 0 0 352 1332
use sky130_osu_sc_18T_hs__decap_1  decap35_0
timestamp 1607194151
transform 1 0 1614 0 1 47492
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_2
timestamp 1607194151
transform 1 0 1064 0 1 47492
box -9 0 553 1341
use sky130_osu_sc_18T_hs__buf_1  delay_2_2
timestamp 1607194151
transform 1 0 2296 0 1 47492
box -9 0 288 1341
use sky130_osu_sc_18T_hs__decap_1  decap35_1
timestamp 1607194151
transform 1 0 2098 0 1 47492
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_2_3
timestamp 1607194151
transform 1 0 1812 0 1 47492
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_131
timestamp 1607194151
transform 1 0 2780 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap35_2
timestamp 1607194151
transform 1 0 2582 0 1 47492
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_132
timestamp 1607194151
transform 1 0 3484 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_133
timestamp 1607194151
transform 1 0 4188 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_134
timestamp 1607194151
transform 1 0 4892 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_135
timestamp 1607194151
transform 1 0 5596 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_136
timestamp 1607194151
transform 1 0 6300 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_137
timestamp 1607194151
transform 1 0 7004 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_138
timestamp 1607194151
transform 1 0 7708 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_139
timestamp 1607194151
transform 1 0 8412 0 1 47492
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_4  FILL_141
timestamp 1607194151
transform 1 0 9468 0 1 47492
box 0 0 88 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_140
timestamp 1607194151
transform 1 0 9116 0 1 47492
box 0 0 352 1332
use sky130_osu_sc_18T_hs__decap_1  decap36_0
timestamp 1607194151
transform 1 0 1614 0 -1 50156
box -9 0 199 1341
use sky130_osu_sc_18T_hs__fill_1  FILL_89
timestamp 1607194151
transform 1 0 1592 0 -1 50156
box 0 0 22 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_88
timestamp 1607194151
transform 1 0 1416 0 -1 50156
box 0 0 176 1332
use sky130_osu_sc_18T_hs__fill_16  FILL_87
timestamp 1607194151
transform 1 0 1064 0 -1 50156
box 0 0 352 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_142
timestamp 1607194151
transform 1 0 2296 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap36_1
timestamp 1607194151
transform 1 0 2098 0 -1 50156
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_1_0
timestamp 1607194151
transform 1 0 1812 0 -1 50156
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_143
timestamp 1607194151
transform 1 0 3000 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_144
timestamp 1607194151
transform 1 0 3704 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_145
timestamp 1607194151
transform 1 0 4408 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_146
timestamp 1607194151
transform 1 0 5112 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_147
timestamp 1607194151
transform 1 0 5816 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_148
timestamp 1607194151
transform 1 0 6520 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_149
timestamp 1607194151
transform 1 0 7224 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_150
timestamp 1607194151
transform 1 0 7928 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_151
timestamp 1607194151
transform 1 0 8632 0 -1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_2  FILL_153 $PDKPATH/libs.ref/sky130_osu_sc_18T_hs/mag
timestamp 1607194151
transform 1 0 9512 0 -1 50156
box 0 0 44 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_152
timestamp 1607194151
transform 1 0 9336 0 -1 50156
box 0 0 176 1332
use sky130_osu_sc_18T_hs__decap_1  decap37_0
timestamp 1607194151
transform 1 0 1614 0 1 50156
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_1
timestamp 1607194151
transform 1 0 1064 0 1 50156
box -9 0 553 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_154
timestamp 1607194151
transform 1 0 2296 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap37_1
timestamp 1607194151
transform 1 0 2098 0 1 50156
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_1_1
timestamp 1607194151
transform 1 0 1812 0 1 50156
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_155
timestamp 1607194151
transform 1 0 3000 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_156
timestamp 1607194151
transform 1 0 3704 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_157
timestamp 1607194151
transform 1 0 4408 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_158
timestamp 1607194151
transform 1 0 5112 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_159
timestamp 1607194151
transform 1 0 5816 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_160
timestamp 1607194151
transform 1 0 6520 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_161
timestamp 1607194151
transform 1 0 7224 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_162
timestamp 1607194151
transform 1 0 7928 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_163
timestamp 1607194151
transform 1 0 8632 0 1 50156
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_2  FILL_165
timestamp 1607194151
transform 1 0 9512 0 1 50156
box 0 0 44 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_164
timestamp 1607194151
transform 1 0 9336 0 1 50156
box 0 0 176 1332
use sky130_osu_sc_18T_hs__decap_1  decap38_0
timestamp 1607194151
transform 1 0 1614 0 -1 52820
box -9 0 199 1341
use sky130_osu_sc_18T_hs__mux2_1  mux_0
timestamp 1607194151
transform 1 0 1064 0 -1 52820
box -9 0 553 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_166
timestamp 1607194151
transform 1 0 2296 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__decap_1  decap38_1
timestamp 1607194151
transform 1 0 2098 0 -1 52820
box -9 0 199 1341
use sky130_osu_sc_18T_hs__buf_1  delay_0_0
timestamp 1607194151
transform 1 0 1812 0 -1 52820
box -9 0 288 1341
use sky130_osu_sc_18T_hs__fill_32  FILL_167
timestamp 1607194151
transform 1 0 3000 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_168
timestamp 1607194151
transform 1 0 3704 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_169
timestamp 1607194151
transform 1 0 4408 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_170
timestamp 1607194151
transform 1 0 5112 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_171
timestamp 1607194151
transform 1 0 5816 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_172
timestamp 1607194151
transform 1 0 6520 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_173
timestamp 1607194151
transform 1 0 7224 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_174
timestamp 1607194151
transform 1 0 7928 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_32  FILL_175
timestamp 1607194151
transform 1 0 8632 0 -1 52820
box 0 0 704 1332
use sky130_osu_sc_18T_hs__fill_2  FILL_177
timestamp 1607194151
transform 1 0 9512 0 -1 52820
box 0 0 44 1332
use sky130_osu_sc_18T_hs__fill_8  FILL_176
timestamp 1607194151
transform 1 0 9336 0 -1 52820
box 0 0 176 1332
<< labels >>
rlabel metal3 s 800 800 920 1056 6 inp_i
port 0 nsew default input
rlabel metal3 s 800 52752 920 53008 6 out_o
port 1 nsew default tristate
rlabel metal3 s 800 20792 920 21048 6 en_i[8]
port 2 nsew default input
rlabel metal3 s 800 31400 920 31656 6 en_i[7]
port 3 nsew default input
rlabel metal3 s 800 36704 920 36960 6 en_i[6]
port 4 nsew default input
rlabel metal3 s 800 39424 920 39680 6 en_i[5]
port 5 nsew default input
rlabel metal3 s 800 42008 920 42264 6 en_i[4]
port 6 nsew default input
rlabel metal3 s 800 44728 920 44984 6 en_i[3]
port 7 nsew default input
rlabel metal3 s 800 47312 920 47568 6 en_i[2]
port 8 nsew default input
rlabel metal3 s 800 50032 920 50288 6 en_i[1]
port 9 nsew default input
rlabel metal3 s 800 51392 920 51648 6 en_i[0]
port 10 nsew default input
rlabel metal5 s 1064 2504 9556 2824 6 VPWR
port 11 nsew default input
rlabel metal5 s 1064 20504 9556 20824 6 VGND
port 12 nsew default input
<< properties >>
string FIXED_BBOX 0 0 10357 53808
<< end >>
